module complete_bipartite_64_64 (
inout input_0,inout input_1,inout input_2,inout input_3,inout input_4,inout input_5,inout input_6,inout input_7,inout input_8,inout input_9,inout input_10,inout input_11,inout input_12,inout input_13,inout input_14,inout input_15,inout input_16,inout input_17,inout input_18,inout input_19,inout input_20,inout input_21,inout input_22,inout input_23,inout input_24,inout input_25,inout input_26,inout input_27,inout input_28,inout input_29,inout input_30,inout input_31,inout input_32,inout input_33,inout input_34,inout input_35,inout input_36,inout input_37,inout input_38,inout input_39,inout input_40,inout input_41,inout input_42,inout input_43,inout input_44,inout input_45,inout input_46,inout input_47,inout input_48,inout input_49,inout input_50,inout input_51,inout input_52,inout input_53,inout input_54,inout input_55,inout input_56,inout input_57,inout input_58,inout input_59,inout input_60,inout input_61,inout input_62,inout input_63,inout output_0,inout output_1,inout output_2,inout output_3,inout output_4,inout output_5,inout output_6,inout output_7,inout output_8,inout output_9,inout output_10,inout output_11,inout output_12,inout output_13,inout output_14,inout output_15,inout output_16,inout output_17,inout output_18,inout output_19,inout output_20,inout output_21,inout output_22,inout output_23,inout output_24,inout output_25,inout output_26,inout output_27,inout output_28,inout output_29,inout output_30,inout output_31,inout output_32,inout output_33,inout output_34,inout output_35,inout output_36,inout output_37,inout output_38,inout output_39,inout output_40,inout output_41,inout output_42,inout output_43,inout output_44,inout output_45,inout output_46,inout output_47,inout output_48,inout output_49,inout output_50,inout output_51,inout output_52,inout output_53,inout output_54,inout output_55,inout output_56,inout output_57,inout output_58,inout output_59,inout output_60,inout output_61,inout output_62,inout output_63
);
assign output_0 = input_0;
assign output_1 = input_0;
assign output_2 = input_0;
assign output_3 = input_0;
assign output_4 = input_0;
assign output_5 = input_0;
assign output_6 = input_0;
assign output_7 = input_0;
assign output_8 = input_0;
assign output_9 = input_0;
assign output_10 = input_0;
assign output_11 = input_0;
assign output_12 = input_0;
assign output_13 = input_0;
assign output_14 = input_0;
assign output_15 = input_0;
assign output_16 = input_0;
assign output_17 = input_0;
assign output_18 = input_0;
assign output_19 = input_0;
assign output_20 = input_0;
assign output_21 = input_0;
assign output_22 = input_0;
assign output_23 = input_0;
assign output_24 = input_0;
assign output_25 = input_0;
assign output_26 = input_0;
assign output_27 = input_0;
assign output_28 = input_0;
assign output_29 = input_0;
assign output_30 = input_0;
assign output_31 = input_0;
assign output_32 = input_0;
assign output_33 = input_0;
assign output_34 = input_0;
assign output_35 = input_0;
assign output_36 = input_0;
assign output_37 = input_0;
assign output_38 = input_0;
assign output_39 = input_0;
assign output_40 = input_0;
assign output_41 = input_0;
assign output_42 = input_0;
assign output_43 = input_0;
assign output_44 = input_0;
assign output_45 = input_0;
assign output_46 = input_0;
assign output_47 = input_0;
assign output_48 = input_0;
assign output_49 = input_0;
assign output_50 = input_0;
assign output_51 = input_0;
assign output_52 = input_0;
assign output_53 = input_0;
assign output_54 = input_0;
assign output_55 = input_0;
assign output_56 = input_0;
assign output_57 = input_0;
assign output_58 = input_0;
assign output_59 = input_0;
assign output_60 = input_0;
assign output_61 = input_0;
assign output_62 = input_0;
assign output_63 = input_0;
assign output_0 = input_1;
assign output_1 = input_1;
assign output_2 = input_1;
assign output_3 = input_1;
assign output_4 = input_1;
assign output_5 = input_1;
assign output_6 = input_1;
assign output_7 = input_1;
assign output_8 = input_1;
assign output_9 = input_1;
assign output_10 = input_1;
assign output_11 = input_1;
assign output_12 = input_1;
assign output_13 = input_1;
assign output_14 = input_1;
assign output_15 = input_1;
assign output_16 = input_1;
assign output_17 = input_1;
assign output_18 = input_1;
assign output_19 = input_1;
assign output_20 = input_1;
assign output_21 = input_1;
assign output_22 = input_1;
assign output_23 = input_1;
assign output_24 = input_1;
assign output_25 = input_1;
assign output_26 = input_1;
assign output_27 = input_1;
assign output_28 = input_1;
assign output_29 = input_1;
assign output_30 = input_1;
assign output_31 = input_1;
assign output_32 = input_1;
assign output_33 = input_1;
assign output_34 = input_1;
assign output_35 = input_1;
assign output_36 = input_1;
assign output_37 = input_1;
assign output_38 = input_1;
assign output_39 = input_1;
assign output_40 = input_1;
assign output_41 = input_1;
assign output_42 = input_1;
assign output_43 = input_1;
assign output_44 = input_1;
assign output_45 = input_1;
assign output_46 = input_1;
assign output_47 = input_1;
assign output_48 = input_1;
assign output_49 = input_1;
assign output_50 = input_1;
assign output_51 = input_1;
assign output_52 = input_1;
assign output_53 = input_1;
assign output_54 = input_1;
assign output_55 = input_1;
assign output_56 = input_1;
assign output_57 = input_1;
assign output_58 = input_1;
assign output_59 = input_1;
assign output_60 = input_1;
assign output_61 = input_1;
assign output_62 = input_1;
assign output_63 = input_1;
assign output_0 = input_2;
assign output_1 = input_2;
assign output_2 = input_2;
assign output_3 = input_2;
assign output_4 = input_2;
assign output_5 = input_2;
assign output_6 = input_2;
assign output_7 = input_2;
assign output_8 = input_2;
assign output_9 = input_2;
assign output_10 = input_2;
assign output_11 = input_2;
assign output_12 = input_2;
assign output_13 = input_2;
assign output_14 = input_2;
assign output_15 = input_2;
assign output_16 = input_2;
assign output_17 = input_2;
assign output_18 = input_2;
assign output_19 = input_2;
assign output_20 = input_2;
assign output_21 = input_2;
assign output_22 = input_2;
assign output_23 = input_2;
assign output_24 = input_2;
assign output_25 = input_2;
assign output_26 = input_2;
assign output_27 = input_2;
assign output_28 = input_2;
assign output_29 = input_2;
assign output_30 = input_2;
assign output_31 = input_2;
assign output_32 = input_2;
assign output_33 = input_2;
assign output_34 = input_2;
assign output_35 = input_2;
assign output_36 = input_2;
assign output_37 = input_2;
assign output_38 = input_2;
assign output_39 = input_2;
assign output_40 = input_2;
assign output_41 = input_2;
assign output_42 = input_2;
assign output_43 = input_2;
assign output_44 = input_2;
assign output_45 = input_2;
assign output_46 = input_2;
assign output_47 = input_2;
assign output_48 = input_2;
assign output_49 = input_2;
assign output_50 = input_2;
assign output_51 = input_2;
assign output_52 = input_2;
assign output_53 = input_2;
assign output_54 = input_2;
assign output_55 = input_2;
assign output_56 = input_2;
assign output_57 = input_2;
assign output_58 = input_2;
assign output_59 = input_2;
assign output_60 = input_2;
assign output_61 = input_2;
assign output_62 = input_2;
assign output_63 = input_2;
assign output_0 = input_3;
assign output_1 = input_3;
assign output_2 = input_3;
assign output_3 = input_3;
assign output_4 = input_3;
assign output_5 = input_3;
assign output_6 = input_3;
assign output_7 = input_3;
assign output_8 = input_3;
assign output_9 = input_3;
assign output_10 = input_3;
assign output_11 = input_3;
assign output_12 = input_3;
assign output_13 = input_3;
assign output_14 = input_3;
assign output_15 = input_3;
assign output_16 = input_3;
assign output_17 = input_3;
assign output_18 = input_3;
assign output_19 = input_3;
assign output_20 = input_3;
assign output_21 = input_3;
assign output_22 = input_3;
assign output_23 = input_3;
assign output_24 = input_3;
assign output_25 = input_3;
assign output_26 = input_3;
assign output_27 = input_3;
assign output_28 = input_3;
assign output_29 = input_3;
assign output_30 = input_3;
assign output_31 = input_3;
assign output_32 = input_3;
assign output_33 = input_3;
assign output_34 = input_3;
assign output_35 = input_3;
assign output_36 = input_3;
assign output_37 = input_3;
assign output_38 = input_3;
assign output_39 = input_3;
assign output_40 = input_3;
assign output_41 = input_3;
assign output_42 = input_3;
assign output_43 = input_3;
assign output_44 = input_3;
assign output_45 = input_3;
assign output_46 = input_3;
assign output_47 = input_3;
assign output_48 = input_3;
assign output_49 = input_3;
assign output_50 = input_3;
assign output_51 = input_3;
assign output_52 = input_3;
assign output_53 = input_3;
assign output_54 = input_3;
assign output_55 = input_3;
assign output_56 = input_3;
assign output_57 = input_3;
assign output_58 = input_3;
assign output_59 = input_3;
assign output_60 = input_3;
assign output_61 = input_3;
assign output_62 = input_3;
assign output_63 = input_3;
assign output_0 = input_4;
assign output_1 = input_4;
assign output_2 = input_4;
assign output_3 = input_4;
assign output_4 = input_4;
assign output_5 = input_4;
assign output_6 = input_4;
assign output_7 = input_4;
assign output_8 = input_4;
assign output_9 = input_4;
assign output_10 = input_4;
assign output_11 = input_4;
assign output_12 = input_4;
assign output_13 = input_4;
assign output_14 = input_4;
assign output_15 = input_4;
assign output_16 = input_4;
assign output_17 = input_4;
assign output_18 = input_4;
assign output_19 = input_4;
assign output_20 = input_4;
assign output_21 = input_4;
assign output_22 = input_4;
assign output_23 = input_4;
assign output_24 = input_4;
assign output_25 = input_4;
assign output_26 = input_4;
assign output_27 = input_4;
assign output_28 = input_4;
assign output_29 = input_4;
assign output_30 = input_4;
assign output_31 = input_4;
assign output_32 = input_4;
assign output_33 = input_4;
assign output_34 = input_4;
assign output_35 = input_4;
assign output_36 = input_4;
assign output_37 = input_4;
assign output_38 = input_4;
assign output_39 = input_4;
assign output_40 = input_4;
assign output_41 = input_4;
assign output_42 = input_4;
assign output_43 = input_4;
assign output_44 = input_4;
assign output_45 = input_4;
assign output_46 = input_4;
assign output_47 = input_4;
assign output_48 = input_4;
assign output_49 = input_4;
assign output_50 = input_4;
assign output_51 = input_4;
assign output_52 = input_4;
assign output_53 = input_4;
assign output_54 = input_4;
assign output_55 = input_4;
assign output_56 = input_4;
assign output_57 = input_4;
assign output_58 = input_4;
assign output_59 = input_4;
assign output_60 = input_4;
assign output_61 = input_4;
assign output_62 = input_4;
assign output_63 = input_4;
assign output_0 = input_5;
assign output_1 = input_5;
assign output_2 = input_5;
assign output_3 = input_5;
assign output_4 = input_5;
assign output_5 = input_5;
assign output_6 = input_5;
assign output_7 = input_5;
assign output_8 = input_5;
assign output_9 = input_5;
assign output_10 = input_5;
assign output_11 = input_5;
assign output_12 = input_5;
assign output_13 = input_5;
assign output_14 = input_5;
assign output_15 = input_5;
assign output_16 = input_5;
assign output_17 = input_5;
assign output_18 = input_5;
assign output_19 = input_5;
assign output_20 = input_5;
assign output_21 = input_5;
assign output_22 = input_5;
assign output_23 = input_5;
assign output_24 = input_5;
assign output_25 = input_5;
assign output_26 = input_5;
assign output_27 = input_5;
assign output_28 = input_5;
assign output_29 = input_5;
assign output_30 = input_5;
assign output_31 = input_5;
assign output_32 = input_5;
assign output_33 = input_5;
assign output_34 = input_5;
assign output_35 = input_5;
assign output_36 = input_5;
assign output_37 = input_5;
assign output_38 = input_5;
assign output_39 = input_5;
assign output_40 = input_5;
assign output_41 = input_5;
assign output_42 = input_5;
assign output_43 = input_5;
assign output_44 = input_5;
assign output_45 = input_5;
assign output_46 = input_5;
assign output_47 = input_5;
assign output_48 = input_5;
assign output_49 = input_5;
assign output_50 = input_5;
assign output_51 = input_5;
assign output_52 = input_5;
assign output_53 = input_5;
assign output_54 = input_5;
assign output_55 = input_5;
assign output_56 = input_5;
assign output_57 = input_5;
assign output_58 = input_5;
assign output_59 = input_5;
assign output_60 = input_5;
assign output_61 = input_5;
assign output_62 = input_5;
assign output_63 = input_5;
assign output_0 = input_6;
assign output_1 = input_6;
assign output_2 = input_6;
assign output_3 = input_6;
assign output_4 = input_6;
assign output_5 = input_6;
assign output_6 = input_6;
assign output_7 = input_6;
assign output_8 = input_6;
assign output_9 = input_6;
assign output_10 = input_6;
assign output_11 = input_6;
assign output_12 = input_6;
assign output_13 = input_6;
assign output_14 = input_6;
assign output_15 = input_6;
assign output_16 = input_6;
assign output_17 = input_6;
assign output_18 = input_6;
assign output_19 = input_6;
assign output_20 = input_6;
assign output_21 = input_6;
assign output_22 = input_6;
assign output_23 = input_6;
assign output_24 = input_6;
assign output_25 = input_6;
assign output_26 = input_6;
assign output_27 = input_6;
assign output_28 = input_6;
assign output_29 = input_6;
assign output_30 = input_6;
assign output_31 = input_6;
assign output_32 = input_6;
assign output_33 = input_6;
assign output_34 = input_6;
assign output_35 = input_6;
assign output_36 = input_6;
assign output_37 = input_6;
assign output_38 = input_6;
assign output_39 = input_6;
assign output_40 = input_6;
assign output_41 = input_6;
assign output_42 = input_6;
assign output_43 = input_6;
assign output_44 = input_6;
assign output_45 = input_6;
assign output_46 = input_6;
assign output_47 = input_6;
assign output_48 = input_6;
assign output_49 = input_6;
assign output_50 = input_6;
assign output_51 = input_6;
assign output_52 = input_6;
assign output_53 = input_6;
assign output_54 = input_6;
assign output_55 = input_6;
assign output_56 = input_6;
assign output_57 = input_6;
assign output_58 = input_6;
assign output_59 = input_6;
assign output_60 = input_6;
assign output_61 = input_6;
assign output_62 = input_6;
assign output_63 = input_6;
assign output_0 = input_7;
assign output_1 = input_7;
assign output_2 = input_7;
assign output_3 = input_7;
assign output_4 = input_7;
assign output_5 = input_7;
assign output_6 = input_7;
assign output_7 = input_7;
assign output_8 = input_7;
assign output_9 = input_7;
assign output_10 = input_7;
assign output_11 = input_7;
assign output_12 = input_7;
assign output_13 = input_7;
assign output_14 = input_7;
assign output_15 = input_7;
assign output_16 = input_7;
assign output_17 = input_7;
assign output_18 = input_7;
assign output_19 = input_7;
assign output_20 = input_7;
assign output_21 = input_7;
assign output_22 = input_7;
assign output_23 = input_7;
assign output_24 = input_7;
assign output_25 = input_7;
assign output_26 = input_7;
assign output_27 = input_7;
assign output_28 = input_7;
assign output_29 = input_7;
assign output_30 = input_7;
assign output_31 = input_7;
assign output_32 = input_7;
assign output_33 = input_7;
assign output_34 = input_7;
assign output_35 = input_7;
assign output_36 = input_7;
assign output_37 = input_7;
assign output_38 = input_7;
assign output_39 = input_7;
assign output_40 = input_7;
assign output_41 = input_7;
assign output_42 = input_7;
assign output_43 = input_7;
assign output_44 = input_7;
assign output_45 = input_7;
assign output_46 = input_7;
assign output_47 = input_7;
assign output_48 = input_7;
assign output_49 = input_7;
assign output_50 = input_7;
assign output_51 = input_7;
assign output_52 = input_7;
assign output_53 = input_7;
assign output_54 = input_7;
assign output_55 = input_7;
assign output_56 = input_7;
assign output_57 = input_7;
assign output_58 = input_7;
assign output_59 = input_7;
assign output_60 = input_7;
assign output_61 = input_7;
assign output_62 = input_7;
assign output_63 = input_7;
assign output_0 = input_8;
assign output_1 = input_8;
assign output_2 = input_8;
assign output_3 = input_8;
assign output_4 = input_8;
assign output_5 = input_8;
assign output_6 = input_8;
assign output_7 = input_8;
assign output_8 = input_8;
assign output_9 = input_8;
assign output_10 = input_8;
assign output_11 = input_8;
assign output_12 = input_8;
assign output_13 = input_8;
assign output_14 = input_8;
assign output_15 = input_8;
assign output_16 = input_8;
assign output_17 = input_8;
assign output_18 = input_8;
assign output_19 = input_8;
assign output_20 = input_8;
assign output_21 = input_8;
assign output_22 = input_8;
assign output_23 = input_8;
assign output_24 = input_8;
assign output_25 = input_8;
assign output_26 = input_8;
assign output_27 = input_8;
assign output_28 = input_8;
assign output_29 = input_8;
assign output_30 = input_8;
assign output_31 = input_8;
assign output_32 = input_8;
assign output_33 = input_8;
assign output_34 = input_8;
assign output_35 = input_8;
assign output_36 = input_8;
assign output_37 = input_8;
assign output_38 = input_8;
assign output_39 = input_8;
assign output_40 = input_8;
assign output_41 = input_8;
assign output_42 = input_8;
assign output_43 = input_8;
assign output_44 = input_8;
assign output_45 = input_8;
assign output_46 = input_8;
assign output_47 = input_8;
assign output_48 = input_8;
assign output_49 = input_8;
assign output_50 = input_8;
assign output_51 = input_8;
assign output_52 = input_8;
assign output_53 = input_8;
assign output_54 = input_8;
assign output_55 = input_8;
assign output_56 = input_8;
assign output_57 = input_8;
assign output_58 = input_8;
assign output_59 = input_8;
assign output_60 = input_8;
assign output_61 = input_8;
assign output_62 = input_8;
assign output_63 = input_8;
assign output_0 = input_9;
assign output_1 = input_9;
assign output_2 = input_9;
assign output_3 = input_9;
assign output_4 = input_9;
assign output_5 = input_9;
assign output_6 = input_9;
assign output_7 = input_9;
assign output_8 = input_9;
assign output_9 = input_9;
assign output_10 = input_9;
assign output_11 = input_9;
assign output_12 = input_9;
assign output_13 = input_9;
assign output_14 = input_9;
assign output_15 = input_9;
assign output_16 = input_9;
assign output_17 = input_9;
assign output_18 = input_9;
assign output_19 = input_9;
assign output_20 = input_9;
assign output_21 = input_9;
assign output_22 = input_9;
assign output_23 = input_9;
assign output_24 = input_9;
assign output_25 = input_9;
assign output_26 = input_9;
assign output_27 = input_9;
assign output_28 = input_9;
assign output_29 = input_9;
assign output_30 = input_9;
assign output_31 = input_9;
assign output_32 = input_9;
assign output_33 = input_9;
assign output_34 = input_9;
assign output_35 = input_9;
assign output_36 = input_9;
assign output_37 = input_9;
assign output_38 = input_9;
assign output_39 = input_9;
assign output_40 = input_9;
assign output_41 = input_9;
assign output_42 = input_9;
assign output_43 = input_9;
assign output_44 = input_9;
assign output_45 = input_9;
assign output_46 = input_9;
assign output_47 = input_9;
assign output_48 = input_9;
assign output_49 = input_9;
assign output_50 = input_9;
assign output_51 = input_9;
assign output_52 = input_9;
assign output_53 = input_9;
assign output_54 = input_9;
assign output_55 = input_9;
assign output_56 = input_9;
assign output_57 = input_9;
assign output_58 = input_9;
assign output_59 = input_9;
assign output_60 = input_9;
assign output_61 = input_9;
assign output_62 = input_9;
assign output_63 = input_9;
assign output_0 = input_10;
assign output_1 = input_10;
assign output_2 = input_10;
assign output_3 = input_10;
assign output_4 = input_10;
assign output_5 = input_10;
assign output_6 = input_10;
assign output_7 = input_10;
assign output_8 = input_10;
assign output_9 = input_10;
assign output_10 = input_10;
assign output_11 = input_10;
assign output_12 = input_10;
assign output_13 = input_10;
assign output_14 = input_10;
assign output_15 = input_10;
assign output_16 = input_10;
assign output_17 = input_10;
assign output_18 = input_10;
assign output_19 = input_10;
assign output_20 = input_10;
assign output_21 = input_10;
assign output_22 = input_10;
assign output_23 = input_10;
assign output_24 = input_10;
assign output_25 = input_10;
assign output_26 = input_10;
assign output_27 = input_10;
assign output_28 = input_10;
assign output_29 = input_10;
assign output_30 = input_10;
assign output_31 = input_10;
assign output_32 = input_10;
assign output_33 = input_10;
assign output_34 = input_10;
assign output_35 = input_10;
assign output_36 = input_10;
assign output_37 = input_10;
assign output_38 = input_10;
assign output_39 = input_10;
assign output_40 = input_10;
assign output_41 = input_10;
assign output_42 = input_10;
assign output_43 = input_10;
assign output_44 = input_10;
assign output_45 = input_10;
assign output_46 = input_10;
assign output_47 = input_10;
assign output_48 = input_10;
assign output_49 = input_10;
assign output_50 = input_10;
assign output_51 = input_10;
assign output_52 = input_10;
assign output_53 = input_10;
assign output_54 = input_10;
assign output_55 = input_10;
assign output_56 = input_10;
assign output_57 = input_10;
assign output_58 = input_10;
assign output_59 = input_10;
assign output_60 = input_10;
assign output_61 = input_10;
assign output_62 = input_10;
assign output_63 = input_10;
assign output_0 = input_11;
assign output_1 = input_11;
assign output_2 = input_11;
assign output_3 = input_11;
assign output_4 = input_11;
assign output_5 = input_11;
assign output_6 = input_11;
assign output_7 = input_11;
assign output_8 = input_11;
assign output_9 = input_11;
assign output_10 = input_11;
assign output_11 = input_11;
assign output_12 = input_11;
assign output_13 = input_11;
assign output_14 = input_11;
assign output_15 = input_11;
assign output_16 = input_11;
assign output_17 = input_11;
assign output_18 = input_11;
assign output_19 = input_11;
assign output_20 = input_11;
assign output_21 = input_11;
assign output_22 = input_11;
assign output_23 = input_11;
assign output_24 = input_11;
assign output_25 = input_11;
assign output_26 = input_11;
assign output_27 = input_11;
assign output_28 = input_11;
assign output_29 = input_11;
assign output_30 = input_11;
assign output_31 = input_11;
assign output_32 = input_11;
assign output_33 = input_11;
assign output_34 = input_11;
assign output_35 = input_11;
assign output_36 = input_11;
assign output_37 = input_11;
assign output_38 = input_11;
assign output_39 = input_11;
assign output_40 = input_11;
assign output_41 = input_11;
assign output_42 = input_11;
assign output_43 = input_11;
assign output_44 = input_11;
assign output_45 = input_11;
assign output_46 = input_11;
assign output_47 = input_11;
assign output_48 = input_11;
assign output_49 = input_11;
assign output_50 = input_11;
assign output_51 = input_11;
assign output_52 = input_11;
assign output_53 = input_11;
assign output_54 = input_11;
assign output_55 = input_11;
assign output_56 = input_11;
assign output_57 = input_11;
assign output_58 = input_11;
assign output_59 = input_11;
assign output_60 = input_11;
assign output_61 = input_11;
assign output_62 = input_11;
assign output_63 = input_11;
assign output_0 = input_12;
assign output_1 = input_12;
assign output_2 = input_12;
assign output_3 = input_12;
assign output_4 = input_12;
assign output_5 = input_12;
assign output_6 = input_12;
assign output_7 = input_12;
assign output_8 = input_12;
assign output_9 = input_12;
assign output_10 = input_12;
assign output_11 = input_12;
assign output_12 = input_12;
assign output_13 = input_12;
assign output_14 = input_12;
assign output_15 = input_12;
assign output_16 = input_12;
assign output_17 = input_12;
assign output_18 = input_12;
assign output_19 = input_12;
assign output_20 = input_12;
assign output_21 = input_12;
assign output_22 = input_12;
assign output_23 = input_12;
assign output_24 = input_12;
assign output_25 = input_12;
assign output_26 = input_12;
assign output_27 = input_12;
assign output_28 = input_12;
assign output_29 = input_12;
assign output_30 = input_12;
assign output_31 = input_12;
assign output_32 = input_12;
assign output_33 = input_12;
assign output_34 = input_12;
assign output_35 = input_12;
assign output_36 = input_12;
assign output_37 = input_12;
assign output_38 = input_12;
assign output_39 = input_12;
assign output_40 = input_12;
assign output_41 = input_12;
assign output_42 = input_12;
assign output_43 = input_12;
assign output_44 = input_12;
assign output_45 = input_12;
assign output_46 = input_12;
assign output_47 = input_12;
assign output_48 = input_12;
assign output_49 = input_12;
assign output_50 = input_12;
assign output_51 = input_12;
assign output_52 = input_12;
assign output_53 = input_12;
assign output_54 = input_12;
assign output_55 = input_12;
assign output_56 = input_12;
assign output_57 = input_12;
assign output_58 = input_12;
assign output_59 = input_12;
assign output_60 = input_12;
assign output_61 = input_12;
assign output_62 = input_12;
assign output_63 = input_12;
assign output_0 = input_13;
assign output_1 = input_13;
assign output_2 = input_13;
assign output_3 = input_13;
assign output_4 = input_13;
assign output_5 = input_13;
assign output_6 = input_13;
assign output_7 = input_13;
assign output_8 = input_13;
assign output_9 = input_13;
assign output_10 = input_13;
assign output_11 = input_13;
assign output_12 = input_13;
assign output_13 = input_13;
assign output_14 = input_13;
assign output_15 = input_13;
assign output_16 = input_13;
assign output_17 = input_13;
assign output_18 = input_13;
assign output_19 = input_13;
assign output_20 = input_13;
assign output_21 = input_13;
assign output_22 = input_13;
assign output_23 = input_13;
assign output_24 = input_13;
assign output_25 = input_13;
assign output_26 = input_13;
assign output_27 = input_13;
assign output_28 = input_13;
assign output_29 = input_13;
assign output_30 = input_13;
assign output_31 = input_13;
assign output_32 = input_13;
assign output_33 = input_13;
assign output_34 = input_13;
assign output_35 = input_13;
assign output_36 = input_13;
assign output_37 = input_13;
assign output_38 = input_13;
assign output_39 = input_13;
assign output_40 = input_13;
assign output_41 = input_13;
assign output_42 = input_13;
assign output_43 = input_13;
assign output_44 = input_13;
assign output_45 = input_13;
assign output_46 = input_13;
assign output_47 = input_13;
assign output_48 = input_13;
assign output_49 = input_13;
assign output_50 = input_13;
assign output_51 = input_13;
assign output_52 = input_13;
assign output_53 = input_13;
assign output_54 = input_13;
assign output_55 = input_13;
assign output_56 = input_13;
assign output_57 = input_13;
assign output_58 = input_13;
assign output_59 = input_13;
assign output_60 = input_13;
assign output_61 = input_13;
assign output_62 = input_13;
assign output_63 = input_13;
assign output_0 = input_14;
assign output_1 = input_14;
assign output_2 = input_14;
assign output_3 = input_14;
assign output_4 = input_14;
assign output_5 = input_14;
assign output_6 = input_14;
assign output_7 = input_14;
assign output_8 = input_14;
assign output_9 = input_14;
assign output_10 = input_14;
assign output_11 = input_14;
assign output_12 = input_14;
assign output_13 = input_14;
assign output_14 = input_14;
assign output_15 = input_14;
assign output_16 = input_14;
assign output_17 = input_14;
assign output_18 = input_14;
assign output_19 = input_14;
assign output_20 = input_14;
assign output_21 = input_14;
assign output_22 = input_14;
assign output_23 = input_14;
assign output_24 = input_14;
assign output_25 = input_14;
assign output_26 = input_14;
assign output_27 = input_14;
assign output_28 = input_14;
assign output_29 = input_14;
assign output_30 = input_14;
assign output_31 = input_14;
assign output_32 = input_14;
assign output_33 = input_14;
assign output_34 = input_14;
assign output_35 = input_14;
assign output_36 = input_14;
assign output_37 = input_14;
assign output_38 = input_14;
assign output_39 = input_14;
assign output_40 = input_14;
assign output_41 = input_14;
assign output_42 = input_14;
assign output_43 = input_14;
assign output_44 = input_14;
assign output_45 = input_14;
assign output_46 = input_14;
assign output_47 = input_14;
assign output_48 = input_14;
assign output_49 = input_14;
assign output_50 = input_14;
assign output_51 = input_14;
assign output_52 = input_14;
assign output_53 = input_14;
assign output_54 = input_14;
assign output_55 = input_14;
assign output_56 = input_14;
assign output_57 = input_14;
assign output_58 = input_14;
assign output_59 = input_14;
assign output_60 = input_14;
assign output_61 = input_14;
assign output_62 = input_14;
assign output_63 = input_14;
assign output_0 = input_15;
assign output_1 = input_15;
assign output_2 = input_15;
assign output_3 = input_15;
assign output_4 = input_15;
assign output_5 = input_15;
assign output_6 = input_15;
assign output_7 = input_15;
assign output_8 = input_15;
assign output_9 = input_15;
assign output_10 = input_15;
assign output_11 = input_15;
assign output_12 = input_15;
assign output_13 = input_15;
assign output_14 = input_15;
assign output_15 = input_15;
assign output_16 = input_15;
assign output_17 = input_15;
assign output_18 = input_15;
assign output_19 = input_15;
assign output_20 = input_15;
assign output_21 = input_15;
assign output_22 = input_15;
assign output_23 = input_15;
assign output_24 = input_15;
assign output_25 = input_15;
assign output_26 = input_15;
assign output_27 = input_15;
assign output_28 = input_15;
assign output_29 = input_15;
assign output_30 = input_15;
assign output_31 = input_15;
assign output_32 = input_15;
assign output_33 = input_15;
assign output_34 = input_15;
assign output_35 = input_15;
assign output_36 = input_15;
assign output_37 = input_15;
assign output_38 = input_15;
assign output_39 = input_15;
assign output_40 = input_15;
assign output_41 = input_15;
assign output_42 = input_15;
assign output_43 = input_15;
assign output_44 = input_15;
assign output_45 = input_15;
assign output_46 = input_15;
assign output_47 = input_15;
assign output_48 = input_15;
assign output_49 = input_15;
assign output_50 = input_15;
assign output_51 = input_15;
assign output_52 = input_15;
assign output_53 = input_15;
assign output_54 = input_15;
assign output_55 = input_15;
assign output_56 = input_15;
assign output_57 = input_15;
assign output_58 = input_15;
assign output_59 = input_15;
assign output_60 = input_15;
assign output_61 = input_15;
assign output_62 = input_15;
assign output_63 = input_15;
assign output_0 = input_16;
assign output_1 = input_16;
assign output_2 = input_16;
assign output_3 = input_16;
assign output_4 = input_16;
assign output_5 = input_16;
assign output_6 = input_16;
assign output_7 = input_16;
assign output_8 = input_16;
assign output_9 = input_16;
assign output_10 = input_16;
assign output_11 = input_16;
assign output_12 = input_16;
assign output_13 = input_16;
assign output_14 = input_16;
assign output_15 = input_16;
assign output_16 = input_16;
assign output_17 = input_16;
assign output_18 = input_16;
assign output_19 = input_16;
assign output_20 = input_16;
assign output_21 = input_16;
assign output_22 = input_16;
assign output_23 = input_16;
assign output_24 = input_16;
assign output_25 = input_16;
assign output_26 = input_16;
assign output_27 = input_16;
assign output_28 = input_16;
assign output_29 = input_16;
assign output_30 = input_16;
assign output_31 = input_16;
assign output_32 = input_16;
assign output_33 = input_16;
assign output_34 = input_16;
assign output_35 = input_16;
assign output_36 = input_16;
assign output_37 = input_16;
assign output_38 = input_16;
assign output_39 = input_16;
assign output_40 = input_16;
assign output_41 = input_16;
assign output_42 = input_16;
assign output_43 = input_16;
assign output_44 = input_16;
assign output_45 = input_16;
assign output_46 = input_16;
assign output_47 = input_16;
assign output_48 = input_16;
assign output_49 = input_16;
assign output_50 = input_16;
assign output_51 = input_16;
assign output_52 = input_16;
assign output_53 = input_16;
assign output_54 = input_16;
assign output_55 = input_16;
assign output_56 = input_16;
assign output_57 = input_16;
assign output_58 = input_16;
assign output_59 = input_16;
assign output_60 = input_16;
assign output_61 = input_16;
assign output_62 = input_16;
assign output_63 = input_16;
assign output_0 = input_17;
assign output_1 = input_17;
assign output_2 = input_17;
assign output_3 = input_17;
assign output_4 = input_17;
assign output_5 = input_17;
assign output_6 = input_17;
assign output_7 = input_17;
assign output_8 = input_17;
assign output_9 = input_17;
assign output_10 = input_17;
assign output_11 = input_17;
assign output_12 = input_17;
assign output_13 = input_17;
assign output_14 = input_17;
assign output_15 = input_17;
assign output_16 = input_17;
assign output_17 = input_17;
assign output_18 = input_17;
assign output_19 = input_17;
assign output_20 = input_17;
assign output_21 = input_17;
assign output_22 = input_17;
assign output_23 = input_17;
assign output_24 = input_17;
assign output_25 = input_17;
assign output_26 = input_17;
assign output_27 = input_17;
assign output_28 = input_17;
assign output_29 = input_17;
assign output_30 = input_17;
assign output_31 = input_17;
assign output_32 = input_17;
assign output_33 = input_17;
assign output_34 = input_17;
assign output_35 = input_17;
assign output_36 = input_17;
assign output_37 = input_17;
assign output_38 = input_17;
assign output_39 = input_17;
assign output_40 = input_17;
assign output_41 = input_17;
assign output_42 = input_17;
assign output_43 = input_17;
assign output_44 = input_17;
assign output_45 = input_17;
assign output_46 = input_17;
assign output_47 = input_17;
assign output_48 = input_17;
assign output_49 = input_17;
assign output_50 = input_17;
assign output_51 = input_17;
assign output_52 = input_17;
assign output_53 = input_17;
assign output_54 = input_17;
assign output_55 = input_17;
assign output_56 = input_17;
assign output_57 = input_17;
assign output_58 = input_17;
assign output_59 = input_17;
assign output_60 = input_17;
assign output_61 = input_17;
assign output_62 = input_17;
assign output_63 = input_17;
assign output_0 = input_18;
assign output_1 = input_18;
assign output_2 = input_18;
assign output_3 = input_18;
assign output_4 = input_18;
assign output_5 = input_18;
assign output_6 = input_18;
assign output_7 = input_18;
assign output_8 = input_18;
assign output_9 = input_18;
assign output_10 = input_18;
assign output_11 = input_18;
assign output_12 = input_18;
assign output_13 = input_18;
assign output_14 = input_18;
assign output_15 = input_18;
assign output_16 = input_18;
assign output_17 = input_18;
assign output_18 = input_18;
assign output_19 = input_18;
assign output_20 = input_18;
assign output_21 = input_18;
assign output_22 = input_18;
assign output_23 = input_18;
assign output_24 = input_18;
assign output_25 = input_18;
assign output_26 = input_18;
assign output_27 = input_18;
assign output_28 = input_18;
assign output_29 = input_18;
assign output_30 = input_18;
assign output_31 = input_18;
assign output_32 = input_18;
assign output_33 = input_18;
assign output_34 = input_18;
assign output_35 = input_18;
assign output_36 = input_18;
assign output_37 = input_18;
assign output_38 = input_18;
assign output_39 = input_18;
assign output_40 = input_18;
assign output_41 = input_18;
assign output_42 = input_18;
assign output_43 = input_18;
assign output_44 = input_18;
assign output_45 = input_18;
assign output_46 = input_18;
assign output_47 = input_18;
assign output_48 = input_18;
assign output_49 = input_18;
assign output_50 = input_18;
assign output_51 = input_18;
assign output_52 = input_18;
assign output_53 = input_18;
assign output_54 = input_18;
assign output_55 = input_18;
assign output_56 = input_18;
assign output_57 = input_18;
assign output_58 = input_18;
assign output_59 = input_18;
assign output_60 = input_18;
assign output_61 = input_18;
assign output_62 = input_18;
assign output_63 = input_18;
assign output_0 = input_19;
assign output_1 = input_19;
assign output_2 = input_19;
assign output_3 = input_19;
assign output_4 = input_19;
assign output_5 = input_19;
assign output_6 = input_19;
assign output_7 = input_19;
assign output_8 = input_19;
assign output_9 = input_19;
assign output_10 = input_19;
assign output_11 = input_19;
assign output_12 = input_19;
assign output_13 = input_19;
assign output_14 = input_19;
assign output_15 = input_19;
assign output_16 = input_19;
assign output_17 = input_19;
assign output_18 = input_19;
assign output_19 = input_19;
assign output_20 = input_19;
assign output_21 = input_19;
assign output_22 = input_19;
assign output_23 = input_19;
assign output_24 = input_19;
assign output_25 = input_19;
assign output_26 = input_19;
assign output_27 = input_19;
assign output_28 = input_19;
assign output_29 = input_19;
assign output_30 = input_19;
assign output_31 = input_19;
assign output_32 = input_19;
assign output_33 = input_19;
assign output_34 = input_19;
assign output_35 = input_19;
assign output_36 = input_19;
assign output_37 = input_19;
assign output_38 = input_19;
assign output_39 = input_19;
assign output_40 = input_19;
assign output_41 = input_19;
assign output_42 = input_19;
assign output_43 = input_19;
assign output_44 = input_19;
assign output_45 = input_19;
assign output_46 = input_19;
assign output_47 = input_19;
assign output_48 = input_19;
assign output_49 = input_19;
assign output_50 = input_19;
assign output_51 = input_19;
assign output_52 = input_19;
assign output_53 = input_19;
assign output_54 = input_19;
assign output_55 = input_19;
assign output_56 = input_19;
assign output_57 = input_19;
assign output_58 = input_19;
assign output_59 = input_19;
assign output_60 = input_19;
assign output_61 = input_19;
assign output_62 = input_19;
assign output_63 = input_19;
assign output_0 = input_20;
assign output_1 = input_20;
assign output_2 = input_20;
assign output_3 = input_20;
assign output_4 = input_20;
assign output_5 = input_20;
assign output_6 = input_20;
assign output_7 = input_20;
assign output_8 = input_20;
assign output_9 = input_20;
assign output_10 = input_20;
assign output_11 = input_20;
assign output_12 = input_20;
assign output_13 = input_20;
assign output_14 = input_20;
assign output_15 = input_20;
assign output_16 = input_20;
assign output_17 = input_20;
assign output_18 = input_20;
assign output_19 = input_20;
assign output_20 = input_20;
assign output_21 = input_20;
assign output_22 = input_20;
assign output_23 = input_20;
assign output_24 = input_20;
assign output_25 = input_20;
assign output_26 = input_20;
assign output_27 = input_20;
assign output_28 = input_20;
assign output_29 = input_20;
assign output_30 = input_20;
assign output_31 = input_20;
assign output_32 = input_20;
assign output_33 = input_20;
assign output_34 = input_20;
assign output_35 = input_20;
assign output_36 = input_20;
assign output_37 = input_20;
assign output_38 = input_20;
assign output_39 = input_20;
assign output_40 = input_20;
assign output_41 = input_20;
assign output_42 = input_20;
assign output_43 = input_20;
assign output_44 = input_20;
assign output_45 = input_20;
assign output_46 = input_20;
assign output_47 = input_20;
assign output_48 = input_20;
assign output_49 = input_20;
assign output_50 = input_20;
assign output_51 = input_20;
assign output_52 = input_20;
assign output_53 = input_20;
assign output_54 = input_20;
assign output_55 = input_20;
assign output_56 = input_20;
assign output_57 = input_20;
assign output_58 = input_20;
assign output_59 = input_20;
assign output_60 = input_20;
assign output_61 = input_20;
assign output_62 = input_20;
assign output_63 = input_20;
assign output_0 = input_21;
assign output_1 = input_21;
assign output_2 = input_21;
assign output_3 = input_21;
assign output_4 = input_21;
assign output_5 = input_21;
assign output_6 = input_21;
assign output_7 = input_21;
assign output_8 = input_21;
assign output_9 = input_21;
assign output_10 = input_21;
assign output_11 = input_21;
assign output_12 = input_21;
assign output_13 = input_21;
assign output_14 = input_21;
assign output_15 = input_21;
assign output_16 = input_21;
assign output_17 = input_21;
assign output_18 = input_21;
assign output_19 = input_21;
assign output_20 = input_21;
assign output_21 = input_21;
assign output_22 = input_21;
assign output_23 = input_21;
assign output_24 = input_21;
assign output_25 = input_21;
assign output_26 = input_21;
assign output_27 = input_21;
assign output_28 = input_21;
assign output_29 = input_21;
assign output_30 = input_21;
assign output_31 = input_21;
assign output_32 = input_21;
assign output_33 = input_21;
assign output_34 = input_21;
assign output_35 = input_21;
assign output_36 = input_21;
assign output_37 = input_21;
assign output_38 = input_21;
assign output_39 = input_21;
assign output_40 = input_21;
assign output_41 = input_21;
assign output_42 = input_21;
assign output_43 = input_21;
assign output_44 = input_21;
assign output_45 = input_21;
assign output_46 = input_21;
assign output_47 = input_21;
assign output_48 = input_21;
assign output_49 = input_21;
assign output_50 = input_21;
assign output_51 = input_21;
assign output_52 = input_21;
assign output_53 = input_21;
assign output_54 = input_21;
assign output_55 = input_21;
assign output_56 = input_21;
assign output_57 = input_21;
assign output_58 = input_21;
assign output_59 = input_21;
assign output_60 = input_21;
assign output_61 = input_21;
assign output_62 = input_21;
assign output_63 = input_21;
assign output_0 = input_22;
assign output_1 = input_22;
assign output_2 = input_22;
assign output_3 = input_22;
assign output_4 = input_22;
assign output_5 = input_22;
assign output_6 = input_22;
assign output_7 = input_22;
assign output_8 = input_22;
assign output_9 = input_22;
assign output_10 = input_22;
assign output_11 = input_22;
assign output_12 = input_22;
assign output_13 = input_22;
assign output_14 = input_22;
assign output_15 = input_22;
assign output_16 = input_22;
assign output_17 = input_22;
assign output_18 = input_22;
assign output_19 = input_22;
assign output_20 = input_22;
assign output_21 = input_22;
assign output_22 = input_22;
assign output_23 = input_22;
assign output_24 = input_22;
assign output_25 = input_22;
assign output_26 = input_22;
assign output_27 = input_22;
assign output_28 = input_22;
assign output_29 = input_22;
assign output_30 = input_22;
assign output_31 = input_22;
assign output_32 = input_22;
assign output_33 = input_22;
assign output_34 = input_22;
assign output_35 = input_22;
assign output_36 = input_22;
assign output_37 = input_22;
assign output_38 = input_22;
assign output_39 = input_22;
assign output_40 = input_22;
assign output_41 = input_22;
assign output_42 = input_22;
assign output_43 = input_22;
assign output_44 = input_22;
assign output_45 = input_22;
assign output_46 = input_22;
assign output_47 = input_22;
assign output_48 = input_22;
assign output_49 = input_22;
assign output_50 = input_22;
assign output_51 = input_22;
assign output_52 = input_22;
assign output_53 = input_22;
assign output_54 = input_22;
assign output_55 = input_22;
assign output_56 = input_22;
assign output_57 = input_22;
assign output_58 = input_22;
assign output_59 = input_22;
assign output_60 = input_22;
assign output_61 = input_22;
assign output_62 = input_22;
assign output_63 = input_22;
assign output_0 = input_23;
assign output_1 = input_23;
assign output_2 = input_23;
assign output_3 = input_23;
assign output_4 = input_23;
assign output_5 = input_23;
assign output_6 = input_23;
assign output_7 = input_23;
assign output_8 = input_23;
assign output_9 = input_23;
assign output_10 = input_23;
assign output_11 = input_23;
assign output_12 = input_23;
assign output_13 = input_23;
assign output_14 = input_23;
assign output_15 = input_23;
assign output_16 = input_23;
assign output_17 = input_23;
assign output_18 = input_23;
assign output_19 = input_23;
assign output_20 = input_23;
assign output_21 = input_23;
assign output_22 = input_23;
assign output_23 = input_23;
assign output_24 = input_23;
assign output_25 = input_23;
assign output_26 = input_23;
assign output_27 = input_23;
assign output_28 = input_23;
assign output_29 = input_23;
assign output_30 = input_23;
assign output_31 = input_23;
assign output_32 = input_23;
assign output_33 = input_23;
assign output_34 = input_23;
assign output_35 = input_23;
assign output_36 = input_23;
assign output_37 = input_23;
assign output_38 = input_23;
assign output_39 = input_23;
assign output_40 = input_23;
assign output_41 = input_23;
assign output_42 = input_23;
assign output_43 = input_23;
assign output_44 = input_23;
assign output_45 = input_23;
assign output_46 = input_23;
assign output_47 = input_23;
assign output_48 = input_23;
assign output_49 = input_23;
assign output_50 = input_23;
assign output_51 = input_23;
assign output_52 = input_23;
assign output_53 = input_23;
assign output_54 = input_23;
assign output_55 = input_23;
assign output_56 = input_23;
assign output_57 = input_23;
assign output_58 = input_23;
assign output_59 = input_23;
assign output_60 = input_23;
assign output_61 = input_23;
assign output_62 = input_23;
assign output_63 = input_23;
assign output_0 = input_24;
assign output_1 = input_24;
assign output_2 = input_24;
assign output_3 = input_24;
assign output_4 = input_24;
assign output_5 = input_24;
assign output_6 = input_24;
assign output_7 = input_24;
assign output_8 = input_24;
assign output_9 = input_24;
assign output_10 = input_24;
assign output_11 = input_24;
assign output_12 = input_24;
assign output_13 = input_24;
assign output_14 = input_24;
assign output_15 = input_24;
assign output_16 = input_24;
assign output_17 = input_24;
assign output_18 = input_24;
assign output_19 = input_24;
assign output_20 = input_24;
assign output_21 = input_24;
assign output_22 = input_24;
assign output_23 = input_24;
assign output_24 = input_24;
assign output_25 = input_24;
assign output_26 = input_24;
assign output_27 = input_24;
assign output_28 = input_24;
assign output_29 = input_24;
assign output_30 = input_24;
assign output_31 = input_24;
assign output_32 = input_24;
assign output_33 = input_24;
assign output_34 = input_24;
assign output_35 = input_24;
assign output_36 = input_24;
assign output_37 = input_24;
assign output_38 = input_24;
assign output_39 = input_24;
assign output_40 = input_24;
assign output_41 = input_24;
assign output_42 = input_24;
assign output_43 = input_24;
assign output_44 = input_24;
assign output_45 = input_24;
assign output_46 = input_24;
assign output_47 = input_24;
assign output_48 = input_24;
assign output_49 = input_24;
assign output_50 = input_24;
assign output_51 = input_24;
assign output_52 = input_24;
assign output_53 = input_24;
assign output_54 = input_24;
assign output_55 = input_24;
assign output_56 = input_24;
assign output_57 = input_24;
assign output_58 = input_24;
assign output_59 = input_24;
assign output_60 = input_24;
assign output_61 = input_24;
assign output_62 = input_24;
assign output_63 = input_24;
assign output_0 = input_25;
assign output_1 = input_25;
assign output_2 = input_25;
assign output_3 = input_25;
assign output_4 = input_25;
assign output_5 = input_25;
assign output_6 = input_25;
assign output_7 = input_25;
assign output_8 = input_25;
assign output_9 = input_25;
assign output_10 = input_25;
assign output_11 = input_25;
assign output_12 = input_25;
assign output_13 = input_25;
assign output_14 = input_25;
assign output_15 = input_25;
assign output_16 = input_25;
assign output_17 = input_25;
assign output_18 = input_25;
assign output_19 = input_25;
assign output_20 = input_25;
assign output_21 = input_25;
assign output_22 = input_25;
assign output_23 = input_25;
assign output_24 = input_25;
assign output_25 = input_25;
assign output_26 = input_25;
assign output_27 = input_25;
assign output_28 = input_25;
assign output_29 = input_25;
assign output_30 = input_25;
assign output_31 = input_25;
assign output_32 = input_25;
assign output_33 = input_25;
assign output_34 = input_25;
assign output_35 = input_25;
assign output_36 = input_25;
assign output_37 = input_25;
assign output_38 = input_25;
assign output_39 = input_25;
assign output_40 = input_25;
assign output_41 = input_25;
assign output_42 = input_25;
assign output_43 = input_25;
assign output_44 = input_25;
assign output_45 = input_25;
assign output_46 = input_25;
assign output_47 = input_25;
assign output_48 = input_25;
assign output_49 = input_25;
assign output_50 = input_25;
assign output_51 = input_25;
assign output_52 = input_25;
assign output_53 = input_25;
assign output_54 = input_25;
assign output_55 = input_25;
assign output_56 = input_25;
assign output_57 = input_25;
assign output_58 = input_25;
assign output_59 = input_25;
assign output_60 = input_25;
assign output_61 = input_25;
assign output_62 = input_25;
assign output_63 = input_25;
assign output_0 = input_26;
assign output_1 = input_26;
assign output_2 = input_26;
assign output_3 = input_26;
assign output_4 = input_26;
assign output_5 = input_26;
assign output_6 = input_26;
assign output_7 = input_26;
assign output_8 = input_26;
assign output_9 = input_26;
assign output_10 = input_26;
assign output_11 = input_26;
assign output_12 = input_26;
assign output_13 = input_26;
assign output_14 = input_26;
assign output_15 = input_26;
assign output_16 = input_26;
assign output_17 = input_26;
assign output_18 = input_26;
assign output_19 = input_26;
assign output_20 = input_26;
assign output_21 = input_26;
assign output_22 = input_26;
assign output_23 = input_26;
assign output_24 = input_26;
assign output_25 = input_26;
assign output_26 = input_26;
assign output_27 = input_26;
assign output_28 = input_26;
assign output_29 = input_26;
assign output_30 = input_26;
assign output_31 = input_26;
assign output_32 = input_26;
assign output_33 = input_26;
assign output_34 = input_26;
assign output_35 = input_26;
assign output_36 = input_26;
assign output_37 = input_26;
assign output_38 = input_26;
assign output_39 = input_26;
assign output_40 = input_26;
assign output_41 = input_26;
assign output_42 = input_26;
assign output_43 = input_26;
assign output_44 = input_26;
assign output_45 = input_26;
assign output_46 = input_26;
assign output_47 = input_26;
assign output_48 = input_26;
assign output_49 = input_26;
assign output_50 = input_26;
assign output_51 = input_26;
assign output_52 = input_26;
assign output_53 = input_26;
assign output_54 = input_26;
assign output_55 = input_26;
assign output_56 = input_26;
assign output_57 = input_26;
assign output_58 = input_26;
assign output_59 = input_26;
assign output_60 = input_26;
assign output_61 = input_26;
assign output_62 = input_26;
assign output_63 = input_26;
assign output_0 = input_27;
assign output_1 = input_27;
assign output_2 = input_27;
assign output_3 = input_27;
assign output_4 = input_27;
assign output_5 = input_27;
assign output_6 = input_27;
assign output_7 = input_27;
assign output_8 = input_27;
assign output_9 = input_27;
assign output_10 = input_27;
assign output_11 = input_27;
assign output_12 = input_27;
assign output_13 = input_27;
assign output_14 = input_27;
assign output_15 = input_27;
assign output_16 = input_27;
assign output_17 = input_27;
assign output_18 = input_27;
assign output_19 = input_27;
assign output_20 = input_27;
assign output_21 = input_27;
assign output_22 = input_27;
assign output_23 = input_27;
assign output_24 = input_27;
assign output_25 = input_27;
assign output_26 = input_27;
assign output_27 = input_27;
assign output_28 = input_27;
assign output_29 = input_27;
assign output_30 = input_27;
assign output_31 = input_27;
assign output_32 = input_27;
assign output_33 = input_27;
assign output_34 = input_27;
assign output_35 = input_27;
assign output_36 = input_27;
assign output_37 = input_27;
assign output_38 = input_27;
assign output_39 = input_27;
assign output_40 = input_27;
assign output_41 = input_27;
assign output_42 = input_27;
assign output_43 = input_27;
assign output_44 = input_27;
assign output_45 = input_27;
assign output_46 = input_27;
assign output_47 = input_27;
assign output_48 = input_27;
assign output_49 = input_27;
assign output_50 = input_27;
assign output_51 = input_27;
assign output_52 = input_27;
assign output_53 = input_27;
assign output_54 = input_27;
assign output_55 = input_27;
assign output_56 = input_27;
assign output_57 = input_27;
assign output_58 = input_27;
assign output_59 = input_27;
assign output_60 = input_27;
assign output_61 = input_27;
assign output_62 = input_27;
assign output_63 = input_27;
assign output_0 = input_28;
assign output_1 = input_28;
assign output_2 = input_28;
assign output_3 = input_28;
assign output_4 = input_28;
assign output_5 = input_28;
assign output_6 = input_28;
assign output_7 = input_28;
assign output_8 = input_28;
assign output_9 = input_28;
assign output_10 = input_28;
assign output_11 = input_28;
assign output_12 = input_28;
assign output_13 = input_28;
assign output_14 = input_28;
assign output_15 = input_28;
assign output_16 = input_28;
assign output_17 = input_28;
assign output_18 = input_28;
assign output_19 = input_28;
assign output_20 = input_28;
assign output_21 = input_28;
assign output_22 = input_28;
assign output_23 = input_28;
assign output_24 = input_28;
assign output_25 = input_28;
assign output_26 = input_28;
assign output_27 = input_28;
assign output_28 = input_28;
assign output_29 = input_28;
assign output_30 = input_28;
assign output_31 = input_28;
assign output_32 = input_28;
assign output_33 = input_28;
assign output_34 = input_28;
assign output_35 = input_28;
assign output_36 = input_28;
assign output_37 = input_28;
assign output_38 = input_28;
assign output_39 = input_28;
assign output_40 = input_28;
assign output_41 = input_28;
assign output_42 = input_28;
assign output_43 = input_28;
assign output_44 = input_28;
assign output_45 = input_28;
assign output_46 = input_28;
assign output_47 = input_28;
assign output_48 = input_28;
assign output_49 = input_28;
assign output_50 = input_28;
assign output_51 = input_28;
assign output_52 = input_28;
assign output_53 = input_28;
assign output_54 = input_28;
assign output_55 = input_28;
assign output_56 = input_28;
assign output_57 = input_28;
assign output_58 = input_28;
assign output_59 = input_28;
assign output_60 = input_28;
assign output_61 = input_28;
assign output_62 = input_28;
assign output_63 = input_28;
assign output_0 = input_29;
assign output_1 = input_29;
assign output_2 = input_29;
assign output_3 = input_29;
assign output_4 = input_29;
assign output_5 = input_29;
assign output_6 = input_29;
assign output_7 = input_29;
assign output_8 = input_29;
assign output_9 = input_29;
assign output_10 = input_29;
assign output_11 = input_29;
assign output_12 = input_29;
assign output_13 = input_29;
assign output_14 = input_29;
assign output_15 = input_29;
assign output_16 = input_29;
assign output_17 = input_29;
assign output_18 = input_29;
assign output_19 = input_29;
assign output_20 = input_29;
assign output_21 = input_29;
assign output_22 = input_29;
assign output_23 = input_29;
assign output_24 = input_29;
assign output_25 = input_29;
assign output_26 = input_29;
assign output_27 = input_29;
assign output_28 = input_29;
assign output_29 = input_29;
assign output_30 = input_29;
assign output_31 = input_29;
assign output_32 = input_29;
assign output_33 = input_29;
assign output_34 = input_29;
assign output_35 = input_29;
assign output_36 = input_29;
assign output_37 = input_29;
assign output_38 = input_29;
assign output_39 = input_29;
assign output_40 = input_29;
assign output_41 = input_29;
assign output_42 = input_29;
assign output_43 = input_29;
assign output_44 = input_29;
assign output_45 = input_29;
assign output_46 = input_29;
assign output_47 = input_29;
assign output_48 = input_29;
assign output_49 = input_29;
assign output_50 = input_29;
assign output_51 = input_29;
assign output_52 = input_29;
assign output_53 = input_29;
assign output_54 = input_29;
assign output_55 = input_29;
assign output_56 = input_29;
assign output_57 = input_29;
assign output_58 = input_29;
assign output_59 = input_29;
assign output_60 = input_29;
assign output_61 = input_29;
assign output_62 = input_29;
assign output_63 = input_29;
assign output_0 = input_30;
assign output_1 = input_30;
assign output_2 = input_30;
assign output_3 = input_30;
assign output_4 = input_30;
assign output_5 = input_30;
assign output_6 = input_30;
assign output_7 = input_30;
assign output_8 = input_30;
assign output_9 = input_30;
assign output_10 = input_30;
assign output_11 = input_30;
assign output_12 = input_30;
assign output_13 = input_30;
assign output_14 = input_30;
assign output_15 = input_30;
assign output_16 = input_30;
assign output_17 = input_30;
assign output_18 = input_30;
assign output_19 = input_30;
assign output_20 = input_30;
assign output_21 = input_30;
assign output_22 = input_30;
assign output_23 = input_30;
assign output_24 = input_30;
assign output_25 = input_30;
assign output_26 = input_30;
assign output_27 = input_30;
assign output_28 = input_30;
assign output_29 = input_30;
assign output_30 = input_30;
assign output_31 = input_30;
assign output_32 = input_30;
assign output_33 = input_30;
assign output_34 = input_30;
assign output_35 = input_30;
assign output_36 = input_30;
assign output_37 = input_30;
assign output_38 = input_30;
assign output_39 = input_30;
assign output_40 = input_30;
assign output_41 = input_30;
assign output_42 = input_30;
assign output_43 = input_30;
assign output_44 = input_30;
assign output_45 = input_30;
assign output_46 = input_30;
assign output_47 = input_30;
assign output_48 = input_30;
assign output_49 = input_30;
assign output_50 = input_30;
assign output_51 = input_30;
assign output_52 = input_30;
assign output_53 = input_30;
assign output_54 = input_30;
assign output_55 = input_30;
assign output_56 = input_30;
assign output_57 = input_30;
assign output_58 = input_30;
assign output_59 = input_30;
assign output_60 = input_30;
assign output_61 = input_30;
assign output_62 = input_30;
assign output_63 = input_30;
assign output_0 = input_31;
assign output_1 = input_31;
assign output_2 = input_31;
assign output_3 = input_31;
assign output_4 = input_31;
assign output_5 = input_31;
assign output_6 = input_31;
assign output_7 = input_31;
assign output_8 = input_31;
assign output_9 = input_31;
assign output_10 = input_31;
assign output_11 = input_31;
assign output_12 = input_31;
assign output_13 = input_31;
assign output_14 = input_31;
assign output_15 = input_31;
assign output_16 = input_31;
assign output_17 = input_31;
assign output_18 = input_31;
assign output_19 = input_31;
assign output_20 = input_31;
assign output_21 = input_31;
assign output_22 = input_31;
assign output_23 = input_31;
assign output_24 = input_31;
assign output_25 = input_31;
assign output_26 = input_31;
assign output_27 = input_31;
assign output_28 = input_31;
assign output_29 = input_31;
assign output_30 = input_31;
assign output_31 = input_31;
assign output_32 = input_31;
assign output_33 = input_31;
assign output_34 = input_31;
assign output_35 = input_31;
assign output_36 = input_31;
assign output_37 = input_31;
assign output_38 = input_31;
assign output_39 = input_31;
assign output_40 = input_31;
assign output_41 = input_31;
assign output_42 = input_31;
assign output_43 = input_31;
assign output_44 = input_31;
assign output_45 = input_31;
assign output_46 = input_31;
assign output_47 = input_31;
assign output_48 = input_31;
assign output_49 = input_31;
assign output_50 = input_31;
assign output_51 = input_31;
assign output_52 = input_31;
assign output_53 = input_31;
assign output_54 = input_31;
assign output_55 = input_31;
assign output_56 = input_31;
assign output_57 = input_31;
assign output_58 = input_31;
assign output_59 = input_31;
assign output_60 = input_31;
assign output_61 = input_31;
assign output_62 = input_31;
assign output_63 = input_31;
assign output_0 = input_32;
assign output_1 = input_32;
assign output_2 = input_32;
assign output_3 = input_32;
assign output_4 = input_32;
assign output_5 = input_32;
assign output_6 = input_32;
assign output_7 = input_32;
assign output_8 = input_32;
assign output_9 = input_32;
assign output_10 = input_32;
assign output_11 = input_32;
assign output_12 = input_32;
assign output_13 = input_32;
assign output_14 = input_32;
assign output_15 = input_32;
assign output_16 = input_32;
assign output_17 = input_32;
assign output_18 = input_32;
assign output_19 = input_32;
assign output_20 = input_32;
assign output_21 = input_32;
assign output_22 = input_32;
assign output_23 = input_32;
assign output_24 = input_32;
assign output_25 = input_32;
assign output_26 = input_32;
assign output_27 = input_32;
assign output_28 = input_32;
assign output_29 = input_32;
assign output_30 = input_32;
assign output_31 = input_32;
assign output_32 = input_32;
assign output_33 = input_32;
assign output_34 = input_32;
assign output_35 = input_32;
assign output_36 = input_32;
assign output_37 = input_32;
assign output_38 = input_32;
assign output_39 = input_32;
assign output_40 = input_32;
assign output_41 = input_32;
assign output_42 = input_32;
assign output_43 = input_32;
assign output_44 = input_32;
assign output_45 = input_32;
assign output_46 = input_32;
assign output_47 = input_32;
assign output_48 = input_32;
assign output_49 = input_32;
assign output_50 = input_32;
assign output_51 = input_32;
assign output_52 = input_32;
assign output_53 = input_32;
assign output_54 = input_32;
assign output_55 = input_32;
assign output_56 = input_32;
assign output_57 = input_32;
assign output_58 = input_32;
assign output_59 = input_32;
assign output_60 = input_32;
assign output_61 = input_32;
assign output_62 = input_32;
assign output_63 = input_32;
assign output_0 = input_33;
assign output_1 = input_33;
assign output_2 = input_33;
assign output_3 = input_33;
assign output_4 = input_33;
assign output_5 = input_33;
assign output_6 = input_33;
assign output_7 = input_33;
assign output_8 = input_33;
assign output_9 = input_33;
assign output_10 = input_33;
assign output_11 = input_33;
assign output_12 = input_33;
assign output_13 = input_33;
assign output_14 = input_33;
assign output_15 = input_33;
assign output_16 = input_33;
assign output_17 = input_33;
assign output_18 = input_33;
assign output_19 = input_33;
assign output_20 = input_33;
assign output_21 = input_33;
assign output_22 = input_33;
assign output_23 = input_33;
assign output_24 = input_33;
assign output_25 = input_33;
assign output_26 = input_33;
assign output_27 = input_33;
assign output_28 = input_33;
assign output_29 = input_33;
assign output_30 = input_33;
assign output_31 = input_33;
assign output_32 = input_33;
assign output_33 = input_33;
assign output_34 = input_33;
assign output_35 = input_33;
assign output_36 = input_33;
assign output_37 = input_33;
assign output_38 = input_33;
assign output_39 = input_33;
assign output_40 = input_33;
assign output_41 = input_33;
assign output_42 = input_33;
assign output_43 = input_33;
assign output_44 = input_33;
assign output_45 = input_33;
assign output_46 = input_33;
assign output_47 = input_33;
assign output_48 = input_33;
assign output_49 = input_33;
assign output_50 = input_33;
assign output_51 = input_33;
assign output_52 = input_33;
assign output_53 = input_33;
assign output_54 = input_33;
assign output_55 = input_33;
assign output_56 = input_33;
assign output_57 = input_33;
assign output_58 = input_33;
assign output_59 = input_33;
assign output_60 = input_33;
assign output_61 = input_33;
assign output_62 = input_33;
assign output_63 = input_33;
assign output_0 = input_34;
assign output_1 = input_34;
assign output_2 = input_34;
assign output_3 = input_34;
assign output_4 = input_34;
assign output_5 = input_34;
assign output_6 = input_34;
assign output_7 = input_34;
assign output_8 = input_34;
assign output_9 = input_34;
assign output_10 = input_34;
assign output_11 = input_34;
assign output_12 = input_34;
assign output_13 = input_34;
assign output_14 = input_34;
assign output_15 = input_34;
assign output_16 = input_34;
assign output_17 = input_34;
assign output_18 = input_34;
assign output_19 = input_34;
assign output_20 = input_34;
assign output_21 = input_34;
assign output_22 = input_34;
assign output_23 = input_34;
assign output_24 = input_34;
assign output_25 = input_34;
assign output_26 = input_34;
assign output_27 = input_34;
assign output_28 = input_34;
assign output_29 = input_34;
assign output_30 = input_34;
assign output_31 = input_34;
assign output_32 = input_34;
assign output_33 = input_34;
assign output_34 = input_34;
assign output_35 = input_34;
assign output_36 = input_34;
assign output_37 = input_34;
assign output_38 = input_34;
assign output_39 = input_34;
assign output_40 = input_34;
assign output_41 = input_34;
assign output_42 = input_34;
assign output_43 = input_34;
assign output_44 = input_34;
assign output_45 = input_34;
assign output_46 = input_34;
assign output_47 = input_34;
assign output_48 = input_34;
assign output_49 = input_34;
assign output_50 = input_34;
assign output_51 = input_34;
assign output_52 = input_34;
assign output_53 = input_34;
assign output_54 = input_34;
assign output_55 = input_34;
assign output_56 = input_34;
assign output_57 = input_34;
assign output_58 = input_34;
assign output_59 = input_34;
assign output_60 = input_34;
assign output_61 = input_34;
assign output_62 = input_34;
assign output_63 = input_34;
assign output_0 = input_35;
assign output_1 = input_35;
assign output_2 = input_35;
assign output_3 = input_35;
assign output_4 = input_35;
assign output_5 = input_35;
assign output_6 = input_35;
assign output_7 = input_35;
assign output_8 = input_35;
assign output_9 = input_35;
assign output_10 = input_35;
assign output_11 = input_35;
assign output_12 = input_35;
assign output_13 = input_35;
assign output_14 = input_35;
assign output_15 = input_35;
assign output_16 = input_35;
assign output_17 = input_35;
assign output_18 = input_35;
assign output_19 = input_35;
assign output_20 = input_35;
assign output_21 = input_35;
assign output_22 = input_35;
assign output_23 = input_35;
assign output_24 = input_35;
assign output_25 = input_35;
assign output_26 = input_35;
assign output_27 = input_35;
assign output_28 = input_35;
assign output_29 = input_35;
assign output_30 = input_35;
assign output_31 = input_35;
assign output_32 = input_35;
assign output_33 = input_35;
assign output_34 = input_35;
assign output_35 = input_35;
assign output_36 = input_35;
assign output_37 = input_35;
assign output_38 = input_35;
assign output_39 = input_35;
assign output_40 = input_35;
assign output_41 = input_35;
assign output_42 = input_35;
assign output_43 = input_35;
assign output_44 = input_35;
assign output_45 = input_35;
assign output_46 = input_35;
assign output_47 = input_35;
assign output_48 = input_35;
assign output_49 = input_35;
assign output_50 = input_35;
assign output_51 = input_35;
assign output_52 = input_35;
assign output_53 = input_35;
assign output_54 = input_35;
assign output_55 = input_35;
assign output_56 = input_35;
assign output_57 = input_35;
assign output_58 = input_35;
assign output_59 = input_35;
assign output_60 = input_35;
assign output_61 = input_35;
assign output_62 = input_35;
assign output_63 = input_35;
assign output_0 = input_36;
assign output_1 = input_36;
assign output_2 = input_36;
assign output_3 = input_36;
assign output_4 = input_36;
assign output_5 = input_36;
assign output_6 = input_36;
assign output_7 = input_36;
assign output_8 = input_36;
assign output_9 = input_36;
assign output_10 = input_36;
assign output_11 = input_36;
assign output_12 = input_36;
assign output_13 = input_36;
assign output_14 = input_36;
assign output_15 = input_36;
assign output_16 = input_36;
assign output_17 = input_36;
assign output_18 = input_36;
assign output_19 = input_36;
assign output_20 = input_36;
assign output_21 = input_36;
assign output_22 = input_36;
assign output_23 = input_36;
assign output_24 = input_36;
assign output_25 = input_36;
assign output_26 = input_36;
assign output_27 = input_36;
assign output_28 = input_36;
assign output_29 = input_36;
assign output_30 = input_36;
assign output_31 = input_36;
assign output_32 = input_36;
assign output_33 = input_36;
assign output_34 = input_36;
assign output_35 = input_36;
assign output_36 = input_36;
assign output_37 = input_36;
assign output_38 = input_36;
assign output_39 = input_36;
assign output_40 = input_36;
assign output_41 = input_36;
assign output_42 = input_36;
assign output_43 = input_36;
assign output_44 = input_36;
assign output_45 = input_36;
assign output_46 = input_36;
assign output_47 = input_36;
assign output_48 = input_36;
assign output_49 = input_36;
assign output_50 = input_36;
assign output_51 = input_36;
assign output_52 = input_36;
assign output_53 = input_36;
assign output_54 = input_36;
assign output_55 = input_36;
assign output_56 = input_36;
assign output_57 = input_36;
assign output_58 = input_36;
assign output_59 = input_36;
assign output_60 = input_36;
assign output_61 = input_36;
assign output_62 = input_36;
assign output_63 = input_36;
assign output_0 = input_37;
assign output_1 = input_37;
assign output_2 = input_37;
assign output_3 = input_37;
assign output_4 = input_37;
assign output_5 = input_37;
assign output_6 = input_37;
assign output_7 = input_37;
assign output_8 = input_37;
assign output_9 = input_37;
assign output_10 = input_37;
assign output_11 = input_37;
assign output_12 = input_37;
assign output_13 = input_37;
assign output_14 = input_37;
assign output_15 = input_37;
assign output_16 = input_37;
assign output_17 = input_37;
assign output_18 = input_37;
assign output_19 = input_37;
assign output_20 = input_37;
assign output_21 = input_37;
assign output_22 = input_37;
assign output_23 = input_37;
assign output_24 = input_37;
assign output_25 = input_37;
assign output_26 = input_37;
assign output_27 = input_37;
assign output_28 = input_37;
assign output_29 = input_37;
assign output_30 = input_37;
assign output_31 = input_37;
assign output_32 = input_37;
assign output_33 = input_37;
assign output_34 = input_37;
assign output_35 = input_37;
assign output_36 = input_37;
assign output_37 = input_37;
assign output_38 = input_37;
assign output_39 = input_37;
assign output_40 = input_37;
assign output_41 = input_37;
assign output_42 = input_37;
assign output_43 = input_37;
assign output_44 = input_37;
assign output_45 = input_37;
assign output_46 = input_37;
assign output_47 = input_37;
assign output_48 = input_37;
assign output_49 = input_37;
assign output_50 = input_37;
assign output_51 = input_37;
assign output_52 = input_37;
assign output_53 = input_37;
assign output_54 = input_37;
assign output_55 = input_37;
assign output_56 = input_37;
assign output_57 = input_37;
assign output_58 = input_37;
assign output_59 = input_37;
assign output_60 = input_37;
assign output_61 = input_37;
assign output_62 = input_37;
assign output_63 = input_37;
assign output_0 = input_38;
assign output_1 = input_38;
assign output_2 = input_38;
assign output_3 = input_38;
assign output_4 = input_38;
assign output_5 = input_38;
assign output_6 = input_38;
assign output_7 = input_38;
assign output_8 = input_38;
assign output_9 = input_38;
assign output_10 = input_38;
assign output_11 = input_38;
assign output_12 = input_38;
assign output_13 = input_38;
assign output_14 = input_38;
assign output_15 = input_38;
assign output_16 = input_38;
assign output_17 = input_38;
assign output_18 = input_38;
assign output_19 = input_38;
assign output_20 = input_38;
assign output_21 = input_38;
assign output_22 = input_38;
assign output_23 = input_38;
assign output_24 = input_38;
assign output_25 = input_38;
assign output_26 = input_38;
assign output_27 = input_38;
assign output_28 = input_38;
assign output_29 = input_38;
assign output_30 = input_38;
assign output_31 = input_38;
assign output_32 = input_38;
assign output_33 = input_38;
assign output_34 = input_38;
assign output_35 = input_38;
assign output_36 = input_38;
assign output_37 = input_38;
assign output_38 = input_38;
assign output_39 = input_38;
assign output_40 = input_38;
assign output_41 = input_38;
assign output_42 = input_38;
assign output_43 = input_38;
assign output_44 = input_38;
assign output_45 = input_38;
assign output_46 = input_38;
assign output_47 = input_38;
assign output_48 = input_38;
assign output_49 = input_38;
assign output_50 = input_38;
assign output_51 = input_38;
assign output_52 = input_38;
assign output_53 = input_38;
assign output_54 = input_38;
assign output_55 = input_38;
assign output_56 = input_38;
assign output_57 = input_38;
assign output_58 = input_38;
assign output_59 = input_38;
assign output_60 = input_38;
assign output_61 = input_38;
assign output_62 = input_38;
assign output_63 = input_38;
assign output_0 = input_39;
assign output_1 = input_39;
assign output_2 = input_39;
assign output_3 = input_39;
assign output_4 = input_39;
assign output_5 = input_39;
assign output_6 = input_39;
assign output_7 = input_39;
assign output_8 = input_39;
assign output_9 = input_39;
assign output_10 = input_39;
assign output_11 = input_39;
assign output_12 = input_39;
assign output_13 = input_39;
assign output_14 = input_39;
assign output_15 = input_39;
assign output_16 = input_39;
assign output_17 = input_39;
assign output_18 = input_39;
assign output_19 = input_39;
assign output_20 = input_39;
assign output_21 = input_39;
assign output_22 = input_39;
assign output_23 = input_39;
assign output_24 = input_39;
assign output_25 = input_39;
assign output_26 = input_39;
assign output_27 = input_39;
assign output_28 = input_39;
assign output_29 = input_39;
assign output_30 = input_39;
assign output_31 = input_39;
assign output_32 = input_39;
assign output_33 = input_39;
assign output_34 = input_39;
assign output_35 = input_39;
assign output_36 = input_39;
assign output_37 = input_39;
assign output_38 = input_39;
assign output_39 = input_39;
assign output_40 = input_39;
assign output_41 = input_39;
assign output_42 = input_39;
assign output_43 = input_39;
assign output_44 = input_39;
assign output_45 = input_39;
assign output_46 = input_39;
assign output_47 = input_39;
assign output_48 = input_39;
assign output_49 = input_39;
assign output_50 = input_39;
assign output_51 = input_39;
assign output_52 = input_39;
assign output_53 = input_39;
assign output_54 = input_39;
assign output_55 = input_39;
assign output_56 = input_39;
assign output_57 = input_39;
assign output_58 = input_39;
assign output_59 = input_39;
assign output_60 = input_39;
assign output_61 = input_39;
assign output_62 = input_39;
assign output_63 = input_39;
assign output_0 = input_40;
assign output_1 = input_40;
assign output_2 = input_40;
assign output_3 = input_40;
assign output_4 = input_40;
assign output_5 = input_40;
assign output_6 = input_40;
assign output_7 = input_40;
assign output_8 = input_40;
assign output_9 = input_40;
assign output_10 = input_40;
assign output_11 = input_40;
assign output_12 = input_40;
assign output_13 = input_40;
assign output_14 = input_40;
assign output_15 = input_40;
assign output_16 = input_40;
assign output_17 = input_40;
assign output_18 = input_40;
assign output_19 = input_40;
assign output_20 = input_40;
assign output_21 = input_40;
assign output_22 = input_40;
assign output_23 = input_40;
assign output_24 = input_40;
assign output_25 = input_40;
assign output_26 = input_40;
assign output_27 = input_40;
assign output_28 = input_40;
assign output_29 = input_40;
assign output_30 = input_40;
assign output_31 = input_40;
assign output_32 = input_40;
assign output_33 = input_40;
assign output_34 = input_40;
assign output_35 = input_40;
assign output_36 = input_40;
assign output_37 = input_40;
assign output_38 = input_40;
assign output_39 = input_40;
assign output_40 = input_40;
assign output_41 = input_40;
assign output_42 = input_40;
assign output_43 = input_40;
assign output_44 = input_40;
assign output_45 = input_40;
assign output_46 = input_40;
assign output_47 = input_40;
assign output_48 = input_40;
assign output_49 = input_40;
assign output_50 = input_40;
assign output_51 = input_40;
assign output_52 = input_40;
assign output_53 = input_40;
assign output_54 = input_40;
assign output_55 = input_40;
assign output_56 = input_40;
assign output_57 = input_40;
assign output_58 = input_40;
assign output_59 = input_40;
assign output_60 = input_40;
assign output_61 = input_40;
assign output_62 = input_40;
assign output_63 = input_40;
assign output_0 = input_41;
assign output_1 = input_41;
assign output_2 = input_41;
assign output_3 = input_41;
assign output_4 = input_41;
assign output_5 = input_41;
assign output_6 = input_41;
assign output_7 = input_41;
assign output_8 = input_41;
assign output_9 = input_41;
assign output_10 = input_41;
assign output_11 = input_41;
assign output_12 = input_41;
assign output_13 = input_41;
assign output_14 = input_41;
assign output_15 = input_41;
assign output_16 = input_41;
assign output_17 = input_41;
assign output_18 = input_41;
assign output_19 = input_41;
assign output_20 = input_41;
assign output_21 = input_41;
assign output_22 = input_41;
assign output_23 = input_41;
assign output_24 = input_41;
assign output_25 = input_41;
assign output_26 = input_41;
assign output_27 = input_41;
assign output_28 = input_41;
assign output_29 = input_41;
assign output_30 = input_41;
assign output_31 = input_41;
assign output_32 = input_41;
assign output_33 = input_41;
assign output_34 = input_41;
assign output_35 = input_41;
assign output_36 = input_41;
assign output_37 = input_41;
assign output_38 = input_41;
assign output_39 = input_41;
assign output_40 = input_41;
assign output_41 = input_41;
assign output_42 = input_41;
assign output_43 = input_41;
assign output_44 = input_41;
assign output_45 = input_41;
assign output_46 = input_41;
assign output_47 = input_41;
assign output_48 = input_41;
assign output_49 = input_41;
assign output_50 = input_41;
assign output_51 = input_41;
assign output_52 = input_41;
assign output_53 = input_41;
assign output_54 = input_41;
assign output_55 = input_41;
assign output_56 = input_41;
assign output_57 = input_41;
assign output_58 = input_41;
assign output_59 = input_41;
assign output_60 = input_41;
assign output_61 = input_41;
assign output_62 = input_41;
assign output_63 = input_41;
assign output_0 = input_42;
assign output_1 = input_42;
assign output_2 = input_42;
assign output_3 = input_42;
assign output_4 = input_42;
assign output_5 = input_42;
assign output_6 = input_42;
assign output_7 = input_42;
assign output_8 = input_42;
assign output_9 = input_42;
assign output_10 = input_42;
assign output_11 = input_42;
assign output_12 = input_42;
assign output_13 = input_42;
assign output_14 = input_42;
assign output_15 = input_42;
assign output_16 = input_42;
assign output_17 = input_42;
assign output_18 = input_42;
assign output_19 = input_42;
assign output_20 = input_42;
assign output_21 = input_42;
assign output_22 = input_42;
assign output_23 = input_42;
assign output_24 = input_42;
assign output_25 = input_42;
assign output_26 = input_42;
assign output_27 = input_42;
assign output_28 = input_42;
assign output_29 = input_42;
assign output_30 = input_42;
assign output_31 = input_42;
assign output_32 = input_42;
assign output_33 = input_42;
assign output_34 = input_42;
assign output_35 = input_42;
assign output_36 = input_42;
assign output_37 = input_42;
assign output_38 = input_42;
assign output_39 = input_42;
assign output_40 = input_42;
assign output_41 = input_42;
assign output_42 = input_42;
assign output_43 = input_42;
assign output_44 = input_42;
assign output_45 = input_42;
assign output_46 = input_42;
assign output_47 = input_42;
assign output_48 = input_42;
assign output_49 = input_42;
assign output_50 = input_42;
assign output_51 = input_42;
assign output_52 = input_42;
assign output_53 = input_42;
assign output_54 = input_42;
assign output_55 = input_42;
assign output_56 = input_42;
assign output_57 = input_42;
assign output_58 = input_42;
assign output_59 = input_42;
assign output_60 = input_42;
assign output_61 = input_42;
assign output_62 = input_42;
assign output_63 = input_42;
assign output_0 = input_43;
assign output_1 = input_43;
assign output_2 = input_43;
assign output_3 = input_43;
assign output_4 = input_43;
assign output_5 = input_43;
assign output_6 = input_43;
assign output_7 = input_43;
assign output_8 = input_43;
assign output_9 = input_43;
assign output_10 = input_43;
assign output_11 = input_43;
assign output_12 = input_43;
assign output_13 = input_43;
assign output_14 = input_43;
assign output_15 = input_43;
assign output_16 = input_43;
assign output_17 = input_43;
assign output_18 = input_43;
assign output_19 = input_43;
assign output_20 = input_43;
assign output_21 = input_43;
assign output_22 = input_43;
assign output_23 = input_43;
assign output_24 = input_43;
assign output_25 = input_43;
assign output_26 = input_43;
assign output_27 = input_43;
assign output_28 = input_43;
assign output_29 = input_43;
assign output_30 = input_43;
assign output_31 = input_43;
assign output_32 = input_43;
assign output_33 = input_43;
assign output_34 = input_43;
assign output_35 = input_43;
assign output_36 = input_43;
assign output_37 = input_43;
assign output_38 = input_43;
assign output_39 = input_43;
assign output_40 = input_43;
assign output_41 = input_43;
assign output_42 = input_43;
assign output_43 = input_43;
assign output_44 = input_43;
assign output_45 = input_43;
assign output_46 = input_43;
assign output_47 = input_43;
assign output_48 = input_43;
assign output_49 = input_43;
assign output_50 = input_43;
assign output_51 = input_43;
assign output_52 = input_43;
assign output_53 = input_43;
assign output_54 = input_43;
assign output_55 = input_43;
assign output_56 = input_43;
assign output_57 = input_43;
assign output_58 = input_43;
assign output_59 = input_43;
assign output_60 = input_43;
assign output_61 = input_43;
assign output_62 = input_43;
assign output_63 = input_43;
assign output_0 = input_44;
assign output_1 = input_44;
assign output_2 = input_44;
assign output_3 = input_44;
assign output_4 = input_44;
assign output_5 = input_44;
assign output_6 = input_44;
assign output_7 = input_44;
assign output_8 = input_44;
assign output_9 = input_44;
assign output_10 = input_44;
assign output_11 = input_44;
assign output_12 = input_44;
assign output_13 = input_44;
assign output_14 = input_44;
assign output_15 = input_44;
assign output_16 = input_44;
assign output_17 = input_44;
assign output_18 = input_44;
assign output_19 = input_44;
assign output_20 = input_44;
assign output_21 = input_44;
assign output_22 = input_44;
assign output_23 = input_44;
assign output_24 = input_44;
assign output_25 = input_44;
assign output_26 = input_44;
assign output_27 = input_44;
assign output_28 = input_44;
assign output_29 = input_44;
assign output_30 = input_44;
assign output_31 = input_44;
assign output_32 = input_44;
assign output_33 = input_44;
assign output_34 = input_44;
assign output_35 = input_44;
assign output_36 = input_44;
assign output_37 = input_44;
assign output_38 = input_44;
assign output_39 = input_44;
assign output_40 = input_44;
assign output_41 = input_44;
assign output_42 = input_44;
assign output_43 = input_44;
assign output_44 = input_44;
assign output_45 = input_44;
assign output_46 = input_44;
assign output_47 = input_44;
assign output_48 = input_44;
assign output_49 = input_44;
assign output_50 = input_44;
assign output_51 = input_44;
assign output_52 = input_44;
assign output_53 = input_44;
assign output_54 = input_44;
assign output_55 = input_44;
assign output_56 = input_44;
assign output_57 = input_44;
assign output_58 = input_44;
assign output_59 = input_44;
assign output_60 = input_44;
assign output_61 = input_44;
assign output_62 = input_44;
assign output_63 = input_44;
assign output_0 = input_45;
assign output_1 = input_45;
assign output_2 = input_45;
assign output_3 = input_45;
assign output_4 = input_45;
assign output_5 = input_45;
assign output_6 = input_45;
assign output_7 = input_45;
assign output_8 = input_45;
assign output_9 = input_45;
assign output_10 = input_45;
assign output_11 = input_45;
assign output_12 = input_45;
assign output_13 = input_45;
assign output_14 = input_45;
assign output_15 = input_45;
assign output_16 = input_45;
assign output_17 = input_45;
assign output_18 = input_45;
assign output_19 = input_45;
assign output_20 = input_45;
assign output_21 = input_45;
assign output_22 = input_45;
assign output_23 = input_45;
assign output_24 = input_45;
assign output_25 = input_45;
assign output_26 = input_45;
assign output_27 = input_45;
assign output_28 = input_45;
assign output_29 = input_45;
assign output_30 = input_45;
assign output_31 = input_45;
assign output_32 = input_45;
assign output_33 = input_45;
assign output_34 = input_45;
assign output_35 = input_45;
assign output_36 = input_45;
assign output_37 = input_45;
assign output_38 = input_45;
assign output_39 = input_45;
assign output_40 = input_45;
assign output_41 = input_45;
assign output_42 = input_45;
assign output_43 = input_45;
assign output_44 = input_45;
assign output_45 = input_45;
assign output_46 = input_45;
assign output_47 = input_45;
assign output_48 = input_45;
assign output_49 = input_45;
assign output_50 = input_45;
assign output_51 = input_45;
assign output_52 = input_45;
assign output_53 = input_45;
assign output_54 = input_45;
assign output_55 = input_45;
assign output_56 = input_45;
assign output_57 = input_45;
assign output_58 = input_45;
assign output_59 = input_45;
assign output_60 = input_45;
assign output_61 = input_45;
assign output_62 = input_45;
assign output_63 = input_45;
assign output_0 = input_46;
assign output_1 = input_46;
assign output_2 = input_46;
assign output_3 = input_46;
assign output_4 = input_46;
assign output_5 = input_46;
assign output_6 = input_46;
assign output_7 = input_46;
assign output_8 = input_46;
assign output_9 = input_46;
assign output_10 = input_46;
assign output_11 = input_46;
assign output_12 = input_46;
assign output_13 = input_46;
assign output_14 = input_46;
assign output_15 = input_46;
assign output_16 = input_46;
assign output_17 = input_46;
assign output_18 = input_46;
assign output_19 = input_46;
assign output_20 = input_46;
assign output_21 = input_46;
assign output_22 = input_46;
assign output_23 = input_46;
assign output_24 = input_46;
assign output_25 = input_46;
assign output_26 = input_46;
assign output_27 = input_46;
assign output_28 = input_46;
assign output_29 = input_46;
assign output_30 = input_46;
assign output_31 = input_46;
assign output_32 = input_46;
assign output_33 = input_46;
assign output_34 = input_46;
assign output_35 = input_46;
assign output_36 = input_46;
assign output_37 = input_46;
assign output_38 = input_46;
assign output_39 = input_46;
assign output_40 = input_46;
assign output_41 = input_46;
assign output_42 = input_46;
assign output_43 = input_46;
assign output_44 = input_46;
assign output_45 = input_46;
assign output_46 = input_46;
assign output_47 = input_46;
assign output_48 = input_46;
assign output_49 = input_46;
assign output_50 = input_46;
assign output_51 = input_46;
assign output_52 = input_46;
assign output_53 = input_46;
assign output_54 = input_46;
assign output_55 = input_46;
assign output_56 = input_46;
assign output_57 = input_46;
assign output_58 = input_46;
assign output_59 = input_46;
assign output_60 = input_46;
assign output_61 = input_46;
assign output_62 = input_46;
assign output_63 = input_46;
assign output_0 = input_47;
assign output_1 = input_47;
assign output_2 = input_47;
assign output_3 = input_47;
assign output_4 = input_47;
assign output_5 = input_47;
assign output_6 = input_47;
assign output_7 = input_47;
assign output_8 = input_47;
assign output_9 = input_47;
assign output_10 = input_47;
assign output_11 = input_47;
assign output_12 = input_47;
assign output_13 = input_47;
assign output_14 = input_47;
assign output_15 = input_47;
assign output_16 = input_47;
assign output_17 = input_47;
assign output_18 = input_47;
assign output_19 = input_47;
assign output_20 = input_47;
assign output_21 = input_47;
assign output_22 = input_47;
assign output_23 = input_47;
assign output_24 = input_47;
assign output_25 = input_47;
assign output_26 = input_47;
assign output_27 = input_47;
assign output_28 = input_47;
assign output_29 = input_47;
assign output_30 = input_47;
assign output_31 = input_47;
assign output_32 = input_47;
assign output_33 = input_47;
assign output_34 = input_47;
assign output_35 = input_47;
assign output_36 = input_47;
assign output_37 = input_47;
assign output_38 = input_47;
assign output_39 = input_47;
assign output_40 = input_47;
assign output_41 = input_47;
assign output_42 = input_47;
assign output_43 = input_47;
assign output_44 = input_47;
assign output_45 = input_47;
assign output_46 = input_47;
assign output_47 = input_47;
assign output_48 = input_47;
assign output_49 = input_47;
assign output_50 = input_47;
assign output_51 = input_47;
assign output_52 = input_47;
assign output_53 = input_47;
assign output_54 = input_47;
assign output_55 = input_47;
assign output_56 = input_47;
assign output_57 = input_47;
assign output_58 = input_47;
assign output_59 = input_47;
assign output_60 = input_47;
assign output_61 = input_47;
assign output_62 = input_47;
assign output_63 = input_47;
assign output_0 = input_48;
assign output_1 = input_48;
assign output_2 = input_48;
assign output_3 = input_48;
assign output_4 = input_48;
assign output_5 = input_48;
assign output_6 = input_48;
assign output_7 = input_48;
assign output_8 = input_48;
assign output_9 = input_48;
assign output_10 = input_48;
assign output_11 = input_48;
assign output_12 = input_48;
assign output_13 = input_48;
assign output_14 = input_48;
assign output_15 = input_48;
assign output_16 = input_48;
assign output_17 = input_48;
assign output_18 = input_48;
assign output_19 = input_48;
assign output_20 = input_48;
assign output_21 = input_48;
assign output_22 = input_48;
assign output_23 = input_48;
assign output_24 = input_48;
assign output_25 = input_48;
assign output_26 = input_48;
assign output_27 = input_48;
assign output_28 = input_48;
assign output_29 = input_48;
assign output_30 = input_48;
assign output_31 = input_48;
assign output_32 = input_48;
assign output_33 = input_48;
assign output_34 = input_48;
assign output_35 = input_48;
assign output_36 = input_48;
assign output_37 = input_48;
assign output_38 = input_48;
assign output_39 = input_48;
assign output_40 = input_48;
assign output_41 = input_48;
assign output_42 = input_48;
assign output_43 = input_48;
assign output_44 = input_48;
assign output_45 = input_48;
assign output_46 = input_48;
assign output_47 = input_48;
assign output_48 = input_48;
assign output_49 = input_48;
assign output_50 = input_48;
assign output_51 = input_48;
assign output_52 = input_48;
assign output_53 = input_48;
assign output_54 = input_48;
assign output_55 = input_48;
assign output_56 = input_48;
assign output_57 = input_48;
assign output_58 = input_48;
assign output_59 = input_48;
assign output_60 = input_48;
assign output_61 = input_48;
assign output_62 = input_48;
assign output_63 = input_48;
assign output_0 = input_49;
assign output_1 = input_49;
assign output_2 = input_49;
assign output_3 = input_49;
assign output_4 = input_49;
assign output_5 = input_49;
assign output_6 = input_49;
assign output_7 = input_49;
assign output_8 = input_49;
assign output_9 = input_49;
assign output_10 = input_49;
assign output_11 = input_49;
assign output_12 = input_49;
assign output_13 = input_49;
assign output_14 = input_49;
assign output_15 = input_49;
assign output_16 = input_49;
assign output_17 = input_49;
assign output_18 = input_49;
assign output_19 = input_49;
assign output_20 = input_49;
assign output_21 = input_49;
assign output_22 = input_49;
assign output_23 = input_49;
assign output_24 = input_49;
assign output_25 = input_49;
assign output_26 = input_49;
assign output_27 = input_49;
assign output_28 = input_49;
assign output_29 = input_49;
assign output_30 = input_49;
assign output_31 = input_49;
assign output_32 = input_49;
assign output_33 = input_49;
assign output_34 = input_49;
assign output_35 = input_49;
assign output_36 = input_49;
assign output_37 = input_49;
assign output_38 = input_49;
assign output_39 = input_49;
assign output_40 = input_49;
assign output_41 = input_49;
assign output_42 = input_49;
assign output_43 = input_49;
assign output_44 = input_49;
assign output_45 = input_49;
assign output_46 = input_49;
assign output_47 = input_49;
assign output_48 = input_49;
assign output_49 = input_49;
assign output_50 = input_49;
assign output_51 = input_49;
assign output_52 = input_49;
assign output_53 = input_49;
assign output_54 = input_49;
assign output_55 = input_49;
assign output_56 = input_49;
assign output_57 = input_49;
assign output_58 = input_49;
assign output_59 = input_49;
assign output_60 = input_49;
assign output_61 = input_49;
assign output_62 = input_49;
assign output_63 = input_49;
assign output_0 = input_50;
assign output_1 = input_50;
assign output_2 = input_50;
assign output_3 = input_50;
assign output_4 = input_50;
assign output_5 = input_50;
assign output_6 = input_50;
assign output_7 = input_50;
assign output_8 = input_50;
assign output_9 = input_50;
assign output_10 = input_50;
assign output_11 = input_50;
assign output_12 = input_50;
assign output_13 = input_50;
assign output_14 = input_50;
assign output_15 = input_50;
assign output_16 = input_50;
assign output_17 = input_50;
assign output_18 = input_50;
assign output_19 = input_50;
assign output_20 = input_50;
assign output_21 = input_50;
assign output_22 = input_50;
assign output_23 = input_50;
assign output_24 = input_50;
assign output_25 = input_50;
assign output_26 = input_50;
assign output_27 = input_50;
assign output_28 = input_50;
assign output_29 = input_50;
assign output_30 = input_50;
assign output_31 = input_50;
assign output_32 = input_50;
assign output_33 = input_50;
assign output_34 = input_50;
assign output_35 = input_50;
assign output_36 = input_50;
assign output_37 = input_50;
assign output_38 = input_50;
assign output_39 = input_50;
assign output_40 = input_50;
assign output_41 = input_50;
assign output_42 = input_50;
assign output_43 = input_50;
assign output_44 = input_50;
assign output_45 = input_50;
assign output_46 = input_50;
assign output_47 = input_50;
assign output_48 = input_50;
assign output_49 = input_50;
assign output_50 = input_50;
assign output_51 = input_50;
assign output_52 = input_50;
assign output_53 = input_50;
assign output_54 = input_50;
assign output_55 = input_50;
assign output_56 = input_50;
assign output_57 = input_50;
assign output_58 = input_50;
assign output_59 = input_50;
assign output_60 = input_50;
assign output_61 = input_50;
assign output_62 = input_50;
assign output_63 = input_50;
assign output_0 = input_51;
assign output_1 = input_51;
assign output_2 = input_51;
assign output_3 = input_51;
assign output_4 = input_51;
assign output_5 = input_51;
assign output_6 = input_51;
assign output_7 = input_51;
assign output_8 = input_51;
assign output_9 = input_51;
assign output_10 = input_51;
assign output_11 = input_51;
assign output_12 = input_51;
assign output_13 = input_51;
assign output_14 = input_51;
assign output_15 = input_51;
assign output_16 = input_51;
assign output_17 = input_51;
assign output_18 = input_51;
assign output_19 = input_51;
assign output_20 = input_51;
assign output_21 = input_51;
assign output_22 = input_51;
assign output_23 = input_51;
assign output_24 = input_51;
assign output_25 = input_51;
assign output_26 = input_51;
assign output_27 = input_51;
assign output_28 = input_51;
assign output_29 = input_51;
assign output_30 = input_51;
assign output_31 = input_51;
assign output_32 = input_51;
assign output_33 = input_51;
assign output_34 = input_51;
assign output_35 = input_51;
assign output_36 = input_51;
assign output_37 = input_51;
assign output_38 = input_51;
assign output_39 = input_51;
assign output_40 = input_51;
assign output_41 = input_51;
assign output_42 = input_51;
assign output_43 = input_51;
assign output_44 = input_51;
assign output_45 = input_51;
assign output_46 = input_51;
assign output_47 = input_51;
assign output_48 = input_51;
assign output_49 = input_51;
assign output_50 = input_51;
assign output_51 = input_51;
assign output_52 = input_51;
assign output_53 = input_51;
assign output_54 = input_51;
assign output_55 = input_51;
assign output_56 = input_51;
assign output_57 = input_51;
assign output_58 = input_51;
assign output_59 = input_51;
assign output_60 = input_51;
assign output_61 = input_51;
assign output_62 = input_51;
assign output_63 = input_51;
assign output_0 = input_52;
assign output_1 = input_52;
assign output_2 = input_52;
assign output_3 = input_52;
assign output_4 = input_52;
assign output_5 = input_52;
assign output_6 = input_52;
assign output_7 = input_52;
assign output_8 = input_52;
assign output_9 = input_52;
assign output_10 = input_52;
assign output_11 = input_52;
assign output_12 = input_52;
assign output_13 = input_52;
assign output_14 = input_52;
assign output_15 = input_52;
assign output_16 = input_52;
assign output_17 = input_52;
assign output_18 = input_52;
assign output_19 = input_52;
assign output_20 = input_52;
assign output_21 = input_52;
assign output_22 = input_52;
assign output_23 = input_52;
assign output_24 = input_52;
assign output_25 = input_52;
assign output_26 = input_52;
assign output_27 = input_52;
assign output_28 = input_52;
assign output_29 = input_52;
assign output_30 = input_52;
assign output_31 = input_52;
assign output_32 = input_52;
assign output_33 = input_52;
assign output_34 = input_52;
assign output_35 = input_52;
assign output_36 = input_52;
assign output_37 = input_52;
assign output_38 = input_52;
assign output_39 = input_52;
assign output_40 = input_52;
assign output_41 = input_52;
assign output_42 = input_52;
assign output_43 = input_52;
assign output_44 = input_52;
assign output_45 = input_52;
assign output_46 = input_52;
assign output_47 = input_52;
assign output_48 = input_52;
assign output_49 = input_52;
assign output_50 = input_52;
assign output_51 = input_52;
assign output_52 = input_52;
assign output_53 = input_52;
assign output_54 = input_52;
assign output_55 = input_52;
assign output_56 = input_52;
assign output_57 = input_52;
assign output_58 = input_52;
assign output_59 = input_52;
assign output_60 = input_52;
assign output_61 = input_52;
assign output_62 = input_52;
assign output_63 = input_52;
assign output_0 = input_53;
assign output_1 = input_53;
assign output_2 = input_53;
assign output_3 = input_53;
assign output_4 = input_53;
assign output_5 = input_53;
assign output_6 = input_53;
assign output_7 = input_53;
assign output_8 = input_53;
assign output_9 = input_53;
assign output_10 = input_53;
assign output_11 = input_53;
assign output_12 = input_53;
assign output_13 = input_53;
assign output_14 = input_53;
assign output_15 = input_53;
assign output_16 = input_53;
assign output_17 = input_53;
assign output_18 = input_53;
assign output_19 = input_53;
assign output_20 = input_53;
assign output_21 = input_53;
assign output_22 = input_53;
assign output_23 = input_53;
assign output_24 = input_53;
assign output_25 = input_53;
assign output_26 = input_53;
assign output_27 = input_53;
assign output_28 = input_53;
assign output_29 = input_53;
assign output_30 = input_53;
assign output_31 = input_53;
assign output_32 = input_53;
assign output_33 = input_53;
assign output_34 = input_53;
assign output_35 = input_53;
assign output_36 = input_53;
assign output_37 = input_53;
assign output_38 = input_53;
assign output_39 = input_53;
assign output_40 = input_53;
assign output_41 = input_53;
assign output_42 = input_53;
assign output_43 = input_53;
assign output_44 = input_53;
assign output_45 = input_53;
assign output_46 = input_53;
assign output_47 = input_53;
assign output_48 = input_53;
assign output_49 = input_53;
assign output_50 = input_53;
assign output_51 = input_53;
assign output_52 = input_53;
assign output_53 = input_53;
assign output_54 = input_53;
assign output_55 = input_53;
assign output_56 = input_53;
assign output_57 = input_53;
assign output_58 = input_53;
assign output_59 = input_53;
assign output_60 = input_53;
assign output_61 = input_53;
assign output_62 = input_53;
assign output_63 = input_53;
assign output_0 = input_54;
assign output_1 = input_54;
assign output_2 = input_54;
assign output_3 = input_54;
assign output_4 = input_54;
assign output_5 = input_54;
assign output_6 = input_54;
assign output_7 = input_54;
assign output_8 = input_54;
assign output_9 = input_54;
assign output_10 = input_54;
assign output_11 = input_54;
assign output_12 = input_54;
assign output_13 = input_54;
assign output_14 = input_54;
assign output_15 = input_54;
assign output_16 = input_54;
assign output_17 = input_54;
assign output_18 = input_54;
assign output_19 = input_54;
assign output_20 = input_54;
assign output_21 = input_54;
assign output_22 = input_54;
assign output_23 = input_54;
assign output_24 = input_54;
assign output_25 = input_54;
assign output_26 = input_54;
assign output_27 = input_54;
assign output_28 = input_54;
assign output_29 = input_54;
assign output_30 = input_54;
assign output_31 = input_54;
assign output_32 = input_54;
assign output_33 = input_54;
assign output_34 = input_54;
assign output_35 = input_54;
assign output_36 = input_54;
assign output_37 = input_54;
assign output_38 = input_54;
assign output_39 = input_54;
assign output_40 = input_54;
assign output_41 = input_54;
assign output_42 = input_54;
assign output_43 = input_54;
assign output_44 = input_54;
assign output_45 = input_54;
assign output_46 = input_54;
assign output_47 = input_54;
assign output_48 = input_54;
assign output_49 = input_54;
assign output_50 = input_54;
assign output_51 = input_54;
assign output_52 = input_54;
assign output_53 = input_54;
assign output_54 = input_54;
assign output_55 = input_54;
assign output_56 = input_54;
assign output_57 = input_54;
assign output_58 = input_54;
assign output_59 = input_54;
assign output_60 = input_54;
assign output_61 = input_54;
assign output_62 = input_54;
assign output_63 = input_54;
assign output_0 = input_55;
assign output_1 = input_55;
assign output_2 = input_55;
assign output_3 = input_55;
assign output_4 = input_55;
assign output_5 = input_55;
assign output_6 = input_55;
assign output_7 = input_55;
assign output_8 = input_55;
assign output_9 = input_55;
assign output_10 = input_55;
assign output_11 = input_55;
assign output_12 = input_55;
assign output_13 = input_55;
assign output_14 = input_55;
assign output_15 = input_55;
assign output_16 = input_55;
assign output_17 = input_55;
assign output_18 = input_55;
assign output_19 = input_55;
assign output_20 = input_55;
assign output_21 = input_55;
assign output_22 = input_55;
assign output_23 = input_55;
assign output_24 = input_55;
assign output_25 = input_55;
assign output_26 = input_55;
assign output_27 = input_55;
assign output_28 = input_55;
assign output_29 = input_55;
assign output_30 = input_55;
assign output_31 = input_55;
assign output_32 = input_55;
assign output_33 = input_55;
assign output_34 = input_55;
assign output_35 = input_55;
assign output_36 = input_55;
assign output_37 = input_55;
assign output_38 = input_55;
assign output_39 = input_55;
assign output_40 = input_55;
assign output_41 = input_55;
assign output_42 = input_55;
assign output_43 = input_55;
assign output_44 = input_55;
assign output_45 = input_55;
assign output_46 = input_55;
assign output_47 = input_55;
assign output_48 = input_55;
assign output_49 = input_55;
assign output_50 = input_55;
assign output_51 = input_55;
assign output_52 = input_55;
assign output_53 = input_55;
assign output_54 = input_55;
assign output_55 = input_55;
assign output_56 = input_55;
assign output_57 = input_55;
assign output_58 = input_55;
assign output_59 = input_55;
assign output_60 = input_55;
assign output_61 = input_55;
assign output_62 = input_55;
assign output_63 = input_55;
assign output_0 = input_56;
assign output_1 = input_56;
assign output_2 = input_56;
assign output_3 = input_56;
assign output_4 = input_56;
assign output_5 = input_56;
assign output_6 = input_56;
assign output_7 = input_56;
assign output_8 = input_56;
assign output_9 = input_56;
assign output_10 = input_56;
assign output_11 = input_56;
assign output_12 = input_56;
assign output_13 = input_56;
assign output_14 = input_56;
assign output_15 = input_56;
assign output_16 = input_56;
assign output_17 = input_56;
assign output_18 = input_56;
assign output_19 = input_56;
assign output_20 = input_56;
assign output_21 = input_56;
assign output_22 = input_56;
assign output_23 = input_56;
assign output_24 = input_56;
assign output_25 = input_56;
assign output_26 = input_56;
assign output_27 = input_56;
assign output_28 = input_56;
assign output_29 = input_56;
assign output_30 = input_56;
assign output_31 = input_56;
assign output_32 = input_56;
assign output_33 = input_56;
assign output_34 = input_56;
assign output_35 = input_56;
assign output_36 = input_56;
assign output_37 = input_56;
assign output_38 = input_56;
assign output_39 = input_56;
assign output_40 = input_56;
assign output_41 = input_56;
assign output_42 = input_56;
assign output_43 = input_56;
assign output_44 = input_56;
assign output_45 = input_56;
assign output_46 = input_56;
assign output_47 = input_56;
assign output_48 = input_56;
assign output_49 = input_56;
assign output_50 = input_56;
assign output_51 = input_56;
assign output_52 = input_56;
assign output_53 = input_56;
assign output_54 = input_56;
assign output_55 = input_56;
assign output_56 = input_56;
assign output_57 = input_56;
assign output_58 = input_56;
assign output_59 = input_56;
assign output_60 = input_56;
assign output_61 = input_56;
assign output_62 = input_56;
assign output_63 = input_56;
assign output_0 = input_57;
assign output_1 = input_57;
assign output_2 = input_57;
assign output_3 = input_57;
assign output_4 = input_57;
assign output_5 = input_57;
assign output_6 = input_57;
assign output_7 = input_57;
assign output_8 = input_57;
assign output_9 = input_57;
assign output_10 = input_57;
assign output_11 = input_57;
assign output_12 = input_57;
assign output_13 = input_57;
assign output_14 = input_57;
assign output_15 = input_57;
assign output_16 = input_57;
assign output_17 = input_57;
assign output_18 = input_57;
assign output_19 = input_57;
assign output_20 = input_57;
assign output_21 = input_57;
assign output_22 = input_57;
assign output_23 = input_57;
assign output_24 = input_57;
assign output_25 = input_57;
assign output_26 = input_57;
assign output_27 = input_57;
assign output_28 = input_57;
assign output_29 = input_57;
assign output_30 = input_57;
assign output_31 = input_57;
assign output_32 = input_57;
assign output_33 = input_57;
assign output_34 = input_57;
assign output_35 = input_57;
assign output_36 = input_57;
assign output_37 = input_57;
assign output_38 = input_57;
assign output_39 = input_57;
assign output_40 = input_57;
assign output_41 = input_57;
assign output_42 = input_57;
assign output_43 = input_57;
assign output_44 = input_57;
assign output_45 = input_57;
assign output_46 = input_57;
assign output_47 = input_57;
assign output_48 = input_57;
assign output_49 = input_57;
assign output_50 = input_57;
assign output_51 = input_57;
assign output_52 = input_57;
assign output_53 = input_57;
assign output_54 = input_57;
assign output_55 = input_57;
assign output_56 = input_57;
assign output_57 = input_57;
assign output_58 = input_57;
assign output_59 = input_57;
assign output_60 = input_57;
assign output_61 = input_57;
assign output_62 = input_57;
assign output_63 = input_57;
assign output_0 = input_58;
assign output_1 = input_58;
assign output_2 = input_58;
assign output_3 = input_58;
assign output_4 = input_58;
assign output_5 = input_58;
assign output_6 = input_58;
assign output_7 = input_58;
assign output_8 = input_58;
assign output_9 = input_58;
assign output_10 = input_58;
assign output_11 = input_58;
assign output_12 = input_58;
assign output_13 = input_58;
assign output_14 = input_58;
assign output_15 = input_58;
assign output_16 = input_58;
assign output_17 = input_58;
assign output_18 = input_58;
assign output_19 = input_58;
assign output_20 = input_58;
assign output_21 = input_58;
assign output_22 = input_58;
assign output_23 = input_58;
assign output_24 = input_58;
assign output_25 = input_58;
assign output_26 = input_58;
assign output_27 = input_58;
assign output_28 = input_58;
assign output_29 = input_58;
assign output_30 = input_58;
assign output_31 = input_58;
assign output_32 = input_58;
assign output_33 = input_58;
assign output_34 = input_58;
assign output_35 = input_58;
assign output_36 = input_58;
assign output_37 = input_58;
assign output_38 = input_58;
assign output_39 = input_58;
assign output_40 = input_58;
assign output_41 = input_58;
assign output_42 = input_58;
assign output_43 = input_58;
assign output_44 = input_58;
assign output_45 = input_58;
assign output_46 = input_58;
assign output_47 = input_58;
assign output_48 = input_58;
assign output_49 = input_58;
assign output_50 = input_58;
assign output_51 = input_58;
assign output_52 = input_58;
assign output_53 = input_58;
assign output_54 = input_58;
assign output_55 = input_58;
assign output_56 = input_58;
assign output_57 = input_58;
assign output_58 = input_58;
assign output_59 = input_58;
assign output_60 = input_58;
assign output_61 = input_58;
assign output_62 = input_58;
assign output_63 = input_58;
assign output_0 = input_59;
assign output_1 = input_59;
assign output_2 = input_59;
assign output_3 = input_59;
assign output_4 = input_59;
assign output_5 = input_59;
assign output_6 = input_59;
assign output_7 = input_59;
assign output_8 = input_59;
assign output_9 = input_59;
assign output_10 = input_59;
assign output_11 = input_59;
assign output_12 = input_59;
assign output_13 = input_59;
assign output_14 = input_59;
assign output_15 = input_59;
assign output_16 = input_59;
assign output_17 = input_59;
assign output_18 = input_59;
assign output_19 = input_59;
assign output_20 = input_59;
assign output_21 = input_59;
assign output_22 = input_59;
assign output_23 = input_59;
assign output_24 = input_59;
assign output_25 = input_59;
assign output_26 = input_59;
assign output_27 = input_59;
assign output_28 = input_59;
assign output_29 = input_59;
assign output_30 = input_59;
assign output_31 = input_59;
assign output_32 = input_59;
assign output_33 = input_59;
assign output_34 = input_59;
assign output_35 = input_59;
assign output_36 = input_59;
assign output_37 = input_59;
assign output_38 = input_59;
assign output_39 = input_59;
assign output_40 = input_59;
assign output_41 = input_59;
assign output_42 = input_59;
assign output_43 = input_59;
assign output_44 = input_59;
assign output_45 = input_59;
assign output_46 = input_59;
assign output_47 = input_59;
assign output_48 = input_59;
assign output_49 = input_59;
assign output_50 = input_59;
assign output_51 = input_59;
assign output_52 = input_59;
assign output_53 = input_59;
assign output_54 = input_59;
assign output_55 = input_59;
assign output_56 = input_59;
assign output_57 = input_59;
assign output_58 = input_59;
assign output_59 = input_59;
assign output_60 = input_59;
assign output_61 = input_59;
assign output_62 = input_59;
assign output_63 = input_59;
assign output_0 = input_60;
assign output_1 = input_60;
assign output_2 = input_60;
assign output_3 = input_60;
assign output_4 = input_60;
assign output_5 = input_60;
assign output_6 = input_60;
assign output_7 = input_60;
assign output_8 = input_60;
assign output_9 = input_60;
assign output_10 = input_60;
assign output_11 = input_60;
assign output_12 = input_60;
assign output_13 = input_60;
assign output_14 = input_60;
assign output_15 = input_60;
assign output_16 = input_60;
assign output_17 = input_60;
assign output_18 = input_60;
assign output_19 = input_60;
assign output_20 = input_60;
assign output_21 = input_60;
assign output_22 = input_60;
assign output_23 = input_60;
assign output_24 = input_60;
assign output_25 = input_60;
assign output_26 = input_60;
assign output_27 = input_60;
assign output_28 = input_60;
assign output_29 = input_60;
assign output_30 = input_60;
assign output_31 = input_60;
assign output_32 = input_60;
assign output_33 = input_60;
assign output_34 = input_60;
assign output_35 = input_60;
assign output_36 = input_60;
assign output_37 = input_60;
assign output_38 = input_60;
assign output_39 = input_60;
assign output_40 = input_60;
assign output_41 = input_60;
assign output_42 = input_60;
assign output_43 = input_60;
assign output_44 = input_60;
assign output_45 = input_60;
assign output_46 = input_60;
assign output_47 = input_60;
assign output_48 = input_60;
assign output_49 = input_60;
assign output_50 = input_60;
assign output_51 = input_60;
assign output_52 = input_60;
assign output_53 = input_60;
assign output_54 = input_60;
assign output_55 = input_60;
assign output_56 = input_60;
assign output_57 = input_60;
assign output_58 = input_60;
assign output_59 = input_60;
assign output_60 = input_60;
assign output_61 = input_60;
assign output_62 = input_60;
assign output_63 = input_60;
assign output_0 = input_61;
assign output_1 = input_61;
assign output_2 = input_61;
assign output_3 = input_61;
assign output_4 = input_61;
assign output_5 = input_61;
assign output_6 = input_61;
assign output_7 = input_61;
assign output_8 = input_61;
assign output_9 = input_61;
assign output_10 = input_61;
assign output_11 = input_61;
assign output_12 = input_61;
assign output_13 = input_61;
assign output_14 = input_61;
assign output_15 = input_61;
assign output_16 = input_61;
assign output_17 = input_61;
assign output_18 = input_61;
assign output_19 = input_61;
assign output_20 = input_61;
assign output_21 = input_61;
assign output_22 = input_61;
assign output_23 = input_61;
assign output_24 = input_61;
assign output_25 = input_61;
assign output_26 = input_61;
assign output_27 = input_61;
assign output_28 = input_61;
assign output_29 = input_61;
assign output_30 = input_61;
assign output_31 = input_61;
assign output_32 = input_61;
assign output_33 = input_61;
assign output_34 = input_61;
assign output_35 = input_61;
assign output_36 = input_61;
assign output_37 = input_61;
assign output_38 = input_61;
assign output_39 = input_61;
assign output_40 = input_61;
assign output_41 = input_61;
assign output_42 = input_61;
assign output_43 = input_61;
assign output_44 = input_61;
assign output_45 = input_61;
assign output_46 = input_61;
assign output_47 = input_61;
assign output_48 = input_61;
assign output_49 = input_61;
assign output_50 = input_61;
assign output_51 = input_61;
assign output_52 = input_61;
assign output_53 = input_61;
assign output_54 = input_61;
assign output_55 = input_61;
assign output_56 = input_61;
assign output_57 = input_61;
assign output_58 = input_61;
assign output_59 = input_61;
assign output_60 = input_61;
assign output_61 = input_61;
assign output_62 = input_61;
assign output_63 = input_61;
assign output_0 = input_62;
assign output_1 = input_62;
assign output_2 = input_62;
assign output_3 = input_62;
assign output_4 = input_62;
assign output_5 = input_62;
assign output_6 = input_62;
assign output_7 = input_62;
assign output_8 = input_62;
assign output_9 = input_62;
assign output_10 = input_62;
assign output_11 = input_62;
assign output_12 = input_62;
assign output_13 = input_62;
assign output_14 = input_62;
assign output_15 = input_62;
assign output_16 = input_62;
assign output_17 = input_62;
assign output_18 = input_62;
assign output_19 = input_62;
assign output_20 = input_62;
assign output_21 = input_62;
assign output_22 = input_62;
assign output_23 = input_62;
assign output_24 = input_62;
assign output_25 = input_62;
assign output_26 = input_62;
assign output_27 = input_62;
assign output_28 = input_62;
assign output_29 = input_62;
assign output_30 = input_62;
assign output_31 = input_62;
assign output_32 = input_62;
assign output_33 = input_62;
assign output_34 = input_62;
assign output_35 = input_62;
assign output_36 = input_62;
assign output_37 = input_62;
assign output_38 = input_62;
assign output_39 = input_62;
assign output_40 = input_62;
assign output_41 = input_62;
assign output_42 = input_62;
assign output_43 = input_62;
assign output_44 = input_62;
assign output_45 = input_62;
assign output_46 = input_62;
assign output_47 = input_62;
assign output_48 = input_62;
assign output_49 = input_62;
assign output_50 = input_62;
assign output_51 = input_62;
assign output_52 = input_62;
assign output_53 = input_62;
assign output_54 = input_62;
assign output_55 = input_62;
assign output_56 = input_62;
assign output_57 = input_62;
assign output_58 = input_62;
assign output_59 = input_62;
assign output_60 = input_62;
assign output_61 = input_62;
assign output_62 = input_62;
assign output_63 = input_62;
assign output_0 = input_63;
assign output_1 = input_63;
assign output_2 = input_63;
assign output_3 = input_63;
assign output_4 = input_63;
assign output_5 = input_63;
assign output_6 = input_63;
assign output_7 = input_63;
assign output_8 = input_63;
assign output_9 = input_63;
assign output_10 = input_63;
assign output_11 = input_63;
assign output_12 = input_63;
assign output_13 = input_63;
assign output_14 = input_63;
assign output_15 = input_63;
assign output_16 = input_63;
assign output_17 = input_63;
assign output_18 = input_63;
assign output_19 = input_63;
assign output_20 = input_63;
assign output_21 = input_63;
assign output_22 = input_63;
assign output_23 = input_63;
assign output_24 = input_63;
assign output_25 = input_63;
assign output_26 = input_63;
assign output_27 = input_63;
assign output_28 = input_63;
assign output_29 = input_63;
assign output_30 = input_63;
assign output_31 = input_63;
assign output_32 = input_63;
assign output_33 = input_63;
assign output_34 = input_63;
assign output_35 = input_63;
assign output_36 = input_63;
assign output_37 = input_63;
assign output_38 = input_63;
assign output_39 = input_63;
assign output_40 = input_63;
assign output_41 = input_63;
assign output_42 = input_63;
assign output_43 = input_63;
assign output_44 = input_63;
assign output_45 = input_63;
assign output_46 = input_63;
assign output_47 = input_63;
assign output_48 = input_63;
assign output_49 = input_63;
assign output_50 = input_63;
assign output_51 = input_63;
assign output_52 = input_63;
assign output_53 = input_63;
assign output_54 = input_63;
assign output_55 = input_63;
assign output_56 = input_63;
assign output_57 = input_63;
assign output_58 = input_63;
assign output_59 = input_63;
assign output_60 = input_63;
assign output_61 = input_63;
assign output_62 = input_63;
assign output_63 = input_63;
endmodule
