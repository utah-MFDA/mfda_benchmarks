module binary_tree_1_12 (
output out_0,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63,input input_64,input input_65,input input_66,input input_67,input input_68,input input_69,input input_70,input input_71,input input_72,input input_73,input input_74,input input_75,input input_76,input input_77,input input_78,input input_79,input input_80,input input_81,input input_82,input input_83,input input_84,input input_85,input input_86,input input_87,input input_88,input input_89,input input_90,input input_91,input input_92,input input_93,input input_94,input input_95,input input_96,input input_97,input input_98,input input_99,input input_100,input input_101,input input_102,input input_103,input input_104,input input_105,input input_106,input input_107,input input_108,input input_109,input input_110,input input_111,input input_112,input input_113,input input_114,input input_115,input input_116,input input_117,input input_118,input input_119,input input_120,input input_121,input input_122,input input_123,input input_124,input input_125,input input_126,input input_127,input input_128,input input_129,input input_130,input input_131,input input_132,input input_133,input input_134,input input_135,input input_136,input input_137,input input_138,input input_139,input input_140,input input_141,input input_142,input input_143,input input_144,input input_145,input input_146,input input_147,input input_148,input input_149,input input_150,input input_151,input input_152,input input_153,input input_154,input input_155,input input_156,input input_157,input input_158,input input_159,input input_160,input input_161,input input_162,input input_163,input input_164,input input_165,input input_166,input input_167,input input_168,input input_169,input input_170,input input_171,input input_172,input input_173,input input_174,input input_175,input input_176,input input_177,input input_178,input input_179,input input_180,input input_181,input input_182,input input_183,input input_184,input input_185,input input_186,input input_187,input input_188,input input_189,input input_190,input input_191,input input_192,input input_193,input input_194,input input_195,input input_196,input input_197,input input_198,input input_199,input input_200,input input_201,input input_202,input input_203,input input_204,input input_205,input input_206,input input_207,input input_208,input input_209,input input_210,input input_211,input input_212,input input_213,input input_214,input input_215,input input_216,input input_217,input input_218,input input_219,input input_220,input input_221,input input_222,input input_223,input input_224,input input_225,input input_226,input input_227,input input_228,input input_229,input input_230,input input_231,input input_232,input input_233,input input_234,input input_235,input input_236,input input_237,input input_238,input input_239,input input_240,input input_241,input input_242,input input_243,input input_244,input input_245,input input_246,input input_247,input input_248,input input_249,input input_250,input input_251,input input_252,input input_253,input input_254,input input_255,input input_256,input input_257,input input_258,input input_259,input input_260,input input_261,input input_262,input input_263,input input_264,input input_265,input input_266,input input_267,input input_268,input input_269,input input_270,input input_271,input input_272,input input_273,input input_274,input input_275,input input_276,input input_277,input input_278,input input_279,input input_280,input input_281,input input_282,input input_283,input input_284,input input_285,input input_286,input input_287,input input_288,input input_289,input input_290,input input_291,input input_292,input input_293,input input_294,input input_295,input input_296,input input_297,input input_298,input input_299,input input_300,input input_301,input input_302,input input_303,input input_304,input input_305,input input_306,input input_307,input input_308,input input_309,input input_310,input input_311,input input_312,input input_313,input input_314,input input_315,input input_316,input input_317,input input_318,input input_319,input input_320,input input_321,input input_322,input input_323,input input_324,input input_325,input input_326,input input_327,input input_328,input input_329,input input_330,input input_331,input input_332,input input_333,input input_334,input input_335,input input_336,input input_337,input input_338,input input_339,input input_340,input input_341,input input_342,input input_343,input input_344,input input_345,input input_346,input input_347,input input_348,input input_349,input input_350,input input_351,input input_352,input input_353,input input_354,input input_355,input input_356,input input_357,input input_358,input input_359,input input_360,input input_361,input input_362,input input_363,input input_364,input input_365,input input_366,input input_367,input input_368,input input_369,input input_370,input input_371,input input_372,input input_373,input input_374,input input_375,input input_376,input input_377,input input_378,input input_379,input input_380,input input_381,input input_382,input input_383,input input_384,input input_385,input input_386,input input_387,input input_388,input input_389,input input_390,input input_391,input input_392,input input_393,input input_394,input input_395,input input_396,input input_397,input input_398,input input_399,input input_400,input input_401,input input_402,input input_403,input input_404,input input_405,input input_406,input input_407,input input_408,input input_409,input input_410,input input_411,input input_412,input input_413,input input_414,input input_415,input input_416,input input_417,input input_418,input input_419,input input_420,input input_421,input input_422,input input_423,input input_424,input input_425,input input_426,input input_427,input input_428,input input_429,input input_430,input input_431,input input_432,input input_433,input input_434,input input_435,input input_436,input input_437,input input_438,input input_439,input input_440,input input_441,input input_442,input input_443,input input_444,input input_445,input input_446,input input_447,input input_448,input input_449,input input_450,input input_451,input input_452,input input_453,input input_454,input input_455,input input_456,input input_457,input input_458,input input_459,input input_460,input input_461,input input_462,input input_463,input input_464,input input_465,input input_466,input input_467,input input_468,input input_469,input input_470,input input_471,input input_472,input input_473,input input_474,input input_475,input input_476,input input_477,input input_478,input input_479,input input_480,input input_481,input input_482,input input_483,input input_484,input input_485,input input_486,input input_487,input input_488,input input_489,input input_490,input input_491,input input_492,input input_493,input input_494,input input_495,input input_496,input input_497,input input_498,input input_499,input input_500,input input_501,input input_502,input input_503,input input_504,input input_505,input input_506,input input_507,input input_508,input input_509,input input_510,input input_511,input input_512,input input_513,input input_514,input input_515,input input_516,input input_517,input input_518,input input_519,input input_520,input input_521,input input_522,input input_523,input input_524,input input_525,input input_526,input input_527,input input_528,input input_529,input input_530,input input_531,input input_532,input input_533,input input_534,input input_535,input input_536,input input_537,input input_538,input input_539,input input_540,input input_541,input input_542,input input_543,input input_544,input input_545,input input_546,input input_547,input input_548,input input_549,input input_550,input input_551,input input_552,input input_553,input input_554,input input_555,input input_556,input input_557,input input_558,input input_559,input input_560,input input_561,input input_562,input input_563,input input_564,input input_565,input input_566,input input_567,input input_568,input input_569,input input_570,input input_571,input input_572,input input_573,input input_574,input input_575,input input_576,input input_577,input input_578,input input_579,input input_580,input input_581,input input_582,input input_583,input input_584,input input_585,input input_586,input input_587,input input_588,input input_589,input input_590,input input_591,input input_592,input input_593,input input_594,input input_595,input input_596,input input_597,input input_598,input input_599,input input_600,input input_601,input input_602,input input_603,input input_604,input input_605,input input_606,input input_607,input input_608,input input_609,input input_610,input input_611,input input_612,input input_613,input input_614,input input_615,input input_616,input input_617,input input_618,input input_619,input input_620,input input_621,input input_622,input input_623,input input_624,input input_625,input input_626,input input_627,input input_628,input input_629,input input_630,input input_631,input input_632,input input_633,input input_634,input input_635,input input_636,input input_637,input input_638,input input_639,input input_640,input input_641,input input_642,input input_643,input input_644,input input_645,input input_646,input input_647,input input_648,input input_649,input input_650,input input_651,input input_652,input input_653,input input_654,input input_655,input input_656,input input_657,input input_658,input input_659,input input_660,input input_661,input input_662,input input_663,input input_664,input input_665,input input_666,input input_667,input input_668,input input_669,input input_670,input input_671,input input_672,input input_673,input input_674,input input_675,input input_676,input input_677,input input_678,input input_679,input input_680,input input_681,input input_682,input input_683,input input_684,input input_685,input input_686,input input_687,input input_688,input input_689,input input_690,input input_691,input input_692,input input_693,input input_694,input input_695,input input_696,input input_697,input input_698,input input_699,input input_700,input input_701,input input_702,input input_703,input input_704,input input_705,input input_706,input input_707,input input_708,input input_709,input input_710,input input_711,input input_712,input input_713,input input_714,input input_715,input input_716,input input_717,input input_718,input input_719,input input_720,input input_721,input input_722,input input_723,input input_724,input input_725,input input_726,input input_727,input input_728,input input_729,input input_730,input input_731,input input_732,input input_733,input input_734,input input_735,input input_736,input input_737,input input_738,input input_739,input input_740,input input_741,input input_742,input input_743,input input_744,input input_745,input input_746,input input_747,input input_748,input input_749,input input_750,input input_751,input input_752,input input_753,input input_754,input input_755,input input_756,input input_757,input input_758,input input_759,input input_760,input input_761,input input_762,input input_763,input input_764,input input_765,input input_766,input input_767,input input_768,input input_769,input input_770,input input_771,input input_772,input input_773,input input_774,input input_775,input input_776,input input_777,input input_778,input input_779,input input_780,input input_781,input input_782,input input_783,input input_784,input input_785,input input_786,input input_787,input input_788,input input_789,input input_790,input input_791,input input_792,input input_793,input input_794,input input_795,input input_796,input input_797,input input_798,input input_799,input input_800,input input_801,input input_802,input input_803,input input_804,input input_805,input input_806,input input_807,input input_808,input input_809,input input_810,input input_811,input input_812,input input_813,input input_814,input input_815,input input_816,input input_817,input input_818,input input_819,input input_820,input input_821,input input_822,input input_823,input input_824,input input_825,input input_826,input input_827,input input_828,input input_829,input input_830,input input_831,input input_832,input input_833,input input_834,input input_835,input input_836,input input_837,input input_838,input input_839,input input_840,input input_841,input input_842,input input_843,input input_844,input input_845,input input_846,input input_847,input input_848,input input_849,input input_850,input input_851,input input_852,input input_853,input input_854,input input_855,input input_856,input input_857,input input_858,input input_859,input input_860,input input_861,input input_862,input input_863,input input_864,input input_865,input input_866,input input_867,input input_868,input input_869,input input_870,input input_871,input input_872,input input_873,input input_874,input input_875,input input_876,input input_877,input input_878,input input_879,input input_880,input input_881,input input_882,input input_883,input input_884,input input_885,input input_886,input input_887,input input_888,input input_889,input input_890,input input_891,input input_892,input input_893,input input_894,input input_895,input input_896,input input_897,input input_898,input input_899,input input_900,input input_901,input input_902,input input_903,input input_904,input input_905,input input_906,input input_907,input input_908,input input_909,input input_910,input input_911,input input_912,input input_913,input input_914,input input_915,input input_916,input input_917,input input_918,input input_919,input input_920,input input_921,input input_922,input input_923,input input_924,input input_925,input input_926,input input_927,input input_928,input input_929,input input_930,input input_931,input input_932,input input_933,input input_934,input input_935,input input_936,input input_937,input input_938,input input_939,input input_940,input input_941,input input_942,input input_943,input input_944,input input_945,input input_946,input input_947,input input_948,input input_949,input input_950,input input_951,input input_952,input input_953,input input_954,input input_955,input input_956,input input_957,input input_958,input input_959,input input_960,input input_961,input input_962,input input_963,input input_964,input input_965,input input_966,input input_967,input input_968,input input_969,input input_970,input input_971,input input_972,input input_973,input input_974,input input_975,input input_976,input input_977,input input_978,input input_979,input input_980,input input_981,input input_982,input input_983,input input_984,input input_985,input input_986,input input_987,input input_988,input input_989,input input_990,input input_991,input input_992,input input_993,input input_994,input input_995,input input_996,input input_997,input input_998,input input_999,input input_1000,input input_1001,input input_1002,input input_1003,input input_1004,input input_1005,input input_1006,input input_1007,input input_1008,input input_1009,input input_1010,input input_1011,input input_1012,input input_1013,input input_1014,input input_1015,input input_1016,input input_1017,input input_1018,input input_1019,input input_1020,input input_1021,input input_1022,input input_1023,input input_1024,input input_1025,input input_1026,input input_1027,input input_1028,input input_1029,input input_1030,input input_1031,input input_1032,input input_1033,input input_1034,input input_1035,input input_1036,input input_1037,input input_1038,input input_1039,input input_1040,input input_1041,input input_1042,input input_1043,input input_1044,input input_1045,input input_1046,input input_1047,input input_1048,input input_1049,input input_1050,input input_1051,input input_1052,input input_1053,input input_1054,input input_1055,input input_1056,input input_1057,input input_1058,input input_1059,input input_1060,input input_1061,input input_1062,input input_1063,input input_1064,input input_1065,input input_1066,input input_1067,input input_1068,input input_1069,input input_1070,input input_1071,input input_1072,input input_1073,input input_1074,input input_1075,input input_1076,input input_1077,input input_1078,input input_1079,input input_1080,input input_1081,input input_1082,input input_1083,input input_1084,input input_1085,input input_1086,input input_1087,input input_1088,input input_1089,input input_1090,input input_1091,input input_1092,input input_1093,input input_1094,input input_1095,input input_1096,input input_1097,input input_1098,input input_1099,input input_1100,input input_1101,input input_1102,input input_1103,input input_1104,input input_1105,input input_1106,input input_1107,input input_1108,input input_1109,input input_1110,input input_1111,input input_1112,input input_1113,input input_1114,input input_1115,input input_1116,input input_1117,input input_1118,input input_1119,input input_1120,input input_1121,input input_1122,input input_1123,input input_1124,input input_1125,input input_1126,input input_1127,input input_1128,input input_1129,input input_1130,input input_1131,input input_1132,input input_1133,input input_1134,input input_1135,input input_1136,input input_1137,input input_1138,input input_1139,input input_1140,input input_1141,input input_1142,input input_1143,input input_1144,input input_1145,input input_1146,input input_1147,input input_1148,input input_1149,input input_1150,input input_1151,input input_1152,input input_1153,input input_1154,input input_1155,input input_1156,input input_1157,input input_1158,input input_1159,input input_1160,input input_1161,input input_1162,input input_1163,input input_1164,input input_1165,input input_1166,input input_1167,input input_1168,input input_1169,input input_1170,input input_1171,input input_1172,input input_1173,input input_1174,input input_1175,input input_1176,input input_1177,input input_1178,input input_1179,input input_1180,input input_1181,input input_1182,input input_1183,input input_1184,input input_1185,input input_1186,input input_1187,input input_1188,input input_1189,input input_1190,input input_1191,input input_1192,input input_1193,input input_1194,input input_1195,input input_1196,input input_1197,input input_1198,input input_1199,input input_1200,input input_1201,input input_1202,input input_1203,input input_1204,input input_1205,input input_1206,input input_1207,input input_1208,input input_1209,input input_1210,input input_1211,input input_1212,input input_1213,input input_1214,input input_1215,input input_1216,input input_1217,input input_1218,input input_1219,input input_1220,input input_1221,input input_1222,input input_1223,input input_1224,input input_1225,input input_1226,input input_1227,input input_1228,input input_1229,input input_1230,input input_1231,input input_1232,input input_1233,input input_1234,input input_1235,input input_1236,input input_1237,input input_1238,input input_1239,input input_1240,input input_1241,input input_1242,input input_1243,input input_1244,input input_1245,input input_1246,input input_1247,input input_1248,input input_1249,input input_1250,input input_1251,input input_1252,input input_1253,input input_1254,input input_1255,input input_1256,input input_1257,input input_1258,input input_1259,input input_1260,input input_1261,input input_1262,input input_1263,input input_1264,input input_1265,input input_1266,input input_1267,input input_1268,input input_1269,input input_1270,input input_1271,input input_1272,input input_1273,input input_1274,input input_1275,input input_1276,input input_1277,input input_1278,input input_1279,input input_1280,input input_1281,input input_1282,input input_1283,input input_1284,input input_1285,input input_1286,input input_1287,input input_1288,input input_1289,input input_1290,input input_1291,input input_1292,input input_1293,input input_1294,input input_1295,input input_1296,input input_1297,input input_1298,input input_1299,input input_1300,input input_1301,input input_1302,input input_1303,input input_1304,input input_1305,input input_1306,input input_1307,input input_1308,input input_1309,input input_1310,input input_1311,input input_1312,input input_1313,input input_1314,input input_1315,input input_1316,input input_1317,input input_1318,input input_1319,input input_1320,input input_1321,input input_1322,input input_1323,input input_1324,input input_1325,input input_1326,input input_1327,input input_1328,input input_1329,input input_1330,input input_1331,input input_1332,input input_1333,input input_1334,input input_1335,input input_1336,input input_1337,input input_1338,input input_1339,input input_1340,input input_1341,input input_1342,input input_1343,input input_1344,input input_1345,input input_1346,input input_1347,input input_1348,input input_1349,input input_1350,input input_1351,input input_1352,input input_1353,input input_1354,input input_1355,input input_1356,input input_1357,input input_1358,input input_1359,input input_1360,input input_1361,input input_1362,input input_1363,input input_1364,input input_1365,input input_1366,input input_1367,input input_1368,input input_1369,input input_1370,input input_1371,input input_1372,input input_1373,input input_1374,input input_1375,input input_1376,input input_1377,input input_1378,input input_1379,input input_1380,input input_1381,input input_1382,input input_1383,input input_1384,input input_1385,input input_1386,input input_1387,input input_1388,input input_1389,input input_1390,input input_1391,input input_1392,input input_1393,input input_1394,input input_1395,input input_1396,input input_1397,input input_1398,input input_1399,input input_1400,input input_1401,input input_1402,input input_1403,input input_1404,input input_1405,input input_1406,input input_1407,input input_1408,input input_1409,input input_1410,input input_1411,input input_1412,input input_1413,input input_1414,input input_1415,input input_1416,input input_1417,input input_1418,input input_1419,input input_1420,input input_1421,input input_1422,input input_1423,input input_1424,input input_1425,input input_1426,input input_1427,input input_1428,input input_1429,input input_1430,input input_1431,input input_1432,input input_1433,input input_1434,input input_1435,input input_1436,input input_1437,input input_1438,input input_1439,input input_1440,input input_1441,input input_1442,input input_1443,input input_1444,input input_1445,input input_1446,input input_1447,input input_1448,input input_1449,input input_1450,input input_1451,input input_1452,input input_1453,input input_1454,input input_1455,input input_1456,input input_1457,input input_1458,input input_1459,input input_1460,input input_1461,input input_1462,input input_1463,input input_1464,input input_1465,input input_1466,input input_1467,input input_1468,input input_1469,input input_1470,input input_1471,input input_1472,input input_1473,input input_1474,input input_1475,input input_1476,input input_1477,input input_1478,input input_1479,input input_1480,input input_1481,input input_1482,input input_1483,input input_1484,input input_1485,input input_1486,input input_1487,input input_1488,input input_1489,input input_1490,input input_1491,input input_1492,input input_1493,input input_1494,input input_1495,input input_1496,input input_1497,input input_1498,input input_1499,input input_1500,input input_1501,input input_1502,input input_1503,input input_1504,input input_1505,input input_1506,input input_1507,input input_1508,input input_1509,input input_1510,input input_1511,input input_1512,input input_1513,input input_1514,input input_1515,input input_1516,input input_1517,input input_1518,input input_1519,input input_1520,input input_1521,input input_1522,input input_1523,input input_1524,input input_1525,input input_1526,input input_1527,input input_1528,input input_1529,input input_1530,input input_1531,input input_1532,input input_1533,input input_1534,input input_1535,input input_1536,input input_1537,input input_1538,input input_1539,input input_1540,input input_1541,input input_1542,input input_1543,input input_1544,input input_1545,input input_1546,input input_1547,input input_1548,input input_1549,input input_1550,input input_1551,input input_1552,input input_1553,input input_1554,input input_1555,input input_1556,input input_1557,input input_1558,input input_1559,input input_1560,input input_1561,input input_1562,input input_1563,input input_1564,input input_1565,input input_1566,input input_1567,input input_1568,input input_1569,input input_1570,input input_1571,input input_1572,input input_1573,input input_1574,input input_1575,input input_1576,input input_1577,input input_1578,input input_1579,input input_1580,input input_1581,input input_1582,input input_1583,input input_1584,input input_1585,input input_1586,input input_1587,input input_1588,input input_1589,input input_1590,input input_1591,input input_1592,input input_1593,input input_1594,input input_1595,input input_1596,input input_1597,input input_1598,input input_1599,input input_1600,input input_1601,input input_1602,input input_1603,input input_1604,input input_1605,input input_1606,input input_1607,input input_1608,input input_1609,input input_1610,input input_1611,input input_1612,input input_1613,input input_1614,input input_1615,input input_1616,input input_1617,input input_1618,input input_1619,input input_1620,input input_1621,input input_1622,input input_1623,input input_1624,input input_1625,input input_1626,input input_1627,input input_1628,input input_1629,input input_1630,input input_1631,input input_1632,input input_1633,input input_1634,input input_1635,input input_1636,input input_1637,input input_1638,input input_1639,input input_1640,input input_1641,input input_1642,input input_1643,input input_1644,input input_1645,input input_1646,input input_1647,input input_1648,input input_1649,input input_1650,input input_1651,input input_1652,input input_1653,input input_1654,input input_1655,input input_1656,input input_1657,input input_1658,input input_1659,input input_1660,input input_1661,input input_1662,input input_1663,input input_1664,input input_1665,input input_1666,input input_1667,input input_1668,input input_1669,input input_1670,input input_1671,input input_1672,input input_1673,input input_1674,input input_1675,input input_1676,input input_1677,input input_1678,input input_1679,input input_1680,input input_1681,input input_1682,input input_1683,input input_1684,input input_1685,input input_1686,input input_1687,input input_1688,input input_1689,input input_1690,input input_1691,input input_1692,input input_1693,input input_1694,input input_1695,input input_1696,input input_1697,input input_1698,input input_1699,input input_1700,input input_1701,input input_1702,input input_1703,input input_1704,input input_1705,input input_1706,input input_1707,input input_1708,input input_1709,input input_1710,input input_1711,input input_1712,input input_1713,input input_1714,input input_1715,input input_1716,input input_1717,input input_1718,input input_1719,input input_1720,input input_1721,input input_1722,input input_1723,input input_1724,input input_1725,input input_1726,input input_1727,input input_1728,input input_1729,input input_1730,input input_1731,input input_1732,input input_1733,input input_1734,input input_1735,input input_1736,input input_1737,input input_1738,input input_1739,input input_1740,input input_1741,input input_1742,input input_1743,input input_1744,input input_1745,input input_1746,input input_1747,input input_1748,input input_1749,input input_1750,input input_1751,input input_1752,input input_1753,input input_1754,input input_1755,input input_1756,input input_1757,input input_1758,input input_1759,input input_1760,input input_1761,input input_1762,input input_1763,input input_1764,input input_1765,input input_1766,input input_1767,input input_1768,input input_1769,input input_1770,input input_1771,input input_1772,input input_1773,input input_1774,input input_1775,input input_1776,input input_1777,input input_1778,input input_1779,input input_1780,input input_1781,input input_1782,input input_1783,input input_1784,input input_1785,input input_1786,input input_1787,input input_1788,input input_1789,input input_1790,input input_1791,input input_1792,input input_1793,input input_1794,input input_1795,input input_1796,input input_1797,input input_1798,input input_1799,input input_1800,input input_1801,input input_1802,input input_1803,input input_1804,input input_1805,input input_1806,input input_1807,input input_1808,input input_1809,input input_1810,input input_1811,input input_1812,input input_1813,input input_1814,input input_1815,input input_1816,input input_1817,input input_1818,input input_1819,input input_1820,input input_1821,input input_1822,input input_1823,input input_1824,input input_1825,input input_1826,input input_1827,input input_1828,input input_1829,input input_1830,input input_1831,input input_1832,input input_1833,input input_1834,input input_1835,input input_1836,input input_1837,input input_1838,input input_1839,input input_1840,input input_1841,input input_1842,input input_1843,input input_1844,input input_1845,input input_1846,input input_1847,input input_1848,input input_1849,input input_1850,input input_1851,input input_1852,input input_1853,input input_1854,input input_1855,input input_1856,input input_1857,input input_1858,input input_1859,input input_1860,input input_1861,input input_1862,input input_1863,input input_1864,input input_1865,input input_1866,input input_1867,input input_1868,input input_1869,input input_1870,input input_1871,input input_1872,input input_1873,input input_1874,input input_1875,input input_1876,input input_1877,input input_1878,input input_1879,input input_1880,input input_1881,input input_1882,input input_1883,input input_1884,input input_1885,input input_1886,input input_1887,input input_1888,input input_1889,input input_1890,input input_1891,input input_1892,input input_1893,input input_1894,input input_1895,input input_1896,input input_1897,input input_1898,input input_1899,input input_1900,input input_1901,input input_1902,input input_1903,input input_1904,input input_1905,input input_1906,input input_1907,input input_1908,input input_1909,input input_1910,input input_1911,input input_1912,input input_1913,input input_1914,input input_1915,input input_1916,input input_1917,input input_1918,input input_1919,input input_1920,input input_1921,input input_1922,input input_1923,input input_1924,input input_1925,input input_1926,input input_1927,input input_1928,input input_1929,input input_1930,input input_1931,input input_1932,input input_1933,input input_1934,input input_1935,input input_1936,input input_1937,input input_1938,input input_1939,input input_1940,input input_1941,input input_1942,input input_1943,input input_1944,input input_1945,input input_1946,input input_1947,input input_1948,input input_1949,input input_1950,input input_1951,input input_1952,input input_1953,input input_1954,input input_1955,input input_1956,input input_1957,input input_1958,input input_1959,input input_1960,input input_1961,input input_1962,input input_1963,input input_1964,input input_1965,input input_1966,input input_1967,input input_1968,input input_1969,input input_1970,input input_1971,input input_1972,input input_1973,input input_1974,input input_1975,input input_1976,input input_1977,input input_1978,input input_1979,input input_1980,input input_1981,input input_1982,input input_1983,input input_1984,input input_1985,input input_1986,input input_1987,input input_1988,input input_1989,input input_1990,input input_1991,input input_1992,input input_1993,input input_1994,input input_1995,input input_1996,input input_1997,input input_1998,input input_1999,input input_2000,input input_2001,input input_2002,input input_2003,input input_2004,input input_2005,input input_2006,input input_2007,input input_2008,input input_2009,input input_2010,input input_2011,input input_2012,input input_2013,input input_2014,input input_2015,input input_2016,input input_2017,input input_2018,input input_2019,input input_2020,input input_2021,input input_2022,input input_2023,input input_2024,input input_2025,input input_2026,input input_2027,input input_2028,input input_2029,input input_2030,input input_2031,input input_2032,input input_2033,input input_2034,input input_2035,input input_2036,input input_2037,input input_2038,input input_2039,input input_2040,input input_2041,input input_2042,input input_2043,input input_2044,input input_2045,input input_2046,input input_2047,input input_2048,input input_2049,input input_2050,input input_2051,input input_2052,input input_2053,input input_2054,input input_2055,input input_2056,input input_2057,input input_2058,input input_2059,input input_2060,input input_2061,input input_2062,input input_2063,input input_2064,input input_2065,input input_2066,input input_2067,input input_2068,input input_2069,input input_2070,input input_2071,input input_2072,input input_2073,input input_2074,input input_2075,input input_2076,input input_2077,input input_2078,input input_2079,input input_2080,input input_2081,input input_2082,input input_2083,input input_2084,input input_2085,input input_2086,input input_2087,input input_2088,input input_2089,input input_2090,input input_2091,input input_2092,input input_2093,input input_2094,input input_2095,input input_2096,input input_2097,input input_2098,input input_2099,input input_2100,input input_2101,input input_2102,input input_2103,input input_2104,input input_2105,input input_2106,input input_2107,input input_2108,input input_2109,input input_2110,input input_2111,input input_2112,input input_2113,input input_2114,input input_2115,input input_2116,input input_2117,input input_2118,input input_2119,input input_2120,input input_2121,input input_2122,input input_2123,input input_2124,input input_2125,input input_2126,input input_2127,input input_2128,input input_2129,input input_2130,input input_2131,input input_2132,input input_2133,input input_2134,input input_2135,input input_2136,input input_2137,input input_2138,input input_2139,input input_2140,input input_2141,input input_2142,input input_2143,input input_2144,input input_2145,input input_2146,input input_2147,input input_2148,input input_2149,input input_2150,input input_2151,input input_2152,input input_2153,input input_2154,input input_2155,input input_2156,input input_2157,input input_2158,input input_2159,input input_2160,input input_2161,input input_2162,input input_2163,input input_2164,input input_2165,input input_2166,input input_2167,input input_2168,input input_2169,input input_2170,input input_2171,input input_2172,input input_2173,input input_2174,input input_2175,input input_2176,input input_2177,input input_2178,input input_2179,input input_2180,input input_2181,input input_2182,input input_2183,input input_2184,input input_2185,input input_2186,input input_2187,input input_2188,input input_2189,input input_2190,input input_2191,input input_2192,input input_2193,input input_2194,input input_2195,input input_2196,input input_2197,input input_2198,input input_2199,input input_2200,input input_2201,input input_2202,input input_2203,input input_2204,input input_2205,input input_2206,input input_2207,input input_2208,input input_2209,input input_2210,input input_2211,input input_2212,input input_2213,input input_2214,input input_2215,input input_2216,input input_2217,input input_2218,input input_2219,input input_2220,input input_2221,input input_2222,input input_2223,input input_2224,input input_2225,input input_2226,input input_2227,input input_2228,input input_2229,input input_2230,input input_2231,input input_2232,input input_2233,input input_2234,input input_2235,input input_2236,input input_2237,input input_2238,input input_2239,input input_2240,input input_2241,input input_2242,input input_2243,input input_2244,input input_2245,input input_2246,input input_2247,input input_2248,input input_2249,input input_2250,input input_2251,input input_2252,input input_2253,input input_2254,input input_2255,input input_2256,input input_2257,input input_2258,input input_2259,input input_2260,input input_2261,input input_2262,input input_2263,input input_2264,input input_2265,input input_2266,input input_2267,input input_2268,input input_2269,input input_2270,input input_2271,input input_2272,input input_2273,input input_2274,input input_2275,input input_2276,input input_2277,input input_2278,input input_2279,input input_2280,input input_2281,input input_2282,input input_2283,input input_2284,input input_2285,input input_2286,input input_2287,input input_2288,input input_2289,input input_2290,input input_2291,input input_2292,input input_2293,input input_2294,input input_2295,input input_2296,input input_2297,input input_2298,input input_2299,input input_2300,input input_2301,input input_2302,input input_2303,input input_2304,input input_2305,input input_2306,input input_2307,input input_2308,input input_2309,input input_2310,input input_2311,input input_2312,input input_2313,input input_2314,input input_2315,input input_2316,input input_2317,input input_2318,input input_2319,input input_2320,input input_2321,input input_2322,input input_2323,input input_2324,input input_2325,input input_2326,input input_2327,input input_2328,input input_2329,input input_2330,input input_2331,input input_2332,input input_2333,input input_2334,input input_2335,input input_2336,input input_2337,input input_2338,input input_2339,input input_2340,input input_2341,input input_2342,input input_2343,input input_2344,input input_2345,input input_2346,input input_2347,input input_2348,input input_2349,input input_2350,input input_2351,input input_2352,input input_2353,input input_2354,input input_2355,input input_2356,input input_2357,input input_2358,input input_2359,input input_2360,input input_2361,input input_2362,input input_2363,input input_2364,input input_2365,input input_2366,input input_2367,input input_2368,input input_2369,input input_2370,input input_2371,input input_2372,input input_2373,input input_2374,input input_2375,input input_2376,input input_2377,input input_2378,input input_2379,input input_2380,input input_2381,input input_2382,input input_2383,input input_2384,input input_2385,input input_2386,input input_2387,input input_2388,input input_2389,input input_2390,input input_2391,input input_2392,input input_2393,input input_2394,input input_2395,input input_2396,input input_2397,input input_2398,input input_2399,input input_2400,input input_2401,input input_2402,input input_2403,input input_2404,input input_2405,input input_2406,input input_2407,input input_2408,input input_2409,input input_2410,input input_2411,input input_2412,input input_2413,input input_2414,input input_2415,input input_2416,input input_2417,input input_2418,input input_2419,input input_2420,input input_2421,input input_2422,input input_2423,input input_2424,input input_2425,input input_2426,input input_2427,input input_2428,input input_2429,input input_2430,input input_2431,input input_2432,input input_2433,input input_2434,input input_2435,input input_2436,input input_2437,input input_2438,input input_2439,input input_2440,input input_2441,input input_2442,input input_2443,input input_2444,input input_2445,input input_2446,input input_2447,input input_2448,input input_2449,input input_2450,input input_2451,input input_2452,input input_2453,input input_2454,input input_2455,input input_2456,input input_2457,input input_2458,input input_2459,input input_2460,input input_2461,input input_2462,input input_2463,input input_2464,input input_2465,input input_2466,input input_2467,input input_2468,input input_2469,input input_2470,input input_2471,input input_2472,input input_2473,input input_2474,input input_2475,input input_2476,input input_2477,input input_2478,input input_2479,input input_2480,input input_2481,input input_2482,input input_2483,input input_2484,input input_2485,input input_2486,input input_2487,input input_2488,input input_2489,input input_2490,input input_2491,input input_2492,input input_2493,input input_2494,input input_2495,input input_2496,input input_2497,input input_2498,input input_2499,input input_2500,input input_2501,input input_2502,input input_2503,input input_2504,input input_2505,input input_2506,input input_2507,input input_2508,input input_2509,input input_2510,input input_2511,input input_2512,input input_2513,input input_2514,input input_2515,input input_2516,input input_2517,input input_2518,input input_2519,input input_2520,input input_2521,input input_2522,input input_2523,input input_2524,input input_2525,input input_2526,input input_2527,input input_2528,input input_2529,input input_2530,input input_2531,input input_2532,input input_2533,input input_2534,input input_2535,input input_2536,input input_2537,input input_2538,input input_2539,input input_2540,input input_2541,input input_2542,input input_2543,input input_2544,input input_2545,input input_2546,input input_2547,input input_2548,input input_2549,input input_2550,input input_2551,input input_2552,input input_2553,input input_2554,input input_2555,input input_2556,input input_2557,input input_2558,input input_2559,input input_2560,input input_2561,input input_2562,input input_2563,input input_2564,input input_2565,input input_2566,input input_2567,input input_2568,input input_2569,input input_2570,input input_2571,input input_2572,input input_2573,input input_2574,input input_2575,input input_2576,input input_2577,input input_2578,input input_2579,input input_2580,input input_2581,input input_2582,input input_2583,input input_2584,input input_2585,input input_2586,input input_2587,input input_2588,input input_2589,input input_2590,input input_2591,input input_2592,input input_2593,input input_2594,input input_2595,input input_2596,input input_2597,input input_2598,input input_2599,input input_2600,input input_2601,input input_2602,input input_2603,input input_2604,input input_2605,input input_2606,input input_2607,input input_2608,input input_2609,input input_2610,input input_2611,input input_2612,input input_2613,input input_2614,input input_2615,input input_2616,input input_2617,input input_2618,input input_2619,input input_2620,input input_2621,input input_2622,input input_2623,input input_2624,input input_2625,input input_2626,input input_2627,input input_2628,input input_2629,input input_2630,input input_2631,input input_2632,input input_2633,input input_2634,input input_2635,input input_2636,input input_2637,input input_2638,input input_2639,input input_2640,input input_2641,input input_2642,input input_2643,input input_2644,input input_2645,input input_2646,input input_2647,input input_2648,input input_2649,input input_2650,input input_2651,input input_2652,input input_2653,input input_2654,input input_2655,input input_2656,input input_2657,input input_2658,input input_2659,input input_2660,input input_2661,input input_2662,input input_2663,input input_2664,input input_2665,input input_2666,input input_2667,input input_2668,input input_2669,input input_2670,input input_2671,input input_2672,input input_2673,input input_2674,input input_2675,input input_2676,input input_2677,input input_2678,input input_2679,input input_2680,input input_2681,input input_2682,input input_2683,input input_2684,input input_2685,input input_2686,input input_2687,input input_2688,input input_2689,input input_2690,input input_2691,input input_2692,input input_2693,input input_2694,input input_2695,input input_2696,input input_2697,input input_2698,input input_2699,input input_2700,input input_2701,input input_2702,input input_2703,input input_2704,input input_2705,input input_2706,input input_2707,input input_2708,input input_2709,input input_2710,input input_2711,input input_2712,input input_2713,input input_2714,input input_2715,input input_2716,input input_2717,input input_2718,input input_2719,input input_2720,input input_2721,input input_2722,input input_2723,input input_2724,input input_2725,input input_2726,input input_2727,input input_2728,input input_2729,input input_2730,input input_2731,input input_2732,input input_2733,input input_2734,input input_2735,input input_2736,input input_2737,input input_2738,input input_2739,input input_2740,input input_2741,input input_2742,input input_2743,input input_2744,input input_2745,input input_2746,input input_2747,input input_2748,input input_2749,input input_2750,input input_2751,input input_2752,input input_2753,input input_2754,input input_2755,input input_2756,input input_2757,input input_2758,input input_2759,input input_2760,input input_2761,input input_2762,input input_2763,input input_2764,input input_2765,input input_2766,input input_2767,input input_2768,input input_2769,input input_2770,input input_2771,input input_2772,input input_2773,input input_2774,input input_2775,input input_2776,input input_2777,input input_2778,input input_2779,input input_2780,input input_2781,input input_2782,input input_2783,input input_2784,input input_2785,input input_2786,input input_2787,input input_2788,input input_2789,input input_2790,input input_2791,input input_2792,input input_2793,input input_2794,input input_2795,input input_2796,input input_2797,input input_2798,input input_2799,input input_2800,input input_2801,input input_2802,input input_2803,input input_2804,input input_2805,input input_2806,input input_2807,input input_2808,input input_2809,input input_2810,input input_2811,input input_2812,input input_2813,input input_2814,input input_2815,input input_2816,input input_2817,input input_2818,input input_2819,input input_2820,input input_2821,input input_2822,input input_2823,input input_2824,input input_2825,input input_2826,input input_2827,input input_2828,input input_2829,input input_2830,input input_2831,input input_2832,input input_2833,input input_2834,input input_2835,input input_2836,input input_2837,input input_2838,input input_2839,input input_2840,input input_2841,input input_2842,input input_2843,input input_2844,input input_2845,input input_2846,input input_2847,input input_2848,input input_2849,input input_2850,input input_2851,input input_2852,input input_2853,input input_2854,input input_2855,input input_2856,input input_2857,input input_2858,input input_2859,input input_2860,input input_2861,input input_2862,input input_2863,input input_2864,input input_2865,input input_2866,input input_2867,input input_2868,input input_2869,input input_2870,input input_2871,input input_2872,input input_2873,input input_2874,input input_2875,input input_2876,input input_2877,input input_2878,input input_2879,input input_2880,input input_2881,input input_2882,input input_2883,input input_2884,input input_2885,input input_2886,input input_2887,input input_2888,input input_2889,input input_2890,input input_2891,input input_2892,input input_2893,input input_2894,input input_2895,input input_2896,input input_2897,input input_2898,input input_2899,input input_2900,input input_2901,input input_2902,input input_2903,input input_2904,input input_2905,input input_2906,input input_2907,input input_2908,input input_2909,input input_2910,input input_2911,input input_2912,input input_2913,input input_2914,input input_2915,input input_2916,input input_2917,input input_2918,input input_2919,input input_2920,input input_2921,input input_2922,input input_2923,input input_2924,input input_2925,input input_2926,input input_2927,input input_2928,input input_2929,input input_2930,input input_2931,input input_2932,input input_2933,input input_2934,input input_2935,input input_2936,input input_2937,input input_2938,input input_2939,input input_2940,input input_2941,input input_2942,input input_2943,input input_2944,input input_2945,input input_2946,input input_2947,input input_2948,input input_2949,input input_2950,input input_2951,input input_2952,input input_2953,input input_2954,input input_2955,input input_2956,input input_2957,input input_2958,input input_2959,input input_2960,input input_2961,input input_2962,input input_2963,input input_2964,input input_2965,input input_2966,input input_2967,input input_2968,input input_2969,input input_2970,input input_2971,input input_2972,input input_2973,input input_2974,input input_2975,input input_2976,input input_2977,input input_2978,input input_2979,input input_2980,input input_2981,input input_2982,input input_2983,input input_2984,input input_2985,input input_2986,input input_2987,input input_2988,input input_2989,input input_2990,input input_2991,input input_2992,input input_2993,input input_2994,input input_2995,input input_2996,input input_2997,input input_2998,input input_2999,input input_3000,input input_3001,input input_3002,input input_3003,input input_3004,input input_3005,input input_3006,input input_3007,input input_3008,input input_3009,input input_3010,input input_3011,input input_3012,input input_3013,input input_3014,input input_3015,input input_3016,input input_3017,input input_3018,input input_3019,input input_3020,input input_3021,input input_3022,input input_3023,input input_3024,input input_3025,input input_3026,input input_3027,input input_3028,input input_3029,input input_3030,input input_3031,input input_3032,input input_3033,input input_3034,input input_3035,input input_3036,input input_3037,input input_3038,input input_3039,input input_3040,input input_3041,input input_3042,input input_3043,input input_3044,input input_3045,input input_3046,input input_3047,input input_3048,input input_3049,input input_3050,input input_3051,input input_3052,input input_3053,input input_3054,input input_3055,input input_3056,input input_3057,input input_3058,input input_3059,input input_3060,input input_3061,input input_3062,input input_3063,input input_3064,input input_3065,input input_3066,input input_3067,input input_3068,input input_3069,input input_3070,input input_3071,input input_3072,input input_3073,input input_3074,input input_3075,input input_3076,input input_3077,input input_3078,input input_3079,input input_3080,input input_3081,input input_3082,input input_3083,input input_3084,input input_3085,input input_3086,input input_3087,input input_3088,input input_3089,input input_3090,input input_3091,input input_3092,input input_3093,input input_3094,input input_3095,input input_3096,input input_3097,input input_3098,input input_3099,input input_3100,input input_3101,input input_3102,input input_3103,input input_3104,input input_3105,input input_3106,input input_3107,input input_3108,input input_3109,input input_3110,input input_3111,input input_3112,input input_3113,input input_3114,input input_3115,input input_3116,input input_3117,input input_3118,input input_3119,input input_3120,input input_3121,input input_3122,input input_3123,input input_3124,input input_3125,input input_3126,input input_3127,input input_3128,input input_3129,input input_3130,input input_3131,input input_3132,input input_3133,input input_3134,input input_3135,input input_3136,input input_3137,input input_3138,input input_3139,input input_3140,input input_3141,input input_3142,input input_3143,input input_3144,input input_3145,input input_3146,input input_3147,input input_3148,input input_3149,input input_3150,input input_3151,input input_3152,input input_3153,input input_3154,input input_3155,input input_3156,input input_3157,input input_3158,input input_3159,input input_3160,input input_3161,input input_3162,input input_3163,input input_3164,input input_3165,input input_3166,input input_3167,input input_3168,input input_3169,input input_3170,input input_3171,input input_3172,input input_3173,input input_3174,input input_3175,input input_3176,input input_3177,input input_3178,input input_3179,input input_3180,input input_3181,input input_3182,input input_3183,input input_3184,input input_3185,input input_3186,input input_3187,input input_3188,input input_3189,input input_3190,input input_3191,input input_3192,input input_3193,input input_3194,input input_3195,input input_3196,input input_3197,input input_3198,input input_3199,input input_3200,input input_3201,input input_3202,input input_3203,input input_3204,input input_3205,input input_3206,input input_3207,input input_3208,input input_3209,input input_3210,input input_3211,input input_3212,input input_3213,input input_3214,input input_3215,input input_3216,input input_3217,input input_3218,input input_3219,input input_3220,input input_3221,input input_3222,input input_3223,input input_3224,input input_3225,input input_3226,input input_3227,input input_3228,input input_3229,input input_3230,input input_3231,input input_3232,input input_3233,input input_3234,input input_3235,input input_3236,input input_3237,input input_3238,input input_3239,input input_3240,input input_3241,input input_3242,input input_3243,input input_3244,input input_3245,input input_3246,input input_3247,input input_3248,input input_3249,input input_3250,input input_3251,input input_3252,input input_3253,input input_3254,input input_3255,input input_3256,input input_3257,input input_3258,input input_3259,input input_3260,input input_3261,input input_3262,input input_3263,input input_3264,input input_3265,input input_3266,input input_3267,input input_3268,input input_3269,input input_3270,input input_3271,input input_3272,input input_3273,input input_3274,input input_3275,input input_3276,input input_3277,input input_3278,input input_3279,input input_3280,input input_3281,input input_3282,input input_3283,input input_3284,input input_3285,input input_3286,input input_3287,input input_3288,input input_3289,input input_3290,input input_3291,input input_3292,input input_3293,input input_3294,input input_3295,input input_3296,input input_3297,input input_3298,input input_3299,input input_3300,input input_3301,input input_3302,input input_3303,input input_3304,input input_3305,input input_3306,input input_3307,input input_3308,input input_3309,input input_3310,input input_3311,input input_3312,input input_3313,input input_3314,input input_3315,input input_3316,input input_3317,input input_3318,input input_3319,input input_3320,input input_3321,input input_3322,input input_3323,input input_3324,input input_3325,input input_3326,input input_3327,input input_3328,input input_3329,input input_3330,input input_3331,input input_3332,input input_3333,input input_3334,input input_3335,input input_3336,input input_3337,input input_3338,input input_3339,input input_3340,input input_3341,input input_3342,input input_3343,input input_3344,input input_3345,input input_3346,input input_3347,input input_3348,input input_3349,input input_3350,input input_3351,input input_3352,input input_3353,input input_3354,input input_3355,input input_3356,input input_3357,input input_3358,input input_3359,input input_3360,input input_3361,input input_3362,input input_3363,input input_3364,input input_3365,input input_3366,input input_3367,input input_3368,input input_3369,input input_3370,input input_3371,input input_3372,input input_3373,input input_3374,input input_3375,input input_3376,input input_3377,input input_3378,input input_3379,input input_3380,input input_3381,input input_3382,input input_3383,input input_3384,input input_3385,input input_3386,input input_3387,input input_3388,input input_3389,input input_3390,input input_3391,input input_3392,input input_3393,input input_3394,input input_3395,input input_3396,input input_3397,input input_3398,input input_3399,input input_3400,input input_3401,input input_3402,input input_3403,input input_3404,input input_3405,input input_3406,input input_3407,input input_3408,input input_3409,input input_3410,input input_3411,input input_3412,input input_3413,input input_3414,input input_3415,input input_3416,input input_3417,input input_3418,input input_3419,input input_3420,input input_3421,input input_3422,input input_3423,input input_3424,input input_3425,input input_3426,input input_3427,input input_3428,input input_3429,input input_3430,input input_3431,input input_3432,input input_3433,input input_3434,input input_3435,input input_3436,input input_3437,input input_3438,input input_3439,input input_3440,input input_3441,input input_3442,input input_3443,input input_3444,input input_3445,input input_3446,input input_3447,input input_3448,input input_3449,input input_3450,input input_3451,input input_3452,input input_3453,input input_3454,input input_3455,input input_3456,input input_3457,input input_3458,input input_3459,input input_3460,input input_3461,input input_3462,input input_3463,input input_3464,input input_3465,input input_3466,input input_3467,input input_3468,input input_3469,input input_3470,input input_3471,input input_3472,input input_3473,input input_3474,input input_3475,input input_3476,input input_3477,input input_3478,input input_3479,input input_3480,input input_3481,input input_3482,input input_3483,input input_3484,input input_3485,input input_3486,input input_3487,input input_3488,input input_3489,input input_3490,input input_3491,input input_3492,input input_3493,input input_3494,input input_3495,input input_3496,input input_3497,input input_3498,input input_3499,input input_3500,input input_3501,input input_3502,input input_3503,input input_3504,input input_3505,input input_3506,input input_3507,input input_3508,input input_3509,input input_3510,input input_3511,input input_3512,input input_3513,input input_3514,input input_3515,input input_3516,input input_3517,input input_3518,input input_3519,input input_3520,input input_3521,input input_3522,input input_3523,input input_3524,input input_3525,input input_3526,input input_3527,input input_3528,input input_3529,input input_3530,input input_3531,input input_3532,input input_3533,input input_3534,input input_3535,input input_3536,input input_3537,input input_3538,input input_3539,input input_3540,input input_3541,input input_3542,input input_3543,input input_3544,input input_3545,input input_3546,input input_3547,input input_3548,input input_3549,input input_3550,input input_3551,input input_3552,input input_3553,input input_3554,input input_3555,input input_3556,input input_3557,input input_3558,input input_3559,input input_3560,input input_3561,input input_3562,input input_3563,input input_3564,input input_3565,input input_3566,input input_3567,input input_3568,input input_3569,input input_3570,input input_3571,input input_3572,input input_3573,input input_3574,input input_3575,input input_3576,input input_3577,input input_3578,input input_3579,input input_3580,input input_3581,input input_3582,input input_3583,input input_3584,input input_3585,input input_3586,input input_3587,input input_3588,input input_3589,input input_3590,input input_3591,input input_3592,input input_3593,input input_3594,input input_3595,input input_3596,input input_3597,input input_3598,input input_3599,input input_3600,input input_3601,input input_3602,input input_3603,input input_3604,input input_3605,input input_3606,input input_3607,input input_3608,input input_3609,input input_3610,input input_3611,input input_3612,input input_3613,input input_3614,input input_3615,input input_3616,input input_3617,input input_3618,input input_3619,input input_3620,input input_3621,input input_3622,input input_3623,input input_3624,input input_3625,input input_3626,input input_3627,input input_3628,input input_3629,input input_3630,input input_3631,input input_3632,input input_3633,input input_3634,input input_3635,input input_3636,input input_3637,input input_3638,input input_3639,input input_3640,input input_3641,input input_3642,input input_3643,input input_3644,input input_3645,input input_3646,input input_3647,input input_3648,input input_3649,input input_3650,input input_3651,input input_3652,input input_3653,input input_3654,input input_3655,input input_3656,input input_3657,input input_3658,input input_3659,input input_3660,input input_3661,input input_3662,input input_3663,input input_3664,input input_3665,input input_3666,input input_3667,input input_3668,input input_3669,input input_3670,input input_3671,input input_3672,input input_3673,input input_3674,input input_3675,input input_3676,input input_3677,input input_3678,input input_3679,input input_3680,input input_3681,input input_3682,input input_3683,input input_3684,input input_3685,input input_3686,input input_3687,input input_3688,input input_3689,input input_3690,input input_3691,input input_3692,input input_3693,input input_3694,input input_3695,input input_3696,input input_3697,input input_3698,input input_3699,input input_3700,input input_3701,input input_3702,input input_3703,input input_3704,input input_3705,input input_3706,input input_3707,input input_3708,input input_3709,input input_3710,input input_3711,input input_3712,input input_3713,input input_3714,input input_3715,input input_3716,input input_3717,input input_3718,input input_3719,input input_3720,input input_3721,input input_3722,input input_3723,input input_3724,input input_3725,input input_3726,input input_3727,input input_3728,input input_3729,input input_3730,input input_3731,input input_3732,input input_3733,input input_3734,input input_3735,input input_3736,input input_3737,input input_3738,input input_3739,input input_3740,input input_3741,input input_3742,input input_3743,input input_3744,input input_3745,input input_3746,input input_3747,input input_3748,input input_3749,input input_3750,input input_3751,input input_3752,input input_3753,input input_3754,input input_3755,input input_3756,input input_3757,input input_3758,input input_3759,input input_3760,input input_3761,input input_3762,input input_3763,input input_3764,input input_3765,input input_3766,input input_3767,input input_3768,input input_3769,input input_3770,input input_3771,input input_3772,input input_3773,input input_3774,input input_3775,input input_3776,input input_3777,input input_3778,input input_3779,input input_3780,input input_3781,input input_3782,input input_3783,input input_3784,input input_3785,input input_3786,input input_3787,input input_3788,input input_3789,input input_3790,input input_3791,input input_3792,input input_3793,input input_3794,input input_3795,input input_3796,input input_3797,input input_3798,input input_3799,input input_3800,input input_3801,input input_3802,input input_3803,input input_3804,input input_3805,input input_3806,input input_3807,input input_3808,input input_3809,input input_3810,input input_3811,input input_3812,input input_3813,input input_3814,input input_3815,input input_3816,input input_3817,input input_3818,input input_3819,input input_3820,input input_3821,input input_3822,input input_3823,input input_3824,input input_3825,input input_3826,input input_3827,input input_3828,input input_3829,input input_3830,input input_3831,input input_3832,input input_3833,input input_3834,input input_3835,input input_3836,input input_3837,input input_3838,input input_3839,input input_3840,input input_3841,input input_3842,input input_3843,input input_3844,input input_3845,input input_3846,input input_3847,input input_3848,input input_3849,input input_3850,input input_3851,input input_3852,input input_3853,input input_3854,input input_3855,input input_3856,input input_3857,input input_3858,input input_3859,input input_3860,input input_3861,input input_3862,input input_3863,input input_3864,input input_3865,input input_3866,input input_3867,input input_3868,input input_3869,input input_3870,input input_3871,input input_3872,input input_3873,input input_3874,input input_3875,input input_3876,input input_3877,input input_3878,input input_3879,input input_3880,input input_3881,input input_3882,input input_3883,input input_3884,input input_3885,input input_3886,input input_3887,input input_3888,input input_3889,input input_3890,input input_3891,input input_3892,input input_3893,input input_3894,input input_3895,input input_3896,input input_3897,input input_3898,input input_3899,input input_3900,input input_3901,input input_3902,input input_3903,input input_3904,input input_3905,input input_3906,input input_3907,input input_3908,input input_3909,input input_3910,input input_3911,input input_3912,input input_3913,input input_3914,input input_3915,input input_3916,input input_3917,input input_3918,input input_3919,input input_3920,input input_3921,input input_3922,input input_3923,input input_3924,input input_3925,input input_3926,input input_3927,input input_3928,input input_3929,input input_3930,input input_3931,input input_3932,input input_3933,input input_3934,input input_3935,input input_3936,input input_3937,input input_3938,input input_3939,input input_3940,input input_3941,input input_3942,input input_3943,input input_3944,input input_3945,input input_3946,input input_3947,input input_3948,input input_3949,input input_3950,input input_3951,input input_3952,input input_3953,input input_3954,input input_3955,input input_3956,input input_3957,input input_3958,input input_3959,input input_3960,input input_3961,input input_3962,input input_3963,input input_3964,input input_3965,input input_3966,input input_3967,input input_3968,input input_3969,input input_3970,input input_3971,input input_3972,input input_3973,input input_3974,input input_3975,input input_3976,input input_3977,input input_3978,input input_3979,input input_3980,input input_3981,input input_3982,input input_3983,input input_3984,input input_3985,input input_3986,input input_3987,input input_3988,input input_3989,input input_3990,input input_3991,input input_3992,input input_3993,input input_3994,input input_3995,input input_3996,input input_3997,input input_3998,input input_3999,input input_4000,input input_4001,input input_4002,input input_4003,input input_4004,input input_4005,input input_4006,input input_4007,input input_4008,input input_4009,input input_4010,input input_4011,input input_4012,input input_4013,input input_4014,input input_4015,input input_4016,input input_4017,input input_4018,input input_4019,input input_4020,input input_4021,input input_4022,input input_4023,input input_4024,input input_4025,input input_4026,input input_4027,input input_4028,input input_4029,input input_4030,input input_4031,input input_4032,input input_4033,input input_4034,input input_4035,input input_4036,input input_4037,input input_4038,input input_4039,input input_4040,input input_4041,input input_4042,input input_4043,input input_4044,input input_4045,input input_4046,input input_4047,input input_4048,input input_4049,input input_4050,input input_4051,input input_4052,input input_4053,input input_4054,input input_4055,input input_4056,input input_4057,input input_4058,input input_4059,input input_4060,input input_4061,input input_4062,input input_4063,input input_4064,input input_4065,input input_4066,input input_4067,input input_4068,input input_4069,input input_4070,input input_4071,input input_4072,input input_4073,input input_4074,input input_4075,input input_4076,input input_4077,input input_4078,input input_4079,input input_4080,input input_4081,input input_4082,input input_4083,input input_4084,input input_4085,input input_4086,input input_4087,input input_4088,input input_4089,input input_4090,input input_4091,input input_4092,input input_4093,input input_4094,input input_4095
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_000000 (.a(t0_0000000), .b(t0_0000001), .y(t0_000000));
wire t0_0000000, t0_0000001;
mixer mix_t0_0000000 (.a(t0_00000000), .b(t0_00000001), .y(t0_0000000));
wire t0_00000000, t0_00000001;
mixer mix_t0_00000000 (.a(t0_000000000), .b(t0_000000001), .y(t0_00000000));
wire t0_000000000, t0_000000001;
mixer mix_t0_000000000 (.a(t0_0000000000), .b(t0_0000000001), .y(t0_000000000));
wire t0_0000000000, t0_0000000001;
mixer mix_t0_0000000000 (.a(t0_00000000000), .b(t0_00000000001), .y(t0_0000000000));
wire t0_00000000000, t0_00000000001;
mixer mix_t0_00000000000 (.a(t0_000000000000), .b(t0_000000000001), .y(t0_00000000000));
wire t0_000000000000, t0_000000000001;
mixer mix_t0_000000000000 (.a(t0_0000000000000), .b(t0_0000000000001), .y(t0_000000000000));
wire t0_0000000000000, t0_0000000000001;
mixer mix_t0_000000000001 (.a(t0_0000000000010), .b(t0_0000000000011), .y(t0_000000000001));
wire t0_0000000000010, t0_0000000000011;
mixer mix_t0_00000000001 (.a(t0_000000000010), .b(t0_000000000011), .y(t0_00000000001));
wire t0_000000000010, t0_000000000011;
mixer mix_t0_000000000010 (.a(t0_0000000000100), .b(t0_0000000000101), .y(t0_000000000010));
wire t0_0000000000100, t0_0000000000101;
mixer mix_t0_000000000011 (.a(t0_0000000000110), .b(t0_0000000000111), .y(t0_000000000011));
wire t0_0000000000110, t0_0000000000111;
mixer mix_t0_0000000001 (.a(t0_00000000010), .b(t0_00000000011), .y(t0_0000000001));
wire t0_00000000010, t0_00000000011;
mixer mix_t0_00000000010 (.a(t0_000000000100), .b(t0_000000000101), .y(t0_00000000010));
wire t0_000000000100, t0_000000000101;
mixer mix_t0_000000000100 (.a(t0_0000000001000), .b(t0_0000000001001), .y(t0_000000000100));
wire t0_0000000001000, t0_0000000001001;
mixer mix_t0_000000000101 (.a(t0_0000000001010), .b(t0_0000000001011), .y(t0_000000000101));
wire t0_0000000001010, t0_0000000001011;
mixer mix_t0_00000000011 (.a(t0_000000000110), .b(t0_000000000111), .y(t0_00000000011));
wire t0_000000000110, t0_000000000111;
mixer mix_t0_000000000110 (.a(t0_0000000001100), .b(t0_0000000001101), .y(t0_000000000110));
wire t0_0000000001100, t0_0000000001101;
mixer mix_t0_000000000111 (.a(t0_0000000001110), .b(t0_0000000001111), .y(t0_000000000111));
wire t0_0000000001110, t0_0000000001111;
mixer mix_t0_000000001 (.a(t0_0000000010), .b(t0_0000000011), .y(t0_000000001));
wire t0_0000000010, t0_0000000011;
mixer mix_t0_0000000010 (.a(t0_00000000100), .b(t0_00000000101), .y(t0_0000000010));
wire t0_00000000100, t0_00000000101;
mixer mix_t0_00000000100 (.a(t0_000000001000), .b(t0_000000001001), .y(t0_00000000100));
wire t0_000000001000, t0_000000001001;
mixer mix_t0_000000001000 (.a(t0_0000000010000), .b(t0_0000000010001), .y(t0_000000001000));
wire t0_0000000010000, t0_0000000010001;
mixer mix_t0_000000001001 (.a(t0_0000000010010), .b(t0_0000000010011), .y(t0_000000001001));
wire t0_0000000010010, t0_0000000010011;
mixer mix_t0_00000000101 (.a(t0_000000001010), .b(t0_000000001011), .y(t0_00000000101));
wire t0_000000001010, t0_000000001011;
mixer mix_t0_000000001010 (.a(t0_0000000010100), .b(t0_0000000010101), .y(t0_000000001010));
wire t0_0000000010100, t0_0000000010101;
mixer mix_t0_000000001011 (.a(t0_0000000010110), .b(t0_0000000010111), .y(t0_000000001011));
wire t0_0000000010110, t0_0000000010111;
mixer mix_t0_0000000011 (.a(t0_00000000110), .b(t0_00000000111), .y(t0_0000000011));
wire t0_00000000110, t0_00000000111;
mixer mix_t0_00000000110 (.a(t0_000000001100), .b(t0_000000001101), .y(t0_00000000110));
wire t0_000000001100, t0_000000001101;
mixer mix_t0_000000001100 (.a(t0_0000000011000), .b(t0_0000000011001), .y(t0_000000001100));
wire t0_0000000011000, t0_0000000011001;
mixer mix_t0_000000001101 (.a(t0_0000000011010), .b(t0_0000000011011), .y(t0_000000001101));
wire t0_0000000011010, t0_0000000011011;
mixer mix_t0_00000000111 (.a(t0_000000001110), .b(t0_000000001111), .y(t0_00000000111));
wire t0_000000001110, t0_000000001111;
mixer mix_t0_000000001110 (.a(t0_0000000011100), .b(t0_0000000011101), .y(t0_000000001110));
wire t0_0000000011100, t0_0000000011101;
mixer mix_t0_000000001111 (.a(t0_0000000011110), .b(t0_0000000011111), .y(t0_000000001111));
wire t0_0000000011110, t0_0000000011111;
mixer mix_t0_00000001 (.a(t0_000000010), .b(t0_000000011), .y(t0_00000001));
wire t0_000000010, t0_000000011;
mixer mix_t0_000000010 (.a(t0_0000000100), .b(t0_0000000101), .y(t0_000000010));
wire t0_0000000100, t0_0000000101;
mixer mix_t0_0000000100 (.a(t0_00000001000), .b(t0_00000001001), .y(t0_0000000100));
wire t0_00000001000, t0_00000001001;
mixer mix_t0_00000001000 (.a(t0_000000010000), .b(t0_000000010001), .y(t0_00000001000));
wire t0_000000010000, t0_000000010001;
mixer mix_t0_000000010000 (.a(t0_0000000100000), .b(t0_0000000100001), .y(t0_000000010000));
wire t0_0000000100000, t0_0000000100001;
mixer mix_t0_000000010001 (.a(t0_0000000100010), .b(t0_0000000100011), .y(t0_000000010001));
wire t0_0000000100010, t0_0000000100011;
mixer mix_t0_00000001001 (.a(t0_000000010010), .b(t0_000000010011), .y(t0_00000001001));
wire t0_000000010010, t0_000000010011;
mixer mix_t0_000000010010 (.a(t0_0000000100100), .b(t0_0000000100101), .y(t0_000000010010));
wire t0_0000000100100, t0_0000000100101;
mixer mix_t0_000000010011 (.a(t0_0000000100110), .b(t0_0000000100111), .y(t0_000000010011));
wire t0_0000000100110, t0_0000000100111;
mixer mix_t0_0000000101 (.a(t0_00000001010), .b(t0_00000001011), .y(t0_0000000101));
wire t0_00000001010, t0_00000001011;
mixer mix_t0_00000001010 (.a(t0_000000010100), .b(t0_000000010101), .y(t0_00000001010));
wire t0_000000010100, t0_000000010101;
mixer mix_t0_000000010100 (.a(t0_0000000101000), .b(t0_0000000101001), .y(t0_000000010100));
wire t0_0000000101000, t0_0000000101001;
mixer mix_t0_000000010101 (.a(t0_0000000101010), .b(t0_0000000101011), .y(t0_000000010101));
wire t0_0000000101010, t0_0000000101011;
mixer mix_t0_00000001011 (.a(t0_000000010110), .b(t0_000000010111), .y(t0_00000001011));
wire t0_000000010110, t0_000000010111;
mixer mix_t0_000000010110 (.a(t0_0000000101100), .b(t0_0000000101101), .y(t0_000000010110));
wire t0_0000000101100, t0_0000000101101;
mixer mix_t0_000000010111 (.a(t0_0000000101110), .b(t0_0000000101111), .y(t0_000000010111));
wire t0_0000000101110, t0_0000000101111;
mixer mix_t0_000000011 (.a(t0_0000000110), .b(t0_0000000111), .y(t0_000000011));
wire t0_0000000110, t0_0000000111;
mixer mix_t0_0000000110 (.a(t0_00000001100), .b(t0_00000001101), .y(t0_0000000110));
wire t0_00000001100, t0_00000001101;
mixer mix_t0_00000001100 (.a(t0_000000011000), .b(t0_000000011001), .y(t0_00000001100));
wire t0_000000011000, t0_000000011001;
mixer mix_t0_000000011000 (.a(t0_0000000110000), .b(t0_0000000110001), .y(t0_000000011000));
wire t0_0000000110000, t0_0000000110001;
mixer mix_t0_000000011001 (.a(t0_0000000110010), .b(t0_0000000110011), .y(t0_000000011001));
wire t0_0000000110010, t0_0000000110011;
mixer mix_t0_00000001101 (.a(t0_000000011010), .b(t0_000000011011), .y(t0_00000001101));
wire t0_000000011010, t0_000000011011;
mixer mix_t0_000000011010 (.a(t0_0000000110100), .b(t0_0000000110101), .y(t0_000000011010));
wire t0_0000000110100, t0_0000000110101;
mixer mix_t0_000000011011 (.a(t0_0000000110110), .b(t0_0000000110111), .y(t0_000000011011));
wire t0_0000000110110, t0_0000000110111;
mixer mix_t0_0000000111 (.a(t0_00000001110), .b(t0_00000001111), .y(t0_0000000111));
wire t0_00000001110, t0_00000001111;
mixer mix_t0_00000001110 (.a(t0_000000011100), .b(t0_000000011101), .y(t0_00000001110));
wire t0_000000011100, t0_000000011101;
mixer mix_t0_000000011100 (.a(t0_0000000111000), .b(t0_0000000111001), .y(t0_000000011100));
wire t0_0000000111000, t0_0000000111001;
mixer mix_t0_000000011101 (.a(t0_0000000111010), .b(t0_0000000111011), .y(t0_000000011101));
wire t0_0000000111010, t0_0000000111011;
mixer mix_t0_00000001111 (.a(t0_000000011110), .b(t0_000000011111), .y(t0_00000001111));
wire t0_000000011110, t0_000000011111;
mixer mix_t0_000000011110 (.a(t0_0000000111100), .b(t0_0000000111101), .y(t0_000000011110));
wire t0_0000000111100, t0_0000000111101;
mixer mix_t0_000000011111 (.a(t0_0000000111110), .b(t0_0000000111111), .y(t0_000000011111));
wire t0_0000000111110, t0_0000000111111;
mixer mix_t0_0000001 (.a(t0_00000010), .b(t0_00000011), .y(t0_0000001));
wire t0_00000010, t0_00000011;
mixer mix_t0_00000010 (.a(t0_000000100), .b(t0_000000101), .y(t0_00000010));
wire t0_000000100, t0_000000101;
mixer mix_t0_000000100 (.a(t0_0000001000), .b(t0_0000001001), .y(t0_000000100));
wire t0_0000001000, t0_0000001001;
mixer mix_t0_0000001000 (.a(t0_00000010000), .b(t0_00000010001), .y(t0_0000001000));
wire t0_00000010000, t0_00000010001;
mixer mix_t0_00000010000 (.a(t0_000000100000), .b(t0_000000100001), .y(t0_00000010000));
wire t0_000000100000, t0_000000100001;
mixer mix_t0_000000100000 (.a(t0_0000001000000), .b(t0_0000001000001), .y(t0_000000100000));
wire t0_0000001000000, t0_0000001000001;
mixer mix_t0_000000100001 (.a(t0_0000001000010), .b(t0_0000001000011), .y(t0_000000100001));
wire t0_0000001000010, t0_0000001000011;
mixer mix_t0_00000010001 (.a(t0_000000100010), .b(t0_000000100011), .y(t0_00000010001));
wire t0_000000100010, t0_000000100011;
mixer mix_t0_000000100010 (.a(t0_0000001000100), .b(t0_0000001000101), .y(t0_000000100010));
wire t0_0000001000100, t0_0000001000101;
mixer mix_t0_000000100011 (.a(t0_0000001000110), .b(t0_0000001000111), .y(t0_000000100011));
wire t0_0000001000110, t0_0000001000111;
mixer mix_t0_0000001001 (.a(t0_00000010010), .b(t0_00000010011), .y(t0_0000001001));
wire t0_00000010010, t0_00000010011;
mixer mix_t0_00000010010 (.a(t0_000000100100), .b(t0_000000100101), .y(t0_00000010010));
wire t0_000000100100, t0_000000100101;
mixer mix_t0_000000100100 (.a(t0_0000001001000), .b(t0_0000001001001), .y(t0_000000100100));
wire t0_0000001001000, t0_0000001001001;
mixer mix_t0_000000100101 (.a(t0_0000001001010), .b(t0_0000001001011), .y(t0_000000100101));
wire t0_0000001001010, t0_0000001001011;
mixer mix_t0_00000010011 (.a(t0_000000100110), .b(t0_000000100111), .y(t0_00000010011));
wire t0_000000100110, t0_000000100111;
mixer mix_t0_000000100110 (.a(t0_0000001001100), .b(t0_0000001001101), .y(t0_000000100110));
wire t0_0000001001100, t0_0000001001101;
mixer mix_t0_000000100111 (.a(t0_0000001001110), .b(t0_0000001001111), .y(t0_000000100111));
wire t0_0000001001110, t0_0000001001111;
mixer mix_t0_000000101 (.a(t0_0000001010), .b(t0_0000001011), .y(t0_000000101));
wire t0_0000001010, t0_0000001011;
mixer mix_t0_0000001010 (.a(t0_00000010100), .b(t0_00000010101), .y(t0_0000001010));
wire t0_00000010100, t0_00000010101;
mixer mix_t0_00000010100 (.a(t0_000000101000), .b(t0_000000101001), .y(t0_00000010100));
wire t0_000000101000, t0_000000101001;
mixer mix_t0_000000101000 (.a(t0_0000001010000), .b(t0_0000001010001), .y(t0_000000101000));
wire t0_0000001010000, t0_0000001010001;
mixer mix_t0_000000101001 (.a(t0_0000001010010), .b(t0_0000001010011), .y(t0_000000101001));
wire t0_0000001010010, t0_0000001010011;
mixer mix_t0_00000010101 (.a(t0_000000101010), .b(t0_000000101011), .y(t0_00000010101));
wire t0_000000101010, t0_000000101011;
mixer mix_t0_000000101010 (.a(t0_0000001010100), .b(t0_0000001010101), .y(t0_000000101010));
wire t0_0000001010100, t0_0000001010101;
mixer mix_t0_000000101011 (.a(t0_0000001010110), .b(t0_0000001010111), .y(t0_000000101011));
wire t0_0000001010110, t0_0000001010111;
mixer mix_t0_0000001011 (.a(t0_00000010110), .b(t0_00000010111), .y(t0_0000001011));
wire t0_00000010110, t0_00000010111;
mixer mix_t0_00000010110 (.a(t0_000000101100), .b(t0_000000101101), .y(t0_00000010110));
wire t0_000000101100, t0_000000101101;
mixer mix_t0_000000101100 (.a(t0_0000001011000), .b(t0_0000001011001), .y(t0_000000101100));
wire t0_0000001011000, t0_0000001011001;
mixer mix_t0_000000101101 (.a(t0_0000001011010), .b(t0_0000001011011), .y(t0_000000101101));
wire t0_0000001011010, t0_0000001011011;
mixer mix_t0_00000010111 (.a(t0_000000101110), .b(t0_000000101111), .y(t0_00000010111));
wire t0_000000101110, t0_000000101111;
mixer mix_t0_000000101110 (.a(t0_0000001011100), .b(t0_0000001011101), .y(t0_000000101110));
wire t0_0000001011100, t0_0000001011101;
mixer mix_t0_000000101111 (.a(t0_0000001011110), .b(t0_0000001011111), .y(t0_000000101111));
wire t0_0000001011110, t0_0000001011111;
mixer mix_t0_00000011 (.a(t0_000000110), .b(t0_000000111), .y(t0_00000011));
wire t0_000000110, t0_000000111;
mixer mix_t0_000000110 (.a(t0_0000001100), .b(t0_0000001101), .y(t0_000000110));
wire t0_0000001100, t0_0000001101;
mixer mix_t0_0000001100 (.a(t0_00000011000), .b(t0_00000011001), .y(t0_0000001100));
wire t0_00000011000, t0_00000011001;
mixer mix_t0_00000011000 (.a(t0_000000110000), .b(t0_000000110001), .y(t0_00000011000));
wire t0_000000110000, t0_000000110001;
mixer mix_t0_000000110000 (.a(t0_0000001100000), .b(t0_0000001100001), .y(t0_000000110000));
wire t0_0000001100000, t0_0000001100001;
mixer mix_t0_000000110001 (.a(t0_0000001100010), .b(t0_0000001100011), .y(t0_000000110001));
wire t0_0000001100010, t0_0000001100011;
mixer mix_t0_00000011001 (.a(t0_000000110010), .b(t0_000000110011), .y(t0_00000011001));
wire t0_000000110010, t0_000000110011;
mixer mix_t0_000000110010 (.a(t0_0000001100100), .b(t0_0000001100101), .y(t0_000000110010));
wire t0_0000001100100, t0_0000001100101;
mixer mix_t0_000000110011 (.a(t0_0000001100110), .b(t0_0000001100111), .y(t0_000000110011));
wire t0_0000001100110, t0_0000001100111;
mixer mix_t0_0000001101 (.a(t0_00000011010), .b(t0_00000011011), .y(t0_0000001101));
wire t0_00000011010, t0_00000011011;
mixer mix_t0_00000011010 (.a(t0_000000110100), .b(t0_000000110101), .y(t0_00000011010));
wire t0_000000110100, t0_000000110101;
mixer mix_t0_000000110100 (.a(t0_0000001101000), .b(t0_0000001101001), .y(t0_000000110100));
wire t0_0000001101000, t0_0000001101001;
mixer mix_t0_000000110101 (.a(t0_0000001101010), .b(t0_0000001101011), .y(t0_000000110101));
wire t0_0000001101010, t0_0000001101011;
mixer mix_t0_00000011011 (.a(t0_000000110110), .b(t0_000000110111), .y(t0_00000011011));
wire t0_000000110110, t0_000000110111;
mixer mix_t0_000000110110 (.a(t0_0000001101100), .b(t0_0000001101101), .y(t0_000000110110));
wire t0_0000001101100, t0_0000001101101;
mixer mix_t0_000000110111 (.a(t0_0000001101110), .b(t0_0000001101111), .y(t0_000000110111));
wire t0_0000001101110, t0_0000001101111;
mixer mix_t0_000000111 (.a(t0_0000001110), .b(t0_0000001111), .y(t0_000000111));
wire t0_0000001110, t0_0000001111;
mixer mix_t0_0000001110 (.a(t0_00000011100), .b(t0_00000011101), .y(t0_0000001110));
wire t0_00000011100, t0_00000011101;
mixer mix_t0_00000011100 (.a(t0_000000111000), .b(t0_000000111001), .y(t0_00000011100));
wire t0_000000111000, t0_000000111001;
mixer mix_t0_000000111000 (.a(t0_0000001110000), .b(t0_0000001110001), .y(t0_000000111000));
wire t0_0000001110000, t0_0000001110001;
mixer mix_t0_000000111001 (.a(t0_0000001110010), .b(t0_0000001110011), .y(t0_000000111001));
wire t0_0000001110010, t0_0000001110011;
mixer mix_t0_00000011101 (.a(t0_000000111010), .b(t0_000000111011), .y(t0_00000011101));
wire t0_000000111010, t0_000000111011;
mixer mix_t0_000000111010 (.a(t0_0000001110100), .b(t0_0000001110101), .y(t0_000000111010));
wire t0_0000001110100, t0_0000001110101;
mixer mix_t0_000000111011 (.a(t0_0000001110110), .b(t0_0000001110111), .y(t0_000000111011));
wire t0_0000001110110, t0_0000001110111;
mixer mix_t0_0000001111 (.a(t0_00000011110), .b(t0_00000011111), .y(t0_0000001111));
wire t0_00000011110, t0_00000011111;
mixer mix_t0_00000011110 (.a(t0_000000111100), .b(t0_000000111101), .y(t0_00000011110));
wire t0_000000111100, t0_000000111101;
mixer mix_t0_000000111100 (.a(t0_0000001111000), .b(t0_0000001111001), .y(t0_000000111100));
wire t0_0000001111000, t0_0000001111001;
mixer mix_t0_000000111101 (.a(t0_0000001111010), .b(t0_0000001111011), .y(t0_000000111101));
wire t0_0000001111010, t0_0000001111011;
mixer mix_t0_00000011111 (.a(t0_000000111110), .b(t0_000000111111), .y(t0_00000011111));
wire t0_000000111110, t0_000000111111;
mixer mix_t0_000000111110 (.a(t0_0000001111100), .b(t0_0000001111101), .y(t0_000000111110));
wire t0_0000001111100, t0_0000001111101;
mixer mix_t0_000000111111 (.a(t0_0000001111110), .b(t0_0000001111111), .y(t0_000000111111));
wire t0_0000001111110, t0_0000001111111;
mixer mix_t0_000001 (.a(t0_0000010), .b(t0_0000011), .y(t0_000001));
wire t0_0000010, t0_0000011;
mixer mix_t0_0000010 (.a(t0_00000100), .b(t0_00000101), .y(t0_0000010));
wire t0_00000100, t0_00000101;
mixer mix_t0_00000100 (.a(t0_000001000), .b(t0_000001001), .y(t0_00000100));
wire t0_000001000, t0_000001001;
mixer mix_t0_000001000 (.a(t0_0000010000), .b(t0_0000010001), .y(t0_000001000));
wire t0_0000010000, t0_0000010001;
mixer mix_t0_0000010000 (.a(t0_00000100000), .b(t0_00000100001), .y(t0_0000010000));
wire t0_00000100000, t0_00000100001;
mixer mix_t0_00000100000 (.a(t0_000001000000), .b(t0_000001000001), .y(t0_00000100000));
wire t0_000001000000, t0_000001000001;
mixer mix_t0_000001000000 (.a(t0_0000010000000), .b(t0_0000010000001), .y(t0_000001000000));
wire t0_0000010000000, t0_0000010000001;
mixer mix_t0_000001000001 (.a(t0_0000010000010), .b(t0_0000010000011), .y(t0_000001000001));
wire t0_0000010000010, t0_0000010000011;
mixer mix_t0_00000100001 (.a(t0_000001000010), .b(t0_000001000011), .y(t0_00000100001));
wire t0_000001000010, t0_000001000011;
mixer mix_t0_000001000010 (.a(t0_0000010000100), .b(t0_0000010000101), .y(t0_000001000010));
wire t0_0000010000100, t0_0000010000101;
mixer mix_t0_000001000011 (.a(t0_0000010000110), .b(t0_0000010000111), .y(t0_000001000011));
wire t0_0000010000110, t0_0000010000111;
mixer mix_t0_0000010001 (.a(t0_00000100010), .b(t0_00000100011), .y(t0_0000010001));
wire t0_00000100010, t0_00000100011;
mixer mix_t0_00000100010 (.a(t0_000001000100), .b(t0_000001000101), .y(t0_00000100010));
wire t0_000001000100, t0_000001000101;
mixer mix_t0_000001000100 (.a(t0_0000010001000), .b(t0_0000010001001), .y(t0_000001000100));
wire t0_0000010001000, t0_0000010001001;
mixer mix_t0_000001000101 (.a(t0_0000010001010), .b(t0_0000010001011), .y(t0_000001000101));
wire t0_0000010001010, t0_0000010001011;
mixer mix_t0_00000100011 (.a(t0_000001000110), .b(t0_000001000111), .y(t0_00000100011));
wire t0_000001000110, t0_000001000111;
mixer mix_t0_000001000110 (.a(t0_0000010001100), .b(t0_0000010001101), .y(t0_000001000110));
wire t0_0000010001100, t0_0000010001101;
mixer mix_t0_000001000111 (.a(t0_0000010001110), .b(t0_0000010001111), .y(t0_000001000111));
wire t0_0000010001110, t0_0000010001111;
mixer mix_t0_000001001 (.a(t0_0000010010), .b(t0_0000010011), .y(t0_000001001));
wire t0_0000010010, t0_0000010011;
mixer mix_t0_0000010010 (.a(t0_00000100100), .b(t0_00000100101), .y(t0_0000010010));
wire t0_00000100100, t0_00000100101;
mixer mix_t0_00000100100 (.a(t0_000001001000), .b(t0_000001001001), .y(t0_00000100100));
wire t0_000001001000, t0_000001001001;
mixer mix_t0_000001001000 (.a(t0_0000010010000), .b(t0_0000010010001), .y(t0_000001001000));
wire t0_0000010010000, t0_0000010010001;
mixer mix_t0_000001001001 (.a(t0_0000010010010), .b(t0_0000010010011), .y(t0_000001001001));
wire t0_0000010010010, t0_0000010010011;
mixer mix_t0_00000100101 (.a(t0_000001001010), .b(t0_000001001011), .y(t0_00000100101));
wire t0_000001001010, t0_000001001011;
mixer mix_t0_000001001010 (.a(t0_0000010010100), .b(t0_0000010010101), .y(t0_000001001010));
wire t0_0000010010100, t0_0000010010101;
mixer mix_t0_000001001011 (.a(t0_0000010010110), .b(t0_0000010010111), .y(t0_000001001011));
wire t0_0000010010110, t0_0000010010111;
mixer mix_t0_0000010011 (.a(t0_00000100110), .b(t0_00000100111), .y(t0_0000010011));
wire t0_00000100110, t0_00000100111;
mixer mix_t0_00000100110 (.a(t0_000001001100), .b(t0_000001001101), .y(t0_00000100110));
wire t0_000001001100, t0_000001001101;
mixer mix_t0_000001001100 (.a(t0_0000010011000), .b(t0_0000010011001), .y(t0_000001001100));
wire t0_0000010011000, t0_0000010011001;
mixer mix_t0_000001001101 (.a(t0_0000010011010), .b(t0_0000010011011), .y(t0_000001001101));
wire t0_0000010011010, t0_0000010011011;
mixer mix_t0_00000100111 (.a(t0_000001001110), .b(t0_000001001111), .y(t0_00000100111));
wire t0_000001001110, t0_000001001111;
mixer mix_t0_000001001110 (.a(t0_0000010011100), .b(t0_0000010011101), .y(t0_000001001110));
wire t0_0000010011100, t0_0000010011101;
mixer mix_t0_000001001111 (.a(t0_0000010011110), .b(t0_0000010011111), .y(t0_000001001111));
wire t0_0000010011110, t0_0000010011111;
mixer mix_t0_00000101 (.a(t0_000001010), .b(t0_000001011), .y(t0_00000101));
wire t0_000001010, t0_000001011;
mixer mix_t0_000001010 (.a(t0_0000010100), .b(t0_0000010101), .y(t0_000001010));
wire t0_0000010100, t0_0000010101;
mixer mix_t0_0000010100 (.a(t0_00000101000), .b(t0_00000101001), .y(t0_0000010100));
wire t0_00000101000, t0_00000101001;
mixer mix_t0_00000101000 (.a(t0_000001010000), .b(t0_000001010001), .y(t0_00000101000));
wire t0_000001010000, t0_000001010001;
mixer mix_t0_000001010000 (.a(t0_0000010100000), .b(t0_0000010100001), .y(t0_000001010000));
wire t0_0000010100000, t0_0000010100001;
mixer mix_t0_000001010001 (.a(t0_0000010100010), .b(t0_0000010100011), .y(t0_000001010001));
wire t0_0000010100010, t0_0000010100011;
mixer mix_t0_00000101001 (.a(t0_000001010010), .b(t0_000001010011), .y(t0_00000101001));
wire t0_000001010010, t0_000001010011;
mixer mix_t0_000001010010 (.a(t0_0000010100100), .b(t0_0000010100101), .y(t0_000001010010));
wire t0_0000010100100, t0_0000010100101;
mixer mix_t0_000001010011 (.a(t0_0000010100110), .b(t0_0000010100111), .y(t0_000001010011));
wire t0_0000010100110, t0_0000010100111;
mixer mix_t0_0000010101 (.a(t0_00000101010), .b(t0_00000101011), .y(t0_0000010101));
wire t0_00000101010, t0_00000101011;
mixer mix_t0_00000101010 (.a(t0_000001010100), .b(t0_000001010101), .y(t0_00000101010));
wire t0_000001010100, t0_000001010101;
mixer mix_t0_000001010100 (.a(t0_0000010101000), .b(t0_0000010101001), .y(t0_000001010100));
wire t0_0000010101000, t0_0000010101001;
mixer mix_t0_000001010101 (.a(t0_0000010101010), .b(t0_0000010101011), .y(t0_000001010101));
wire t0_0000010101010, t0_0000010101011;
mixer mix_t0_00000101011 (.a(t0_000001010110), .b(t0_000001010111), .y(t0_00000101011));
wire t0_000001010110, t0_000001010111;
mixer mix_t0_000001010110 (.a(t0_0000010101100), .b(t0_0000010101101), .y(t0_000001010110));
wire t0_0000010101100, t0_0000010101101;
mixer mix_t0_000001010111 (.a(t0_0000010101110), .b(t0_0000010101111), .y(t0_000001010111));
wire t0_0000010101110, t0_0000010101111;
mixer mix_t0_000001011 (.a(t0_0000010110), .b(t0_0000010111), .y(t0_000001011));
wire t0_0000010110, t0_0000010111;
mixer mix_t0_0000010110 (.a(t0_00000101100), .b(t0_00000101101), .y(t0_0000010110));
wire t0_00000101100, t0_00000101101;
mixer mix_t0_00000101100 (.a(t0_000001011000), .b(t0_000001011001), .y(t0_00000101100));
wire t0_000001011000, t0_000001011001;
mixer mix_t0_000001011000 (.a(t0_0000010110000), .b(t0_0000010110001), .y(t0_000001011000));
wire t0_0000010110000, t0_0000010110001;
mixer mix_t0_000001011001 (.a(t0_0000010110010), .b(t0_0000010110011), .y(t0_000001011001));
wire t0_0000010110010, t0_0000010110011;
mixer mix_t0_00000101101 (.a(t0_000001011010), .b(t0_000001011011), .y(t0_00000101101));
wire t0_000001011010, t0_000001011011;
mixer mix_t0_000001011010 (.a(t0_0000010110100), .b(t0_0000010110101), .y(t0_000001011010));
wire t0_0000010110100, t0_0000010110101;
mixer mix_t0_000001011011 (.a(t0_0000010110110), .b(t0_0000010110111), .y(t0_000001011011));
wire t0_0000010110110, t0_0000010110111;
mixer mix_t0_0000010111 (.a(t0_00000101110), .b(t0_00000101111), .y(t0_0000010111));
wire t0_00000101110, t0_00000101111;
mixer mix_t0_00000101110 (.a(t0_000001011100), .b(t0_000001011101), .y(t0_00000101110));
wire t0_000001011100, t0_000001011101;
mixer mix_t0_000001011100 (.a(t0_0000010111000), .b(t0_0000010111001), .y(t0_000001011100));
wire t0_0000010111000, t0_0000010111001;
mixer mix_t0_000001011101 (.a(t0_0000010111010), .b(t0_0000010111011), .y(t0_000001011101));
wire t0_0000010111010, t0_0000010111011;
mixer mix_t0_00000101111 (.a(t0_000001011110), .b(t0_000001011111), .y(t0_00000101111));
wire t0_000001011110, t0_000001011111;
mixer mix_t0_000001011110 (.a(t0_0000010111100), .b(t0_0000010111101), .y(t0_000001011110));
wire t0_0000010111100, t0_0000010111101;
mixer mix_t0_000001011111 (.a(t0_0000010111110), .b(t0_0000010111111), .y(t0_000001011111));
wire t0_0000010111110, t0_0000010111111;
mixer mix_t0_0000011 (.a(t0_00000110), .b(t0_00000111), .y(t0_0000011));
wire t0_00000110, t0_00000111;
mixer mix_t0_00000110 (.a(t0_000001100), .b(t0_000001101), .y(t0_00000110));
wire t0_000001100, t0_000001101;
mixer mix_t0_000001100 (.a(t0_0000011000), .b(t0_0000011001), .y(t0_000001100));
wire t0_0000011000, t0_0000011001;
mixer mix_t0_0000011000 (.a(t0_00000110000), .b(t0_00000110001), .y(t0_0000011000));
wire t0_00000110000, t0_00000110001;
mixer mix_t0_00000110000 (.a(t0_000001100000), .b(t0_000001100001), .y(t0_00000110000));
wire t0_000001100000, t0_000001100001;
mixer mix_t0_000001100000 (.a(t0_0000011000000), .b(t0_0000011000001), .y(t0_000001100000));
wire t0_0000011000000, t0_0000011000001;
mixer mix_t0_000001100001 (.a(t0_0000011000010), .b(t0_0000011000011), .y(t0_000001100001));
wire t0_0000011000010, t0_0000011000011;
mixer mix_t0_00000110001 (.a(t0_000001100010), .b(t0_000001100011), .y(t0_00000110001));
wire t0_000001100010, t0_000001100011;
mixer mix_t0_000001100010 (.a(t0_0000011000100), .b(t0_0000011000101), .y(t0_000001100010));
wire t0_0000011000100, t0_0000011000101;
mixer mix_t0_000001100011 (.a(t0_0000011000110), .b(t0_0000011000111), .y(t0_000001100011));
wire t0_0000011000110, t0_0000011000111;
mixer mix_t0_0000011001 (.a(t0_00000110010), .b(t0_00000110011), .y(t0_0000011001));
wire t0_00000110010, t0_00000110011;
mixer mix_t0_00000110010 (.a(t0_000001100100), .b(t0_000001100101), .y(t0_00000110010));
wire t0_000001100100, t0_000001100101;
mixer mix_t0_000001100100 (.a(t0_0000011001000), .b(t0_0000011001001), .y(t0_000001100100));
wire t0_0000011001000, t0_0000011001001;
mixer mix_t0_000001100101 (.a(t0_0000011001010), .b(t0_0000011001011), .y(t0_000001100101));
wire t0_0000011001010, t0_0000011001011;
mixer mix_t0_00000110011 (.a(t0_000001100110), .b(t0_000001100111), .y(t0_00000110011));
wire t0_000001100110, t0_000001100111;
mixer mix_t0_000001100110 (.a(t0_0000011001100), .b(t0_0000011001101), .y(t0_000001100110));
wire t0_0000011001100, t0_0000011001101;
mixer mix_t0_000001100111 (.a(t0_0000011001110), .b(t0_0000011001111), .y(t0_000001100111));
wire t0_0000011001110, t0_0000011001111;
mixer mix_t0_000001101 (.a(t0_0000011010), .b(t0_0000011011), .y(t0_000001101));
wire t0_0000011010, t0_0000011011;
mixer mix_t0_0000011010 (.a(t0_00000110100), .b(t0_00000110101), .y(t0_0000011010));
wire t0_00000110100, t0_00000110101;
mixer mix_t0_00000110100 (.a(t0_000001101000), .b(t0_000001101001), .y(t0_00000110100));
wire t0_000001101000, t0_000001101001;
mixer mix_t0_000001101000 (.a(t0_0000011010000), .b(t0_0000011010001), .y(t0_000001101000));
wire t0_0000011010000, t0_0000011010001;
mixer mix_t0_000001101001 (.a(t0_0000011010010), .b(t0_0000011010011), .y(t0_000001101001));
wire t0_0000011010010, t0_0000011010011;
mixer mix_t0_00000110101 (.a(t0_000001101010), .b(t0_000001101011), .y(t0_00000110101));
wire t0_000001101010, t0_000001101011;
mixer mix_t0_000001101010 (.a(t0_0000011010100), .b(t0_0000011010101), .y(t0_000001101010));
wire t0_0000011010100, t0_0000011010101;
mixer mix_t0_000001101011 (.a(t0_0000011010110), .b(t0_0000011010111), .y(t0_000001101011));
wire t0_0000011010110, t0_0000011010111;
mixer mix_t0_0000011011 (.a(t0_00000110110), .b(t0_00000110111), .y(t0_0000011011));
wire t0_00000110110, t0_00000110111;
mixer mix_t0_00000110110 (.a(t0_000001101100), .b(t0_000001101101), .y(t0_00000110110));
wire t0_000001101100, t0_000001101101;
mixer mix_t0_000001101100 (.a(t0_0000011011000), .b(t0_0000011011001), .y(t0_000001101100));
wire t0_0000011011000, t0_0000011011001;
mixer mix_t0_000001101101 (.a(t0_0000011011010), .b(t0_0000011011011), .y(t0_000001101101));
wire t0_0000011011010, t0_0000011011011;
mixer mix_t0_00000110111 (.a(t0_000001101110), .b(t0_000001101111), .y(t0_00000110111));
wire t0_000001101110, t0_000001101111;
mixer mix_t0_000001101110 (.a(t0_0000011011100), .b(t0_0000011011101), .y(t0_000001101110));
wire t0_0000011011100, t0_0000011011101;
mixer mix_t0_000001101111 (.a(t0_0000011011110), .b(t0_0000011011111), .y(t0_000001101111));
wire t0_0000011011110, t0_0000011011111;
mixer mix_t0_00000111 (.a(t0_000001110), .b(t0_000001111), .y(t0_00000111));
wire t0_000001110, t0_000001111;
mixer mix_t0_000001110 (.a(t0_0000011100), .b(t0_0000011101), .y(t0_000001110));
wire t0_0000011100, t0_0000011101;
mixer mix_t0_0000011100 (.a(t0_00000111000), .b(t0_00000111001), .y(t0_0000011100));
wire t0_00000111000, t0_00000111001;
mixer mix_t0_00000111000 (.a(t0_000001110000), .b(t0_000001110001), .y(t0_00000111000));
wire t0_000001110000, t0_000001110001;
mixer mix_t0_000001110000 (.a(t0_0000011100000), .b(t0_0000011100001), .y(t0_000001110000));
wire t0_0000011100000, t0_0000011100001;
mixer mix_t0_000001110001 (.a(t0_0000011100010), .b(t0_0000011100011), .y(t0_000001110001));
wire t0_0000011100010, t0_0000011100011;
mixer mix_t0_00000111001 (.a(t0_000001110010), .b(t0_000001110011), .y(t0_00000111001));
wire t0_000001110010, t0_000001110011;
mixer mix_t0_000001110010 (.a(t0_0000011100100), .b(t0_0000011100101), .y(t0_000001110010));
wire t0_0000011100100, t0_0000011100101;
mixer mix_t0_000001110011 (.a(t0_0000011100110), .b(t0_0000011100111), .y(t0_000001110011));
wire t0_0000011100110, t0_0000011100111;
mixer mix_t0_0000011101 (.a(t0_00000111010), .b(t0_00000111011), .y(t0_0000011101));
wire t0_00000111010, t0_00000111011;
mixer mix_t0_00000111010 (.a(t0_000001110100), .b(t0_000001110101), .y(t0_00000111010));
wire t0_000001110100, t0_000001110101;
mixer mix_t0_000001110100 (.a(t0_0000011101000), .b(t0_0000011101001), .y(t0_000001110100));
wire t0_0000011101000, t0_0000011101001;
mixer mix_t0_000001110101 (.a(t0_0000011101010), .b(t0_0000011101011), .y(t0_000001110101));
wire t0_0000011101010, t0_0000011101011;
mixer mix_t0_00000111011 (.a(t0_000001110110), .b(t0_000001110111), .y(t0_00000111011));
wire t0_000001110110, t0_000001110111;
mixer mix_t0_000001110110 (.a(t0_0000011101100), .b(t0_0000011101101), .y(t0_000001110110));
wire t0_0000011101100, t0_0000011101101;
mixer mix_t0_000001110111 (.a(t0_0000011101110), .b(t0_0000011101111), .y(t0_000001110111));
wire t0_0000011101110, t0_0000011101111;
mixer mix_t0_000001111 (.a(t0_0000011110), .b(t0_0000011111), .y(t0_000001111));
wire t0_0000011110, t0_0000011111;
mixer mix_t0_0000011110 (.a(t0_00000111100), .b(t0_00000111101), .y(t0_0000011110));
wire t0_00000111100, t0_00000111101;
mixer mix_t0_00000111100 (.a(t0_000001111000), .b(t0_000001111001), .y(t0_00000111100));
wire t0_000001111000, t0_000001111001;
mixer mix_t0_000001111000 (.a(t0_0000011110000), .b(t0_0000011110001), .y(t0_000001111000));
wire t0_0000011110000, t0_0000011110001;
mixer mix_t0_000001111001 (.a(t0_0000011110010), .b(t0_0000011110011), .y(t0_000001111001));
wire t0_0000011110010, t0_0000011110011;
mixer mix_t0_00000111101 (.a(t0_000001111010), .b(t0_000001111011), .y(t0_00000111101));
wire t0_000001111010, t0_000001111011;
mixer mix_t0_000001111010 (.a(t0_0000011110100), .b(t0_0000011110101), .y(t0_000001111010));
wire t0_0000011110100, t0_0000011110101;
mixer mix_t0_000001111011 (.a(t0_0000011110110), .b(t0_0000011110111), .y(t0_000001111011));
wire t0_0000011110110, t0_0000011110111;
mixer mix_t0_0000011111 (.a(t0_00000111110), .b(t0_00000111111), .y(t0_0000011111));
wire t0_00000111110, t0_00000111111;
mixer mix_t0_00000111110 (.a(t0_000001111100), .b(t0_000001111101), .y(t0_00000111110));
wire t0_000001111100, t0_000001111101;
mixer mix_t0_000001111100 (.a(t0_0000011111000), .b(t0_0000011111001), .y(t0_000001111100));
wire t0_0000011111000, t0_0000011111001;
mixer mix_t0_000001111101 (.a(t0_0000011111010), .b(t0_0000011111011), .y(t0_000001111101));
wire t0_0000011111010, t0_0000011111011;
mixer mix_t0_00000111111 (.a(t0_000001111110), .b(t0_000001111111), .y(t0_00000111111));
wire t0_000001111110, t0_000001111111;
mixer mix_t0_000001111110 (.a(t0_0000011111100), .b(t0_0000011111101), .y(t0_000001111110));
wire t0_0000011111100, t0_0000011111101;
mixer mix_t0_000001111111 (.a(t0_0000011111110), .b(t0_0000011111111), .y(t0_000001111111));
wire t0_0000011111110, t0_0000011111111;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_000010 (.a(t0_0000100), .b(t0_0000101), .y(t0_000010));
wire t0_0000100, t0_0000101;
mixer mix_t0_0000100 (.a(t0_00001000), .b(t0_00001001), .y(t0_0000100));
wire t0_00001000, t0_00001001;
mixer mix_t0_00001000 (.a(t0_000010000), .b(t0_000010001), .y(t0_00001000));
wire t0_000010000, t0_000010001;
mixer mix_t0_000010000 (.a(t0_0000100000), .b(t0_0000100001), .y(t0_000010000));
wire t0_0000100000, t0_0000100001;
mixer mix_t0_0000100000 (.a(t0_00001000000), .b(t0_00001000001), .y(t0_0000100000));
wire t0_00001000000, t0_00001000001;
mixer mix_t0_00001000000 (.a(t0_000010000000), .b(t0_000010000001), .y(t0_00001000000));
wire t0_000010000000, t0_000010000001;
mixer mix_t0_000010000000 (.a(t0_0000100000000), .b(t0_0000100000001), .y(t0_000010000000));
wire t0_0000100000000, t0_0000100000001;
mixer mix_t0_000010000001 (.a(t0_0000100000010), .b(t0_0000100000011), .y(t0_000010000001));
wire t0_0000100000010, t0_0000100000011;
mixer mix_t0_00001000001 (.a(t0_000010000010), .b(t0_000010000011), .y(t0_00001000001));
wire t0_000010000010, t0_000010000011;
mixer mix_t0_000010000010 (.a(t0_0000100000100), .b(t0_0000100000101), .y(t0_000010000010));
wire t0_0000100000100, t0_0000100000101;
mixer mix_t0_000010000011 (.a(t0_0000100000110), .b(t0_0000100000111), .y(t0_000010000011));
wire t0_0000100000110, t0_0000100000111;
mixer mix_t0_0000100001 (.a(t0_00001000010), .b(t0_00001000011), .y(t0_0000100001));
wire t0_00001000010, t0_00001000011;
mixer mix_t0_00001000010 (.a(t0_000010000100), .b(t0_000010000101), .y(t0_00001000010));
wire t0_000010000100, t0_000010000101;
mixer mix_t0_000010000100 (.a(t0_0000100001000), .b(t0_0000100001001), .y(t0_000010000100));
wire t0_0000100001000, t0_0000100001001;
mixer mix_t0_000010000101 (.a(t0_0000100001010), .b(t0_0000100001011), .y(t0_000010000101));
wire t0_0000100001010, t0_0000100001011;
mixer mix_t0_00001000011 (.a(t0_000010000110), .b(t0_000010000111), .y(t0_00001000011));
wire t0_000010000110, t0_000010000111;
mixer mix_t0_000010000110 (.a(t0_0000100001100), .b(t0_0000100001101), .y(t0_000010000110));
wire t0_0000100001100, t0_0000100001101;
mixer mix_t0_000010000111 (.a(t0_0000100001110), .b(t0_0000100001111), .y(t0_000010000111));
wire t0_0000100001110, t0_0000100001111;
mixer mix_t0_000010001 (.a(t0_0000100010), .b(t0_0000100011), .y(t0_000010001));
wire t0_0000100010, t0_0000100011;
mixer mix_t0_0000100010 (.a(t0_00001000100), .b(t0_00001000101), .y(t0_0000100010));
wire t0_00001000100, t0_00001000101;
mixer mix_t0_00001000100 (.a(t0_000010001000), .b(t0_000010001001), .y(t0_00001000100));
wire t0_000010001000, t0_000010001001;
mixer mix_t0_000010001000 (.a(t0_0000100010000), .b(t0_0000100010001), .y(t0_000010001000));
wire t0_0000100010000, t0_0000100010001;
mixer mix_t0_000010001001 (.a(t0_0000100010010), .b(t0_0000100010011), .y(t0_000010001001));
wire t0_0000100010010, t0_0000100010011;
mixer mix_t0_00001000101 (.a(t0_000010001010), .b(t0_000010001011), .y(t0_00001000101));
wire t0_000010001010, t0_000010001011;
mixer mix_t0_000010001010 (.a(t0_0000100010100), .b(t0_0000100010101), .y(t0_000010001010));
wire t0_0000100010100, t0_0000100010101;
mixer mix_t0_000010001011 (.a(t0_0000100010110), .b(t0_0000100010111), .y(t0_000010001011));
wire t0_0000100010110, t0_0000100010111;
mixer mix_t0_0000100011 (.a(t0_00001000110), .b(t0_00001000111), .y(t0_0000100011));
wire t0_00001000110, t0_00001000111;
mixer mix_t0_00001000110 (.a(t0_000010001100), .b(t0_000010001101), .y(t0_00001000110));
wire t0_000010001100, t0_000010001101;
mixer mix_t0_000010001100 (.a(t0_0000100011000), .b(t0_0000100011001), .y(t0_000010001100));
wire t0_0000100011000, t0_0000100011001;
mixer mix_t0_000010001101 (.a(t0_0000100011010), .b(t0_0000100011011), .y(t0_000010001101));
wire t0_0000100011010, t0_0000100011011;
mixer mix_t0_00001000111 (.a(t0_000010001110), .b(t0_000010001111), .y(t0_00001000111));
wire t0_000010001110, t0_000010001111;
mixer mix_t0_000010001110 (.a(t0_0000100011100), .b(t0_0000100011101), .y(t0_000010001110));
wire t0_0000100011100, t0_0000100011101;
mixer mix_t0_000010001111 (.a(t0_0000100011110), .b(t0_0000100011111), .y(t0_000010001111));
wire t0_0000100011110, t0_0000100011111;
mixer mix_t0_00001001 (.a(t0_000010010), .b(t0_000010011), .y(t0_00001001));
wire t0_000010010, t0_000010011;
mixer mix_t0_000010010 (.a(t0_0000100100), .b(t0_0000100101), .y(t0_000010010));
wire t0_0000100100, t0_0000100101;
mixer mix_t0_0000100100 (.a(t0_00001001000), .b(t0_00001001001), .y(t0_0000100100));
wire t0_00001001000, t0_00001001001;
mixer mix_t0_00001001000 (.a(t0_000010010000), .b(t0_000010010001), .y(t0_00001001000));
wire t0_000010010000, t0_000010010001;
mixer mix_t0_000010010000 (.a(t0_0000100100000), .b(t0_0000100100001), .y(t0_000010010000));
wire t0_0000100100000, t0_0000100100001;
mixer mix_t0_000010010001 (.a(t0_0000100100010), .b(t0_0000100100011), .y(t0_000010010001));
wire t0_0000100100010, t0_0000100100011;
mixer mix_t0_00001001001 (.a(t0_000010010010), .b(t0_000010010011), .y(t0_00001001001));
wire t0_000010010010, t0_000010010011;
mixer mix_t0_000010010010 (.a(t0_0000100100100), .b(t0_0000100100101), .y(t0_000010010010));
wire t0_0000100100100, t0_0000100100101;
mixer mix_t0_000010010011 (.a(t0_0000100100110), .b(t0_0000100100111), .y(t0_000010010011));
wire t0_0000100100110, t0_0000100100111;
mixer mix_t0_0000100101 (.a(t0_00001001010), .b(t0_00001001011), .y(t0_0000100101));
wire t0_00001001010, t0_00001001011;
mixer mix_t0_00001001010 (.a(t0_000010010100), .b(t0_000010010101), .y(t0_00001001010));
wire t0_000010010100, t0_000010010101;
mixer mix_t0_000010010100 (.a(t0_0000100101000), .b(t0_0000100101001), .y(t0_000010010100));
wire t0_0000100101000, t0_0000100101001;
mixer mix_t0_000010010101 (.a(t0_0000100101010), .b(t0_0000100101011), .y(t0_000010010101));
wire t0_0000100101010, t0_0000100101011;
mixer mix_t0_00001001011 (.a(t0_000010010110), .b(t0_000010010111), .y(t0_00001001011));
wire t0_000010010110, t0_000010010111;
mixer mix_t0_000010010110 (.a(t0_0000100101100), .b(t0_0000100101101), .y(t0_000010010110));
wire t0_0000100101100, t0_0000100101101;
mixer mix_t0_000010010111 (.a(t0_0000100101110), .b(t0_0000100101111), .y(t0_000010010111));
wire t0_0000100101110, t0_0000100101111;
mixer mix_t0_000010011 (.a(t0_0000100110), .b(t0_0000100111), .y(t0_000010011));
wire t0_0000100110, t0_0000100111;
mixer mix_t0_0000100110 (.a(t0_00001001100), .b(t0_00001001101), .y(t0_0000100110));
wire t0_00001001100, t0_00001001101;
mixer mix_t0_00001001100 (.a(t0_000010011000), .b(t0_000010011001), .y(t0_00001001100));
wire t0_000010011000, t0_000010011001;
mixer mix_t0_000010011000 (.a(t0_0000100110000), .b(t0_0000100110001), .y(t0_000010011000));
wire t0_0000100110000, t0_0000100110001;
mixer mix_t0_000010011001 (.a(t0_0000100110010), .b(t0_0000100110011), .y(t0_000010011001));
wire t0_0000100110010, t0_0000100110011;
mixer mix_t0_00001001101 (.a(t0_000010011010), .b(t0_000010011011), .y(t0_00001001101));
wire t0_000010011010, t0_000010011011;
mixer mix_t0_000010011010 (.a(t0_0000100110100), .b(t0_0000100110101), .y(t0_000010011010));
wire t0_0000100110100, t0_0000100110101;
mixer mix_t0_000010011011 (.a(t0_0000100110110), .b(t0_0000100110111), .y(t0_000010011011));
wire t0_0000100110110, t0_0000100110111;
mixer mix_t0_0000100111 (.a(t0_00001001110), .b(t0_00001001111), .y(t0_0000100111));
wire t0_00001001110, t0_00001001111;
mixer mix_t0_00001001110 (.a(t0_000010011100), .b(t0_000010011101), .y(t0_00001001110));
wire t0_000010011100, t0_000010011101;
mixer mix_t0_000010011100 (.a(t0_0000100111000), .b(t0_0000100111001), .y(t0_000010011100));
wire t0_0000100111000, t0_0000100111001;
mixer mix_t0_000010011101 (.a(t0_0000100111010), .b(t0_0000100111011), .y(t0_000010011101));
wire t0_0000100111010, t0_0000100111011;
mixer mix_t0_00001001111 (.a(t0_000010011110), .b(t0_000010011111), .y(t0_00001001111));
wire t0_000010011110, t0_000010011111;
mixer mix_t0_000010011110 (.a(t0_0000100111100), .b(t0_0000100111101), .y(t0_000010011110));
wire t0_0000100111100, t0_0000100111101;
mixer mix_t0_000010011111 (.a(t0_0000100111110), .b(t0_0000100111111), .y(t0_000010011111));
wire t0_0000100111110, t0_0000100111111;
mixer mix_t0_0000101 (.a(t0_00001010), .b(t0_00001011), .y(t0_0000101));
wire t0_00001010, t0_00001011;
mixer mix_t0_00001010 (.a(t0_000010100), .b(t0_000010101), .y(t0_00001010));
wire t0_000010100, t0_000010101;
mixer mix_t0_000010100 (.a(t0_0000101000), .b(t0_0000101001), .y(t0_000010100));
wire t0_0000101000, t0_0000101001;
mixer mix_t0_0000101000 (.a(t0_00001010000), .b(t0_00001010001), .y(t0_0000101000));
wire t0_00001010000, t0_00001010001;
mixer mix_t0_00001010000 (.a(t0_000010100000), .b(t0_000010100001), .y(t0_00001010000));
wire t0_000010100000, t0_000010100001;
mixer mix_t0_000010100000 (.a(t0_0000101000000), .b(t0_0000101000001), .y(t0_000010100000));
wire t0_0000101000000, t0_0000101000001;
mixer mix_t0_000010100001 (.a(t0_0000101000010), .b(t0_0000101000011), .y(t0_000010100001));
wire t0_0000101000010, t0_0000101000011;
mixer mix_t0_00001010001 (.a(t0_000010100010), .b(t0_000010100011), .y(t0_00001010001));
wire t0_000010100010, t0_000010100011;
mixer mix_t0_000010100010 (.a(t0_0000101000100), .b(t0_0000101000101), .y(t0_000010100010));
wire t0_0000101000100, t0_0000101000101;
mixer mix_t0_000010100011 (.a(t0_0000101000110), .b(t0_0000101000111), .y(t0_000010100011));
wire t0_0000101000110, t0_0000101000111;
mixer mix_t0_0000101001 (.a(t0_00001010010), .b(t0_00001010011), .y(t0_0000101001));
wire t0_00001010010, t0_00001010011;
mixer mix_t0_00001010010 (.a(t0_000010100100), .b(t0_000010100101), .y(t0_00001010010));
wire t0_000010100100, t0_000010100101;
mixer mix_t0_000010100100 (.a(t0_0000101001000), .b(t0_0000101001001), .y(t0_000010100100));
wire t0_0000101001000, t0_0000101001001;
mixer mix_t0_000010100101 (.a(t0_0000101001010), .b(t0_0000101001011), .y(t0_000010100101));
wire t0_0000101001010, t0_0000101001011;
mixer mix_t0_00001010011 (.a(t0_000010100110), .b(t0_000010100111), .y(t0_00001010011));
wire t0_000010100110, t0_000010100111;
mixer mix_t0_000010100110 (.a(t0_0000101001100), .b(t0_0000101001101), .y(t0_000010100110));
wire t0_0000101001100, t0_0000101001101;
mixer mix_t0_000010100111 (.a(t0_0000101001110), .b(t0_0000101001111), .y(t0_000010100111));
wire t0_0000101001110, t0_0000101001111;
mixer mix_t0_000010101 (.a(t0_0000101010), .b(t0_0000101011), .y(t0_000010101));
wire t0_0000101010, t0_0000101011;
mixer mix_t0_0000101010 (.a(t0_00001010100), .b(t0_00001010101), .y(t0_0000101010));
wire t0_00001010100, t0_00001010101;
mixer mix_t0_00001010100 (.a(t0_000010101000), .b(t0_000010101001), .y(t0_00001010100));
wire t0_000010101000, t0_000010101001;
mixer mix_t0_000010101000 (.a(t0_0000101010000), .b(t0_0000101010001), .y(t0_000010101000));
wire t0_0000101010000, t0_0000101010001;
mixer mix_t0_000010101001 (.a(t0_0000101010010), .b(t0_0000101010011), .y(t0_000010101001));
wire t0_0000101010010, t0_0000101010011;
mixer mix_t0_00001010101 (.a(t0_000010101010), .b(t0_000010101011), .y(t0_00001010101));
wire t0_000010101010, t0_000010101011;
mixer mix_t0_000010101010 (.a(t0_0000101010100), .b(t0_0000101010101), .y(t0_000010101010));
wire t0_0000101010100, t0_0000101010101;
mixer mix_t0_000010101011 (.a(t0_0000101010110), .b(t0_0000101010111), .y(t0_000010101011));
wire t0_0000101010110, t0_0000101010111;
mixer mix_t0_0000101011 (.a(t0_00001010110), .b(t0_00001010111), .y(t0_0000101011));
wire t0_00001010110, t0_00001010111;
mixer mix_t0_00001010110 (.a(t0_000010101100), .b(t0_000010101101), .y(t0_00001010110));
wire t0_000010101100, t0_000010101101;
mixer mix_t0_000010101100 (.a(t0_0000101011000), .b(t0_0000101011001), .y(t0_000010101100));
wire t0_0000101011000, t0_0000101011001;
mixer mix_t0_000010101101 (.a(t0_0000101011010), .b(t0_0000101011011), .y(t0_000010101101));
wire t0_0000101011010, t0_0000101011011;
mixer mix_t0_00001010111 (.a(t0_000010101110), .b(t0_000010101111), .y(t0_00001010111));
wire t0_000010101110, t0_000010101111;
mixer mix_t0_000010101110 (.a(t0_0000101011100), .b(t0_0000101011101), .y(t0_000010101110));
wire t0_0000101011100, t0_0000101011101;
mixer mix_t0_000010101111 (.a(t0_0000101011110), .b(t0_0000101011111), .y(t0_000010101111));
wire t0_0000101011110, t0_0000101011111;
mixer mix_t0_00001011 (.a(t0_000010110), .b(t0_000010111), .y(t0_00001011));
wire t0_000010110, t0_000010111;
mixer mix_t0_000010110 (.a(t0_0000101100), .b(t0_0000101101), .y(t0_000010110));
wire t0_0000101100, t0_0000101101;
mixer mix_t0_0000101100 (.a(t0_00001011000), .b(t0_00001011001), .y(t0_0000101100));
wire t0_00001011000, t0_00001011001;
mixer mix_t0_00001011000 (.a(t0_000010110000), .b(t0_000010110001), .y(t0_00001011000));
wire t0_000010110000, t0_000010110001;
mixer mix_t0_000010110000 (.a(t0_0000101100000), .b(t0_0000101100001), .y(t0_000010110000));
wire t0_0000101100000, t0_0000101100001;
mixer mix_t0_000010110001 (.a(t0_0000101100010), .b(t0_0000101100011), .y(t0_000010110001));
wire t0_0000101100010, t0_0000101100011;
mixer mix_t0_00001011001 (.a(t0_000010110010), .b(t0_000010110011), .y(t0_00001011001));
wire t0_000010110010, t0_000010110011;
mixer mix_t0_000010110010 (.a(t0_0000101100100), .b(t0_0000101100101), .y(t0_000010110010));
wire t0_0000101100100, t0_0000101100101;
mixer mix_t0_000010110011 (.a(t0_0000101100110), .b(t0_0000101100111), .y(t0_000010110011));
wire t0_0000101100110, t0_0000101100111;
mixer mix_t0_0000101101 (.a(t0_00001011010), .b(t0_00001011011), .y(t0_0000101101));
wire t0_00001011010, t0_00001011011;
mixer mix_t0_00001011010 (.a(t0_000010110100), .b(t0_000010110101), .y(t0_00001011010));
wire t0_000010110100, t0_000010110101;
mixer mix_t0_000010110100 (.a(t0_0000101101000), .b(t0_0000101101001), .y(t0_000010110100));
wire t0_0000101101000, t0_0000101101001;
mixer mix_t0_000010110101 (.a(t0_0000101101010), .b(t0_0000101101011), .y(t0_000010110101));
wire t0_0000101101010, t0_0000101101011;
mixer mix_t0_00001011011 (.a(t0_000010110110), .b(t0_000010110111), .y(t0_00001011011));
wire t0_000010110110, t0_000010110111;
mixer mix_t0_000010110110 (.a(t0_0000101101100), .b(t0_0000101101101), .y(t0_000010110110));
wire t0_0000101101100, t0_0000101101101;
mixer mix_t0_000010110111 (.a(t0_0000101101110), .b(t0_0000101101111), .y(t0_000010110111));
wire t0_0000101101110, t0_0000101101111;
mixer mix_t0_000010111 (.a(t0_0000101110), .b(t0_0000101111), .y(t0_000010111));
wire t0_0000101110, t0_0000101111;
mixer mix_t0_0000101110 (.a(t0_00001011100), .b(t0_00001011101), .y(t0_0000101110));
wire t0_00001011100, t0_00001011101;
mixer mix_t0_00001011100 (.a(t0_000010111000), .b(t0_000010111001), .y(t0_00001011100));
wire t0_000010111000, t0_000010111001;
mixer mix_t0_000010111000 (.a(t0_0000101110000), .b(t0_0000101110001), .y(t0_000010111000));
wire t0_0000101110000, t0_0000101110001;
mixer mix_t0_000010111001 (.a(t0_0000101110010), .b(t0_0000101110011), .y(t0_000010111001));
wire t0_0000101110010, t0_0000101110011;
mixer mix_t0_00001011101 (.a(t0_000010111010), .b(t0_000010111011), .y(t0_00001011101));
wire t0_000010111010, t0_000010111011;
mixer mix_t0_000010111010 (.a(t0_0000101110100), .b(t0_0000101110101), .y(t0_000010111010));
wire t0_0000101110100, t0_0000101110101;
mixer mix_t0_000010111011 (.a(t0_0000101110110), .b(t0_0000101110111), .y(t0_000010111011));
wire t0_0000101110110, t0_0000101110111;
mixer mix_t0_0000101111 (.a(t0_00001011110), .b(t0_00001011111), .y(t0_0000101111));
wire t0_00001011110, t0_00001011111;
mixer mix_t0_00001011110 (.a(t0_000010111100), .b(t0_000010111101), .y(t0_00001011110));
wire t0_000010111100, t0_000010111101;
mixer mix_t0_000010111100 (.a(t0_0000101111000), .b(t0_0000101111001), .y(t0_000010111100));
wire t0_0000101111000, t0_0000101111001;
mixer mix_t0_000010111101 (.a(t0_0000101111010), .b(t0_0000101111011), .y(t0_000010111101));
wire t0_0000101111010, t0_0000101111011;
mixer mix_t0_00001011111 (.a(t0_000010111110), .b(t0_000010111111), .y(t0_00001011111));
wire t0_000010111110, t0_000010111111;
mixer mix_t0_000010111110 (.a(t0_0000101111100), .b(t0_0000101111101), .y(t0_000010111110));
wire t0_0000101111100, t0_0000101111101;
mixer mix_t0_000010111111 (.a(t0_0000101111110), .b(t0_0000101111111), .y(t0_000010111111));
wire t0_0000101111110, t0_0000101111111;
mixer mix_t0_000011 (.a(t0_0000110), .b(t0_0000111), .y(t0_000011));
wire t0_0000110, t0_0000111;
mixer mix_t0_0000110 (.a(t0_00001100), .b(t0_00001101), .y(t0_0000110));
wire t0_00001100, t0_00001101;
mixer mix_t0_00001100 (.a(t0_000011000), .b(t0_000011001), .y(t0_00001100));
wire t0_000011000, t0_000011001;
mixer mix_t0_000011000 (.a(t0_0000110000), .b(t0_0000110001), .y(t0_000011000));
wire t0_0000110000, t0_0000110001;
mixer mix_t0_0000110000 (.a(t0_00001100000), .b(t0_00001100001), .y(t0_0000110000));
wire t0_00001100000, t0_00001100001;
mixer mix_t0_00001100000 (.a(t0_000011000000), .b(t0_000011000001), .y(t0_00001100000));
wire t0_000011000000, t0_000011000001;
mixer mix_t0_000011000000 (.a(t0_0000110000000), .b(t0_0000110000001), .y(t0_000011000000));
wire t0_0000110000000, t0_0000110000001;
mixer mix_t0_000011000001 (.a(t0_0000110000010), .b(t0_0000110000011), .y(t0_000011000001));
wire t0_0000110000010, t0_0000110000011;
mixer mix_t0_00001100001 (.a(t0_000011000010), .b(t0_000011000011), .y(t0_00001100001));
wire t0_000011000010, t0_000011000011;
mixer mix_t0_000011000010 (.a(t0_0000110000100), .b(t0_0000110000101), .y(t0_000011000010));
wire t0_0000110000100, t0_0000110000101;
mixer mix_t0_000011000011 (.a(t0_0000110000110), .b(t0_0000110000111), .y(t0_000011000011));
wire t0_0000110000110, t0_0000110000111;
mixer mix_t0_0000110001 (.a(t0_00001100010), .b(t0_00001100011), .y(t0_0000110001));
wire t0_00001100010, t0_00001100011;
mixer mix_t0_00001100010 (.a(t0_000011000100), .b(t0_000011000101), .y(t0_00001100010));
wire t0_000011000100, t0_000011000101;
mixer mix_t0_000011000100 (.a(t0_0000110001000), .b(t0_0000110001001), .y(t0_000011000100));
wire t0_0000110001000, t0_0000110001001;
mixer mix_t0_000011000101 (.a(t0_0000110001010), .b(t0_0000110001011), .y(t0_000011000101));
wire t0_0000110001010, t0_0000110001011;
mixer mix_t0_00001100011 (.a(t0_000011000110), .b(t0_000011000111), .y(t0_00001100011));
wire t0_000011000110, t0_000011000111;
mixer mix_t0_000011000110 (.a(t0_0000110001100), .b(t0_0000110001101), .y(t0_000011000110));
wire t0_0000110001100, t0_0000110001101;
mixer mix_t0_000011000111 (.a(t0_0000110001110), .b(t0_0000110001111), .y(t0_000011000111));
wire t0_0000110001110, t0_0000110001111;
mixer mix_t0_000011001 (.a(t0_0000110010), .b(t0_0000110011), .y(t0_000011001));
wire t0_0000110010, t0_0000110011;
mixer mix_t0_0000110010 (.a(t0_00001100100), .b(t0_00001100101), .y(t0_0000110010));
wire t0_00001100100, t0_00001100101;
mixer mix_t0_00001100100 (.a(t0_000011001000), .b(t0_000011001001), .y(t0_00001100100));
wire t0_000011001000, t0_000011001001;
mixer mix_t0_000011001000 (.a(t0_0000110010000), .b(t0_0000110010001), .y(t0_000011001000));
wire t0_0000110010000, t0_0000110010001;
mixer mix_t0_000011001001 (.a(t0_0000110010010), .b(t0_0000110010011), .y(t0_000011001001));
wire t0_0000110010010, t0_0000110010011;
mixer mix_t0_00001100101 (.a(t0_000011001010), .b(t0_000011001011), .y(t0_00001100101));
wire t0_000011001010, t0_000011001011;
mixer mix_t0_000011001010 (.a(t0_0000110010100), .b(t0_0000110010101), .y(t0_000011001010));
wire t0_0000110010100, t0_0000110010101;
mixer mix_t0_000011001011 (.a(t0_0000110010110), .b(t0_0000110010111), .y(t0_000011001011));
wire t0_0000110010110, t0_0000110010111;
mixer mix_t0_0000110011 (.a(t0_00001100110), .b(t0_00001100111), .y(t0_0000110011));
wire t0_00001100110, t0_00001100111;
mixer mix_t0_00001100110 (.a(t0_000011001100), .b(t0_000011001101), .y(t0_00001100110));
wire t0_000011001100, t0_000011001101;
mixer mix_t0_000011001100 (.a(t0_0000110011000), .b(t0_0000110011001), .y(t0_000011001100));
wire t0_0000110011000, t0_0000110011001;
mixer mix_t0_000011001101 (.a(t0_0000110011010), .b(t0_0000110011011), .y(t0_000011001101));
wire t0_0000110011010, t0_0000110011011;
mixer mix_t0_00001100111 (.a(t0_000011001110), .b(t0_000011001111), .y(t0_00001100111));
wire t0_000011001110, t0_000011001111;
mixer mix_t0_000011001110 (.a(t0_0000110011100), .b(t0_0000110011101), .y(t0_000011001110));
wire t0_0000110011100, t0_0000110011101;
mixer mix_t0_000011001111 (.a(t0_0000110011110), .b(t0_0000110011111), .y(t0_000011001111));
wire t0_0000110011110, t0_0000110011111;
mixer mix_t0_00001101 (.a(t0_000011010), .b(t0_000011011), .y(t0_00001101));
wire t0_000011010, t0_000011011;
mixer mix_t0_000011010 (.a(t0_0000110100), .b(t0_0000110101), .y(t0_000011010));
wire t0_0000110100, t0_0000110101;
mixer mix_t0_0000110100 (.a(t0_00001101000), .b(t0_00001101001), .y(t0_0000110100));
wire t0_00001101000, t0_00001101001;
mixer mix_t0_00001101000 (.a(t0_000011010000), .b(t0_000011010001), .y(t0_00001101000));
wire t0_000011010000, t0_000011010001;
mixer mix_t0_000011010000 (.a(t0_0000110100000), .b(t0_0000110100001), .y(t0_000011010000));
wire t0_0000110100000, t0_0000110100001;
mixer mix_t0_000011010001 (.a(t0_0000110100010), .b(t0_0000110100011), .y(t0_000011010001));
wire t0_0000110100010, t0_0000110100011;
mixer mix_t0_00001101001 (.a(t0_000011010010), .b(t0_000011010011), .y(t0_00001101001));
wire t0_000011010010, t0_000011010011;
mixer mix_t0_000011010010 (.a(t0_0000110100100), .b(t0_0000110100101), .y(t0_000011010010));
wire t0_0000110100100, t0_0000110100101;
mixer mix_t0_000011010011 (.a(t0_0000110100110), .b(t0_0000110100111), .y(t0_000011010011));
wire t0_0000110100110, t0_0000110100111;
mixer mix_t0_0000110101 (.a(t0_00001101010), .b(t0_00001101011), .y(t0_0000110101));
wire t0_00001101010, t0_00001101011;
mixer mix_t0_00001101010 (.a(t0_000011010100), .b(t0_000011010101), .y(t0_00001101010));
wire t0_000011010100, t0_000011010101;
mixer mix_t0_000011010100 (.a(t0_0000110101000), .b(t0_0000110101001), .y(t0_000011010100));
wire t0_0000110101000, t0_0000110101001;
mixer mix_t0_000011010101 (.a(t0_0000110101010), .b(t0_0000110101011), .y(t0_000011010101));
wire t0_0000110101010, t0_0000110101011;
mixer mix_t0_00001101011 (.a(t0_000011010110), .b(t0_000011010111), .y(t0_00001101011));
wire t0_000011010110, t0_000011010111;
mixer mix_t0_000011010110 (.a(t0_0000110101100), .b(t0_0000110101101), .y(t0_000011010110));
wire t0_0000110101100, t0_0000110101101;
mixer mix_t0_000011010111 (.a(t0_0000110101110), .b(t0_0000110101111), .y(t0_000011010111));
wire t0_0000110101110, t0_0000110101111;
mixer mix_t0_000011011 (.a(t0_0000110110), .b(t0_0000110111), .y(t0_000011011));
wire t0_0000110110, t0_0000110111;
mixer mix_t0_0000110110 (.a(t0_00001101100), .b(t0_00001101101), .y(t0_0000110110));
wire t0_00001101100, t0_00001101101;
mixer mix_t0_00001101100 (.a(t0_000011011000), .b(t0_000011011001), .y(t0_00001101100));
wire t0_000011011000, t0_000011011001;
mixer mix_t0_000011011000 (.a(t0_0000110110000), .b(t0_0000110110001), .y(t0_000011011000));
wire t0_0000110110000, t0_0000110110001;
mixer mix_t0_000011011001 (.a(t0_0000110110010), .b(t0_0000110110011), .y(t0_000011011001));
wire t0_0000110110010, t0_0000110110011;
mixer mix_t0_00001101101 (.a(t0_000011011010), .b(t0_000011011011), .y(t0_00001101101));
wire t0_000011011010, t0_000011011011;
mixer mix_t0_000011011010 (.a(t0_0000110110100), .b(t0_0000110110101), .y(t0_000011011010));
wire t0_0000110110100, t0_0000110110101;
mixer mix_t0_000011011011 (.a(t0_0000110110110), .b(t0_0000110110111), .y(t0_000011011011));
wire t0_0000110110110, t0_0000110110111;
mixer mix_t0_0000110111 (.a(t0_00001101110), .b(t0_00001101111), .y(t0_0000110111));
wire t0_00001101110, t0_00001101111;
mixer mix_t0_00001101110 (.a(t0_000011011100), .b(t0_000011011101), .y(t0_00001101110));
wire t0_000011011100, t0_000011011101;
mixer mix_t0_000011011100 (.a(t0_0000110111000), .b(t0_0000110111001), .y(t0_000011011100));
wire t0_0000110111000, t0_0000110111001;
mixer mix_t0_000011011101 (.a(t0_0000110111010), .b(t0_0000110111011), .y(t0_000011011101));
wire t0_0000110111010, t0_0000110111011;
mixer mix_t0_00001101111 (.a(t0_000011011110), .b(t0_000011011111), .y(t0_00001101111));
wire t0_000011011110, t0_000011011111;
mixer mix_t0_000011011110 (.a(t0_0000110111100), .b(t0_0000110111101), .y(t0_000011011110));
wire t0_0000110111100, t0_0000110111101;
mixer mix_t0_000011011111 (.a(t0_0000110111110), .b(t0_0000110111111), .y(t0_000011011111));
wire t0_0000110111110, t0_0000110111111;
mixer mix_t0_0000111 (.a(t0_00001110), .b(t0_00001111), .y(t0_0000111));
wire t0_00001110, t0_00001111;
mixer mix_t0_00001110 (.a(t0_000011100), .b(t0_000011101), .y(t0_00001110));
wire t0_000011100, t0_000011101;
mixer mix_t0_000011100 (.a(t0_0000111000), .b(t0_0000111001), .y(t0_000011100));
wire t0_0000111000, t0_0000111001;
mixer mix_t0_0000111000 (.a(t0_00001110000), .b(t0_00001110001), .y(t0_0000111000));
wire t0_00001110000, t0_00001110001;
mixer mix_t0_00001110000 (.a(t0_000011100000), .b(t0_000011100001), .y(t0_00001110000));
wire t0_000011100000, t0_000011100001;
mixer mix_t0_000011100000 (.a(t0_0000111000000), .b(t0_0000111000001), .y(t0_000011100000));
wire t0_0000111000000, t0_0000111000001;
mixer mix_t0_000011100001 (.a(t0_0000111000010), .b(t0_0000111000011), .y(t0_000011100001));
wire t0_0000111000010, t0_0000111000011;
mixer mix_t0_00001110001 (.a(t0_000011100010), .b(t0_000011100011), .y(t0_00001110001));
wire t0_000011100010, t0_000011100011;
mixer mix_t0_000011100010 (.a(t0_0000111000100), .b(t0_0000111000101), .y(t0_000011100010));
wire t0_0000111000100, t0_0000111000101;
mixer mix_t0_000011100011 (.a(t0_0000111000110), .b(t0_0000111000111), .y(t0_000011100011));
wire t0_0000111000110, t0_0000111000111;
mixer mix_t0_0000111001 (.a(t0_00001110010), .b(t0_00001110011), .y(t0_0000111001));
wire t0_00001110010, t0_00001110011;
mixer mix_t0_00001110010 (.a(t0_000011100100), .b(t0_000011100101), .y(t0_00001110010));
wire t0_000011100100, t0_000011100101;
mixer mix_t0_000011100100 (.a(t0_0000111001000), .b(t0_0000111001001), .y(t0_000011100100));
wire t0_0000111001000, t0_0000111001001;
mixer mix_t0_000011100101 (.a(t0_0000111001010), .b(t0_0000111001011), .y(t0_000011100101));
wire t0_0000111001010, t0_0000111001011;
mixer mix_t0_00001110011 (.a(t0_000011100110), .b(t0_000011100111), .y(t0_00001110011));
wire t0_000011100110, t0_000011100111;
mixer mix_t0_000011100110 (.a(t0_0000111001100), .b(t0_0000111001101), .y(t0_000011100110));
wire t0_0000111001100, t0_0000111001101;
mixer mix_t0_000011100111 (.a(t0_0000111001110), .b(t0_0000111001111), .y(t0_000011100111));
wire t0_0000111001110, t0_0000111001111;
mixer mix_t0_000011101 (.a(t0_0000111010), .b(t0_0000111011), .y(t0_000011101));
wire t0_0000111010, t0_0000111011;
mixer mix_t0_0000111010 (.a(t0_00001110100), .b(t0_00001110101), .y(t0_0000111010));
wire t0_00001110100, t0_00001110101;
mixer mix_t0_00001110100 (.a(t0_000011101000), .b(t0_000011101001), .y(t0_00001110100));
wire t0_000011101000, t0_000011101001;
mixer mix_t0_000011101000 (.a(t0_0000111010000), .b(t0_0000111010001), .y(t0_000011101000));
wire t0_0000111010000, t0_0000111010001;
mixer mix_t0_000011101001 (.a(t0_0000111010010), .b(t0_0000111010011), .y(t0_000011101001));
wire t0_0000111010010, t0_0000111010011;
mixer mix_t0_00001110101 (.a(t0_000011101010), .b(t0_000011101011), .y(t0_00001110101));
wire t0_000011101010, t0_000011101011;
mixer mix_t0_000011101010 (.a(t0_0000111010100), .b(t0_0000111010101), .y(t0_000011101010));
wire t0_0000111010100, t0_0000111010101;
mixer mix_t0_000011101011 (.a(t0_0000111010110), .b(t0_0000111010111), .y(t0_000011101011));
wire t0_0000111010110, t0_0000111010111;
mixer mix_t0_0000111011 (.a(t0_00001110110), .b(t0_00001110111), .y(t0_0000111011));
wire t0_00001110110, t0_00001110111;
mixer mix_t0_00001110110 (.a(t0_000011101100), .b(t0_000011101101), .y(t0_00001110110));
wire t0_000011101100, t0_000011101101;
mixer mix_t0_000011101100 (.a(t0_0000111011000), .b(t0_0000111011001), .y(t0_000011101100));
wire t0_0000111011000, t0_0000111011001;
mixer mix_t0_000011101101 (.a(t0_0000111011010), .b(t0_0000111011011), .y(t0_000011101101));
wire t0_0000111011010, t0_0000111011011;
mixer mix_t0_00001110111 (.a(t0_000011101110), .b(t0_000011101111), .y(t0_00001110111));
wire t0_000011101110, t0_000011101111;
mixer mix_t0_000011101110 (.a(t0_0000111011100), .b(t0_0000111011101), .y(t0_000011101110));
wire t0_0000111011100, t0_0000111011101;
mixer mix_t0_000011101111 (.a(t0_0000111011110), .b(t0_0000111011111), .y(t0_000011101111));
wire t0_0000111011110, t0_0000111011111;
mixer mix_t0_00001111 (.a(t0_000011110), .b(t0_000011111), .y(t0_00001111));
wire t0_000011110, t0_000011111;
mixer mix_t0_000011110 (.a(t0_0000111100), .b(t0_0000111101), .y(t0_000011110));
wire t0_0000111100, t0_0000111101;
mixer mix_t0_0000111100 (.a(t0_00001111000), .b(t0_00001111001), .y(t0_0000111100));
wire t0_00001111000, t0_00001111001;
mixer mix_t0_00001111000 (.a(t0_000011110000), .b(t0_000011110001), .y(t0_00001111000));
wire t0_000011110000, t0_000011110001;
mixer mix_t0_000011110000 (.a(t0_0000111100000), .b(t0_0000111100001), .y(t0_000011110000));
wire t0_0000111100000, t0_0000111100001;
mixer mix_t0_000011110001 (.a(t0_0000111100010), .b(t0_0000111100011), .y(t0_000011110001));
wire t0_0000111100010, t0_0000111100011;
mixer mix_t0_00001111001 (.a(t0_000011110010), .b(t0_000011110011), .y(t0_00001111001));
wire t0_000011110010, t0_000011110011;
mixer mix_t0_000011110010 (.a(t0_0000111100100), .b(t0_0000111100101), .y(t0_000011110010));
wire t0_0000111100100, t0_0000111100101;
mixer mix_t0_000011110011 (.a(t0_0000111100110), .b(t0_0000111100111), .y(t0_000011110011));
wire t0_0000111100110, t0_0000111100111;
mixer mix_t0_0000111101 (.a(t0_00001111010), .b(t0_00001111011), .y(t0_0000111101));
wire t0_00001111010, t0_00001111011;
mixer mix_t0_00001111010 (.a(t0_000011110100), .b(t0_000011110101), .y(t0_00001111010));
wire t0_000011110100, t0_000011110101;
mixer mix_t0_000011110100 (.a(t0_0000111101000), .b(t0_0000111101001), .y(t0_000011110100));
wire t0_0000111101000, t0_0000111101001;
mixer mix_t0_000011110101 (.a(t0_0000111101010), .b(t0_0000111101011), .y(t0_000011110101));
wire t0_0000111101010, t0_0000111101011;
mixer mix_t0_00001111011 (.a(t0_000011110110), .b(t0_000011110111), .y(t0_00001111011));
wire t0_000011110110, t0_000011110111;
mixer mix_t0_000011110110 (.a(t0_0000111101100), .b(t0_0000111101101), .y(t0_000011110110));
wire t0_0000111101100, t0_0000111101101;
mixer mix_t0_000011110111 (.a(t0_0000111101110), .b(t0_0000111101111), .y(t0_000011110111));
wire t0_0000111101110, t0_0000111101111;
mixer mix_t0_000011111 (.a(t0_0000111110), .b(t0_0000111111), .y(t0_000011111));
wire t0_0000111110, t0_0000111111;
mixer mix_t0_0000111110 (.a(t0_00001111100), .b(t0_00001111101), .y(t0_0000111110));
wire t0_00001111100, t0_00001111101;
mixer mix_t0_00001111100 (.a(t0_000011111000), .b(t0_000011111001), .y(t0_00001111100));
wire t0_000011111000, t0_000011111001;
mixer mix_t0_000011111000 (.a(t0_0000111110000), .b(t0_0000111110001), .y(t0_000011111000));
wire t0_0000111110000, t0_0000111110001;
mixer mix_t0_000011111001 (.a(t0_0000111110010), .b(t0_0000111110011), .y(t0_000011111001));
wire t0_0000111110010, t0_0000111110011;
mixer mix_t0_00001111101 (.a(t0_000011111010), .b(t0_000011111011), .y(t0_00001111101));
wire t0_000011111010, t0_000011111011;
mixer mix_t0_000011111010 (.a(t0_0000111110100), .b(t0_0000111110101), .y(t0_000011111010));
wire t0_0000111110100, t0_0000111110101;
mixer mix_t0_000011111011 (.a(t0_0000111110110), .b(t0_0000111110111), .y(t0_000011111011));
wire t0_0000111110110, t0_0000111110111;
mixer mix_t0_0000111111 (.a(t0_00001111110), .b(t0_00001111111), .y(t0_0000111111));
wire t0_00001111110, t0_00001111111;
mixer mix_t0_00001111110 (.a(t0_000011111100), .b(t0_000011111101), .y(t0_00001111110));
wire t0_000011111100, t0_000011111101;
mixer mix_t0_000011111100 (.a(t0_0000111111000), .b(t0_0000111111001), .y(t0_000011111100));
wire t0_0000111111000, t0_0000111111001;
mixer mix_t0_000011111101 (.a(t0_0000111111010), .b(t0_0000111111011), .y(t0_000011111101));
wire t0_0000111111010, t0_0000111111011;
mixer mix_t0_00001111111 (.a(t0_000011111110), .b(t0_000011111111), .y(t0_00001111111));
wire t0_000011111110, t0_000011111111;
mixer mix_t0_000011111110 (.a(t0_0000111111100), .b(t0_0000111111101), .y(t0_000011111110));
wire t0_0000111111100, t0_0000111111101;
mixer mix_t0_000011111111 (.a(t0_0000111111110), .b(t0_0000111111111), .y(t0_000011111111));
wire t0_0000111111110, t0_0000111111111;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_000100 (.a(t0_0001000), .b(t0_0001001), .y(t0_000100));
wire t0_0001000, t0_0001001;
mixer mix_t0_0001000 (.a(t0_00010000), .b(t0_00010001), .y(t0_0001000));
wire t0_00010000, t0_00010001;
mixer mix_t0_00010000 (.a(t0_000100000), .b(t0_000100001), .y(t0_00010000));
wire t0_000100000, t0_000100001;
mixer mix_t0_000100000 (.a(t0_0001000000), .b(t0_0001000001), .y(t0_000100000));
wire t0_0001000000, t0_0001000001;
mixer mix_t0_0001000000 (.a(t0_00010000000), .b(t0_00010000001), .y(t0_0001000000));
wire t0_00010000000, t0_00010000001;
mixer mix_t0_00010000000 (.a(t0_000100000000), .b(t0_000100000001), .y(t0_00010000000));
wire t0_000100000000, t0_000100000001;
mixer mix_t0_000100000000 (.a(t0_0001000000000), .b(t0_0001000000001), .y(t0_000100000000));
wire t0_0001000000000, t0_0001000000001;
mixer mix_t0_000100000001 (.a(t0_0001000000010), .b(t0_0001000000011), .y(t0_000100000001));
wire t0_0001000000010, t0_0001000000011;
mixer mix_t0_00010000001 (.a(t0_000100000010), .b(t0_000100000011), .y(t0_00010000001));
wire t0_000100000010, t0_000100000011;
mixer mix_t0_000100000010 (.a(t0_0001000000100), .b(t0_0001000000101), .y(t0_000100000010));
wire t0_0001000000100, t0_0001000000101;
mixer mix_t0_000100000011 (.a(t0_0001000000110), .b(t0_0001000000111), .y(t0_000100000011));
wire t0_0001000000110, t0_0001000000111;
mixer mix_t0_0001000001 (.a(t0_00010000010), .b(t0_00010000011), .y(t0_0001000001));
wire t0_00010000010, t0_00010000011;
mixer mix_t0_00010000010 (.a(t0_000100000100), .b(t0_000100000101), .y(t0_00010000010));
wire t0_000100000100, t0_000100000101;
mixer mix_t0_000100000100 (.a(t0_0001000001000), .b(t0_0001000001001), .y(t0_000100000100));
wire t0_0001000001000, t0_0001000001001;
mixer mix_t0_000100000101 (.a(t0_0001000001010), .b(t0_0001000001011), .y(t0_000100000101));
wire t0_0001000001010, t0_0001000001011;
mixer mix_t0_00010000011 (.a(t0_000100000110), .b(t0_000100000111), .y(t0_00010000011));
wire t0_000100000110, t0_000100000111;
mixer mix_t0_000100000110 (.a(t0_0001000001100), .b(t0_0001000001101), .y(t0_000100000110));
wire t0_0001000001100, t0_0001000001101;
mixer mix_t0_000100000111 (.a(t0_0001000001110), .b(t0_0001000001111), .y(t0_000100000111));
wire t0_0001000001110, t0_0001000001111;
mixer mix_t0_000100001 (.a(t0_0001000010), .b(t0_0001000011), .y(t0_000100001));
wire t0_0001000010, t0_0001000011;
mixer mix_t0_0001000010 (.a(t0_00010000100), .b(t0_00010000101), .y(t0_0001000010));
wire t0_00010000100, t0_00010000101;
mixer mix_t0_00010000100 (.a(t0_000100001000), .b(t0_000100001001), .y(t0_00010000100));
wire t0_000100001000, t0_000100001001;
mixer mix_t0_000100001000 (.a(t0_0001000010000), .b(t0_0001000010001), .y(t0_000100001000));
wire t0_0001000010000, t0_0001000010001;
mixer mix_t0_000100001001 (.a(t0_0001000010010), .b(t0_0001000010011), .y(t0_000100001001));
wire t0_0001000010010, t0_0001000010011;
mixer mix_t0_00010000101 (.a(t0_000100001010), .b(t0_000100001011), .y(t0_00010000101));
wire t0_000100001010, t0_000100001011;
mixer mix_t0_000100001010 (.a(t0_0001000010100), .b(t0_0001000010101), .y(t0_000100001010));
wire t0_0001000010100, t0_0001000010101;
mixer mix_t0_000100001011 (.a(t0_0001000010110), .b(t0_0001000010111), .y(t0_000100001011));
wire t0_0001000010110, t0_0001000010111;
mixer mix_t0_0001000011 (.a(t0_00010000110), .b(t0_00010000111), .y(t0_0001000011));
wire t0_00010000110, t0_00010000111;
mixer mix_t0_00010000110 (.a(t0_000100001100), .b(t0_000100001101), .y(t0_00010000110));
wire t0_000100001100, t0_000100001101;
mixer mix_t0_000100001100 (.a(t0_0001000011000), .b(t0_0001000011001), .y(t0_000100001100));
wire t0_0001000011000, t0_0001000011001;
mixer mix_t0_000100001101 (.a(t0_0001000011010), .b(t0_0001000011011), .y(t0_000100001101));
wire t0_0001000011010, t0_0001000011011;
mixer mix_t0_00010000111 (.a(t0_000100001110), .b(t0_000100001111), .y(t0_00010000111));
wire t0_000100001110, t0_000100001111;
mixer mix_t0_000100001110 (.a(t0_0001000011100), .b(t0_0001000011101), .y(t0_000100001110));
wire t0_0001000011100, t0_0001000011101;
mixer mix_t0_000100001111 (.a(t0_0001000011110), .b(t0_0001000011111), .y(t0_000100001111));
wire t0_0001000011110, t0_0001000011111;
mixer mix_t0_00010001 (.a(t0_000100010), .b(t0_000100011), .y(t0_00010001));
wire t0_000100010, t0_000100011;
mixer mix_t0_000100010 (.a(t0_0001000100), .b(t0_0001000101), .y(t0_000100010));
wire t0_0001000100, t0_0001000101;
mixer mix_t0_0001000100 (.a(t0_00010001000), .b(t0_00010001001), .y(t0_0001000100));
wire t0_00010001000, t0_00010001001;
mixer mix_t0_00010001000 (.a(t0_000100010000), .b(t0_000100010001), .y(t0_00010001000));
wire t0_000100010000, t0_000100010001;
mixer mix_t0_000100010000 (.a(t0_0001000100000), .b(t0_0001000100001), .y(t0_000100010000));
wire t0_0001000100000, t0_0001000100001;
mixer mix_t0_000100010001 (.a(t0_0001000100010), .b(t0_0001000100011), .y(t0_000100010001));
wire t0_0001000100010, t0_0001000100011;
mixer mix_t0_00010001001 (.a(t0_000100010010), .b(t0_000100010011), .y(t0_00010001001));
wire t0_000100010010, t0_000100010011;
mixer mix_t0_000100010010 (.a(t0_0001000100100), .b(t0_0001000100101), .y(t0_000100010010));
wire t0_0001000100100, t0_0001000100101;
mixer mix_t0_000100010011 (.a(t0_0001000100110), .b(t0_0001000100111), .y(t0_000100010011));
wire t0_0001000100110, t0_0001000100111;
mixer mix_t0_0001000101 (.a(t0_00010001010), .b(t0_00010001011), .y(t0_0001000101));
wire t0_00010001010, t0_00010001011;
mixer mix_t0_00010001010 (.a(t0_000100010100), .b(t0_000100010101), .y(t0_00010001010));
wire t0_000100010100, t0_000100010101;
mixer mix_t0_000100010100 (.a(t0_0001000101000), .b(t0_0001000101001), .y(t0_000100010100));
wire t0_0001000101000, t0_0001000101001;
mixer mix_t0_000100010101 (.a(t0_0001000101010), .b(t0_0001000101011), .y(t0_000100010101));
wire t0_0001000101010, t0_0001000101011;
mixer mix_t0_00010001011 (.a(t0_000100010110), .b(t0_000100010111), .y(t0_00010001011));
wire t0_000100010110, t0_000100010111;
mixer mix_t0_000100010110 (.a(t0_0001000101100), .b(t0_0001000101101), .y(t0_000100010110));
wire t0_0001000101100, t0_0001000101101;
mixer mix_t0_000100010111 (.a(t0_0001000101110), .b(t0_0001000101111), .y(t0_000100010111));
wire t0_0001000101110, t0_0001000101111;
mixer mix_t0_000100011 (.a(t0_0001000110), .b(t0_0001000111), .y(t0_000100011));
wire t0_0001000110, t0_0001000111;
mixer mix_t0_0001000110 (.a(t0_00010001100), .b(t0_00010001101), .y(t0_0001000110));
wire t0_00010001100, t0_00010001101;
mixer mix_t0_00010001100 (.a(t0_000100011000), .b(t0_000100011001), .y(t0_00010001100));
wire t0_000100011000, t0_000100011001;
mixer mix_t0_000100011000 (.a(t0_0001000110000), .b(t0_0001000110001), .y(t0_000100011000));
wire t0_0001000110000, t0_0001000110001;
mixer mix_t0_000100011001 (.a(t0_0001000110010), .b(t0_0001000110011), .y(t0_000100011001));
wire t0_0001000110010, t0_0001000110011;
mixer mix_t0_00010001101 (.a(t0_000100011010), .b(t0_000100011011), .y(t0_00010001101));
wire t0_000100011010, t0_000100011011;
mixer mix_t0_000100011010 (.a(t0_0001000110100), .b(t0_0001000110101), .y(t0_000100011010));
wire t0_0001000110100, t0_0001000110101;
mixer mix_t0_000100011011 (.a(t0_0001000110110), .b(t0_0001000110111), .y(t0_000100011011));
wire t0_0001000110110, t0_0001000110111;
mixer mix_t0_0001000111 (.a(t0_00010001110), .b(t0_00010001111), .y(t0_0001000111));
wire t0_00010001110, t0_00010001111;
mixer mix_t0_00010001110 (.a(t0_000100011100), .b(t0_000100011101), .y(t0_00010001110));
wire t0_000100011100, t0_000100011101;
mixer mix_t0_000100011100 (.a(t0_0001000111000), .b(t0_0001000111001), .y(t0_000100011100));
wire t0_0001000111000, t0_0001000111001;
mixer mix_t0_000100011101 (.a(t0_0001000111010), .b(t0_0001000111011), .y(t0_000100011101));
wire t0_0001000111010, t0_0001000111011;
mixer mix_t0_00010001111 (.a(t0_000100011110), .b(t0_000100011111), .y(t0_00010001111));
wire t0_000100011110, t0_000100011111;
mixer mix_t0_000100011110 (.a(t0_0001000111100), .b(t0_0001000111101), .y(t0_000100011110));
wire t0_0001000111100, t0_0001000111101;
mixer mix_t0_000100011111 (.a(t0_0001000111110), .b(t0_0001000111111), .y(t0_000100011111));
wire t0_0001000111110, t0_0001000111111;
mixer mix_t0_0001001 (.a(t0_00010010), .b(t0_00010011), .y(t0_0001001));
wire t0_00010010, t0_00010011;
mixer mix_t0_00010010 (.a(t0_000100100), .b(t0_000100101), .y(t0_00010010));
wire t0_000100100, t0_000100101;
mixer mix_t0_000100100 (.a(t0_0001001000), .b(t0_0001001001), .y(t0_000100100));
wire t0_0001001000, t0_0001001001;
mixer mix_t0_0001001000 (.a(t0_00010010000), .b(t0_00010010001), .y(t0_0001001000));
wire t0_00010010000, t0_00010010001;
mixer mix_t0_00010010000 (.a(t0_000100100000), .b(t0_000100100001), .y(t0_00010010000));
wire t0_000100100000, t0_000100100001;
mixer mix_t0_000100100000 (.a(t0_0001001000000), .b(t0_0001001000001), .y(t0_000100100000));
wire t0_0001001000000, t0_0001001000001;
mixer mix_t0_000100100001 (.a(t0_0001001000010), .b(t0_0001001000011), .y(t0_000100100001));
wire t0_0001001000010, t0_0001001000011;
mixer mix_t0_00010010001 (.a(t0_000100100010), .b(t0_000100100011), .y(t0_00010010001));
wire t0_000100100010, t0_000100100011;
mixer mix_t0_000100100010 (.a(t0_0001001000100), .b(t0_0001001000101), .y(t0_000100100010));
wire t0_0001001000100, t0_0001001000101;
mixer mix_t0_000100100011 (.a(t0_0001001000110), .b(t0_0001001000111), .y(t0_000100100011));
wire t0_0001001000110, t0_0001001000111;
mixer mix_t0_0001001001 (.a(t0_00010010010), .b(t0_00010010011), .y(t0_0001001001));
wire t0_00010010010, t0_00010010011;
mixer mix_t0_00010010010 (.a(t0_000100100100), .b(t0_000100100101), .y(t0_00010010010));
wire t0_000100100100, t0_000100100101;
mixer mix_t0_000100100100 (.a(t0_0001001001000), .b(t0_0001001001001), .y(t0_000100100100));
wire t0_0001001001000, t0_0001001001001;
mixer mix_t0_000100100101 (.a(t0_0001001001010), .b(t0_0001001001011), .y(t0_000100100101));
wire t0_0001001001010, t0_0001001001011;
mixer mix_t0_00010010011 (.a(t0_000100100110), .b(t0_000100100111), .y(t0_00010010011));
wire t0_000100100110, t0_000100100111;
mixer mix_t0_000100100110 (.a(t0_0001001001100), .b(t0_0001001001101), .y(t0_000100100110));
wire t0_0001001001100, t0_0001001001101;
mixer mix_t0_000100100111 (.a(t0_0001001001110), .b(t0_0001001001111), .y(t0_000100100111));
wire t0_0001001001110, t0_0001001001111;
mixer mix_t0_000100101 (.a(t0_0001001010), .b(t0_0001001011), .y(t0_000100101));
wire t0_0001001010, t0_0001001011;
mixer mix_t0_0001001010 (.a(t0_00010010100), .b(t0_00010010101), .y(t0_0001001010));
wire t0_00010010100, t0_00010010101;
mixer mix_t0_00010010100 (.a(t0_000100101000), .b(t0_000100101001), .y(t0_00010010100));
wire t0_000100101000, t0_000100101001;
mixer mix_t0_000100101000 (.a(t0_0001001010000), .b(t0_0001001010001), .y(t0_000100101000));
wire t0_0001001010000, t0_0001001010001;
mixer mix_t0_000100101001 (.a(t0_0001001010010), .b(t0_0001001010011), .y(t0_000100101001));
wire t0_0001001010010, t0_0001001010011;
mixer mix_t0_00010010101 (.a(t0_000100101010), .b(t0_000100101011), .y(t0_00010010101));
wire t0_000100101010, t0_000100101011;
mixer mix_t0_000100101010 (.a(t0_0001001010100), .b(t0_0001001010101), .y(t0_000100101010));
wire t0_0001001010100, t0_0001001010101;
mixer mix_t0_000100101011 (.a(t0_0001001010110), .b(t0_0001001010111), .y(t0_000100101011));
wire t0_0001001010110, t0_0001001010111;
mixer mix_t0_0001001011 (.a(t0_00010010110), .b(t0_00010010111), .y(t0_0001001011));
wire t0_00010010110, t0_00010010111;
mixer mix_t0_00010010110 (.a(t0_000100101100), .b(t0_000100101101), .y(t0_00010010110));
wire t0_000100101100, t0_000100101101;
mixer mix_t0_000100101100 (.a(t0_0001001011000), .b(t0_0001001011001), .y(t0_000100101100));
wire t0_0001001011000, t0_0001001011001;
mixer mix_t0_000100101101 (.a(t0_0001001011010), .b(t0_0001001011011), .y(t0_000100101101));
wire t0_0001001011010, t0_0001001011011;
mixer mix_t0_00010010111 (.a(t0_000100101110), .b(t0_000100101111), .y(t0_00010010111));
wire t0_000100101110, t0_000100101111;
mixer mix_t0_000100101110 (.a(t0_0001001011100), .b(t0_0001001011101), .y(t0_000100101110));
wire t0_0001001011100, t0_0001001011101;
mixer mix_t0_000100101111 (.a(t0_0001001011110), .b(t0_0001001011111), .y(t0_000100101111));
wire t0_0001001011110, t0_0001001011111;
mixer mix_t0_00010011 (.a(t0_000100110), .b(t0_000100111), .y(t0_00010011));
wire t0_000100110, t0_000100111;
mixer mix_t0_000100110 (.a(t0_0001001100), .b(t0_0001001101), .y(t0_000100110));
wire t0_0001001100, t0_0001001101;
mixer mix_t0_0001001100 (.a(t0_00010011000), .b(t0_00010011001), .y(t0_0001001100));
wire t0_00010011000, t0_00010011001;
mixer mix_t0_00010011000 (.a(t0_000100110000), .b(t0_000100110001), .y(t0_00010011000));
wire t0_000100110000, t0_000100110001;
mixer mix_t0_000100110000 (.a(t0_0001001100000), .b(t0_0001001100001), .y(t0_000100110000));
wire t0_0001001100000, t0_0001001100001;
mixer mix_t0_000100110001 (.a(t0_0001001100010), .b(t0_0001001100011), .y(t0_000100110001));
wire t0_0001001100010, t0_0001001100011;
mixer mix_t0_00010011001 (.a(t0_000100110010), .b(t0_000100110011), .y(t0_00010011001));
wire t0_000100110010, t0_000100110011;
mixer mix_t0_000100110010 (.a(t0_0001001100100), .b(t0_0001001100101), .y(t0_000100110010));
wire t0_0001001100100, t0_0001001100101;
mixer mix_t0_000100110011 (.a(t0_0001001100110), .b(t0_0001001100111), .y(t0_000100110011));
wire t0_0001001100110, t0_0001001100111;
mixer mix_t0_0001001101 (.a(t0_00010011010), .b(t0_00010011011), .y(t0_0001001101));
wire t0_00010011010, t0_00010011011;
mixer mix_t0_00010011010 (.a(t0_000100110100), .b(t0_000100110101), .y(t0_00010011010));
wire t0_000100110100, t0_000100110101;
mixer mix_t0_000100110100 (.a(t0_0001001101000), .b(t0_0001001101001), .y(t0_000100110100));
wire t0_0001001101000, t0_0001001101001;
mixer mix_t0_000100110101 (.a(t0_0001001101010), .b(t0_0001001101011), .y(t0_000100110101));
wire t0_0001001101010, t0_0001001101011;
mixer mix_t0_00010011011 (.a(t0_000100110110), .b(t0_000100110111), .y(t0_00010011011));
wire t0_000100110110, t0_000100110111;
mixer mix_t0_000100110110 (.a(t0_0001001101100), .b(t0_0001001101101), .y(t0_000100110110));
wire t0_0001001101100, t0_0001001101101;
mixer mix_t0_000100110111 (.a(t0_0001001101110), .b(t0_0001001101111), .y(t0_000100110111));
wire t0_0001001101110, t0_0001001101111;
mixer mix_t0_000100111 (.a(t0_0001001110), .b(t0_0001001111), .y(t0_000100111));
wire t0_0001001110, t0_0001001111;
mixer mix_t0_0001001110 (.a(t0_00010011100), .b(t0_00010011101), .y(t0_0001001110));
wire t0_00010011100, t0_00010011101;
mixer mix_t0_00010011100 (.a(t0_000100111000), .b(t0_000100111001), .y(t0_00010011100));
wire t0_000100111000, t0_000100111001;
mixer mix_t0_000100111000 (.a(t0_0001001110000), .b(t0_0001001110001), .y(t0_000100111000));
wire t0_0001001110000, t0_0001001110001;
mixer mix_t0_000100111001 (.a(t0_0001001110010), .b(t0_0001001110011), .y(t0_000100111001));
wire t0_0001001110010, t0_0001001110011;
mixer mix_t0_00010011101 (.a(t0_000100111010), .b(t0_000100111011), .y(t0_00010011101));
wire t0_000100111010, t0_000100111011;
mixer mix_t0_000100111010 (.a(t0_0001001110100), .b(t0_0001001110101), .y(t0_000100111010));
wire t0_0001001110100, t0_0001001110101;
mixer mix_t0_000100111011 (.a(t0_0001001110110), .b(t0_0001001110111), .y(t0_000100111011));
wire t0_0001001110110, t0_0001001110111;
mixer mix_t0_0001001111 (.a(t0_00010011110), .b(t0_00010011111), .y(t0_0001001111));
wire t0_00010011110, t0_00010011111;
mixer mix_t0_00010011110 (.a(t0_000100111100), .b(t0_000100111101), .y(t0_00010011110));
wire t0_000100111100, t0_000100111101;
mixer mix_t0_000100111100 (.a(t0_0001001111000), .b(t0_0001001111001), .y(t0_000100111100));
wire t0_0001001111000, t0_0001001111001;
mixer mix_t0_000100111101 (.a(t0_0001001111010), .b(t0_0001001111011), .y(t0_000100111101));
wire t0_0001001111010, t0_0001001111011;
mixer mix_t0_00010011111 (.a(t0_000100111110), .b(t0_000100111111), .y(t0_00010011111));
wire t0_000100111110, t0_000100111111;
mixer mix_t0_000100111110 (.a(t0_0001001111100), .b(t0_0001001111101), .y(t0_000100111110));
wire t0_0001001111100, t0_0001001111101;
mixer mix_t0_000100111111 (.a(t0_0001001111110), .b(t0_0001001111111), .y(t0_000100111111));
wire t0_0001001111110, t0_0001001111111;
mixer mix_t0_000101 (.a(t0_0001010), .b(t0_0001011), .y(t0_000101));
wire t0_0001010, t0_0001011;
mixer mix_t0_0001010 (.a(t0_00010100), .b(t0_00010101), .y(t0_0001010));
wire t0_00010100, t0_00010101;
mixer mix_t0_00010100 (.a(t0_000101000), .b(t0_000101001), .y(t0_00010100));
wire t0_000101000, t0_000101001;
mixer mix_t0_000101000 (.a(t0_0001010000), .b(t0_0001010001), .y(t0_000101000));
wire t0_0001010000, t0_0001010001;
mixer mix_t0_0001010000 (.a(t0_00010100000), .b(t0_00010100001), .y(t0_0001010000));
wire t0_00010100000, t0_00010100001;
mixer mix_t0_00010100000 (.a(t0_000101000000), .b(t0_000101000001), .y(t0_00010100000));
wire t0_000101000000, t0_000101000001;
mixer mix_t0_000101000000 (.a(t0_0001010000000), .b(t0_0001010000001), .y(t0_000101000000));
wire t0_0001010000000, t0_0001010000001;
mixer mix_t0_000101000001 (.a(t0_0001010000010), .b(t0_0001010000011), .y(t0_000101000001));
wire t0_0001010000010, t0_0001010000011;
mixer mix_t0_00010100001 (.a(t0_000101000010), .b(t0_000101000011), .y(t0_00010100001));
wire t0_000101000010, t0_000101000011;
mixer mix_t0_000101000010 (.a(t0_0001010000100), .b(t0_0001010000101), .y(t0_000101000010));
wire t0_0001010000100, t0_0001010000101;
mixer mix_t0_000101000011 (.a(t0_0001010000110), .b(t0_0001010000111), .y(t0_000101000011));
wire t0_0001010000110, t0_0001010000111;
mixer mix_t0_0001010001 (.a(t0_00010100010), .b(t0_00010100011), .y(t0_0001010001));
wire t0_00010100010, t0_00010100011;
mixer mix_t0_00010100010 (.a(t0_000101000100), .b(t0_000101000101), .y(t0_00010100010));
wire t0_000101000100, t0_000101000101;
mixer mix_t0_000101000100 (.a(t0_0001010001000), .b(t0_0001010001001), .y(t0_000101000100));
wire t0_0001010001000, t0_0001010001001;
mixer mix_t0_000101000101 (.a(t0_0001010001010), .b(t0_0001010001011), .y(t0_000101000101));
wire t0_0001010001010, t0_0001010001011;
mixer mix_t0_00010100011 (.a(t0_000101000110), .b(t0_000101000111), .y(t0_00010100011));
wire t0_000101000110, t0_000101000111;
mixer mix_t0_000101000110 (.a(t0_0001010001100), .b(t0_0001010001101), .y(t0_000101000110));
wire t0_0001010001100, t0_0001010001101;
mixer mix_t0_000101000111 (.a(t0_0001010001110), .b(t0_0001010001111), .y(t0_000101000111));
wire t0_0001010001110, t0_0001010001111;
mixer mix_t0_000101001 (.a(t0_0001010010), .b(t0_0001010011), .y(t0_000101001));
wire t0_0001010010, t0_0001010011;
mixer mix_t0_0001010010 (.a(t0_00010100100), .b(t0_00010100101), .y(t0_0001010010));
wire t0_00010100100, t0_00010100101;
mixer mix_t0_00010100100 (.a(t0_000101001000), .b(t0_000101001001), .y(t0_00010100100));
wire t0_000101001000, t0_000101001001;
mixer mix_t0_000101001000 (.a(t0_0001010010000), .b(t0_0001010010001), .y(t0_000101001000));
wire t0_0001010010000, t0_0001010010001;
mixer mix_t0_000101001001 (.a(t0_0001010010010), .b(t0_0001010010011), .y(t0_000101001001));
wire t0_0001010010010, t0_0001010010011;
mixer mix_t0_00010100101 (.a(t0_000101001010), .b(t0_000101001011), .y(t0_00010100101));
wire t0_000101001010, t0_000101001011;
mixer mix_t0_000101001010 (.a(t0_0001010010100), .b(t0_0001010010101), .y(t0_000101001010));
wire t0_0001010010100, t0_0001010010101;
mixer mix_t0_000101001011 (.a(t0_0001010010110), .b(t0_0001010010111), .y(t0_000101001011));
wire t0_0001010010110, t0_0001010010111;
mixer mix_t0_0001010011 (.a(t0_00010100110), .b(t0_00010100111), .y(t0_0001010011));
wire t0_00010100110, t0_00010100111;
mixer mix_t0_00010100110 (.a(t0_000101001100), .b(t0_000101001101), .y(t0_00010100110));
wire t0_000101001100, t0_000101001101;
mixer mix_t0_000101001100 (.a(t0_0001010011000), .b(t0_0001010011001), .y(t0_000101001100));
wire t0_0001010011000, t0_0001010011001;
mixer mix_t0_000101001101 (.a(t0_0001010011010), .b(t0_0001010011011), .y(t0_000101001101));
wire t0_0001010011010, t0_0001010011011;
mixer mix_t0_00010100111 (.a(t0_000101001110), .b(t0_000101001111), .y(t0_00010100111));
wire t0_000101001110, t0_000101001111;
mixer mix_t0_000101001110 (.a(t0_0001010011100), .b(t0_0001010011101), .y(t0_000101001110));
wire t0_0001010011100, t0_0001010011101;
mixer mix_t0_000101001111 (.a(t0_0001010011110), .b(t0_0001010011111), .y(t0_000101001111));
wire t0_0001010011110, t0_0001010011111;
mixer mix_t0_00010101 (.a(t0_000101010), .b(t0_000101011), .y(t0_00010101));
wire t0_000101010, t0_000101011;
mixer mix_t0_000101010 (.a(t0_0001010100), .b(t0_0001010101), .y(t0_000101010));
wire t0_0001010100, t0_0001010101;
mixer mix_t0_0001010100 (.a(t0_00010101000), .b(t0_00010101001), .y(t0_0001010100));
wire t0_00010101000, t0_00010101001;
mixer mix_t0_00010101000 (.a(t0_000101010000), .b(t0_000101010001), .y(t0_00010101000));
wire t0_000101010000, t0_000101010001;
mixer mix_t0_000101010000 (.a(t0_0001010100000), .b(t0_0001010100001), .y(t0_000101010000));
wire t0_0001010100000, t0_0001010100001;
mixer mix_t0_000101010001 (.a(t0_0001010100010), .b(t0_0001010100011), .y(t0_000101010001));
wire t0_0001010100010, t0_0001010100011;
mixer mix_t0_00010101001 (.a(t0_000101010010), .b(t0_000101010011), .y(t0_00010101001));
wire t0_000101010010, t0_000101010011;
mixer mix_t0_000101010010 (.a(t0_0001010100100), .b(t0_0001010100101), .y(t0_000101010010));
wire t0_0001010100100, t0_0001010100101;
mixer mix_t0_000101010011 (.a(t0_0001010100110), .b(t0_0001010100111), .y(t0_000101010011));
wire t0_0001010100110, t0_0001010100111;
mixer mix_t0_0001010101 (.a(t0_00010101010), .b(t0_00010101011), .y(t0_0001010101));
wire t0_00010101010, t0_00010101011;
mixer mix_t0_00010101010 (.a(t0_000101010100), .b(t0_000101010101), .y(t0_00010101010));
wire t0_000101010100, t0_000101010101;
mixer mix_t0_000101010100 (.a(t0_0001010101000), .b(t0_0001010101001), .y(t0_000101010100));
wire t0_0001010101000, t0_0001010101001;
mixer mix_t0_000101010101 (.a(t0_0001010101010), .b(t0_0001010101011), .y(t0_000101010101));
wire t0_0001010101010, t0_0001010101011;
mixer mix_t0_00010101011 (.a(t0_000101010110), .b(t0_000101010111), .y(t0_00010101011));
wire t0_000101010110, t0_000101010111;
mixer mix_t0_000101010110 (.a(t0_0001010101100), .b(t0_0001010101101), .y(t0_000101010110));
wire t0_0001010101100, t0_0001010101101;
mixer mix_t0_000101010111 (.a(t0_0001010101110), .b(t0_0001010101111), .y(t0_000101010111));
wire t0_0001010101110, t0_0001010101111;
mixer mix_t0_000101011 (.a(t0_0001010110), .b(t0_0001010111), .y(t0_000101011));
wire t0_0001010110, t0_0001010111;
mixer mix_t0_0001010110 (.a(t0_00010101100), .b(t0_00010101101), .y(t0_0001010110));
wire t0_00010101100, t0_00010101101;
mixer mix_t0_00010101100 (.a(t0_000101011000), .b(t0_000101011001), .y(t0_00010101100));
wire t0_000101011000, t0_000101011001;
mixer mix_t0_000101011000 (.a(t0_0001010110000), .b(t0_0001010110001), .y(t0_000101011000));
wire t0_0001010110000, t0_0001010110001;
mixer mix_t0_000101011001 (.a(t0_0001010110010), .b(t0_0001010110011), .y(t0_000101011001));
wire t0_0001010110010, t0_0001010110011;
mixer mix_t0_00010101101 (.a(t0_000101011010), .b(t0_000101011011), .y(t0_00010101101));
wire t0_000101011010, t0_000101011011;
mixer mix_t0_000101011010 (.a(t0_0001010110100), .b(t0_0001010110101), .y(t0_000101011010));
wire t0_0001010110100, t0_0001010110101;
mixer mix_t0_000101011011 (.a(t0_0001010110110), .b(t0_0001010110111), .y(t0_000101011011));
wire t0_0001010110110, t0_0001010110111;
mixer mix_t0_0001010111 (.a(t0_00010101110), .b(t0_00010101111), .y(t0_0001010111));
wire t0_00010101110, t0_00010101111;
mixer mix_t0_00010101110 (.a(t0_000101011100), .b(t0_000101011101), .y(t0_00010101110));
wire t0_000101011100, t0_000101011101;
mixer mix_t0_000101011100 (.a(t0_0001010111000), .b(t0_0001010111001), .y(t0_000101011100));
wire t0_0001010111000, t0_0001010111001;
mixer mix_t0_000101011101 (.a(t0_0001010111010), .b(t0_0001010111011), .y(t0_000101011101));
wire t0_0001010111010, t0_0001010111011;
mixer mix_t0_00010101111 (.a(t0_000101011110), .b(t0_000101011111), .y(t0_00010101111));
wire t0_000101011110, t0_000101011111;
mixer mix_t0_000101011110 (.a(t0_0001010111100), .b(t0_0001010111101), .y(t0_000101011110));
wire t0_0001010111100, t0_0001010111101;
mixer mix_t0_000101011111 (.a(t0_0001010111110), .b(t0_0001010111111), .y(t0_000101011111));
wire t0_0001010111110, t0_0001010111111;
mixer mix_t0_0001011 (.a(t0_00010110), .b(t0_00010111), .y(t0_0001011));
wire t0_00010110, t0_00010111;
mixer mix_t0_00010110 (.a(t0_000101100), .b(t0_000101101), .y(t0_00010110));
wire t0_000101100, t0_000101101;
mixer mix_t0_000101100 (.a(t0_0001011000), .b(t0_0001011001), .y(t0_000101100));
wire t0_0001011000, t0_0001011001;
mixer mix_t0_0001011000 (.a(t0_00010110000), .b(t0_00010110001), .y(t0_0001011000));
wire t0_00010110000, t0_00010110001;
mixer mix_t0_00010110000 (.a(t0_000101100000), .b(t0_000101100001), .y(t0_00010110000));
wire t0_000101100000, t0_000101100001;
mixer mix_t0_000101100000 (.a(t0_0001011000000), .b(t0_0001011000001), .y(t0_000101100000));
wire t0_0001011000000, t0_0001011000001;
mixer mix_t0_000101100001 (.a(t0_0001011000010), .b(t0_0001011000011), .y(t0_000101100001));
wire t0_0001011000010, t0_0001011000011;
mixer mix_t0_00010110001 (.a(t0_000101100010), .b(t0_000101100011), .y(t0_00010110001));
wire t0_000101100010, t0_000101100011;
mixer mix_t0_000101100010 (.a(t0_0001011000100), .b(t0_0001011000101), .y(t0_000101100010));
wire t0_0001011000100, t0_0001011000101;
mixer mix_t0_000101100011 (.a(t0_0001011000110), .b(t0_0001011000111), .y(t0_000101100011));
wire t0_0001011000110, t0_0001011000111;
mixer mix_t0_0001011001 (.a(t0_00010110010), .b(t0_00010110011), .y(t0_0001011001));
wire t0_00010110010, t0_00010110011;
mixer mix_t0_00010110010 (.a(t0_000101100100), .b(t0_000101100101), .y(t0_00010110010));
wire t0_000101100100, t0_000101100101;
mixer mix_t0_000101100100 (.a(t0_0001011001000), .b(t0_0001011001001), .y(t0_000101100100));
wire t0_0001011001000, t0_0001011001001;
mixer mix_t0_000101100101 (.a(t0_0001011001010), .b(t0_0001011001011), .y(t0_000101100101));
wire t0_0001011001010, t0_0001011001011;
mixer mix_t0_00010110011 (.a(t0_000101100110), .b(t0_000101100111), .y(t0_00010110011));
wire t0_000101100110, t0_000101100111;
mixer mix_t0_000101100110 (.a(t0_0001011001100), .b(t0_0001011001101), .y(t0_000101100110));
wire t0_0001011001100, t0_0001011001101;
mixer mix_t0_000101100111 (.a(t0_0001011001110), .b(t0_0001011001111), .y(t0_000101100111));
wire t0_0001011001110, t0_0001011001111;
mixer mix_t0_000101101 (.a(t0_0001011010), .b(t0_0001011011), .y(t0_000101101));
wire t0_0001011010, t0_0001011011;
mixer mix_t0_0001011010 (.a(t0_00010110100), .b(t0_00010110101), .y(t0_0001011010));
wire t0_00010110100, t0_00010110101;
mixer mix_t0_00010110100 (.a(t0_000101101000), .b(t0_000101101001), .y(t0_00010110100));
wire t0_000101101000, t0_000101101001;
mixer mix_t0_000101101000 (.a(t0_0001011010000), .b(t0_0001011010001), .y(t0_000101101000));
wire t0_0001011010000, t0_0001011010001;
mixer mix_t0_000101101001 (.a(t0_0001011010010), .b(t0_0001011010011), .y(t0_000101101001));
wire t0_0001011010010, t0_0001011010011;
mixer mix_t0_00010110101 (.a(t0_000101101010), .b(t0_000101101011), .y(t0_00010110101));
wire t0_000101101010, t0_000101101011;
mixer mix_t0_000101101010 (.a(t0_0001011010100), .b(t0_0001011010101), .y(t0_000101101010));
wire t0_0001011010100, t0_0001011010101;
mixer mix_t0_000101101011 (.a(t0_0001011010110), .b(t0_0001011010111), .y(t0_000101101011));
wire t0_0001011010110, t0_0001011010111;
mixer mix_t0_0001011011 (.a(t0_00010110110), .b(t0_00010110111), .y(t0_0001011011));
wire t0_00010110110, t0_00010110111;
mixer mix_t0_00010110110 (.a(t0_000101101100), .b(t0_000101101101), .y(t0_00010110110));
wire t0_000101101100, t0_000101101101;
mixer mix_t0_000101101100 (.a(t0_0001011011000), .b(t0_0001011011001), .y(t0_000101101100));
wire t0_0001011011000, t0_0001011011001;
mixer mix_t0_000101101101 (.a(t0_0001011011010), .b(t0_0001011011011), .y(t0_000101101101));
wire t0_0001011011010, t0_0001011011011;
mixer mix_t0_00010110111 (.a(t0_000101101110), .b(t0_000101101111), .y(t0_00010110111));
wire t0_000101101110, t0_000101101111;
mixer mix_t0_000101101110 (.a(t0_0001011011100), .b(t0_0001011011101), .y(t0_000101101110));
wire t0_0001011011100, t0_0001011011101;
mixer mix_t0_000101101111 (.a(t0_0001011011110), .b(t0_0001011011111), .y(t0_000101101111));
wire t0_0001011011110, t0_0001011011111;
mixer mix_t0_00010111 (.a(t0_000101110), .b(t0_000101111), .y(t0_00010111));
wire t0_000101110, t0_000101111;
mixer mix_t0_000101110 (.a(t0_0001011100), .b(t0_0001011101), .y(t0_000101110));
wire t0_0001011100, t0_0001011101;
mixer mix_t0_0001011100 (.a(t0_00010111000), .b(t0_00010111001), .y(t0_0001011100));
wire t0_00010111000, t0_00010111001;
mixer mix_t0_00010111000 (.a(t0_000101110000), .b(t0_000101110001), .y(t0_00010111000));
wire t0_000101110000, t0_000101110001;
mixer mix_t0_000101110000 (.a(t0_0001011100000), .b(t0_0001011100001), .y(t0_000101110000));
wire t0_0001011100000, t0_0001011100001;
mixer mix_t0_000101110001 (.a(t0_0001011100010), .b(t0_0001011100011), .y(t0_000101110001));
wire t0_0001011100010, t0_0001011100011;
mixer mix_t0_00010111001 (.a(t0_000101110010), .b(t0_000101110011), .y(t0_00010111001));
wire t0_000101110010, t0_000101110011;
mixer mix_t0_000101110010 (.a(t0_0001011100100), .b(t0_0001011100101), .y(t0_000101110010));
wire t0_0001011100100, t0_0001011100101;
mixer mix_t0_000101110011 (.a(t0_0001011100110), .b(t0_0001011100111), .y(t0_000101110011));
wire t0_0001011100110, t0_0001011100111;
mixer mix_t0_0001011101 (.a(t0_00010111010), .b(t0_00010111011), .y(t0_0001011101));
wire t0_00010111010, t0_00010111011;
mixer mix_t0_00010111010 (.a(t0_000101110100), .b(t0_000101110101), .y(t0_00010111010));
wire t0_000101110100, t0_000101110101;
mixer mix_t0_000101110100 (.a(t0_0001011101000), .b(t0_0001011101001), .y(t0_000101110100));
wire t0_0001011101000, t0_0001011101001;
mixer mix_t0_000101110101 (.a(t0_0001011101010), .b(t0_0001011101011), .y(t0_000101110101));
wire t0_0001011101010, t0_0001011101011;
mixer mix_t0_00010111011 (.a(t0_000101110110), .b(t0_000101110111), .y(t0_00010111011));
wire t0_000101110110, t0_000101110111;
mixer mix_t0_000101110110 (.a(t0_0001011101100), .b(t0_0001011101101), .y(t0_000101110110));
wire t0_0001011101100, t0_0001011101101;
mixer mix_t0_000101110111 (.a(t0_0001011101110), .b(t0_0001011101111), .y(t0_000101110111));
wire t0_0001011101110, t0_0001011101111;
mixer mix_t0_000101111 (.a(t0_0001011110), .b(t0_0001011111), .y(t0_000101111));
wire t0_0001011110, t0_0001011111;
mixer mix_t0_0001011110 (.a(t0_00010111100), .b(t0_00010111101), .y(t0_0001011110));
wire t0_00010111100, t0_00010111101;
mixer mix_t0_00010111100 (.a(t0_000101111000), .b(t0_000101111001), .y(t0_00010111100));
wire t0_000101111000, t0_000101111001;
mixer mix_t0_000101111000 (.a(t0_0001011110000), .b(t0_0001011110001), .y(t0_000101111000));
wire t0_0001011110000, t0_0001011110001;
mixer mix_t0_000101111001 (.a(t0_0001011110010), .b(t0_0001011110011), .y(t0_000101111001));
wire t0_0001011110010, t0_0001011110011;
mixer mix_t0_00010111101 (.a(t0_000101111010), .b(t0_000101111011), .y(t0_00010111101));
wire t0_000101111010, t0_000101111011;
mixer mix_t0_000101111010 (.a(t0_0001011110100), .b(t0_0001011110101), .y(t0_000101111010));
wire t0_0001011110100, t0_0001011110101;
mixer mix_t0_000101111011 (.a(t0_0001011110110), .b(t0_0001011110111), .y(t0_000101111011));
wire t0_0001011110110, t0_0001011110111;
mixer mix_t0_0001011111 (.a(t0_00010111110), .b(t0_00010111111), .y(t0_0001011111));
wire t0_00010111110, t0_00010111111;
mixer mix_t0_00010111110 (.a(t0_000101111100), .b(t0_000101111101), .y(t0_00010111110));
wire t0_000101111100, t0_000101111101;
mixer mix_t0_000101111100 (.a(t0_0001011111000), .b(t0_0001011111001), .y(t0_000101111100));
wire t0_0001011111000, t0_0001011111001;
mixer mix_t0_000101111101 (.a(t0_0001011111010), .b(t0_0001011111011), .y(t0_000101111101));
wire t0_0001011111010, t0_0001011111011;
mixer mix_t0_00010111111 (.a(t0_000101111110), .b(t0_000101111111), .y(t0_00010111111));
wire t0_000101111110, t0_000101111111;
mixer mix_t0_000101111110 (.a(t0_0001011111100), .b(t0_0001011111101), .y(t0_000101111110));
wire t0_0001011111100, t0_0001011111101;
mixer mix_t0_000101111111 (.a(t0_0001011111110), .b(t0_0001011111111), .y(t0_000101111111));
wire t0_0001011111110, t0_0001011111111;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_000110 (.a(t0_0001100), .b(t0_0001101), .y(t0_000110));
wire t0_0001100, t0_0001101;
mixer mix_t0_0001100 (.a(t0_00011000), .b(t0_00011001), .y(t0_0001100));
wire t0_00011000, t0_00011001;
mixer mix_t0_00011000 (.a(t0_000110000), .b(t0_000110001), .y(t0_00011000));
wire t0_000110000, t0_000110001;
mixer mix_t0_000110000 (.a(t0_0001100000), .b(t0_0001100001), .y(t0_000110000));
wire t0_0001100000, t0_0001100001;
mixer mix_t0_0001100000 (.a(t0_00011000000), .b(t0_00011000001), .y(t0_0001100000));
wire t0_00011000000, t0_00011000001;
mixer mix_t0_00011000000 (.a(t0_000110000000), .b(t0_000110000001), .y(t0_00011000000));
wire t0_000110000000, t0_000110000001;
mixer mix_t0_000110000000 (.a(t0_0001100000000), .b(t0_0001100000001), .y(t0_000110000000));
wire t0_0001100000000, t0_0001100000001;
mixer mix_t0_000110000001 (.a(t0_0001100000010), .b(t0_0001100000011), .y(t0_000110000001));
wire t0_0001100000010, t0_0001100000011;
mixer mix_t0_00011000001 (.a(t0_000110000010), .b(t0_000110000011), .y(t0_00011000001));
wire t0_000110000010, t0_000110000011;
mixer mix_t0_000110000010 (.a(t0_0001100000100), .b(t0_0001100000101), .y(t0_000110000010));
wire t0_0001100000100, t0_0001100000101;
mixer mix_t0_000110000011 (.a(t0_0001100000110), .b(t0_0001100000111), .y(t0_000110000011));
wire t0_0001100000110, t0_0001100000111;
mixer mix_t0_0001100001 (.a(t0_00011000010), .b(t0_00011000011), .y(t0_0001100001));
wire t0_00011000010, t0_00011000011;
mixer mix_t0_00011000010 (.a(t0_000110000100), .b(t0_000110000101), .y(t0_00011000010));
wire t0_000110000100, t0_000110000101;
mixer mix_t0_000110000100 (.a(t0_0001100001000), .b(t0_0001100001001), .y(t0_000110000100));
wire t0_0001100001000, t0_0001100001001;
mixer mix_t0_000110000101 (.a(t0_0001100001010), .b(t0_0001100001011), .y(t0_000110000101));
wire t0_0001100001010, t0_0001100001011;
mixer mix_t0_00011000011 (.a(t0_000110000110), .b(t0_000110000111), .y(t0_00011000011));
wire t0_000110000110, t0_000110000111;
mixer mix_t0_000110000110 (.a(t0_0001100001100), .b(t0_0001100001101), .y(t0_000110000110));
wire t0_0001100001100, t0_0001100001101;
mixer mix_t0_000110000111 (.a(t0_0001100001110), .b(t0_0001100001111), .y(t0_000110000111));
wire t0_0001100001110, t0_0001100001111;
mixer mix_t0_000110001 (.a(t0_0001100010), .b(t0_0001100011), .y(t0_000110001));
wire t0_0001100010, t0_0001100011;
mixer mix_t0_0001100010 (.a(t0_00011000100), .b(t0_00011000101), .y(t0_0001100010));
wire t0_00011000100, t0_00011000101;
mixer mix_t0_00011000100 (.a(t0_000110001000), .b(t0_000110001001), .y(t0_00011000100));
wire t0_000110001000, t0_000110001001;
mixer mix_t0_000110001000 (.a(t0_0001100010000), .b(t0_0001100010001), .y(t0_000110001000));
wire t0_0001100010000, t0_0001100010001;
mixer mix_t0_000110001001 (.a(t0_0001100010010), .b(t0_0001100010011), .y(t0_000110001001));
wire t0_0001100010010, t0_0001100010011;
mixer mix_t0_00011000101 (.a(t0_000110001010), .b(t0_000110001011), .y(t0_00011000101));
wire t0_000110001010, t0_000110001011;
mixer mix_t0_000110001010 (.a(t0_0001100010100), .b(t0_0001100010101), .y(t0_000110001010));
wire t0_0001100010100, t0_0001100010101;
mixer mix_t0_000110001011 (.a(t0_0001100010110), .b(t0_0001100010111), .y(t0_000110001011));
wire t0_0001100010110, t0_0001100010111;
mixer mix_t0_0001100011 (.a(t0_00011000110), .b(t0_00011000111), .y(t0_0001100011));
wire t0_00011000110, t0_00011000111;
mixer mix_t0_00011000110 (.a(t0_000110001100), .b(t0_000110001101), .y(t0_00011000110));
wire t0_000110001100, t0_000110001101;
mixer mix_t0_000110001100 (.a(t0_0001100011000), .b(t0_0001100011001), .y(t0_000110001100));
wire t0_0001100011000, t0_0001100011001;
mixer mix_t0_000110001101 (.a(t0_0001100011010), .b(t0_0001100011011), .y(t0_000110001101));
wire t0_0001100011010, t0_0001100011011;
mixer mix_t0_00011000111 (.a(t0_000110001110), .b(t0_000110001111), .y(t0_00011000111));
wire t0_000110001110, t0_000110001111;
mixer mix_t0_000110001110 (.a(t0_0001100011100), .b(t0_0001100011101), .y(t0_000110001110));
wire t0_0001100011100, t0_0001100011101;
mixer mix_t0_000110001111 (.a(t0_0001100011110), .b(t0_0001100011111), .y(t0_000110001111));
wire t0_0001100011110, t0_0001100011111;
mixer mix_t0_00011001 (.a(t0_000110010), .b(t0_000110011), .y(t0_00011001));
wire t0_000110010, t0_000110011;
mixer mix_t0_000110010 (.a(t0_0001100100), .b(t0_0001100101), .y(t0_000110010));
wire t0_0001100100, t0_0001100101;
mixer mix_t0_0001100100 (.a(t0_00011001000), .b(t0_00011001001), .y(t0_0001100100));
wire t0_00011001000, t0_00011001001;
mixer mix_t0_00011001000 (.a(t0_000110010000), .b(t0_000110010001), .y(t0_00011001000));
wire t0_000110010000, t0_000110010001;
mixer mix_t0_000110010000 (.a(t0_0001100100000), .b(t0_0001100100001), .y(t0_000110010000));
wire t0_0001100100000, t0_0001100100001;
mixer mix_t0_000110010001 (.a(t0_0001100100010), .b(t0_0001100100011), .y(t0_000110010001));
wire t0_0001100100010, t0_0001100100011;
mixer mix_t0_00011001001 (.a(t0_000110010010), .b(t0_000110010011), .y(t0_00011001001));
wire t0_000110010010, t0_000110010011;
mixer mix_t0_000110010010 (.a(t0_0001100100100), .b(t0_0001100100101), .y(t0_000110010010));
wire t0_0001100100100, t0_0001100100101;
mixer mix_t0_000110010011 (.a(t0_0001100100110), .b(t0_0001100100111), .y(t0_000110010011));
wire t0_0001100100110, t0_0001100100111;
mixer mix_t0_0001100101 (.a(t0_00011001010), .b(t0_00011001011), .y(t0_0001100101));
wire t0_00011001010, t0_00011001011;
mixer mix_t0_00011001010 (.a(t0_000110010100), .b(t0_000110010101), .y(t0_00011001010));
wire t0_000110010100, t0_000110010101;
mixer mix_t0_000110010100 (.a(t0_0001100101000), .b(t0_0001100101001), .y(t0_000110010100));
wire t0_0001100101000, t0_0001100101001;
mixer mix_t0_000110010101 (.a(t0_0001100101010), .b(t0_0001100101011), .y(t0_000110010101));
wire t0_0001100101010, t0_0001100101011;
mixer mix_t0_00011001011 (.a(t0_000110010110), .b(t0_000110010111), .y(t0_00011001011));
wire t0_000110010110, t0_000110010111;
mixer mix_t0_000110010110 (.a(t0_0001100101100), .b(t0_0001100101101), .y(t0_000110010110));
wire t0_0001100101100, t0_0001100101101;
mixer mix_t0_000110010111 (.a(t0_0001100101110), .b(t0_0001100101111), .y(t0_000110010111));
wire t0_0001100101110, t0_0001100101111;
mixer mix_t0_000110011 (.a(t0_0001100110), .b(t0_0001100111), .y(t0_000110011));
wire t0_0001100110, t0_0001100111;
mixer mix_t0_0001100110 (.a(t0_00011001100), .b(t0_00011001101), .y(t0_0001100110));
wire t0_00011001100, t0_00011001101;
mixer mix_t0_00011001100 (.a(t0_000110011000), .b(t0_000110011001), .y(t0_00011001100));
wire t0_000110011000, t0_000110011001;
mixer mix_t0_000110011000 (.a(t0_0001100110000), .b(t0_0001100110001), .y(t0_000110011000));
wire t0_0001100110000, t0_0001100110001;
mixer mix_t0_000110011001 (.a(t0_0001100110010), .b(t0_0001100110011), .y(t0_000110011001));
wire t0_0001100110010, t0_0001100110011;
mixer mix_t0_00011001101 (.a(t0_000110011010), .b(t0_000110011011), .y(t0_00011001101));
wire t0_000110011010, t0_000110011011;
mixer mix_t0_000110011010 (.a(t0_0001100110100), .b(t0_0001100110101), .y(t0_000110011010));
wire t0_0001100110100, t0_0001100110101;
mixer mix_t0_000110011011 (.a(t0_0001100110110), .b(t0_0001100110111), .y(t0_000110011011));
wire t0_0001100110110, t0_0001100110111;
mixer mix_t0_0001100111 (.a(t0_00011001110), .b(t0_00011001111), .y(t0_0001100111));
wire t0_00011001110, t0_00011001111;
mixer mix_t0_00011001110 (.a(t0_000110011100), .b(t0_000110011101), .y(t0_00011001110));
wire t0_000110011100, t0_000110011101;
mixer mix_t0_000110011100 (.a(t0_0001100111000), .b(t0_0001100111001), .y(t0_000110011100));
wire t0_0001100111000, t0_0001100111001;
mixer mix_t0_000110011101 (.a(t0_0001100111010), .b(t0_0001100111011), .y(t0_000110011101));
wire t0_0001100111010, t0_0001100111011;
mixer mix_t0_00011001111 (.a(t0_000110011110), .b(t0_000110011111), .y(t0_00011001111));
wire t0_000110011110, t0_000110011111;
mixer mix_t0_000110011110 (.a(t0_0001100111100), .b(t0_0001100111101), .y(t0_000110011110));
wire t0_0001100111100, t0_0001100111101;
mixer mix_t0_000110011111 (.a(t0_0001100111110), .b(t0_0001100111111), .y(t0_000110011111));
wire t0_0001100111110, t0_0001100111111;
mixer mix_t0_0001101 (.a(t0_00011010), .b(t0_00011011), .y(t0_0001101));
wire t0_00011010, t0_00011011;
mixer mix_t0_00011010 (.a(t0_000110100), .b(t0_000110101), .y(t0_00011010));
wire t0_000110100, t0_000110101;
mixer mix_t0_000110100 (.a(t0_0001101000), .b(t0_0001101001), .y(t0_000110100));
wire t0_0001101000, t0_0001101001;
mixer mix_t0_0001101000 (.a(t0_00011010000), .b(t0_00011010001), .y(t0_0001101000));
wire t0_00011010000, t0_00011010001;
mixer mix_t0_00011010000 (.a(t0_000110100000), .b(t0_000110100001), .y(t0_00011010000));
wire t0_000110100000, t0_000110100001;
mixer mix_t0_000110100000 (.a(t0_0001101000000), .b(t0_0001101000001), .y(t0_000110100000));
wire t0_0001101000000, t0_0001101000001;
mixer mix_t0_000110100001 (.a(t0_0001101000010), .b(t0_0001101000011), .y(t0_000110100001));
wire t0_0001101000010, t0_0001101000011;
mixer mix_t0_00011010001 (.a(t0_000110100010), .b(t0_000110100011), .y(t0_00011010001));
wire t0_000110100010, t0_000110100011;
mixer mix_t0_000110100010 (.a(t0_0001101000100), .b(t0_0001101000101), .y(t0_000110100010));
wire t0_0001101000100, t0_0001101000101;
mixer mix_t0_000110100011 (.a(t0_0001101000110), .b(t0_0001101000111), .y(t0_000110100011));
wire t0_0001101000110, t0_0001101000111;
mixer mix_t0_0001101001 (.a(t0_00011010010), .b(t0_00011010011), .y(t0_0001101001));
wire t0_00011010010, t0_00011010011;
mixer mix_t0_00011010010 (.a(t0_000110100100), .b(t0_000110100101), .y(t0_00011010010));
wire t0_000110100100, t0_000110100101;
mixer mix_t0_000110100100 (.a(t0_0001101001000), .b(t0_0001101001001), .y(t0_000110100100));
wire t0_0001101001000, t0_0001101001001;
mixer mix_t0_000110100101 (.a(t0_0001101001010), .b(t0_0001101001011), .y(t0_000110100101));
wire t0_0001101001010, t0_0001101001011;
mixer mix_t0_00011010011 (.a(t0_000110100110), .b(t0_000110100111), .y(t0_00011010011));
wire t0_000110100110, t0_000110100111;
mixer mix_t0_000110100110 (.a(t0_0001101001100), .b(t0_0001101001101), .y(t0_000110100110));
wire t0_0001101001100, t0_0001101001101;
mixer mix_t0_000110100111 (.a(t0_0001101001110), .b(t0_0001101001111), .y(t0_000110100111));
wire t0_0001101001110, t0_0001101001111;
mixer mix_t0_000110101 (.a(t0_0001101010), .b(t0_0001101011), .y(t0_000110101));
wire t0_0001101010, t0_0001101011;
mixer mix_t0_0001101010 (.a(t0_00011010100), .b(t0_00011010101), .y(t0_0001101010));
wire t0_00011010100, t0_00011010101;
mixer mix_t0_00011010100 (.a(t0_000110101000), .b(t0_000110101001), .y(t0_00011010100));
wire t0_000110101000, t0_000110101001;
mixer mix_t0_000110101000 (.a(t0_0001101010000), .b(t0_0001101010001), .y(t0_000110101000));
wire t0_0001101010000, t0_0001101010001;
mixer mix_t0_000110101001 (.a(t0_0001101010010), .b(t0_0001101010011), .y(t0_000110101001));
wire t0_0001101010010, t0_0001101010011;
mixer mix_t0_00011010101 (.a(t0_000110101010), .b(t0_000110101011), .y(t0_00011010101));
wire t0_000110101010, t0_000110101011;
mixer mix_t0_000110101010 (.a(t0_0001101010100), .b(t0_0001101010101), .y(t0_000110101010));
wire t0_0001101010100, t0_0001101010101;
mixer mix_t0_000110101011 (.a(t0_0001101010110), .b(t0_0001101010111), .y(t0_000110101011));
wire t0_0001101010110, t0_0001101010111;
mixer mix_t0_0001101011 (.a(t0_00011010110), .b(t0_00011010111), .y(t0_0001101011));
wire t0_00011010110, t0_00011010111;
mixer mix_t0_00011010110 (.a(t0_000110101100), .b(t0_000110101101), .y(t0_00011010110));
wire t0_000110101100, t0_000110101101;
mixer mix_t0_000110101100 (.a(t0_0001101011000), .b(t0_0001101011001), .y(t0_000110101100));
wire t0_0001101011000, t0_0001101011001;
mixer mix_t0_000110101101 (.a(t0_0001101011010), .b(t0_0001101011011), .y(t0_000110101101));
wire t0_0001101011010, t0_0001101011011;
mixer mix_t0_00011010111 (.a(t0_000110101110), .b(t0_000110101111), .y(t0_00011010111));
wire t0_000110101110, t0_000110101111;
mixer mix_t0_000110101110 (.a(t0_0001101011100), .b(t0_0001101011101), .y(t0_000110101110));
wire t0_0001101011100, t0_0001101011101;
mixer mix_t0_000110101111 (.a(t0_0001101011110), .b(t0_0001101011111), .y(t0_000110101111));
wire t0_0001101011110, t0_0001101011111;
mixer mix_t0_00011011 (.a(t0_000110110), .b(t0_000110111), .y(t0_00011011));
wire t0_000110110, t0_000110111;
mixer mix_t0_000110110 (.a(t0_0001101100), .b(t0_0001101101), .y(t0_000110110));
wire t0_0001101100, t0_0001101101;
mixer mix_t0_0001101100 (.a(t0_00011011000), .b(t0_00011011001), .y(t0_0001101100));
wire t0_00011011000, t0_00011011001;
mixer mix_t0_00011011000 (.a(t0_000110110000), .b(t0_000110110001), .y(t0_00011011000));
wire t0_000110110000, t0_000110110001;
mixer mix_t0_000110110000 (.a(t0_0001101100000), .b(t0_0001101100001), .y(t0_000110110000));
wire t0_0001101100000, t0_0001101100001;
mixer mix_t0_000110110001 (.a(t0_0001101100010), .b(t0_0001101100011), .y(t0_000110110001));
wire t0_0001101100010, t0_0001101100011;
mixer mix_t0_00011011001 (.a(t0_000110110010), .b(t0_000110110011), .y(t0_00011011001));
wire t0_000110110010, t0_000110110011;
mixer mix_t0_000110110010 (.a(t0_0001101100100), .b(t0_0001101100101), .y(t0_000110110010));
wire t0_0001101100100, t0_0001101100101;
mixer mix_t0_000110110011 (.a(t0_0001101100110), .b(t0_0001101100111), .y(t0_000110110011));
wire t0_0001101100110, t0_0001101100111;
mixer mix_t0_0001101101 (.a(t0_00011011010), .b(t0_00011011011), .y(t0_0001101101));
wire t0_00011011010, t0_00011011011;
mixer mix_t0_00011011010 (.a(t0_000110110100), .b(t0_000110110101), .y(t0_00011011010));
wire t0_000110110100, t0_000110110101;
mixer mix_t0_000110110100 (.a(t0_0001101101000), .b(t0_0001101101001), .y(t0_000110110100));
wire t0_0001101101000, t0_0001101101001;
mixer mix_t0_000110110101 (.a(t0_0001101101010), .b(t0_0001101101011), .y(t0_000110110101));
wire t0_0001101101010, t0_0001101101011;
mixer mix_t0_00011011011 (.a(t0_000110110110), .b(t0_000110110111), .y(t0_00011011011));
wire t0_000110110110, t0_000110110111;
mixer mix_t0_000110110110 (.a(t0_0001101101100), .b(t0_0001101101101), .y(t0_000110110110));
wire t0_0001101101100, t0_0001101101101;
mixer mix_t0_000110110111 (.a(t0_0001101101110), .b(t0_0001101101111), .y(t0_000110110111));
wire t0_0001101101110, t0_0001101101111;
mixer mix_t0_000110111 (.a(t0_0001101110), .b(t0_0001101111), .y(t0_000110111));
wire t0_0001101110, t0_0001101111;
mixer mix_t0_0001101110 (.a(t0_00011011100), .b(t0_00011011101), .y(t0_0001101110));
wire t0_00011011100, t0_00011011101;
mixer mix_t0_00011011100 (.a(t0_000110111000), .b(t0_000110111001), .y(t0_00011011100));
wire t0_000110111000, t0_000110111001;
mixer mix_t0_000110111000 (.a(t0_0001101110000), .b(t0_0001101110001), .y(t0_000110111000));
wire t0_0001101110000, t0_0001101110001;
mixer mix_t0_000110111001 (.a(t0_0001101110010), .b(t0_0001101110011), .y(t0_000110111001));
wire t0_0001101110010, t0_0001101110011;
mixer mix_t0_00011011101 (.a(t0_000110111010), .b(t0_000110111011), .y(t0_00011011101));
wire t0_000110111010, t0_000110111011;
mixer mix_t0_000110111010 (.a(t0_0001101110100), .b(t0_0001101110101), .y(t0_000110111010));
wire t0_0001101110100, t0_0001101110101;
mixer mix_t0_000110111011 (.a(t0_0001101110110), .b(t0_0001101110111), .y(t0_000110111011));
wire t0_0001101110110, t0_0001101110111;
mixer mix_t0_0001101111 (.a(t0_00011011110), .b(t0_00011011111), .y(t0_0001101111));
wire t0_00011011110, t0_00011011111;
mixer mix_t0_00011011110 (.a(t0_000110111100), .b(t0_000110111101), .y(t0_00011011110));
wire t0_000110111100, t0_000110111101;
mixer mix_t0_000110111100 (.a(t0_0001101111000), .b(t0_0001101111001), .y(t0_000110111100));
wire t0_0001101111000, t0_0001101111001;
mixer mix_t0_000110111101 (.a(t0_0001101111010), .b(t0_0001101111011), .y(t0_000110111101));
wire t0_0001101111010, t0_0001101111011;
mixer mix_t0_00011011111 (.a(t0_000110111110), .b(t0_000110111111), .y(t0_00011011111));
wire t0_000110111110, t0_000110111111;
mixer mix_t0_000110111110 (.a(t0_0001101111100), .b(t0_0001101111101), .y(t0_000110111110));
wire t0_0001101111100, t0_0001101111101;
mixer mix_t0_000110111111 (.a(t0_0001101111110), .b(t0_0001101111111), .y(t0_000110111111));
wire t0_0001101111110, t0_0001101111111;
mixer mix_t0_000111 (.a(t0_0001110), .b(t0_0001111), .y(t0_000111));
wire t0_0001110, t0_0001111;
mixer mix_t0_0001110 (.a(t0_00011100), .b(t0_00011101), .y(t0_0001110));
wire t0_00011100, t0_00011101;
mixer mix_t0_00011100 (.a(t0_000111000), .b(t0_000111001), .y(t0_00011100));
wire t0_000111000, t0_000111001;
mixer mix_t0_000111000 (.a(t0_0001110000), .b(t0_0001110001), .y(t0_000111000));
wire t0_0001110000, t0_0001110001;
mixer mix_t0_0001110000 (.a(t0_00011100000), .b(t0_00011100001), .y(t0_0001110000));
wire t0_00011100000, t0_00011100001;
mixer mix_t0_00011100000 (.a(t0_000111000000), .b(t0_000111000001), .y(t0_00011100000));
wire t0_000111000000, t0_000111000001;
mixer mix_t0_000111000000 (.a(t0_0001110000000), .b(t0_0001110000001), .y(t0_000111000000));
wire t0_0001110000000, t0_0001110000001;
mixer mix_t0_000111000001 (.a(t0_0001110000010), .b(t0_0001110000011), .y(t0_000111000001));
wire t0_0001110000010, t0_0001110000011;
mixer mix_t0_00011100001 (.a(t0_000111000010), .b(t0_000111000011), .y(t0_00011100001));
wire t0_000111000010, t0_000111000011;
mixer mix_t0_000111000010 (.a(t0_0001110000100), .b(t0_0001110000101), .y(t0_000111000010));
wire t0_0001110000100, t0_0001110000101;
mixer mix_t0_000111000011 (.a(t0_0001110000110), .b(t0_0001110000111), .y(t0_000111000011));
wire t0_0001110000110, t0_0001110000111;
mixer mix_t0_0001110001 (.a(t0_00011100010), .b(t0_00011100011), .y(t0_0001110001));
wire t0_00011100010, t0_00011100011;
mixer mix_t0_00011100010 (.a(t0_000111000100), .b(t0_000111000101), .y(t0_00011100010));
wire t0_000111000100, t0_000111000101;
mixer mix_t0_000111000100 (.a(t0_0001110001000), .b(t0_0001110001001), .y(t0_000111000100));
wire t0_0001110001000, t0_0001110001001;
mixer mix_t0_000111000101 (.a(t0_0001110001010), .b(t0_0001110001011), .y(t0_000111000101));
wire t0_0001110001010, t0_0001110001011;
mixer mix_t0_00011100011 (.a(t0_000111000110), .b(t0_000111000111), .y(t0_00011100011));
wire t0_000111000110, t0_000111000111;
mixer mix_t0_000111000110 (.a(t0_0001110001100), .b(t0_0001110001101), .y(t0_000111000110));
wire t0_0001110001100, t0_0001110001101;
mixer mix_t0_000111000111 (.a(t0_0001110001110), .b(t0_0001110001111), .y(t0_000111000111));
wire t0_0001110001110, t0_0001110001111;
mixer mix_t0_000111001 (.a(t0_0001110010), .b(t0_0001110011), .y(t0_000111001));
wire t0_0001110010, t0_0001110011;
mixer mix_t0_0001110010 (.a(t0_00011100100), .b(t0_00011100101), .y(t0_0001110010));
wire t0_00011100100, t0_00011100101;
mixer mix_t0_00011100100 (.a(t0_000111001000), .b(t0_000111001001), .y(t0_00011100100));
wire t0_000111001000, t0_000111001001;
mixer mix_t0_000111001000 (.a(t0_0001110010000), .b(t0_0001110010001), .y(t0_000111001000));
wire t0_0001110010000, t0_0001110010001;
mixer mix_t0_000111001001 (.a(t0_0001110010010), .b(t0_0001110010011), .y(t0_000111001001));
wire t0_0001110010010, t0_0001110010011;
mixer mix_t0_00011100101 (.a(t0_000111001010), .b(t0_000111001011), .y(t0_00011100101));
wire t0_000111001010, t0_000111001011;
mixer mix_t0_000111001010 (.a(t0_0001110010100), .b(t0_0001110010101), .y(t0_000111001010));
wire t0_0001110010100, t0_0001110010101;
mixer mix_t0_000111001011 (.a(t0_0001110010110), .b(t0_0001110010111), .y(t0_000111001011));
wire t0_0001110010110, t0_0001110010111;
mixer mix_t0_0001110011 (.a(t0_00011100110), .b(t0_00011100111), .y(t0_0001110011));
wire t0_00011100110, t0_00011100111;
mixer mix_t0_00011100110 (.a(t0_000111001100), .b(t0_000111001101), .y(t0_00011100110));
wire t0_000111001100, t0_000111001101;
mixer mix_t0_000111001100 (.a(t0_0001110011000), .b(t0_0001110011001), .y(t0_000111001100));
wire t0_0001110011000, t0_0001110011001;
mixer mix_t0_000111001101 (.a(t0_0001110011010), .b(t0_0001110011011), .y(t0_000111001101));
wire t0_0001110011010, t0_0001110011011;
mixer mix_t0_00011100111 (.a(t0_000111001110), .b(t0_000111001111), .y(t0_00011100111));
wire t0_000111001110, t0_000111001111;
mixer mix_t0_000111001110 (.a(t0_0001110011100), .b(t0_0001110011101), .y(t0_000111001110));
wire t0_0001110011100, t0_0001110011101;
mixer mix_t0_000111001111 (.a(t0_0001110011110), .b(t0_0001110011111), .y(t0_000111001111));
wire t0_0001110011110, t0_0001110011111;
mixer mix_t0_00011101 (.a(t0_000111010), .b(t0_000111011), .y(t0_00011101));
wire t0_000111010, t0_000111011;
mixer mix_t0_000111010 (.a(t0_0001110100), .b(t0_0001110101), .y(t0_000111010));
wire t0_0001110100, t0_0001110101;
mixer mix_t0_0001110100 (.a(t0_00011101000), .b(t0_00011101001), .y(t0_0001110100));
wire t0_00011101000, t0_00011101001;
mixer mix_t0_00011101000 (.a(t0_000111010000), .b(t0_000111010001), .y(t0_00011101000));
wire t0_000111010000, t0_000111010001;
mixer mix_t0_000111010000 (.a(t0_0001110100000), .b(t0_0001110100001), .y(t0_000111010000));
wire t0_0001110100000, t0_0001110100001;
mixer mix_t0_000111010001 (.a(t0_0001110100010), .b(t0_0001110100011), .y(t0_000111010001));
wire t0_0001110100010, t0_0001110100011;
mixer mix_t0_00011101001 (.a(t0_000111010010), .b(t0_000111010011), .y(t0_00011101001));
wire t0_000111010010, t0_000111010011;
mixer mix_t0_000111010010 (.a(t0_0001110100100), .b(t0_0001110100101), .y(t0_000111010010));
wire t0_0001110100100, t0_0001110100101;
mixer mix_t0_000111010011 (.a(t0_0001110100110), .b(t0_0001110100111), .y(t0_000111010011));
wire t0_0001110100110, t0_0001110100111;
mixer mix_t0_0001110101 (.a(t0_00011101010), .b(t0_00011101011), .y(t0_0001110101));
wire t0_00011101010, t0_00011101011;
mixer mix_t0_00011101010 (.a(t0_000111010100), .b(t0_000111010101), .y(t0_00011101010));
wire t0_000111010100, t0_000111010101;
mixer mix_t0_000111010100 (.a(t0_0001110101000), .b(t0_0001110101001), .y(t0_000111010100));
wire t0_0001110101000, t0_0001110101001;
mixer mix_t0_000111010101 (.a(t0_0001110101010), .b(t0_0001110101011), .y(t0_000111010101));
wire t0_0001110101010, t0_0001110101011;
mixer mix_t0_00011101011 (.a(t0_000111010110), .b(t0_000111010111), .y(t0_00011101011));
wire t0_000111010110, t0_000111010111;
mixer mix_t0_000111010110 (.a(t0_0001110101100), .b(t0_0001110101101), .y(t0_000111010110));
wire t0_0001110101100, t0_0001110101101;
mixer mix_t0_000111010111 (.a(t0_0001110101110), .b(t0_0001110101111), .y(t0_000111010111));
wire t0_0001110101110, t0_0001110101111;
mixer mix_t0_000111011 (.a(t0_0001110110), .b(t0_0001110111), .y(t0_000111011));
wire t0_0001110110, t0_0001110111;
mixer mix_t0_0001110110 (.a(t0_00011101100), .b(t0_00011101101), .y(t0_0001110110));
wire t0_00011101100, t0_00011101101;
mixer mix_t0_00011101100 (.a(t0_000111011000), .b(t0_000111011001), .y(t0_00011101100));
wire t0_000111011000, t0_000111011001;
mixer mix_t0_000111011000 (.a(t0_0001110110000), .b(t0_0001110110001), .y(t0_000111011000));
wire t0_0001110110000, t0_0001110110001;
mixer mix_t0_000111011001 (.a(t0_0001110110010), .b(t0_0001110110011), .y(t0_000111011001));
wire t0_0001110110010, t0_0001110110011;
mixer mix_t0_00011101101 (.a(t0_000111011010), .b(t0_000111011011), .y(t0_00011101101));
wire t0_000111011010, t0_000111011011;
mixer mix_t0_000111011010 (.a(t0_0001110110100), .b(t0_0001110110101), .y(t0_000111011010));
wire t0_0001110110100, t0_0001110110101;
mixer mix_t0_000111011011 (.a(t0_0001110110110), .b(t0_0001110110111), .y(t0_000111011011));
wire t0_0001110110110, t0_0001110110111;
mixer mix_t0_0001110111 (.a(t0_00011101110), .b(t0_00011101111), .y(t0_0001110111));
wire t0_00011101110, t0_00011101111;
mixer mix_t0_00011101110 (.a(t0_000111011100), .b(t0_000111011101), .y(t0_00011101110));
wire t0_000111011100, t0_000111011101;
mixer mix_t0_000111011100 (.a(t0_0001110111000), .b(t0_0001110111001), .y(t0_000111011100));
wire t0_0001110111000, t0_0001110111001;
mixer mix_t0_000111011101 (.a(t0_0001110111010), .b(t0_0001110111011), .y(t0_000111011101));
wire t0_0001110111010, t0_0001110111011;
mixer mix_t0_00011101111 (.a(t0_000111011110), .b(t0_000111011111), .y(t0_00011101111));
wire t0_000111011110, t0_000111011111;
mixer mix_t0_000111011110 (.a(t0_0001110111100), .b(t0_0001110111101), .y(t0_000111011110));
wire t0_0001110111100, t0_0001110111101;
mixer mix_t0_000111011111 (.a(t0_0001110111110), .b(t0_0001110111111), .y(t0_000111011111));
wire t0_0001110111110, t0_0001110111111;
mixer mix_t0_0001111 (.a(t0_00011110), .b(t0_00011111), .y(t0_0001111));
wire t0_00011110, t0_00011111;
mixer mix_t0_00011110 (.a(t0_000111100), .b(t0_000111101), .y(t0_00011110));
wire t0_000111100, t0_000111101;
mixer mix_t0_000111100 (.a(t0_0001111000), .b(t0_0001111001), .y(t0_000111100));
wire t0_0001111000, t0_0001111001;
mixer mix_t0_0001111000 (.a(t0_00011110000), .b(t0_00011110001), .y(t0_0001111000));
wire t0_00011110000, t0_00011110001;
mixer mix_t0_00011110000 (.a(t0_000111100000), .b(t0_000111100001), .y(t0_00011110000));
wire t0_000111100000, t0_000111100001;
mixer mix_t0_000111100000 (.a(t0_0001111000000), .b(t0_0001111000001), .y(t0_000111100000));
wire t0_0001111000000, t0_0001111000001;
mixer mix_t0_000111100001 (.a(t0_0001111000010), .b(t0_0001111000011), .y(t0_000111100001));
wire t0_0001111000010, t0_0001111000011;
mixer mix_t0_00011110001 (.a(t0_000111100010), .b(t0_000111100011), .y(t0_00011110001));
wire t0_000111100010, t0_000111100011;
mixer mix_t0_000111100010 (.a(t0_0001111000100), .b(t0_0001111000101), .y(t0_000111100010));
wire t0_0001111000100, t0_0001111000101;
mixer mix_t0_000111100011 (.a(t0_0001111000110), .b(t0_0001111000111), .y(t0_000111100011));
wire t0_0001111000110, t0_0001111000111;
mixer mix_t0_0001111001 (.a(t0_00011110010), .b(t0_00011110011), .y(t0_0001111001));
wire t0_00011110010, t0_00011110011;
mixer mix_t0_00011110010 (.a(t0_000111100100), .b(t0_000111100101), .y(t0_00011110010));
wire t0_000111100100, t0_000111100101;
mixer mix_t0_000111100100 (.a(t0_0001111001000), .b(t0_0001111001001), .y(t0_000111100100));
wire t0_0001111001000, t0_0001111001001;
mixer mix_t0_000111100101 (.a(t0_0001111001010), .b(t0_0001111001011), .y(t0_000111100101));
wire t0_0001111001010, t0_0001111001011;
mixer mix_t0_00011110011 (.a(t0_000111100110), .b(t0_000111100111), .y(t0_00011110011));
wire t0_000111100110, t0_000111100111;
mixer mix_t0_000111100110 (.a(t0_0001111001100), .b(t0_0001111001101), .y(t0_000111100110));
wire t0_0001111001100, t0_0001111001101;
mixer mix_t0_000111100111 (.a(t0_0001111001110), .b(t0_0001111001111), .y(t0_000111100111));
wire t0_0001111001110, t0_0001111001111;
mixer mix_t0_000111101 (.a(t0_0001111010), .b(t0_0001111011), .y(t0_000111101));
wire t0_0001111010, t0_0001111011;
mixer mix_t0_0001111010 (.a(t0_00011110100), .b(t0_00011110101), .y(t0_0001111010));
wire t0_00011110100, t0_00011110101;
mixer mix_t0_00011110100 (.a(t0_000111101000), .b(t0_000111101001), .y(t0_00011110100));
wire t0_000111101000, t0_000111101001;
mixer mix_t0_000111101000 (.a(t0_0001111010000), .b(t0_0001111010001), .y(t0_000111101000));
wire t0_0001111010000, t0_0001111010001;
mixer mix_t0_000111101001 (.a(t0_0001111010010), .b(t0_0001111010011), .y(t0_000111101001));
wire t0_0001111010010, t0_0001111010011;
mixer mix_t0_00011110101 (.a(t0_000111101010), .b(t0_000111101011), .y(t0_00011110101));
wire t0_000111101010, t0_000111101011;
mixer mix_t0_000111101010 (.a(t0_0001111010100), .b(t0_0001111010101), .y(t0_000111101010));
wire t0_0001111010100, t0_0001111010101;
mixer mix_t0_000111101011 (.a(t0_0001111010110), .b(t0_0001111010111), .y(t0_000111101011));
wire t0_0001111010110, t0_0001111010111;
mixer mix_t0_0001111011 (.a(t0_00011110110), .b(t0_00011110111), .y(t0_0001111011));
wire t0_00011110110, t0_00011110111;
mixer mix_t0_00011110110 (.a(t0_000111101100), .b(t0_000111101101), .y(t0_00011110110));
wire t0_000111101100, t0_000111101101;
mixer mix_t0_000111101100 (.a(t0_0001111011000), .b(t0_0001111011001), .y(t0_000111101100));
wire t0_0001111011000, t0_0001111011001;
mixer mix_t0_000111101101 (.a(t0_0001111011010), .b(t0_0001111011011), .y(t0_000111101101));
wire t0_0001111011010, t0_0001111011011;
mixer mix_t0_00011110111 (.a(t0_000111101110), .b(t0_000111101111), .y(t0_00011110111));
wire t0_000111101110, t0_000111101111;
mixer mix_t0_000111101110 (.a(t0_0001111011100), .b(t0_0001111011101), .y(t0_000111101110));
wire t0_0001111011100, t0_0001111011101;
mixer mix_t0_000111101111 (.a(t0_0001111011110), .b(t0_0001111011111), .y(t0_000111101111));
wire t0_0001111011110, t0_0001111011111;
mixer mix_t0_00011111 (.a(t0_000111110), .b(t0_000111111), .y(t0_00011111));
wire t0_000111110, t0_000111111;
mixer mix_t0_000111110 (.a(t0_0001111100), .b(t0_0001111101), .y(t0_000111110));
wire t0_0001111100, t0_0001111101;
mixer mix_t0_0001111100 (.a(t0_00011111000), .b(t0_00011111001), .y(t0_0001111100));
wire t0_00011111000, t0_00011111001;
mixer mix_t0_00011111000 (.a(t0_000111110000), .b(t0_000111110001), .y(t0_00011111000));
wire t0_000111110000, t0_000111110001;
mixer mix_t0_000111110000 (.a(t0_0001111100000), .b(t0_0001111100001), .y(t0_000111110000));
wire t0_0001111100000, t0_0001111100001;
mixer mix_t0_000111110001 (.a(t0_0001111100010), .b(t0_0001111100011), .y(t0_000111110001));
wire t0_0001111100010, t0_0001111100011;
mixer mix_t0_00011111001 (.a(t0_000111110010), .b(t0_000111110011), .y(t0_00011111001));
wire t0_000111110010, t0_000111110011;
mixer mix_t0_000111110010 (.a(t0_0001111100100), .b(t0_0001111100101), .y(t0_000111110010));
wire t0_0001111100100, t0_0001111100101;
mixer mix_t0_000111110011 (.a(t0_0001111100110), .b(t0_0001111100111), .y(t0_000111110011));
wire t0_0001111100110, t0_0001111100111;
mixer mix_t0_0001111101 (.a(t0_00011111010), .b(t0_00011111011), .y(t0_0001111101));
wire t0_00011111010, t0_00011111011;
mixer mix_t0_00011111010 (.a(t0_000111110100), .b(t0_000111110101), .y(t0_00011111010));
wire t0_000111110100, t0_000111110101;
mixer mix_t0_000111110100 (.a(t0_0001111101000), .b(t0_0001111101001), .y(t0_000111110100));
wire t0_0001111101000, t0_0001111101001;
mixer mix_t0_000111110101 (.a(t0_0001111101010), .b(t0_0001111101011), .y(t0_000111110101));
wire t0_0001111101010, t0_0001111101011;
mixer mix_t0_00011111011 (.a(t0_000111110110), .b(t0_000111110111), .y(t0_00011111011));
wire t0_000111110110, t0_000111110111;
mixer mix_t0_000111110110 (.a(t0_0001111101100), .b(t0_0001111101101), .y(t0_000111110110));
wire t0_0001111101100, t0_0001111101101;
mixer mix_t0_000111110111 (.a(t0_0001111101110), .b(t0_0001111101111), .y(t0_000111110111));
wire t0_0001111101110, t0_0001111101111;
mixer mix_t0_000111111 (.a(t0_0001111110), .b(t0_0001111111), .y(t0_000111111));
wire t0_0001111110, t0_0001111111;
mixer mix_t0_0001111110 (.a(t0_00011111100), .b(t0_00011111101), .y(t0_0001111110));
wire t0_00011111100, t0_00011111101;
mixer mix_t0_00011111100 (.a(t0_000111111000), .b(t0_000111111001), .y(t0_00011111100));
wire t0_000111111000, t0_000111111001;
mixer mix_t0_000111111000 (.a(t0_0001111110000), .b(t0_0001111110001), .y(t0_000111111000));
wire t0_0001111110000, t0_0001111110001;
mixer mix_t0_000111111001 (.a(t0_0001111110010), .b(t0_0001111110011), .y(t0_000111111001));
wire t0_0001111110010, t0_0001111110011;
mixer mix_t0_00011111101 (.a(t0_000111111010), .b(t0_000111111011), .y(t0_00011111101));
wire t0_000111111010, t0_000111111011;
mixer mix_t0_000111111010 (.a(t0_0001111110100), .b(t0_0001111110101), .y(t0_000111111010));
wire t0_0001111110100, t0_0001111110101;
mixer mix_t0_000111111011 (.a(t0_0001111110110), .b(t0_0001111110111), .y(t0_000111111011));
wire t0_0001111110110, t0_0001111110111;
mixer mix_t0_0001111111 (.a(t0_00011111110), .b(t0_00011111111), .y(t0_0001111111));
wire t0_00011111110, t0_00011111111;
mixer mix_t0_00011111110 (.a(t0_000111111100), .b(t0_000111111101), .y(t0_00011111110));
wire t0_000111111100, t0_000111111101;
mixer mix_t0_000111111100 (.a(t0_0001111111000), .b(t0_0001111111001), .y(t0_000111111100));
wire t0_0001111111000, t0_0001111111001;
mixer mix_t0_000111111101 (.a(t0_0001111111010), .b(t0_0001111111011), .y(t0_000111111101));
wire t0_0001111111010, t0_0001111111011;
mixer mix_t0_00011111111 (.a(t0_000111111110), .b(t0_000111111111), .y(t0_00011111111));
wire t0_000111111110, t0_000111111111;
mixer mix_t0_000111111110 (.a(t0_0001111111100), .b(t0_0001111111101), .y(t0_000111111110));
wire t0_0001111111100, t0_0001111111101;
mixer mix_t0_000111111111 (.a(t0_0001111111110), .b(t0_0001111111111), .y(t0_000111111111));
wire t0_0001111111110, t0_0001111111111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_001000 (.a(t0_0010000), .b(t0_0010001), .y(t0_001000));
wire t0_0010000, t0_0010001;
mixer mix_t0_0010000 (.a(t0_00100000), .b(t0_00100001), .y(t0_0010000));
wire t0_00100000, t0_00100001;
mixer mix_t0_00100000 (.a(t0_001000000), .b(t0_001000001), .y(t0_00100000));
wire t0_001000000, t0_001000001;
mixer mix_t0_001000000 (.a(t0_0010000000), .b(t0_0010000001), .y(t0_001000000));
wire t0_0010000000, t0_0010000001;
mixer mix_t0_0010000000 (.a(t0_00100000000), .b(t0_00100000001), .y(t0_0010000000));
wire t0_00100000000, t0_00100000001;
mixer mix_t0_00100000000 (.a(t0_001000000000), .b(t0_001000000001), .y(t0_00100000000));
wire t0_001000000000, t0_001000000001;
mixer mix_t0_001000000000 (.a(t0_0010000000000), .b(t0_0010000000001), .y(t0_001000000000));
wire t0_0010000000000, t0_0010000000001;
mixer mix_t0_001000000001 (.a(t0_0010000000010), .b(t0_0010000000011), .y(t0_001000000001));
wire t0_0010000000010, t0_0010000000011;
mixer mix_t0_00100000001 (.a(t0_001000000010), .b(t0_001000000011), .y(t0_00100000001));
wire t0_001000000010, t0_001000000011;
mixer mix_t0_001000000010 (.a(t0_0010000000100), .b(t0_0010000000101), .y(t0_001000000010));
wire t0_0010000000100, t0_0010000000101;
mixer mix_t0_001000000011 (.a(t0_0010000000110), .b(t0_0010000000111), .y(t0_001000000011));
wire t0_0010000000110, t0_0010000000111;
mixer mix_t0_0010000001 (.a(t0_00100000010), .b(t0_00100000011), .y(t0_0010000001));
wire t0_00100000010, t0_00100000011;
mixer mix_t0_00100000010 (.a(t0_001000000100), .b(t0_001000000101), .y(t0_00100000010));
wire t0_001000000100, t0_001000000101;
mixer mix_t0_001000000100 (.a(t0_0010000001000), .b(t0_0010000001001), .y(t0_001000000100));
wire t0_0010000001000, t0_0010000001001;
mixer mix_t0_001000000101 (.a(t0_0010000001010), .b(t0_0010000001011), .y(t0_001000000101));
wire t0_0010000001010, t0_0010000001011;
mixer mix_t0_00100000011 (.a(t0_001000000110), .b(t0_001000000111), .y(t0_00100000011));
wire t0_001000000110, t0_001000000111;
mixer mix_t0_001000000110 (.a(t0_0010000001100), .b(t0_0010000001101), .y(t0_001000000110));
wire t0_0010000001100, t0_0010000001101;
mixer mix_t0_001000000111 (.a(t0_0010000001110), .b(t0_0010000001111), .y(t0_001000000111));
wire t0_0010000001110, t0_0010000001111;
mixer mix_t0_001000001 (.a(t0_0010000010), .b(t0_0010000011), .y(t0_001000001));
wire t0_0010000010, t0_0010000011;
mixer mix_t0_0010000010 (.a(t0_00100000100), .b(t0_00100000101), .y(t0_0010000010));
wire t0_00100000100, t0_00100000101;
mixer mix_t0_00100000100 (.a(t0_001000001000), .b(t0_001000001001), .y(t0_00100000100));
wire t0_001000001000, t0_001000001001;
mixer mix_t0_001000001000 (.a(t0_0010000010000), .b(t0_0010000010001), .y(t0_001000001000));
wire t0_0010000010000, t0_0010000010001;
mixer mix_t0_001000001001 (.a(t0_0010000010010), .b(t0_0010000010011), .y(t0_001000001001));
wire t0_0010000010010, t0_0010000010011;
mixer mix_t0_00100000101 (.a(t0_001000001010), .b(t0_001000001011), .y(t0_00100000101));
wire t0_001000001010, t0_001000001011;
mixer mix_t0_001000001010 (.a(t0_0010000010100), .b(t0_0010000010101), .y(t0_001000001010));
wire t0_0010000010100, t0_0010000010101;
mixer mix_t0_001000001011 (.a(t0_0010000010110), .b(t0_0010000010111), .y(t0_001000001011));
wire t0_0010000010110, t0_0010000010111;
mixer mix_t0_0010000011 (.a(t0_00100000110), .b(t0_00100000111), .y(t0_0010000011));
wire t0_00100000110, t0_00100000111;
mixer mix_t0_00100000110 (.a(t0_001000001100), .b(t0_001000001101), .y(t0_00100000110));
wire t0_001000001100, t0_001000001101;
mixer mix_t0_001000001100 (.a(t0_0010000011000), .b(t0_0010000011001), .y(t0_001000001100));
wire t0_0010000011000, t0_0010000011001;
mixer mix_t0_001000001101 (.a(t0_0010000011010), .b(t0_0010000011011), .y(t0_001000001101));
wire t0_0010000011010, t0_0010000011011;
mixer mix_t0_00100000111 (.a(t0_001000001110), .b(t0_001000001111), .y(t0_00100000111));
wire t0_001000001110, t0_001000001111;
mixer mix_t0_001000001110 (.a(t0_0010000011100), .b(t0_0010000011101), .y(t0_001000001110));
wire t0_0010000011100, t0_0010000011101;
mixer mix_t0_001000001111 (.a(t0_0010000011110), .b(t0_0010000011111), .y(t0_001000001111));
wire t0_0010000011110, t0_0010000011111;
mixer mix_t0_00100001 (.a(t0_001000010), .b(t0_001000011), .y(t0_00100001));
wire t0_001000010, t0_001000011;
mixer mix_t0_001000010 (.a(t0_0010000100), .b(t0_0010000101), .y(t0_001000010));
wire t0_0010000100, t0_0010000101;
mixer mix_t0_0010000100 (.a(t0_00100001000), .b(t0_00100001001), .y(t0_0010000100));
wire t0_00100001000, t0_00100001001;
mixer mix_t0_00100001000 (.a(t0_001000010000), .b(t0_001000010001), .y(t0_00100001000));
wire t0_001000010000, t0_001000010001;
mixer mix_t0_001000010000 (.a(t0_0010000100000), .b(t0_0010000100001), .y(t0_001000010000));
wire t0_0010000100000, t0_0010000100001;
mixer mix_t0_001000010001 (.a(t0_0010000100010), .b(t0_0010000100011), .y(t0_001000010001));
wire t0_0010000100010, t0_0010000100011;
mixer mix_t0_00100001001 (.a(t0_001000010010), .b(t0_001000010011), .y(t0_00100001001));
wire t0_001000010010, t0_001000010011;
mixer mix_t0_001000010010 (.a(t0_0010000100100), .b(t0_0010000100101), .y(t0_001000010010));
wire t0_0010000100100, t0_0010000100101;
mixer mix_t0_001000010011 (.a(t0_0010000100110), .b(t0_0010000100111), .y(t0_001000010011));
wire t0_0010000100110, t0_0010000100111;
mixer mix_t0_0010000101 (.a(t0_00100001010), .b(t0_00100001011), .y(t0_0010000101));
wire t0_00100001010, t0_00100001011;
mixer mix_t0_00100001010 (.a(t0_001000010100), .b(t0_001000010101), .y(t0_00100001010));
wire t0_001000010100, t0_001000010101;
mixer mix_t0_001000010100 (.a(t0_0010000101000), .b(t0_0010000101001), .y(t0_001000010100));
wire t0_0010000101000, t0_0010000101001;
mixer mix_t0_001000010101 (.a(t0_0010000101010), .b(t0_0010000101011), .y(t0_001000010101));
wire t0_0010000101010, t0_0010000101011;
mixer mix_t0_00100001011 (.a(t0_001000010110), .b(t0_001000010111), .y(t0_00100001011));
wire t0_001000010110, t0_001000010111;
mixer mix_t0_001000010110 (.a(t0_0010000101100), .b(t0_0010000101101), .y(t0_001000010110));
wire t0_0010000101100, t0_0010000101101;
mixer mix_t0_001000010111 (.a(t0_0010000101110), .b(t0_0010000101111), .y(t0_001000010111));
wire t0_0010000101110, t0_0010000101111;
mixer mix_t0_001000011 (.a(t0_0010000110), .b(t0_0010000111), .y(t0_001000011));
wire t0_0010000110, t0_0010000111;
mixer mix_t0_0010000110 (.a(t0_00100001100), .b(t0_00100001101), .y(t0_0010000110));
wire t0_00100001100, t0_00100001101;
mixer mix_t0_00100001100 (.a(t0_001000011000), .b(t0_001000011001), .y(t0_00100001100));
wire t0_001000011000, t0_001000011001;
mixer mix_t0_001000011000 (.a(t0_0010000110000), .b(t0_0010000110001), .y(t0_001000011000));
wire t0_0010000110000, t0_0010000110001;
mixer mix_t0_001000011001 (.a(t0_0010000110010), .b(t0_0010000110011), .y(t0_001000011001));
wire t0_0010000110010, t0_0010000110011;
mixer mix_t0_00100001101 (.a(t0_001000011010), .b(t0_001000011011), .y(t0_00100001101));
wire t0_001000011010, t0_001000011011;
mixer mix_t0_001000011010 (.a(t0_0010000110100), .b(t0_0010000110101), .y(t0_001000011010));
wire t0_0010000110100, t0_0010000110101;
mixer mix_t0_001000011011 (.a(t0_0010000110110), .b(t0_0010000110111), .y(t0_001000011011));
wire t0_0010000110110, t0_0010000110111;
mixer mix_t0_0010000111 (.a(t0_00100001110), .b(t0_00100001111), .y(t0_0010000111));
wire t0_00100001110, t0_00100001111;
mixer mix_t0_00100001110 (.a(t0_001000011100), .b(t0_001000011101), .y(t0_00100001110));
wire t0_001000011100, t0_001000011101;
mixer mix_t0_001000011100 (.a(t0_0010000111000), .b(t0_0010000111001), .y(t0_001000011100));
wire t0_0010000111000, t0_0010000111001;
mixer mix_t0_001000011101 (.a(t0_0010000111010), .b(t0_0010000111011), .y(t0_001000011101));
wire t0_0010000111010, t0_0010000111011;
mixer mix_t0_00100001111 (.a(t0_001000011110), .b(t0_001000011111), .y(t0_00100001111));
wire t0_001000011110, t0_001000011111;
mixer mix_t0_001000011110 (.a(t0_0010000111100), .b(t0_0010000111101), .y(t0_001000011110));
wire t0_0010000111100, t0_0010000111101;
mixer mix_t0_001000011111 (.a(t0_0010000111110), .b(t0_0010000111111), .y(t0_001000011111));
wire t0_0010000111110, t0_0010000111111;
mixer mix_t0_0010001 (.a(t0_00100010), .b(t0_00100011), .y(t0_0010001));
wire t0_00100010, t0_00100011;
mixer mix_t0_00100010 (.a(t0_001000100), .b(t0_001000101), .y(t0_00100010));
wire t0_001000100, t0_001000101;
mixer mix_t0_001000100 (.a(t0_0010001000), .b(t0_0010001001), .y(t0_001000100));
wire t0_0010001000, t0_0010001001;
mixer mix_t0_0010001000 (.a(t0_00100010000), .b(t0_00100010001), .y(t0_0010001000));
wire t0_00100010000, t0_00100010001;
mixer mix_t0_00100010000 (.a(t0_001000100000), .b(t0_001000100001), .y(t0_00100010000));
wire t0_001000100000, t0_001000100001;
mixer mix_t0_001000100000 (.a(t0_0010001000000), .b(t0_0010001000001), .y(t0_001000100000));
wire t0_0010001000000, t0_0010001000001;
mixer mix_t0_001000100001 (.a(t0_0010001000010), .b(t0_0010001000011), .y(t0_001000100001));
wire t0_0010001000010, t0_0010001000011;
mixer mix_t0_00100010001 (.a(t0_001000100010), .b(t0_001000100011), .y(t0_00100010001));
wire t0_001000100010, t0_001000100011;
mixer mix_t0_001000100010 (.a(t0_0010001000100), .b(t0_0010001000101), .y(t0_001000100010));
wire t0_0010001000100, t0_0010001000101;
mixer mix_t0_001000100011 (.a(t0_0010001000110), .b(t0_0010001000111), .y(t0_001000100011));
wire t0_0010001000110, t0_0010001000111;
mixer mix_t0_0010001001 (.a(t0_00100010010), .b(t0_00100010011), .y(t0_0010001001));
wire t0_00100010010, t0_00100010011;
mixer mix_t0_00100010010 (.a(t0_001000100100), .b(t0_001000100101), .y(t0_00100010010));
wire t0_001000100100, t0_001000100101;
mixer mix_t0_001000100100 (.a(t0_0010001001000), .b(t0_0010001001001), .y(t0_001000100100));
wire t0_0010001001000, t0_0010001001001;
mixer mix_t0_001000100101 (.a(t0_0010001001010), .b(t0_0010001001011), .y(t0_001000100101));
wire t0_0010001001010, t0_0010001001011;
mixer mix_t0_00100010011 (.a(t0_001000100110), .b(t0_001000100111), .y(t0_00100010011));
wire t0_001000100110, t0_001000100111;
mixer mix_t0_001000100110 (.a(t0_0010001001100), .b(t0_0010001001101), .y(t0_001000100110));
wire t0_0010001001100, t0_0010001001101;
mixer mix_t0_001000100111 (.a(t0_0010001001110), .b(t0_0010001001111), .y(t0_001000100111));
wire t0_0010001001110, t0_0010001001111;
mixer mix_t0_001000101 (.a(t0_0010001010), .b(t0_0010001011), .y(t0_001000101));
wire t0_0010001010, t0_0010001011;
mixer mix_t0_0010001010 (.a(t0_00100010100), .b(t0_00100010101), .y(t0_0010001010));
wire t0_00100010100, t0_00100010101;
mixer mix_t0_00100010100 (.a(t0_001000101000), .b(t0_001000101001), .y(t0_00100010100));
wire t0_001000101000, t0_001000101001;
mixer mix_t0_001000101000 (.a(t0_0010001010000), .b(t0_0010001010001), .y(t0_001000101000));
wire t0_0010001010000, t0_0010001010001;
mixer mix_t0_001000101001 (.a(t0_0010001010010), .b(t0_0010001010011), .y(t0_001000101001));
wire t0_0010001010010, t0_0010001010011;
mixer mix_t0_00100010101 (.a(t0_001000101010), .b(t0_001000101011), .y(t0_00100010101));
wire t0_001000101010, t0_001000101011;
mixer mix_t0_001000101010 (.a(t0_0010001010100), .b(t0_0010001010101), .y(t0_001000101010));
wire t0_0010001010100, t0_0010001010101;
mixer mix_t0_001000101011 (.a(t0_0010001010110), .b(t0_0010001010111), .y(t0_001000101011));
wire t0_0010001010110, t0_0010001010111;
mixer mix_t0_0010001011 (.a(t0_00100010110), .b(t0_00100010111), .y(t0_0010001011));
wire t0_00100010110, t0_00100010111;
mixer mix_t0_00100010110 (.a(t0_001000101100), .b(t0_001000101101), .y(t0_00100010110));
wire t0_001000101100, t0_001000101101;
mixer mix_t0_001000101100 (.a(t0_0010001011000), .b(t0_0010001011001), .y(t0_001000101100));
wire t0_0010001011000, t0_0010001011001;
mixer mix_t0_001000101101 (.a(t0_0010001011010), .b(t0_0010001011011), .y(t0_001000101101));
wire t0_0010001011010, t0_0010001011011;
mixer mix_t0_00100010111 (.a(t0_001000101110), .b(t0_001000101111), .y(t0_00100010111));
wire t0_001000101110, t0_001000101111;
mixer mix_t0_001000101110 (.a(t0_0010001011100), .b(t0_0010001011101), .y(t0_001000101110));
wire t0_0010001011100, t0_0010001011101;
mixer mix_t0_001000101111 (.a(t0_0010001011110), .b(t0_0010001011111), .y(t0_001000101111));
wire t0_0010001011110, t0_0010001011111;
mixer mix_t0_00100011 (.a(t0_001000110), .b(t0_001000111), .y(t0_00100011));
wire t0_001000110, t0_001000111;
mixer mix_t0_001000110 (.a(t0_0010001100), .b(t0_0010001101), .y(t0_001000110));
wire t0_0010001100, t0_0010001101;
mixer mix_t0_0010001100 (.a(t0_00100011000), .b(t0_00100011001), .y(t0_0010001100));
wire t0_00100011000, t0_00100011001;
mixer mix_t0_00100011000 (.a(t0_001000110000), .b(t0_001000110001), .y(t0_00100011000));
wire t0_001000110000, t0_001000110001;
mixer mix_t0_001000110000 (.a(t0_0010001100000), .b(t0_0010001100001), .y(t0_001000110000));
wire t0_0010001100000, t0_0010001100001;
mixer mix_t0_001000110001 (.a(t0_0010001100010), .b(t0_0010001100011), .y(t0_001000110001));
wire t0_0010001100010, t0_0010001100011;
mixer mix_t0_00100011001 (.a(t0_001000110010), .b(t0_001000110011), .y(t0_00100011001));
wire t0_001000110010, t0_001000110011;
mixer mix_t0_001000110010 (.a(t0_0010001100100), .b(t0_0010001100101), .y(t0_001000110010));
wire t0_0010001100100, t0_0010001100101;
mixer mix_t0_001000110011 (.a(t0_0010001100110), .b(t0_0010001100111), .y(t0_001000110011));
wire t0_0010001100110, t0_0010001100111;
mixer mix_t0_0010001101 (.a(t0_00100011010), .b(t0_00100011011), .y(t0_0010001101));
wire t0_00100011010, t0_00100011011;
mixer mix_t0_00100011010 (.a(t0_001000110100), .b(t0_001000110101), .y(t0_00100011010));
wire t0_001000110100, t0_001000110101;
mixer mix_t0_001000110100 (.a(t0_0010001101000), .b(t0_0010001101001), .y(t0_001000110100));
wire t0_0010001101000, t0_0010001101001;
mixer mix_t0_001000110101 (.a(t0_0010001101010), .b(t0_0010001101011), .y(t0_001000110101));
wire t0_0010001101010, t0_0010001101011;
mixer mix_t0_00100011011 (.a(t0_001000110110), .b(t0_001000110111), .y(t0_00100011011));
wire t0_001000110110, t0_001000110111;
mixer mix_t0_001000110110 (.a(t0_0010001101100), .b(t0_0010001101101), .y(t0_001000110110));
wire t0_0010001101100, t0_0010001101101;
mixer mix_t0_001000110111 (.a(t0_0010001101110), .b(t0_0010001101111), .y(t0_001000110111));
wire t0_0010001101110, t0_0010001101111;
mixer mix_t0_001000111 (.a(t0_0010001110), .b(t0_0010001111), .y(t0_001000111));
wire t0_0010001110, t0_0010001111;
mixer mix_t0_0010001110 (.a(t0_00100011100), .b(t0_00100011101), .y(t0_0010001110));
wire t0_00100011100, t0_00100011101;
mixer mix_t0_00100011100 (.a(t0_001000111000), .b(t0_001000111001), .y(t0_00100011100));
wire t0_001000111000, t0_001000111001;
mixer mix_t0_001000111000 (.a(t0_0010001110000), .b(t0_0010001110001), .y(t0_001000111000));
wire t0_0010001110000, t0_0010001110001;
mixer mix_t0_001000111001 (.a(t0_0010001110010), .b(t0_0010001110011), .y(t0_001000111001));
wire t0_0010001110010, t0_0010001110011;
mixer mix_t0_00100011101 (.a(t0_001000111010), .b(t0_001000111011), .y(t0_00100011101));
wire t0_001000111010, t0_001000111011;
mixer mix_t0_001000111010 (.a(t0_0010001110100), .b(t0_0010001110101), .y(t0_001000111010));
wire t0_0010001110100, t0_0010001110101;
mixer mix_t0_001000111011 (.a(t0_0010001110110), .b(t0_0010001110111), .y(t0_001000111011));
wire t0_0010001110110, t0_0010001110111;
mixer mix_t0_0010001111 (.a(t0_00100011110), .b(t0_00100011111), .y(t0_0010001111));
wire t0_00100011110, t0_00100011111;
mixer mix_t0_00100011110 (.a(t0_001000111100), .b(t0_001000111101), .y(t0_00100011110));
wire t0_001000111100, t0_001000111101;
mixer mix_t0_001000111100 (.a(t0_0010001111000), .b(t0_0010001111001), .y(t0_001000111100));
wire t0_0010001111000, t0_0010001111001;
mixer mix_t0_001000111101 (.a(t0_0010001111010), .b(t0_0010001111011), .y(t0_001000111101));
wire t0_0010001111010, t0_0010001111011;
mixer mix_t0_00100011111 (.a(t0_001000111110), .b(t0_001000111111), .y(t0_00100011111));
wire t0_001000111110, t0_001000111111;
mixer mix_t0_001000111110 (.a(t0_0010001111100), .b(t0_0010001111101), .y(t0_001000111110));
wire t0_0010001111100, t0_0010001111101;
mixer mix_t0_001000111111 (.a(t0_0010001111110), .b(t0_0010001111111), .y(t0_001000111111));
wire t0_0010001111110, t0_0010001111111;
mixer mix_t0_001001 (.a(t0_0010010), .b(t0_0010011), .y(t0_001001));
wire t0_0010010, t0_0010011;
mixer mix_t0_0010010 (.a(t0_00100100), .b(t0_00100101), .y(t0_0010010));
wire t0_00100100, t0_00100101;
mixer mix_t0_00100100 (.a(t0_001001000), .b(t0_001001001), .y(t0_00100100));
wire t0_001001000, t0_001001001;
mixer mix_t0_001001000 (.a(t0_0010010000), .b(t0_0010010001), .y(t0_001001000));
wire t0_0010010000, t0_0010010001;
mixer mix_t0_0010010000 (.a(t0_00100100000), .b(t0_00100100001), .y(t0_0010010000));
wire t0_00100100000, t0_00100100001;
mixer mix_t0_00100100000 (.a(t0_001001000000), .b(t0_001001000001), .y(t0_00100100000));
wire t0_001001000000, t0_001001000001;
mixer mix_t0_001001000000 (.a(t0_0010010000000), .b(t0_0010010000001), .y(t0_001001000000));
wire t0_0010010000000, t0_0010010000001;
mixer mix_t0_001001000001 (.a(t0_0010010000010), .b(t0_0010010000011), .y(t0_001001000001));
wire t0_0010010000010, t0_0010010000011;
mixer mix_t0_00100100001 (.a(t0_001001000010), .b(t0_001001000011), .y(t0_00100100001));
wire t0_001001000010, t0_001001000011;
mixer mix_t0_001001000010 (.a(t0_0010010000100), .b(t0_0010010000101), .y(t0_001001000010));
wire t0_0010010000100, t0_0010010000101;
mixer mix_t0_001001000011 (.a(t0_0010010000110), .b(t0_0010010000111), .y(t0_001001000011));
wire t0_0010010000110, t0_0010010000111;
mixer mix_t0_0010010001 (.a(t0_00100100010), .b(t0_00100100011), .y(t0_0010010001));
wire t0_00100100010, t0_00100100011;
mixer mix_t0_00100100010 (.a(t0_001001000100), .b(t0_001001000101), .y(t0_00100100010));
wire t0_001001000100, t0_001001000101;
mixer mix_t0_001001000100 (.a(t0_0010010001000), .b(t0_0010010001001), .y(t0_001001000100));
wire t0_0010010001000, t0_0010010001001;
mixer mix_t0_001001000101 (.a(t0_0010010001010), .b(t0_0010010001011), .y(t0_001001000101));
wire t0_0010010001010, t0_0010010001011;
mixer mix_t0_00100100011 (.a(t0_001001000110), .b(t0_001001000111), .y(t0_00100100011));
wire t0_001001000110, t0_001001000111;
mixer mix_t0_001001000110 (.a(t0_0010010001100), .b(t0_0010010001101), .y(t0_001001000110));
wire t0_0010010001100, t0_0010010001101;
mixer mix_t0_001001000111 (.a(t0_0010010001110), .b(t0_0010010001111), .y(t0_001001000111));
wire t0_0010010001110, t0_0010010001111;
mixer mix_t0_001001001 (.a(t0_0010010010), .b(t0_0010010011), .y(t0_001001001));
wire t0_0010010010, t0_0010010011;
mixer mix_t0_0010010010 (.a(t0_00100100100), .b(t0_00100100101), .y(t0_0010010010));
wire t0_00100100100, t0_00100100101;
mixer mix_t0_00100100100 (.a(t0_001001001000), .b(t0_001001001001), .y(t0_00100100100));
wire t0_001001001000, t0_001001001001;
mixer mix_t0_001001001000 (.a(t0_0010010010000), .b(t0_0010010010001), .y(t0_001001001000));
wire t0_0010010010000, t0_0010010010001;
mixer mix_t0_001001001001 (.a(t0_0010010010010), .b(t0_0010010010011), .y(t0_001001001001));
wire t0_0010010010010, t0_0010010010011;
mixer mix_t0_00100100101 (.a(t0_001001001010), .b(t0_001001001011), .y(t0_00100100101));
wire t0_001001001010, t0_001001001011;
mixer mix_t0_001001001010 (.a(t0_0010010010100), .b(t0_0010010010101), .y(t0_001001001010));
wire t0_0010010010100, t0_0010010010101;
mixer mix_t0_001001001011 (.a(t0_0010010010110), .b(t0_0010010010111), .y(t0_001001001011));
wire t0_0010010010110, t0_0010010010111;
mixer mix_t0_0010010011 (.a(t0_00100100110), .b(t0_00100100111), .y(t0_0010010011));
wire t0_00100100110, t0_00100100111;
mixer mix_t0_00100100110 (.a(t0_001001001100), .b(t0_001001001101), .y(t0_00100100110));
wire t0_001001001100, t0_001001001101;
mixer mix_t0_001001001100 (.a(t0_0010010011000), .b(t0_0010010011001), .y(t0_001001001100));
wire t0_0010010011000, t0_0010010011001;
mixer mix_t0_001001001101 (.a(t0_0010010011010), .b(t0_0010010011011), .y(t0_001001001101));
wire t0_0010010011010, t0_0010010011011;
mixer mix_t0_00100100111 (.a(t0_001001001110), .b(t0_001001001111), .y(t0_00100100111));
wire t0_001001001110, t0_001001001111;
mixer mix_t0_001001001110 (.a(t0_0010010011100), .b(t0_0010010011101), .y(t0_001001001110));
wire t0_0010010011100, t0_0010010011101;
mixer mix_t0_001001001111 (.a(t0_0010010011110), .b(t0_0010010011111), .y(t0_001001001111));
wire t0_0010010011110, t0_0010010011111;
mixer mix_t0_00100101 (.a(t0_001001010), .b(t0_001001011), .y(t0_00100101));
wire t0_001001010, t0_001001011;
mixer mix_t0_001001010 (.a(t0_0010010100), .b(t0_0010010101), .y(t0_001001010));
wire t0_0010010100, t0_0010010101;
mixer mix_t0_0010010100 (.a(t0_00100101000), .b(t0_00100101001), .y(t0_0010010100));
wire t0_00100101000, t0_00100101001;
mixer mix_t0_00100101000 (.a(t0_001001010000), .b(t0_001001010001), .y(t0_00100101000));
wire t0_001001010000, t0_001001010001;
mixer mix_t0_001001010000 (.a(t0_0010010100000), .b(t0_0010010100001), .y(t0_001001010000));
wire t0_0010010100000, t0_0010010100001;
mixer mix_t0_001001010001 (.a(t0_0010010100010), .b(t0_0010010100011), .y(t0_001001010001));
wire t0_0010010100010, t0_0010010100011;
mixer mix_t0_00100101001 (.a(t0_001001010010), .b(t0_001001010011), .y(t0_00100101001));
wire t0_001001010010, t0_001001010011;
mixer mix_t0_001001010010 (.a(t0_0010010100100), .b(t0_0010010100101), .y(t0_001001010010));
wire t0_0010010100100, t0_0010010100101;
mixer mix_t0_001001010011 (.a(t0_0010010100110), .b(t0_0010010100111), .y(t0_001001010011));
wire t0_0010010100110, t0_0010010100111;
mixer mix_t0_0010010101 (.a(t0_00100101010), .b(t0_00100101011), .y(t0_0010010101));
wire t0_00100101010, t0_00100101011;
mixer mix_t0_00100101010 (.a(t0_001001010100), .b(t0_001001010101), .y(t0_00100101010));
wire t0_001001010100, t0_001001010101;
mixer mix_t0_001001010100 (.a(t0_0010010101000), .b(t0_0010010101001), .y(t0_001001010100));
wire t0_0010010101000, t0_0010010101001;
mixer mix_t0_001001010101 (.a(t0_0010010101010), .b(t0_0010010101011), .y(t0_001001010101));
wire t0_0010010101010, t0_0010010101011;
mixer mix_t0_00100101011 (.a(t0_001001010110), .b(t0_001001010111), .y(t0_00100101011));
wire t0_001001010110, t0_001001010111;
mixer mix_t0_001001010110 (.a(t0_0010010101100), .b(t0_0010010101101), .y(t0_001001010110));
wire t0_0010010101100, t0_0010010101101;
mixer mix_t0_001001010111 (.a(t0_0010010101110), .b(t0_0010010101111), .y(t0_001001010111));
wire t0_0010010101110, t0_0010010101111;
mixer mix_t0_001001011 (.a(t0_0010010110), .b(t0_0010010111), .y(t0_001001011));
wire t0_0010010110, t0_0010010111;
mixer mix_t0_0010010110 (.a(t0_00100101100), .b(t0_00100101101), .y(t0_0010010110));
wire t0_00100101100, t0_00100101101;
mixer mix_t0_00100101100 (.a(t0_001001011000), .b(t0_001001011001), .y(t0_00100101100));
wire t0_001001011000, t0_001001011001;
mixer mix_t0_001001011000 (.a(t0_0010010110000), .b(t0_0010010110001), .y(t0_001001011000));
wire t0_0010010110000, t0_0010010110001;
mixer mix_t0_001001011001 (.a(t0_0010010110010), .b(t0_0010010110011), .y(t0_001001011001));
wire t0_0010010110010, t0_0010010110011;
mixer mix_t0_00100101101 (.a(t0_001001011010), .b(t0_001001011011), .y(t0_00100101101));
wire t0_001001011010, t0_001001011011;
mixer mix_t0_001001011010 (.a(t0_0010010110100), .b(t0_0010010110101), .y(t0_001001011010));
wire t0_0010010110100, t0_0010010110101;
mixer mix_t0_001001011011 (.a(t0_0010010110110), .b(t0_0010010110111), .y(t0_001001011011));
wire t0_0010010110110, t0_0010010110111;
mixer mix_t0_0010010111 (.a(t0_00100101110), .b(t0_00100101111), .y(t0_0010010111));
wire t0_00100101110, t0_00100101111;
mixer mix_t0_00100101110 (.a(t0_001001011100), .b(t0_001001011101), .y(t0_00100101110));
wire t0_001001011100, t0_001001011101;
mixer mix_t0_001001011100 (.a(t0_0010010111000), .b(t0_0010010111001), .y(t0_001001011100));
wire t0_0010010111000, t0_0010010111001;
mixer mix_t0_001001011101 (.a(t0_0010010111010), .b(t0_0010010111011), .y(t0_001001011101));
wire t0_0010010111010, t0_0010010111011;
mixer mix_t0_00100101111 (.a(t0_001001011110), .b(t0_001001011111), .y(t0_00100101111));
wire t0_001001011110, t0_001001011111;
mixer mix_t0_001001011110 (.a(t0_0010010111100), .b(t0_0010010111101), .y(t0_001001011110));
wire t0_0010010111100, t0_0010010111101;
mixer mix_t0_001001011111 (.a(t0_0010010111110), .b(t0_0010010111111), .y(t0_001001011111));
wire t0_0010010111110, t0_0010010111111;
mixer mix_t0_0010011 (.a(t0_00100110), .b(t0_00100111), .y(t0_0010011));
wire t0_00100110, t0_00100111;
mixer mix_t0_00100110 (.a(t0_001001100), .b(t0_001001101), .y(t0_00100110));
wire t0_001001100, t0_001001101;
mixer mix_t0_001001100 (.a(t0_0010011000), .b(t0_0010011001), .y(t0_001001100));
wire t0_0010011000, t0_0010011001;
mixer mix_t0_0010011000 (.a(t0_00100110000), .b(t0_00100110001), .y(t0_0010011000));
wire t0_00100110000, t0_00100110001;
mixer mix_t0_00100110000 (.a(t0_001001100000), .b(t0_001001100001), .y(t0_00100110000));
wire t0_001001100000, t0_001001100001;
mixer mix_t0_001001100000 (.a(t0_0010011000000), .b(t0_0010011000001), .y(t0_001001100000));
wire t0_0010011000000, t0_0010011000001;
mixer mix_t0_001001100001 (.a(t0_0010011000010), .b(t0_0010011000011), .y(t0_001001100001));
wire t0_0010011000010, t0_0010011000011;
mixer mix_t0_00100110001 (.a(t0_001001100010), .b(t0_001001100011), .y(t0_00100110001));
wire t0_001001100010, t0_001001100011;
mixer mix_t0_001001100010 (.a(t0_0010011000100), .b(t0_0010011000101), .y(t0_001001100010));
wire t0_0010011000100, t0_0010011000101;
mixer mix_t0_001001100011 (.a(t0_0010011000110), .b(t0_0010011000111), .y(t0_001001100011));
wire t0_0010011000110, t0_0010011000111;
mixer mix_t0_0010011001 (.a(t0_00100110010), .b(t0_00100110011), .y(t0_0010011001));
wire t0_00100110010, t0_00100110011;
mixer mix_t0_00100110010 (.a(t0_001001100100), .b(t0_001001100101), .y(t0_00100110010));
wire t0_001001100100, t0_001001100101;
mixer mix_t0_001001100100 (.a(t0_0010011001000), .b(t0_0010011001001), .y(t0_001001100100));
wire t0_0010011001000, t0_0010011001001;
mixer mix_t0_001001100101 (.a(t0_0010011001010), .b(t0_0010011001011), .y(t0_001001100101));
wire t0_0010011001010, t0_0010011001011;
mixer mix_t0_00100110011 (.a(t0_001001100110), .b(t0_001001100111), .y(t0_00100110011));
wire t0_001001100110, t0_001001100111;
mixer mix_t0_001001100110 (.a(t0_0010011001100), .b(t0_0010011001101), .y(t0_001001100110));
wire t0_0010011001100, t0_0010011001101;
mixer mix_t0_001001100111 (.a(t0_0010011001110), .b(t0_0010011001111), .y(t0_001001100111));
wire t0_0010011001110, t0_0010011001111;
mixer mix_t0_001001101 (.a(t0_0010011010), .b(t0_0010011011), .y(t0_001001101));
wire t0_0010011010, t0_0010011011;
mixer mix_t0_0010011010 (.a(t0_00100110100), .b(t0_00100110101), .y(t0_0010011010));
wire t0_00100110100, t0_00100110101;
mixer mix_t0_00100110100 (.a(t0_001001101000), .b(t0_001001101001), .y(t0_00100110100));
wire t0_001001101000, t0_001001101001;
mixer mix_t0_001001101000 (.a(t0_0010011010000), .b(t0_0010011010001), .y(t0_001001101000));
wire t0_0010011010000, t0_0010011010001;
mixer mix_t0_001001101001 (.a(t0_0010011010010), .b(t0_0010011010011), .y(t0_001001101001));
wire t0_0010011010010, t0_0010011010011;
mixer mix_t0_00100110101 (.a(t0_001001101010), .b(t0_001001101011), .y(t0_00100110101));
wire t0_001001101010, t0_001001101011;
mixer mix_t0_001001101010 (.a(t0_0010011010100), .b(t0_0010011010101), .y(t0_001001101010));
wire t0_0010011010100, t0_0010011010101;
mixer mix_t0_001001101011 (.a(t0_0010011010110), .b(t0_0010011010111), .y(t0_001001101011));
wire t0_0010011010110, t0_0010011010111;
mixer mix_t0_0010011011 (.a(t0_00100110110), .b(t0_00100110111), .y(t0_0010011011));
wire t0_00100110110, t0_00100110111;
mixer mix_t0_00100110110 (.a(t0_001001101100), .b(t0_001001101101), .y(t0_00100110110));
wire t0_001001101100, t0_001001101101;
mixer mix_t0_001001101100 (.a(t0_0010011011000), .b(t0_0010011011001), .y(t0_001001101100));
wire t0_0010011011000, t0_0010011011001;
mixer mix_t0_001001101101 (.a(t0_0010011011010), .b(t0_0010011011011), .y(t0_001001101101));
wire t0_0010011011010, t0_0010011011011;
mixer mix_t0_00100110111 (.a(t0_001001101110), .b(t0_001001101111), .y(t0_00100110111));
wire t0_001001101110, t0_001001101111;
mixer mix_t0_001001101110 (.a(t0_0010011011100), .b(t0_0010011011101), .y(t0_001001101110));
wire t0_0010011011100, t0_0010011011101;
mixer mix_t0_001001101111 (.a(t0_0010011011110), .b(t0_0010011011111), .y(t0_001001101111));
wire t0_0010011011110, t0_0010011011111;
mixer mix_t0_00100111 (.a(t0_001001110), .b(t0_001001111), .y(t0_00100111));
wire t0_001001110, t0_001001111;
mixer mix_t0_001001110 (.a(t0_0010011100), .b(t0_0010011101), .y(t0_001001110));
wire t0_0010011100, t0_0010011101;
mixer mix_t0_0010011100 (.a(t0_00100111000), .b(t0_00100111001), .y(t0_0010011100));
wire t0_00100111000, t0_00100111001;
mixer mix_t0_00100111000 (.a(t0_001001110000), .b(t0_001001110001), .y(t0_00100111000));
wire t0_001001110000, t0_001001110001;
mixer mix_t0_001001110000 (.a(t0_0010011100000), .b(t0_0010011100001), .y(t0_001001110000));
wire t0_0010011100000, t0_0010011100001;
mixer mix_t0_001001110001 (.a(t0_0010011100010), .b(t0_0010011100011), .y(t0_001001110001));
wire t0_0010011100010, t0_0010011100011;
mixer mix_t0_00100111001 (.a(t0_001001110010), .b(t0_001001110011), .y(t0_00100111001));
wire t0_001001110010, t0_001001110011;
mixer mix_t0_001001110010 (.a(t0_0010011100100), .b(t0_0010011100101), .y(t0_001001110010));
wire t0_0010011100100, t0_0010011100101;
mixer mix_t0_001001110011 (.a(t0_0010011100110), .b(t0_0010011100111), .y(t0_001001110011));
wire t0_0010011100110, t0_0010011100111;
mixer mix_t0_0010011101 (.a(t0_00100111010), .b(t0_00100111011), .y(t0_0010011101));
wire t0_00100111010, t0_00100111011;
mixer mix_t0_00100111010 (.a(t0_001001110100), .b(t0_001001110101), .y(t0_00100111010));
wire t0_001001110100, t0_001001110101;
mixer mix_t0_001001110100 (.a(t0_0010011101000), .b(t0_0010011101001), .y(t0_001001110100));
wire t0_0010011101000, t0_0010011101001;
mixer mix_t0_001001110101 (.a(t0_0010011101010), .b(t0_0010011101011), .y(t0_001001110101));
wire t0_0010011101010, t0_0010011101011;
mixer mix_t0_00100111011 (.a(t0_001001110110), .b(t0_001001110111), .y(t0_00100111011));
wire t0_001001110110, t0_001001110111;
mixer mix_t0_001001110110 (.a(t0_0010011101100), .b(t0_0010011101101), .y(t0_001001110110));
wire t0_0010011101100, t0_0010011101101;
mixer mix_t0_001001110111 (.a(t0_0010011101110), .b(t0_0010011101111), .y(t0_001001110111));
wire t0_0010011101110, t0_0010011101111;
mixer mix_t0_001001111 (.a(t0_0010011110), .b(t0_0010011111), .y(t0_001001111));
wire t0_0010011110, t0_0010011111;
mixer mix_t0_0010011110 (.a(t0_00100111100), .b(t0_00100111101), .y(t0_0010011110));
wire t0_00100111100, t0_00100111101;
mixer mix_t0_00100111100 (.a(t0_001001111000), .b(t0_001001111001), .y(t0_00100111100));
wire t0_001001111000, t0_001001111001;
mixer mix_t0_001001111000 (.a(t0_0010011110000), .b(t0_0010011110001), .y(t0_001001111000));
wire t0_0010011110000, t0_0010011110001;
mixer mix_t0_001001111001 (.a(t0_0010011110010), .b(t0_0010011110011), .y(t0_001001111001));
wire t0_0010011110010, t0_0010011110011;
mixer mix_t0_00100111101 (.a(t0_001001111010), .b(t0_001001111011), .y(t0_00100111101));
wire t0_001001111010, t0_001001111011;
mixer mix_t0_001001111010 (.a(t0_0010011110100), .b(t0_0010011110101), .y(t0_001001111010));
wire t0_0010011110100, t0_0010011110101;
mixer mix_t0_001001111011 (.a(t0_0010011110110), .b(t0_0010011110111), .y(t0_001001111011));
wire t0_0010011110110, t0_0010011110111;
mixer mix_t0_0010011111 (.a(t0_00100111110), .b(t0_00100111111), .y(t0_0010011111));
wire t0_00100111110, t0_00100111111;
mixer mix_t0_00100111110 (.a(t0_001001111100), .b(t0_001001111101), .y(t0_00100111110));
wire t0_001001111100, t0_001001111101;
mixer mix_t0_001001111100 (.a(t0_0010011111000), .b(t0_0010011111001), .y(t0_001001111100));
wire t0_0010011111000, t0_0010011111001;
mixer mix_t0_001001111101 (.a(t0_0010011111010), .b(t0_0010011111011), .y(t0_001001111101));
wire t0_0010011111010, t0_0010011111011;
mixer mix_t0_00100111111 (.a(t0_001001111110), .b(t0_001001111111), .y(t0_00100111111));
wire t0_001001111110, t0_001001111111;
mixer mix_t0_001001111110 (.a(t0_0010011111100), .b(t0_0010011111101), .y(t0_001001111110));
wire t0_0010011111100, t0_0010011111101;
mixer mix_t0_001001111111 (.a(t0_0010011111110), .b(t0_0010011111111), .y(t0_001001111111));
wire t0_0010011111110, t0_0010011111111;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_001010 (.a(t0_0010100), .b(t0_0010101), .y(t0_001010));
wire t0_0010100, t0_0010101;
mixer mix_t0_0010100 (.a(t0_00101000), .b(t0_00101001), .y(t0_0010100));
wire t0_00101000, t0_00101001;
mixer mix_t0_00101000 (.a(t0_001010000), .b(t0_001010001), .y(t0_00101000));
wire t0_001010000, t0_001010001;
mixer mix_t0_001010000 (.a(t0_0010100000), .b(t0_0010100001), .y(t0_001010000));
wire t0_0010100000, t0_0010100001;
mixer mix_t0_0010100000 (.a(t0_00101000000), .b(t0_00101000001), .y(t0_0010100000));
wire t0_00101000000, t0_00101000001;
mixer mix_t0_00101000000 (.a(t0_001010000000), .b(t0_001010000001), .y(t0_00101000000));
wire t0_001010000000, t0_001010000001;
mixer mix_t0_001010000000 (.a(t0_0010100000000), .b(t0_0010100000001), .y(t0_001010000000));
wire t0_0010100000000, t0_0010100000001;
mixer mix_t0_001010000001 (.a(t0_0010100000010), .b(t0_0010100000011), .y(t0_001010000001));
wire t0_0010100000010, t0_0010100000011;
mixer mix_t0_00101000001 (.a(t0_001010000010), .b(t0_001010000011), .y(t0_00101000001));
wire t0_001010000010, t0_001010000011;
mixer mix_t0_001010000010 (.a(t0_0010100000100), .b(t0_0010100000101), .y(t0_001010000010));
wire t0_0010100000100, t0_0010100000101;
mixer mix_t0_001010000011 (.a(t0_0010100000110), .b(t0_0010100000111), .y(t0_001010000011));
wire t0_0010100000110, t0_0010100000111;
mixer mix_t0_0010100001 (.a(t0_00101000010), .b(t0_00101000011), .y(t0_0010100001));
wire t0_00101000010, t0_00101000011;
mixer mix_t0_00101000010 (.a(t0_001010000100), .b(t0_001010000101), .y(t0_00101000010));
wire t0_001010000100, t0_001010000101;
mixer mix_t0_001010000100 (.a(t0_0010100001000), .b(t0_0010100001001), .y(t0_001010000100));
wire t0_0010100001000, t0_0010100001001;
mixer mix_t0_001010000101 (.a(t0_0010100001010), .b(t0_0010100001011), .y(t0_001010000101));
wire t0_0010100001010, t0_0010100001011;
mixer mix_t0_00101000011 (.a(t0_001010000110), .b(t0_001010000111), .y(t0_00101000011));
wire t0_001010000110, t0_001010000111;
mixer mix_t0_001010000110 (.a(t0_0010100001100), .b(t0_0010100001101), .y(t0_001010000110));
wire t0_0010100001100, t0_0010100001101;
mixer mix_t0_001010000111 (.a(t0_0010100001110), .b(t0_0010100001111), .y(t0_001010000111));
wire t0_0010100001110, t0_0010100001111;
mixer mix_t0_001010001 (.a(t0_0010100010), .b(t0_0010100011), .y(t0_001010001));
wire t0_0010100010, t0_0010100011;
mixer mix_t0_0010100010 (.a(t0_00101000100), .b(t0_00101000101), .y(t0_0010100010));
wire t0_00101000100, t0_00101000101;
mixer mix_t0_00101000100 (.a(t0_001010001000), .b(t0_001010001001), .y(t0_00101000100));
wire t0_001010001000, t0_001010001001;
mixer mix_t0_001010001000 (.a(t0_0010100010000), .b(t0_0010100010001), .y(t0_001010001000));
wire t0_0010100010000, t0_0010100010001;
mixer mix_t0_001010001001 (.a(t0_0010100010010), .b(t0_0010100010011), .y(t0_001010001001));
wire t0_0010100010010, t0_0010100010011;
mixer mix_t0_00101000101 (.a(t0_001010001010), .b(t0_001010001011), .y(t0_00101000101));
wire t0_001010001010, t0_001010001011;
mixer mix_t0_001010001010 (.a(t0_0010100010100), .b(t0_0010100010101), .y(t0_001010001010));
wire t0_0010100010100, t0_0010100010101;
mixer mix_t0_001010001011 (.a(t0_0010100010110), .b(t0_0010100010111), .y(t0_001010001011));
wire t0_0010100010110, t0_0010100010111;
mixer mix_t0_0010100011 (.a(t0_00101000110), .b(t0_00101000111), .y(t0_0010100011));
wire t0_00101000110, t0_00101000111;
mixer mix_t0_00101000110 (.a(t0_001010001100), .b(t0_001010001101), .y(t0_00101000110));
wire t0_001010001100, t0_001010001101;
mixer mix_t0_001010001100 (.a(t0_0010100011000), .b(t0_0010100011001), .y(t0_001010001100));
wire t0_0010100011000, t0_0010100011001;
mixer mix_t0_001010001101 (.a(t0_0010100011010), .b(t0_0010100011011), .y(t0_001010001101));
wire t0_0010100011010, t0_0010100011011;
mixer mix_t0_00101000111 (.a(t0_001010001110), .b(t0_001010001111), .y(t0_00101000111));
wire t0_001010001110, t0_001010001111;
mixer mix_t0_001010001110 (.a(t0_0010100011100), .b(t0_0010100011101), .y(t0_001010001110));
wire t0_0010100011100, t0_0010100011101;
mixer mix_t0_001010001111 (.a(t0_0010100011110), .b(t0_0010100011111), .y(t0_001010001111));
wire t0_0010100011110, t0_0010100011111;
mixer mix_t0_00101001 (.a(t0_001010010), .b(t0_001010011), .y(t0_00101001));
wire t0_001010010, t0_001010011;
mixer mix_t0_001010010 (.a(t0_0010100100), .b(t0_0010100101), .y(t0_001010010));
wire t0_0010100100, t0_0010100101;
mixer mix_t0_0010100100 (.a(t0_00101001000), .b(t0_00101001001), .y(t0_0010100100));
wire t0_00101001000, t0_00101001001;
mixer mix_t0_00101001000 (.a(t0_001010010000), .b(t0_001010010001), .y(t0_00101001000));
wire t0_001010010000, t0_001010010001;
mixer mix_t0_001010010000 (.a(t0_0010100100000), .b(t0_0010100100001), .y(t0_001010010000));
wire t0_0010100100000, t0_0010100100001;
mixer mix_t0_001010010001 (.a(t0_0010100100010), .b(t0_0010100100011), .y(t0_001010010001));
wire t0_0010100100010, t0_0010100100011;
mixer mix_t0_00101001001 (.a(t0_001010010010), .b(t0_001010010011), .y(t0_00101001001));
wire t0_001010010010, t0_001010010011;
mixer mix_t0_001010010010 (.a(t0_0010100100100), .b(t0_0010100100101), .y(t0_001010010010));
wire t0_0010100100100, t0_0010100100101;
mixer mix_t0_001010010011 (.a(t0_0010100100110), .b(t0_0010100100111), .y(t0_001010010011));
wire t0_0010100100110, t0_0010100100111;
mixer mix_t0_0010100101 (.a(t0_00101001010), .b(t0_00101001011), .y(t0_0010100101));
wire t0_00101001010, t0_00101001011;
mixer mix_t0_00101001010 (.a(t0_001010010100), .b(t0_001010010101), .y(t0_00101001010));
wire t0_001010010100, t0_001010010101;
mixer mix_t0_001010010100 (.a(t0_0010100101000), .b(t0_0010100101001), .y(t0_001010010100));
wire t0_0010100101000, t0_0010100101001;
mixer mix_t0_001010010101 (.a(t0_0010100101010), .b(t0_0010100101011), .y(t0_001010010101));
wire t0_0010100101010, t0_0010100101011;
mixer mix_t0_00101001011 (.a(t0_001010010110), .b(t0_001010010111), .y(t0_00101001011));
wire t0_001010010110, t0_001010010111;
mixer mix_t0_001010010110 (.a(t0_0010100101100), .b(t0_0010100101101), .y(t0_001010010110));
wire t0_0010100101100, t0_0010100101101;
mixer mix_t0_001010010111 (.a(t0_0010100101110), .b(t0_0010100101111), .y(t0_001010010111));
wire t0_0010100101110, t0_0010100101111;
mixer mix_t0_001010011 (.a(t0_0010100110), .b(t0_0010100111), .y(t0_001010011));
wire t0_0010100110, t0_0010100111;
mixer mix_t0_0010100110 (.a(t0_00101001100), .b(t0_00101001101), .y(t0_0010100110));
wire t0_00101001100, t0_00101001101;
mixer mix_t0_00101001100 (.a(t0_001010011000), .b(t0_001010011001), .y(t0_00101001100));
wire t0_001010011000, t0_001010011001;
mixer mix_t0_001010011000 (.a(t0_0010100110000), .b(t0_0010100110001), .y(t0_001010011000));
wire t0_0010100110000, t0_0010100110001;
mixer mix_t0_001010011001 (.a(t0_0010100110010), .b(t0_0010100110011), .y(t0_001010011001));
wire t0_0010100110010, t0_0010100110011;
mixer mix_t0_00101001101 (.a(t0_001010011010), .b(t0_001010011011), .y(t0_00101001101));
wire t0_001010011010, t0_001010011011;
mixer mix_t0_001010011010 (.a(t0_0010100110100), .b(t0_0010100110101), .y(t0_001010011010));
wire t0_0010100110100, t0_0010100110101;
mixer mix_t0_001010011011 (.a(t0_0010100110110), .b(t0_0010100110111), .y(t0_001010011011));
wire t0_0010100110110, t0_0010100110111;
mixer mix_t0_0010100111 (.a(t0_00101001110), .b(t0_00101001111), .y(t0_0010100111));
wire t0_00101001110, t0_00101001111;
mixer mix_t0_00101001110 (.a(t0_001010011100), .b(t0_001010011101), .y(t0_00101001110));
wire t0_001010011100, t0_001010011101;
mixer mix_t0_001010011100 (.a(t0_0010100111000), .b(t0_0010100111001), .y(t0_001010011100));
wire t0_0010100111000, t0_0010100111001;
mixer mix_t0_001010011101 (.a(t0_0010100111010), .b(t0_0010100111011), .y(t0_001010011101));
wire t0_0010100111010, t0_0010100111011;
mixer mix_t0_00101001111 (.a(t0_001010011110), .b(t0_001010011111), .y(t0_00101001111));
wire t0_001010011110, t0_001010011111;
mixer mix_t0_001010011110 (.a(t0_0010100111100), .b(t0_0010100111101), .y(t0_001010011110));
wire t0_0010100111100, t0_0010100111101;
mixer mix_t0_001010011111 (.a(t0_0010100111110), .b(t0_0010100111111), .y(t0_001010011111));
wire t0_0010100111110, t0_0010100111111;
mixer mix_t0_0010101 (.a(t0_00101010), .b(t0_00101011), .y(t0_0010101));
wire t0_00101010, t0_00101011;
mixer mix_t0_00101010 (.a(t0_001010100), .b(t0_001010101), .y(t0_00101010));
wire t0_001010100, t0_001010101;
mixer mix_t0_001010100 (.a(t0_0010101000), .b(t0_0010101001), .y(t0_001010100));
wire t0_0010101000, t0_0010101001;
mixer mix_t0_0010101000 (.a(t0_00101010000), .b(t0_00101010001), .y(t0_0010101000));
wire t0_00101010000, t0_00101010001;
mixer mix_t0_00101010000 (.a(t0_001010100000), .b(t0_001010100001), .y(t0_00101010000));
wire t0_001010100000, t0_001010100001;
mixer mix_t0_001010100000 (.a(t0_0010101000000), .b(t0_0010101000001), .y(t0_001010100000));
wire t0_0010101000000, t0_0010101000001;
mixer mix_t0_001010100001 (.a(t0_0010101000010), .b(t0_0010101000011), .y(t0_001010100001));
wire t0_0010101000010, t0_0010101000011;
mixer mix_t0_00101010001 (.a(t0_001010100010), .b(t0_001010100011), .y(t0_00101010001));
wire t0_001010100010, t0_001010100011;
mixer mix_t0_001010100010 (.a(t0_0010101000100), .b(t0_0010101000101), .y(t0_001010100010));
wire t0_0010101000100, t0_0010101000101;
mixer mix_t0_001010100011 (.a(t0_0010101000110), .b(t0_0010101000111), .y(t0_001010100011));
wire t0_0010101000110, t0_0010101000111;
mixer mix_t0_0010101001 (.a(t0_00101010010), .b(t0_00101010011), .y(t0_0010101001));
wire t0_00101010010, t0_00101010011;
mixer mix_t0_00101010010 (.a(t0_001010100100), .b(t0_001010100101), .y(t0_00101010010));
wire t0_001010100100, t0_001010100101;
mixer mix_t0_001010100100 (.a(t0_0010101001000), .b(t0_0010101001001), .y(t0_001010100100));
wire t0_0010101001000, t0_0010101001001;
mixer mix_t0_001010100101 (.a(t0_0010101001010), .b(t0_0010101001011), .y(t0_001010100101));
wire t0_0010101001010, t0_0010101001011;
mixer mix_t0_00101010011 (.a(t0_001010100110), .b(t0_001010100111), .y(t0_00101010011));
wire t0_001010100110, t0_001010100111;
mixer mix_t0_001010100110 (.a(t0_0010101001100), .b(t0_0010101001101), .y(t0_001010100110));
wire t0_0010101001100, t0_0010101001101;
mixer mix_t0_001010100111 (.a(t0_0010101001110), .b(t0_0010101001111), .y(t0_001010100111));
wire t0_0010101001110, t0_0010101001111;
mixer mix_t0_001010101 (.a(t0_0010101010), .b(t0_0010101011), .y(t0_001010101));
wire t0_0010101010, t0_0010101011;
mixer mix_t0_0010101010 (.a(t0_00101010100), .b(t0_00101010101), .y(t0_0010101010));
wire t0_00101010100, t0_00101010101;
mixer mix_t0_00101010100 (.a(t0_001010101000), .b(t0_001010101001), .y(t0_00101010100));
wire t0_001010101000, t0_001010101001;
mixer mix_t0_001010101000 (.a(t0_0010101010000), .b(t0_0010101010001), .y(t0_001010101000));
wire t0_0010101010000, t0_0010101010001;
mixer mix_t0_001010101001 (.a(t0_0010101010010), .b(t0_0010101010011), .y(t0_001010101001));
wire t0_0010101010010, t0_0010101010011;
mixer mix_t0_00101010101 (.a(t0_001010101010), .b(t0_001010101011), .y(t0_00101010101));
wire t0_001010101010, t0_001010101011;
mixer mix_t0_001010101010 (.a(t0_0010101010100), .b(t0_0010101010101), .y(t0_001010101010));
wire t0_0010101010100, t0_0010101010101;
mixer mix_t0_001010101011 (.a(t0_0010101010110), .b(t0_0010101010111), .y(t0_001010101011));
wire t0_0010101010110, t0_0010101010111;
mixer mix_t0_0010101011 (.a(t0_00101010110), .b(t0_00101010111), .y(t0_0010101011));
wire t0_00101010110, t0_00101010111;
mixer mix_t0_00101010110 (.a(t0_001010101100), .b(t0_001010101101), .y(t0_00101010110));
wire t0_001010101100, t0_001010101101;
mixer mix_t0_001010101100 (.a(t0_0010101011000), .b(t0_0010101011001), .y(t0_001010101100));
wire t0_0010101011000, t0_0010101011001;
mixer mix_t0_001010101101 (.a(t0_0010101011010), .b(t0_0010101011011), .y(t0_001010101101));
wire t0_0010101011010, t0_0010101011011;
mixer mix_t0_00101010111 (.a(t0_001010101110), .b(t0_001010101111), .y(t0_00101010111));
wire t0_001010101110, t0_001010101111;
mixer mix_t0_001010101110 (.a(t0_0010101011100), .b(t0_0010101011101), .y(t0_001010101110));
wire t0_0010101011100, t0_0010101011101;
mixer mix_t0_001010101111 (.a(t0_0010101011110), .b(t0_0010101011111), .y(t0_001010101111));
wire t0_0010101011110, t0_0010101011111;
mixer mix_t0_00101011 (.a(t0_001010110), .b(t0_001010111), .y(t0_00101011));
wire t0_001010110, t0_001010111;
mixer mix_t0_001010110 (.a(t0_0010101100), .b(t0_0010101101), .y(t0_001010110));
wire t0_0010101100, t0_0010101101;
mixer mix_t0_0010101100 (.a(t0_00101011000), .b(t0_00101011001), .y(t0_0010101100));
wire t0_00101011000, t0_00101011001;
mixer mix_t0_00101011000 (.a(t0_001010110000), .b(t0_001010110001), .y(t0_00101011000));
wire t0_001010110000, t0_001010110001;
mixer mix_t0_001010110000 (.a(t0_0010101100000), .b(t0_0010101100001), .y(t0_001010110000));
wire t0_0010101100000, t0_0010101100001;
mixer mix_t0_001010110001 (.a(t0_0010101100010), .b(t0_0010101100011), .y(t0_001010110001));
wire t0_0010101100010, t0_0010101100011;
mixer mix_t0_00101011001 (.a(t0_001010110010), .b(t0_001010110011), .y(t0_00101011001));
wire t0_001010110010, t0_001010110011;
mixer mix_t0_001010110010 (.a(t0_0010101100100), .b(t0_0010101100101), .y(t0_001010110010));
wire t0_0010101100100, t0_0010101100101;
mixer mix_t0_001010110011 (.a(t0_0010101100110), .b(t0_0010101100111), .y(t0_001010110011));
wire t0_0010101100110, t0_0010101100111;
mixer mix_t0_0010101101 (.a(t0_00101011010), .b(t0_00101011011), .y(t0_0010101101));
wire t0_00101011010, t0_00101011011;
mixer mix_t0_00101011010 (.a(t0_001010110100), .b(t0_001010110101), .y(t0_00101011010));
wire t0_001010110100, t0_001010110101;
mixer mix_t0_001010110100 (.a(t0_0010101101000), .b(t0_0010101101001), .y(t0_001010110100));
wire t0_0010101101000, t0_0010101101001;
mixer mix_t0_001010110101 (.a(t0_0010101101010), .b(t0_0010101101011), .y(t0_001010110101));
wire t0_0010101101010, t0_0010101101011;
mixer mix_t0_00101011011 (.a(t0_001010110110), .b(t0_001010110111), .y(t0_00101011011));
wire t0_001010110110, t0_001010110111;
mixer mix_t0_001010110110 (.a(t0_0010101101100), .b(t0_0010101101101), .y(t0_001010110110));
wire t0_0010101101100, t0_0010101101101;
mixer mix_t0_001010110111 (.a(t0_0010101101110), .b(t0_0010101101111), .y(t0_001010110111));
wire t0_0010101101110, t0_0010101101111;
mixer mix_t0_001010111 (.a(t0_0010101110), .b(t0_0010101111), .y(t0_001010111));
wire t0_0010101110, t0_0010101111;
mixer mix_t0_0010101110 (.a(t0_00101011100), .b(t0_00101011101), .y(t0_0010101110));
wire t0_00101011100, t0_00101011101;
mixer mix_t0_00101011100 (.a(t0_001010111000), .b(t0_001010111001), .y(t0_00101011100));
wire t0_001010111000, t0_001010111001;
mixer mix_t0_001010111000 (.a(t0_0010101110000), .b(t0_0010101110001), .y(t0_001010111000));
wire t0_0010101110000, t0_0010101110001;
mixer mix_t0_001010111001 (.a(t0_0010101110010), .b(t0_0010101110011), .y(t0_001010111001));
wire t0_0010101110010, t0_0010101110011;
mixer mix_t0_00101011101 (.a(t0_001010111010), .b(t0_001010111011), .y(t0_00101011101));
wire t0_001010111010, t0_001010111011;
mixer mix_t0_001010111010 (.a(t0_0010101110100), .b(t0_0010101110101), .y(t0_001010111010));
wire t0_0010101110100, t0_0010101110101;
mixer mix_t0_001010111011 (.a(t0_0010101110110), .b(t0_0010101110111), .y(t0_001010111011));
wire t0_0010101110110, t0_0010101110111;
mixer mix_t0_0010101111 (.a(t0_00101011110), .b(t0_00101011111), .y(t0_0010101111));
wire t0_00101011110, t0_00101011111;
mixer mix_t0_00101011110 (.a(t0_001010111100), .b(t0_001010111101), .y(t0_00101011110));
wire t0_001010111100, t0_001010111101;
mixer mix_t0_001010111100 (.a(t0_0010101111000), .b(t0_0010101111001), .y(t0_001010111100));
wire t0_0010101111000, t0_0010101111001;
mixer mix_t0_001010111101 (.a(t0_0010101111010), .b(t0_0010101111011), .y(t0_001010111101));
wire t0_0010101111010, t0_0010101111011;
mixer mix_t0_00101011111 (.a(t0_001010111110), .b(t0_001010111111), .y(t0_00101011111));
wire t0_001010111110, t0_001010111111;
mixer mix_t0_001010111110 (.a(t0_0010101111100), .b(t0_0010101111101), .y(t0_001010111110));
wire t0_0010101111100, t0_0010101111101;
mixer mix_t0_001010111111 (.a(t0_0010101111110), .b(t0_0010101111111), .y(t0_001010111111));
wire t0_0010101111110, t0_0010101111111;
mixer mix_t0_001011 (.a(t0_0010110), .b(t0_0010111), .y(t0_001011));
wire t0_0010110, t0_0010111;
mixer mix_t0_0010110 (.a(t0_00101100), .b(t0_00101101), .y(t0_0010110));
wire t0_00101100, t0_00101101;
mixer mix_t0_00101100 (.a(t0_001011000), .b(t0_001011001), .y(t0_00101100));
wire t0_001011000, t0_001011001;
mixer mix_t0_001011000 (.a(t0_0010110000), .b(t0_0010110001), .y(t0_001011000));
wire t0_0010110000, t0_0010110001;
mixer mix_t0_0010110000 (.a(t0_00101100000), .b(t0_00101100001), .y(t0_0010110000));
wire t0_00101100000, t0_00101100001;
mixer mix_t0_00101100000 (.a(t0_001011000000), .b(t0_001011000001), .y(t0_00101100000));
wire t0_001011000000, t0_001011000001;
mixer mix_t0_001011000000 (.a(t0_0010110000000), .b(t0_0010110000001), .y(t0_001011000000));
wire t0_0010110000000, t0_0010110000001;
mixer mix_t0_001011000001 (.a(t0_0010110000010), .b(t0_0010110000011), .y(t0_001011000001));
wire t0_0010110000010, t0_0010110000011;
mixer mix_t0_00101100001 (.a(t0_001011000010), .b(t0_001011000011), .y(t0_00101100001));
wire t0_001011000010, t0_001011000011;
mixer mix_t0_001011000010 (.a(t0_0010110000100), .b(t0_0010110000101), .y(t0_001011000010));
wire t0_0010110000100, t0_0010110000101;
mixer mix_t0_001011000011 (.a(t0_0010110000110), .b(t0_0010110000111), .y(t0_001011000011));
wire t0_0010110000110, t0_0010110000111;
mixer mix_t0_0010110001 (.a(t0_00101100010), .b(t0_00101100011), .y(t0_0010110001));
wire t0_00101100010, t0_00101100011;
mixer mix_t0_00101100010 (.a(t0_001011000100), .b(t0_001011000101), .y(t0_00101100010));
wire t0_001011000100, t0_001011000101;
mixer mix_t0_001011000100 (.a(t0_0010110001000), .b(t0_0010110001001), .y(t0_001011000100));
wire t0_0010110001000, t0_0010110001001;
mixer mix_t0_001011000101 (.a(t0_0010110001010), .b(t0_0010110001011), .y(t0_001011000101));
wire t0_0010110001010, t0_0010110001011;
mixer mix_t0_00101100011 (.a(t0_001011000110), .b(t0_001011000111), .y(t0_00101100011));
wire t0_001011000110, t0_001011000111;
mixer mix_t0_001011000110 (.a(t0_0010110001100), .b(t0_0010110001101), .y(t0_001011000110));
wire t0_0010110001100, t0_0010110001101;
mixer mix_t0_001011000111 (.a(t0_0010110001110), .b(t0_0010110001111), .y(t0_001011000111));
wire t0_0010110001110, t0_0010110001111;
mixer mix_t0_001011001 (.a(t0_0010110010), .b(t0_0010110011), .y(t0_001011001));
wire t0_0010110010, t0_0010110011;
mixer mix_t0_0010110010 (.a(t0_00101100100), .b(t0_00101100101), .y(t0_0010110010));
wire t0_00101100100, t0_00101100101;
mixer mix_t0_00101100100 (.a(t0_001011001000), .b(t0_001011001001), .y(t0_00101100100));
wire t0_001011001000, t0_001011001001;
mixer mix_t0_001011001000 (.a(t0_0010110010000), .b(t0_0010110010001), .y(t0_001011001000));
wire t0_0010110010000, t0_0010110010001;
mixer mix_t0_001011001001 (.a(t0_0010110010010), .b(t0_0010110010011), .y(t0_001011001001));
wire t0_0010110010010, t0_0010110010011;
mixer mix_t0_00101100101 (.a(t0_001011001010), .b(t0_001011001011), .y(t0_00101100101));
wire t0_001011001010, t0_001011001011;
mixer mix_t0_001011001010 (.a(t0_0010110010100), .b(t0_0010110010101), .y(t0_001011001010));
wire t0_0010110010100, t0_0010110010101;
mixer mix_t0_001011001011 (.a(t0_0010110010110), .b(t0_0010110010111), .y(t0_001011001011));
wire t0_0010110010110, t0_0010110010111;
mixer mix_t0_0010110011 (.a(t0_00101100110), .b(t0_00101100111), .y(t0_0010110011));
wire t0_00101100110, t0_00101100111;
mixer mix_t0_00101100110 (.a(t0_001011001100), .b(t0_001011001101), .y(t0_00101100110));
wire t0_001011001100, t0_001011001101;
mixer mix_t0_001011001100 (.a(t0_0010110011000), .b(t0_0010110011001), .y(t0_001011001100));
wire t0_0010110011000, t0_0010110011001;
mixer mix_t0_001011001101 (.a(t0_0010110011010), .b(t0_0010110011011), .y(t0_001011001101));
wire t0_0010110011010, t0_0010110011011;
mixer mix_t0_00101100111 (.a(t0_001011001110), .b(t0_001011001111), .y(t0_00101100111));
wire t0_001011001110, t0_001011001111;
mixer mix_t0_001011001110 (.a(t0_0010110011100), .b(t0_0010110011101), .y(t0_001011001110));
wire t0_0010110011100, t0_0010110011101;
mixer mix_t0_001011001111 (.a(t0_0010110011110), .b(t0_0010110011111), .y(t0_001011001111));
wire t0_0010110011110, t0_0010110011111;
mixer mix_t0_00101101 (.a(t0_001011010), .b(t0_001011011), .y(t0_00101101));
wire t0_001011010, t0_001011011;
mixer mix_t0_001011010 (.a(t0_0010110100), .b(t0_0010110101), .y(t0_001011010));
wire t0_0010110100, t0_0010110101;
mixer mix_t0_0010110100 (.a(t0_00101101000), .b(t0_00101101001), .y(t0_0010110100));
wire t0_00101101000, t0_00101101001;
mixer mix_t0_00101101000 (.a(t0_001011010000), .b(t0_001011010001), .y(t0_00101101000));
wire t0_001011010000, t0_001011010001;
mixer mix_t0_001011010000 (.a(t0_0010110100000), .b(t0_0010110100001), .y(t0_001011010000));
wire t0_0010110100000, t0_0010110100001;
mixer mix_t0_001011010001 (.a(t0_0010110100010), .b(t0_0010110100011), .y(t0_001011010001));
wire t0_0010110100010, t0_0010110100011;
mixer mix_t0_00101101001 (.a(t0_001011010010), .b(t0_001011010011), .y(t0_00101101001));
wire t0_001011010010, t0_001011010011;
mixer mix_t0_001011010010 (.a(t0_0010110100100), .b(t0_0010110100101), .y(t0_001011010010));
wire t0_0010110100100, t0_0010110100101;
mixer mix_t0_001011010011 (.a(t0_0010110100110), .b(t0_0010110100111), .y(t0_001011010011));
wire t0_0010110100110, t0_0010110100111;
mixer mix_t0_0010110101 (.a(t0_00101101010), .b(t0_00101101011), .y(t0_0010110101));
wire t0_00101101010, t0_00101101011;
mixer mix_t0_00101101010 (.a(t0_001011010100), .b(t0_001011010101), .y(t0_00101101010));
wire t0_001011010100, t0_001011010101;
mixer mix_t0_001011010100 (.a(t0_0010110101000), .b(t0_0010110101001), .y(t0_001011010100));
wire t0_0010110101000, t0_0010110101001;
mixer mix_t0_001011010101 (.a(t0_0010110101010), .b(t0_0010110101011), .y(t0_001011010101));
wire t0_0010110101010, t0_0010110101011;
mixer mix_t0_00101101011 (.a(t0_001011010110), .b(t0_001011010111), .y(t0_00101101011));
wire t0_001011010110, t0_001011010111;
mixer mix_t0_001011010110 (.a(t0_0010110101100), .b(t0_0010110101101), .y(t0_001011010110));
wire t0_0010110101100, t0_0010110101101;
mixer mix_t0_001011010111 (.a(t0_0010110101110), .b(t0_0010110101111), .y(t0_001011010111));
wire t0_0010110101110, t0_0010110101111;
mixer mix_t0_001011011 (.a(t0_0010110110), .b(t0_0010110111), .y(t0_001011011));
wire t0_0010110110, t0_0010110111;
mixer mix_t0_0010110110 (.a(t0_00101101100), .b(t0_00101101101), .y(t0_0010110110));
wire t0_00101101100, t0_00101101101;
mixer mix_t0_00101101100 (.a(t0_001011011000), .b(t0_001011011001), .y(t0_00101101100));
wire t0_001011011000, t0_001011011001;
mixer mix_t0_001011011000 (.a(t0_0010110110000), .b(t0_0010110110001), .y(t0_001011011000));
wire t0_0010110110000, t0_0010110110001;
mixer mix_t0_001011011001 (.a(t0_0010110110010), .b(t0_0010110110011), .y(t0_001011011001));
wire t0_0010110110010, t0_0010110110011;
mixer mix_t0_00101101101 (.a(t0_001011011010), .b(t0_001011011011), .y(t0_00101101101));
wire t0_001011011010, t0_001011011011;
mixer mix_t0_001011011010 (.a(t0_0010110110100), .b(t0_0010110110101), .y(t0_001011011010));
wire t0_0010110110100, t0_0010110110101;
mixer mix_t0_001011011011 (.a(t0_0010110110110), .b(t0_0010110110111), .y(t0_001011011011));
wire t0_0010110110110, t0_0010110110111;
mixer mix_t0_0010110111 (.a(t0_00101101110), .b(t0_00101101111), .y(t0_0010110111));
wire t0_00101101110, t0_00101101111;
mixer mix_t0_00101101110 (.a(t0_001011011100), .b(t0_001011011101), .y(t0_00101101110));
wire t0_001011011100, t0_001011011101;
mixer mix_t0_001011011100 (.a(t0_0010110111000), .b(t0_0010110111001), .y(t0_001011011100));
wire t0_0010110111000, t0_0010110111001;
mixer mix_t0_001011011101 (.a(t0_0010110111010), .b(t0_0010110111011), .y(t0_001011011101));
wire t0_0010110111010, t0_0010110111011;
mixer mix_t0_00101101111 (.a(t0_001011011110), .b(t0_001011011111), .y(t0_00101101111));
wire t0_001011011110, t0_001011011111;
mixer mix_t0_001011011110 (.a(t0_0010110111100), .b(t0_0010110111101), .y(t0_001011011110));
wire t0_0010110111100, t0_0010110111101;
mixer mix_t0_001011011111 (.a(t0_0010110111110), .b(t0_0010110111111), .y(t0_001011011111));
wire t0_0010110111110, t0_0010110111111;
mixer mix_t0_0010111 (.a(t0_00101110), .b(t0_00101111), .y(t0_0010111));
wire t0_00101110, t0_00101111;
mixer mix_t0_00101110 (.a(t0_001011100), .b(t0_001011101), .y(t0_00101110));
wire t0_001011100, t0_001011101;
mixer mix_t0_001011100 (.a(t0_0010111000), .b(t0_0010111001), .y(t0_001011100));
wire t0_0010111000, t0_0010111001;
mixer mix_t0_0010111000 (.a(t0_00101110000), .b(t0_00101110001), .y(t0_0010111000));
wire t0_00101110000, t0_00101110001;
mixer mix_t0_00101110000 (.a(t0_001011100000), .b(t0_001011100001), .y(t0_00101110000));
wire t0_001011100000, t0_001011100001;
mixer mix_t0_001011100000 (.a(t0_0010111000000), .b(t0_0010111000001), .y(t0_001011100000));
wire t0_0010111000000, t0_0010111000001;
mixer mix_t0_001011100001 (.a(t0_0010111000010), .b(t0_0010111000011), .y(t0_001011100001));
wire t0_0010111000010, t0_0010111000011;
mixer mix_t0_00101110001 (.a(t0_001011100010), .b(t0_001011100011), .y(t0_00101110001));
wire t0_001011100010, t0_001011100011;
mixer mix_t0_001011100010 (.a(t0_0010111000100), .b(t0_0010111000101), .y(t0_001011100010));
wire t0_0010111000100, t0_0010111000101;
mixer mix_t0_001011100011 (.a(t0_0010111000110), .b(t0_0010111000111), .y(t0_001011100011));
wire t0_0010111000110, t0_0010111000111;
mixer mix_t0_0010111001 (.a(t0_00101110010), .b(t0_00101110011), .y(t0_0010111001));
wire t0_00101110010, t0_00101110011;
mixer mix_t0_00101110010 (.a(t0_001011100100), .b(t0_001011100101), .y(t0_00101110010));
wire t0_001011100100, t0_001011100101;
mixer mix_t0_001011100100 (.a(t0_0010111001000), .b(t0_0010111001001), .y(t0_001011100100));
wire t0_0010111001000, t0_0010111001001;
mixer mix_t0_001011100101 (.a(t0_0010111001010), .b(t0_0010111001011), .y(t0_001011100101));
wire t0_0010111001010, t0_0010111001011;
mixer mix_t0_00101110011 (.a(t0_001011100110), .b(t0_001011100111), .y(t0_00101110011));
wire t0_001011100110, t0_001011100111;
mixer mix_t0_001011100110 (.a(t0_0010111001100), .b(t0_0010111001101), .y(t0_001011100110));
wire t0_0010111001100, t0_0010111001101;
mixer mix_t0_001011100111 (.a(t0_0010111001110), .b(t0_0010111001111), .y(t0_001011100111));
wire t0_0010111001110, t0_0010111001111;
mixer mix_t0_001011101 (.a(t0_0010111010), .b(t0_0010111011), .y(t0_001011101));
wire t0_0010111010, t0_0010111011;
mixer mix_t0_0010111010 (.a(t0_00101110100), .b(t0_00101110101), .y(t0_0010111010));
wire t0_00101110100, t0_00101110101;
mixer mix_t0_00101110100 (.a(t0_001011101000), .b(t0_001011101001), .y(t0_00101110100));
wire t0_001011101000, t0_001011101001;
mixer mix_t0_001011101000 (.a(t0_0010111010000), .b(t0_0010111010001), .y(t0_001011101000));
wire t0_0010111010000, t0_0010111010001;
mixer mix_t0_001011101001 (.a(t0_0010111010010), .b(t0_0010111010011), .y(t0_001011101001));
wire t0_0010111010010, t0_0010111010011;
mixer mix_t0_00101110101 (.a(t0_001011101010), .b(t0_001011101011), .y(t0_00101110101));
wire t0_001011101010, t0_001011101011;
mixer mix_t0_001011101010 (.a(t0_0010111010100), .b(t0_0010111010101), .y(t0_001011101010));
wire t0_0010111010100, t0_0010111010101;
mixer mix_t0_001011101011 (.a(t0_0010111010110), .b(t0_0010111010111), .y(t0_001011101011));
wire t0_0010111010110, t0_0010111010111;
mixer mix_t0_0010111011 (.a(t0_00101110110), .b(t0_00101110111), .y(t0_0010111011));
wire t0_00101110110, t0_00101110111;
mixer mix_t0_00101110110 (.a(t0_001011101100), .b(t0_001011101101), .y(t0_00101110110));
wire t0_001011101100, t0_001011101101;
mixer mix_t0_001011101100 (.a(t0_0010111011000), .b(t0_0010111011001), .y(t0_001011101100));
wire t0_0010111011000, t0_0010111011001;
mixer mix_t0_001011101101 (.a(t0_0010111011010), .b(t0_0010111011011), .y(t0_001011101101));
wire t0_0010111011010, t0_0010111011011;
mixer mix_t0_00101110111 (.a(t0_001011101110), .b(t0_001011101111), .y(t0_00101110111));
wire t0_001011101110, t0_001011101111;
mixer mix_t0_001011101110 (.a(t0_0010111011100), .b(t0_0010111011101), .y(t0_001011101110));
wire t0_0010111011100, t0_0010111011101;
mixer mix_t0_001011101111 (.a(t0_0010111011110), .b(t0_0010111011111), .y(t0_001011101111));
wire t0_0010111011110, t0_0010111011111;
mixer mix_t0_00101111 (.a(t0_001011110), .b(t0_001011111), .y(t0_00101111));
wire t0_001011110, t0_001011111;
mixer mix_t0_001011110 (.a(t0_0010111100), .b(t0_0010111101), .y(t0_001011110));
wire t0_0010111100, t0_0010111101;
mixer mix_t0_0010111100 (.a(t0_00101111000), .b(t0_00101111001), .y(t0_0010111100));
wire t0_00101111000, t0_00101111001;
mixer mix_t0_00101111000 (.a(t0_001011110000), .b(t0_001011110001), .y(t0_00101111000));
wire t0_001011110000, t0_001011110001;
mixer mix_t0_001011110000 (.a(t0_0010111100000), .b(t0_0010111100001), .y(t0_001011110000));
wire t0_0010111100000, t0_0010111100001;
mixer mix_t0_001011110001 (.a(t0_0010111100010), .b(t0_0010111100011), .y(t0_001011110001));
wire t0_0010111100010, t0_0010111100011;
mixer mix_t0_00101111001 (.a(t0_001011110010), .b(t0_001011110011), .y(t0_00101111001));
wire t0_001011110010, t0_001011110011;
mixer mix_t0_001011110010 (.a(t0_0010111100100), .b(t0_0010111100101), .y(t0_001011110010));
wire t0_0010111100100, t0_0010111100101;
mixer mix_t0_001011110011 (.a(t0_0010111100110), .b(t0_0010111100111), .y(t0_001011110011));
wire t0_0010111100110, t0_0010111100111;
mixer mix_t0_0010111101 (.a(t0_00101111010), .b(t0_00101111011), .y(t0_0010111101));
wire t0_00101111010, t0_00101111011;
mixer mix_t0_00101111010 (.a(t0_001011110100), .b(t0_001011110101), .y(t0_00101111010));
wire t0_001011110100, t0_001011110101;
mixer mix_t0_001011110100 (.a(t0_0010111101000), .b(t0_0010111101001), .y(t0_001011110100));
wire t0_0010111101000, t0_0010111101001;
mixer mix_t0_001011110101 (.a(t0_0010111101010), .b(t0_0010111101011), .y(t0_001011110101));
wire t0_0010111101010, t0_0010111101011;
mixer mix_t0_00101111011 (.a(t0_001011110110), .b(t0_001011110111), .y(t0_00101111011));
wire t0_001011110110, t0_001011110111;
mixer mix_t0_001011110110 (.a(t0_0010111101100), .b(t0_0010111101101), .y(t0_001011110110));
wire t0_0010111101100, t0_0010111101101;
mixer mix_t0_001011110111 (.a(t0_0010111101110), .b(t0_0010111101111), .y(t0_001011110111));
wire t0_0010111101110, t0_0010111101111;
mixer mix_t0_001011111 (.a(t0_0010111110), .b(t0_0010111111), .y(t0_001011111));
wire t0_0010111110, t0_0010111111;
mixer mix_t0_0010111110 (.a(t0_00101111100), .b(t0_00101111101), .y(t0_0010111110));
wire t0_00101111100, t0_00101111101;
mixer mix_t0_00101111100 (.a(t0_001011111000), .b(t0_001011111001), .y(t0_00101111100));
wire t0_001011111000, t0_001011111001;
mixer mix_t0_001011111000 (.a(t0_0010111110000), .b(t0_0010111110001), .y(t0_001011111000));
wire t0_0010111110000, t0_0010111110001;
mixer mix_t0_001011111001 (.a(t0_0010111110010), .b(t0_0010111110011), .y(t0_001011111001));
wire t0_0010111110010, t0_0010111110011;
mixer mix_t0_00101111101 (.a(t0_001011111010), .b(t0_001011111011), .y(t0_00101111101));
wire t0_001011111010, t0_001011111011;
mixer mix_t0_001011111010 (.a(t0_0010111110100), .b(t0_0010111110101), .y(t0_001011111010));
wire t0_0010111110100, t0_0010111110101;
mixer mix_t0_001011111011 (.a(t0_0010111110110), .b(t0_0010111110111), .y(t0_001011111011));
wire t0_0010111110110, t0_0010111110111;
mixer mix_t0_0010111111 (.a(t0_00101111110), .b(t0_00101111111), .y(t0_0010111111));
wire t0_00101111110, t0_00101111111;
mixer mix_t0_00101111110 (.a(t0_001011111100), .b(t0_001011111101), .y(t0_00101111110));
wire t0_001011111100, t0_001011111101;
mixer mix_t0_001011111100 (.a(t0_0010111111000), .b(t0_0010111111001), .y(t0_001011111100));
wire t0_0010111111000, t0_0010111111001;
mixer mix_t0_001011111101 (.a(t0_0010111111010), .b(t0_0010111111011), .y(t0_001011111101));
wire t0_0010111111010, t0_0010111111011;
mixer mix_t0_00101111111 (.a(t0_001011111110), .b(t0_001011111111), .y(t0_00101111111));
wire t0_001011111110, t0_001011111111;
mixer mix_t0_001011111110 (.a(t0_0010111111100), .b(t0_0010111111101), .y(t0_001011111110));
wire t0_0010111111100, t0_0010111111101;
mixer mix_t0_001011111111 (.a(t0_0010111111110), .b(t0_0010111111111), .y(t0_001011111111));
wire t0_0010111111110, t0_0010111111111;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_001100 (.a(t0_0011000), .b(t0_0011001), .y(t0_001100));
wire t0_0011000, t0_0011001;
mixer mix_t0_0011000 (.a(t0_00110000), .b(t0_00110001), .y(t0_0011000));
wire t0_00110000, t0_00110001;
mixer mix_t0_00110000 (.a(t0_001100000), .b(t0_001100001), .y(t0_00110000));
wire t0_001100000, t0_001100001;
mixer mix_t0_001100000 (.a(t0_0011000000), .b(t0_0011000001), .y(t0_001100000));
wire t0_0011000000, t0_0011000001;
mixer mix_t0_0011000000 (.a(t0_00110000000), .b(t0_00110000001), .y(t0_0011000000));
wire t0_00110000000, t0_00110000001;
mixer mix_t0_00110000000 (.a(t0_001100000000), .b(t0_001100000001), .y(t0_00110000000));
wire t0_001100000000, t0_001100000001;
mixer mix_t0_001100000000 (.a(t0_0011000000000), .b(t0_0011000000001), .y(t0_001100000000));
wire t0_0011000000000, t0_0011000000001;
mixer mix_t0_001100000001 (.a(t0_0011000000010), .b(t0_0011000000011), .y(t0_001100000001));
wire t0_0011000000010, t0_0011000000011;
mixer mix_t0_00110000001 (.a(t0_001100000010), .b(t0_001100000011), .y(t0_00110000001));
wire t0_001100000010, t0_001100000011;
mixer mix_t0_001100000010 (.a(t0_0011000000100), .b(t0_0011000000101), .y(t0_001100000010));
wire t0_0011000000100, t0_0011000000101;
mixer mix_t0_001100000011 (.a(t0_0011000000110), .b(t0_0011000000111), .y(t0_001100000011));
wire t0_0011000000110, t0_0011000000111;
mixer mix_t0_0011000001 (.a(t0_00110000010), .b(t0_00110000011), .y(t0_0011000001));
wire t0_00110000010, t0_00110000011;
mixer mix_t0_00110000010 (.a(t0_001100000100), .b(t0_001100000101), .y(t0_00110000010));
wire t0_001100000100, t0_001100000101;
mixer mix_t0_001100000100 (.a(t0_0011000001000), .b(t0_0011000001001), .y(t0_001100000100));
wire t0_0011000001000, t0_0011000001001;
mixer mix_t0_001100000101 (.a(t0_0011000001010), .b(t0_0011000001011), .y(t0_001100000101));
wire t0_0011000001010, t0_0011000001011;
mixer mix_t0_00110000011 (.a(t0_001100000110), .b(t0_001100000111), .y(t0_00110000011));
wire t0_001100000110, t0_001100000111;
mixer mix_t0_001100000110 (.a(t0_0011000001100), .b(t0_0011000001101), .y(t0_001100000110));
wire t0_0011000001100, t0_0011000001101;
mixer mix_t0_001100000111 (.a(t0_0011000001110), .b(t0_0011000001111), .y(t0_001100000111));
wire t0_0011000001110, t0_0011000001111;
mixer mix_t0_001100001 (.a(t0_0011000010), .b(t0_0011000011), .y(t0_001100001));
wire t0_0011000010, t0_0011000011;
mixer mix_t0_0011000010 (.a(t0_00110000100), .b(t0_00110000101), .y(t0_0011000010));
wire t0_00110000100, t0_00110000101;
mixer mix_t0_00110000100 (.a(t0_001100001000), .b(t0_001100001001), .y(t0_00110000100));
wire t0_001100001000, t0_001100001001;
mixer mix_t0_001100001000 (.a(t0_0011000010000), .b(t0_0011000010001), .y(t0_001100001000));
wire t0_0011000010000, t0_0011000010001;
mixer mix_t0_001100001001 (.a(t0_0011000010010), .b(t0_0011000010011), .y(t0_001100001001));
wire t0_0011000010010, t0_0011000010011;
mixer mix_t0_00110000101 (.a(t0_001100001010), .b(t0_001100001011), .y(t0_00110000101));
wire t0_001100001010, t0_001100001011;
mixer mix_t0_001100001010 (.a(t0_0011000010100), .b(t0_0011000010101), .y(t0_001100001010));
wire t0_0011000010100, t0_0011000010101;
mixer mix_t0_001100001011 (.a(t0_0011000010110), .b(t0_0011000010111), .y(t0_001100001011));
wire t0_0011000010110, t0_0011000010111;
mixer mix_t0_0011000011 (.a(t0_00110000110), .b(t0_00110000111), .y(t0_0011000011));
wire t0_00110000110, t0_00110000111;
mixer mix_t0_00110000110 (.a(t0_001100001100), .b(t0_001100001101), .y(t0_00110000110));
wire t0_001100001100, t0_001100001101;
mixer mix_t0_001100001100 (.a(t0_0011000011000), .b(t0_0011000011001), .y(t0_001100001100));
wire t0_0011000011000, t0_0011000011001;
mixer mix_t0_001100001101 (.a(t0_0011000011010), .b(t0_0011000011011), .y(t0_001100001101));
wire t0_0011000011010, t0_0011000011011;
mixer mix_t0_00110000111 (.a(t0_001100001110), .b(t0_001100001111), .y(t0_00110000111));
wire t0_001100001110, t0_001100001111;
mixer mix_t0_001100001110 (.a(t0_0011000011100), .b(t0_0011000011101), .y(t0_001100001110));
wire t0_0011000011100, t0_0011000011101;
mixer mix_t0_001100001111 (.a(t0_0011000011110), .b(t0_0011000011111), .y(t0_001100001111));
wire t0_0011000011110, t0_0011000011111;
mixer mix_t0_00110001 (.a(t0_001100010), .b(t0_001100011), .y(t0_00110001));
wire t0_001100010, t0_001100011;
mixer mix_t0_001100010 (.a(t0_0011000100), .b(t0_0011000101), .y(t0_001100010));
wire t0_0011000100, t0_0011000101;
mixer mix_t0_0011000100 (.a(t0_00110001000), .b(t0_00110001001), .y(t0_0011000100));
wire t0_00110001000, t0_00110001001;
mixer mix_t0_00110001000 (.a(t0_001100010000), .b(t0_001100010001), .y(t0_00110001000));
wire t0_001100010000, t0_001100010001;
mixer mix_t0_001100010000 (.a(t0_0011000100000), .b(t0_0011000100001), .y(t0_001100010000));
wire t0_0011000100000, t0_0011000100001;
mixer mix_t0_001100010001 (.a(t0_0011000100010), .b(t0_0011000100011), .y(t0_001100010001));
wire t0_0011000100010, t0_0011000100011;
mixer mix_t0_00110001001 (.a(t0_001100010010), .b(t0_001100010011), .y(t0_00110001001));
wire t0_001100010010, t0_001100010011;
mixer mix_t0_001100010010 (.a(t0_0011000100100), .b(t0_0011000100101), .y(t0_001100010010));
wire t0_0011000100100, t0_0011000100101;
mixer mix_t0_001100010011 (.a(t0_0011000100110), .b(t0_0011000100111), .y(t0_001100010011));
wire t0_0011000100110, t0_0011000100111;
mixer mix_t0_0011000101 (.a(t0_00110001010), .b(t0_00110001011), .y(t0_0011000101));
wire t0_00110001010, t0_00110001011;
mixer mix_t0_00110001010 (.a(t0_001100010100), .b(t0_001100010101), .y(t0_00110001010));
wire t0_001100010100, t0_001100010101;
mixer mix_t0_001100010100 (.a(t0_0011000101000), .b(t0_0011000101001), .y(t0_001100010100));
wire t0_0011000101000, t0_0011000101001;
mixer mix_t0_001100010101 (.a(t0_0011000101010), .b(t0_0011000101011), .y(t0_001100010101));
wire t0_0011000101010, t0_0011000101011;
mixer mix_t0_00110001011 (.a(t0_001100010110), .b(t0_001100010111), .y(t0_00110001011));
wire t0_001100010110, t0_001100010111;
mixer mix_t0_001100010110 (.a(t0_0011000101100), .b(t0_0011000101101), .y(t0_001100010110));
wire t0_0011000101100, t0_0011000101101;
mixer mix_t0_001100010111 (.a(t0_0011000101110), .b(t0_0011000101111), .y(t0_001100010111));
wire t0_0011000101110, t0_0011000101111;
mixer mix_t0_001100011 (.a(t0_0011000110), .b(t0_0011000111), .y(t0_001100011));
wire t0_0011000110, t0_0011000111;
mixer mix_t0_0011000110 (.a(t0_00110001100), .b(t0_00110001101), .y(t0_0011000110));
wire t0_00110001100, t0_00110001101;
mixer mix_t0_00110001100 (.a(t0_001100011000), .b(t0_001100011001), .y(t0_00110001100));
wire t0_001100011000, t0_001100011001;
mixer mix_t0_001100011000 (.a(t0_0011000110000), .b(t0_0011000110001), .y(t0_001100011000));
wire t0_0011000110000, t0_0011000110001;
mixer mix_t0_001100011001 (.a(t0_0011000110010), .b(t0_0011000110011), .y(t0_001100011001));
wire t0_0011000110010, t0_0011000110011;
mixer mix_t0_00110001101 (.a(t0_001100011010), .b(t0_001100011011), .y(t0_00110001101));
wire t0_001100011010, t0_001100011011;
mixer mix_t0_001100011010 (.a(t0_0011000110100), .b(t0_0011000110101), .y(t0_001100011010));
wire t0_0011000110100, t0_0011000110101;
mixer mix_t0_001100011011 (.a(t0_0011000110110), .b(t0_0011000110111), .y(t0_001100011011));
wire t0_0011000110110, t0_0011000110111;
mixer mix_t0_0011000111 (.a(t0_00110001110), .b(t0_00110001111), .y(t0_0011000111));
wire t0_00110001110, t0_00110001111;
mixer mix_t0_00110001110 (.a(t0_001100011100), .b(t0_001100011101), .y(t0_00110001110));
wire t0_001100011100, t0_001100011101;
mixer mix_t0_001100011100 (.a(t0_0011000111000), .b(t0_0011000111001), .y(t0_001100011100));
wire t0_0011000111000, t0_0011000111001;
mixer mix_t0_001100011101 (.a(t0_0011000111010), .b(t0_0011000111011), .y(t0_001100011101));
wire t0_0011000111010, t0_0011000111011;
mixer mix_t0_00110001111 (.a(t0_001100011110), .b(t0_001100011111), .y(t0_00110001111));
wire t0_001100011110, t0_001100011111;
mixer mix_t0_001100011110 (.a(t0_0011000111100), .b(t0_0011000111101), .y(t0_001100011110));
wire t0_0011000111100, t0_0011000111101;
mixer mix_t0_001100011111 (.a(t0_0011000111110), .b(t0_0011000111111), .y(t0_001100011111));
wire t0_0011000111110, t0_0011000111111;
mixer mix_t0_0011001 (.a(t0_00110010), .b(t0_00110011), .y(t0_0011001));
wire t0_00110010, t0_00110011;
mixer mix_t0_00110010 (.a(t0_001100100), .b(t0_001100101), .y(t0_00110010));
wire t0_001100100, t0_001100101;
mixer mix_t0_001100100 (.a(t0_0011001000), .b(t0_0011001001), .y(t0_001100100));
wire t0_0011001000, t0_0011001001;
mixer mix_t0_0011001000 (.a(t0_00110010000), .b(t0_00110010001), .y(t0_0011001000));
wire t0_00110010000, t0_00110010001;
mixer mix_t0_00110010000 (.a(t0_001100100000), .b(t0_001100100001), .y(t0_00110010000));
wire t0_001100100000, t0_001100100001;
mixer mix_t0_001100100000 (.a(t0_0011001000000), .b(t0_0011001000001), .y(t0_001100100000));
wire t0_0011001000000, t0_0011001000001;
mixer mix_t0_001100100001 (.a(t0_0011001000010), .b(t0_0011001000011), .y(t0_001100100001));
wire t0_0011001000010, t0_0011001000011;
mixer mix_t0_00110010001 (.a(t0_001100100010), .b(t0_001100100011), .y(t0_00110010001));
wire t0_001100100010, t0_001100100011;
mixer mix_t0_001100100010 (.a(t0_0011001000100), .b(t0_0011001000101), .y(t0_001100100010));
wire t0_0011001000100, t0_0011001000101;
mixer mix_t0_001100100011 (.a(t0_0011001000110), .b(t0_0011001000111), .y(t0_001100100011));
wire t0_0011001000110, t0_0011001000111;
mixer mix_t0_0011001001 (.a(t0_00110010010), .b(t0_00110010011), .y(t0_0011001001));
wire t0_00110010010, t0_00110010011;
mixer mix_t0_00110010010 (.a(t0_001100100100), .b(t0_001100100101), .y(t0_00110010010));
wire t0_001100100100, t0_001100100101;
mixer mix_t0_001100100100 (.a(t0_0011001001000), .b(t0_0011001001001), .y(t0_001100100100));
wire t0_0011001001000, t0_0011001001001;
mixer mix_t0_001100100101 (.a(t0_0011001001010), .b(t0_0011001001011), .y(t0_001100100101));
wire t0_0011001001010, t0_0011001001011;
mixer mix_t0_00110010011 (.a(t0_001100100110), .b(t0_001100100111), .y(t0_00110010011));
wire t0_001100100110, t0_001100100111;
mixer mix_t0_001100100110 (.a(t0_0011001001100), .b(t0_0011001001101), .y(t0_001100100110));
wire t0_0011001001100, t0_0011001001101;
mixer mix_t0_001100100111 (.a(t0_0011001001110), .b(t0_0011001001111), .y(t0_001100100111));
wire t0_0011001001110, t0_0011001001111;
mixer mix_t0_001100101 (.a(t0_0011001010), .b(t0_0011001011), .y(t0_001100101));
wire t0_0011001010, t0_0011001011;
mixer mix_t0_0011001010 (.a(t0_00110010100), .b(t0_00110010101), .y(t0_0011001010));
wire t0_00110010100, t0_00110010101;
mixer mix_t0_00110010100 (.a(t0_001100101000), .b(t0_001100101001), .y(t0_00110010100));
wire t0_001100101000, t0_001100101001;
mixer mix_t0_001100101000 (.a(t0_0011001010000), .b(t0_0011001010001), .y(t0_001100101000));
wire t0_0011001010000, t0_0011001010001;
mixer mix_t0_001100101001 (.a(t0_0011001010010), .b(t0_0011001010011), .y(t0_001100101001));
wire t0_0011001010010, t0_0011001010011;
mixer mix_t0_00110010101 (.a(t0_001100101010), .b(t0_001100101011), .y(t0_00110010101));
wire t0_001100101010, t0_001100101011;
mixer mix_t0_001100101010 (.a(t0_0011001010100), .b(t0_0011001010101), .y(t0_001100101010));
wire t0_0011001010100, t0_0011001010101;
mixer mix_t0_001100101011 (.a(t0_0011001010110), .b(t0_0011001010111), .y(t0_001100101011));
wire t0_0011001010110, t0_0011001010111;
mixer mix_t0_0011001011 (.a(t0_00110010110), .b(t0_00110010111), .y(t0_0011001011));
wire t0_00110010110, t0_00110010111;
mixer mix_t0_00110010110 (.a(t0_001100101100), .b(t0_001100101101), .y(t0_00110010110));
wire t0_001100101100, t0_001100101101;
mixer mix_t0_001100101100 (.a(t0_0011001011000), .b(t0_0011001011001), .y(t0_001100101100));
wire t0_0011001011000, t0_0011001011001;
mixer mix_t0_001100101101 (.a(t0_0011001011010), .b(t0_0011001011011), .y(t0_001100101101));
wire t0_0011001011010, t0_0011001011011;
mixer mix_t0_00110010111 (.a(t0_001100101110), .b(t0_001100101111), .y(t0_00110010111));
wire t0_001100101110, t0_001100101111;
mixer mix_t0_001100101110 (.a(t0_0011001011100), .b(t0_0011001011101), .y(t0_001100101110));
wire t0_0011001011100, t0_0011001011101;
mixer mix_t0_001100101111 (.a(t0_0011001011110), .b(t0_0011001011111), .y(t0_001100101111));
wire t0_0011001011110, t0_0011001011111;
mixer mix_t0_00110011 (.a(t0_001100110), .b(t0_001100111), .y(t0_00110011));
wire t0_001100110, t0_001100111;
mixer mix_t0_001100110 (.a(t0_0011001100), .b(t0_0011001101), .y(t0_001100110));
wire t0_0011001100, t0_0011001101;
mixer mix_t0_0011001100 (.a(t0_00110011000), .b(t0_00110011001), .y(t0_0011001100));
wire t0_00110011000, t0_00110011001;
mixer mix_t0_00110011000 (.a(t0_001100110000), .b(t0_001100110001), .y(t0_00110011000));
wire t0_001100110000, t0_001100110001;
mixer mix_t0_001100110000 (.a(t0_0011001100000), .b(t0_0011001100001), .y(t0_001100110000));
wire t0_0011001100000, t0_0011001100001;
mixer mix_t0_001100110001 (.a(t0_0011001100010), .b(t0_0011001100011), .y(t0_001100110001));
wire t0_0011001100010, t0_0011001100011;
mixer mix_t0_00110011001 (.a(t0_001100110010), .b(t0_001100110011), .y(t0_00110011001));
wire t0_001100110010, t0_001100110011;
mixer mix_t0_001100110010 (.a(t0_0011001100100), .b(t0_0011001100101), .y(t0_001100110010));
wire t0_0011001100100, t0_0011001100101;
mixer mix_t0_001100110011 (.a(t0_0011001100110), .b(t0_0011001100111), .y(t0_001100110011));
wire t0_0011001100110, t0_0011001100111;
mixer mix_t0_0011001101 (.a(t0_00110011010), .b(t0_00110011011), .y(t0_0011001101));
wire t0_00110011010, t0_00110011011;
mixer mix_t0_00110011010 (.a(t0_001100110100), .b(t0_001100110101), .y(t0_00110011010));
wire t0_001100110100, t0_001100110101;
mixer mix_t0_001100110100 (.a(t0_0011001101000), .b(t0_0011001101001), .y(t0_001100110100));
wire t0_0011001101000, t0_0011001101001;
mixer mix_t0_001100110101 (.a(t0_0011001101010), .b(t0_0011001101011), .y(t0_001100110101));
wire t0_0011001101010, t0_0011001101011;
mixer mix_t0_00110011011 (.a(t0_001100110110), .b(t0_001100110111), .y(t0_00110011011));
wire t0_001100110110, t0_001100110111;
mixer mix_t0_001100110110 (.a(t0_0011001101100), .b(t0_0011001101101), .y(t0_001100110110));
wire t0_0011001101100, t0_0011001101101;
mixer mix_t0_001100110111 (.a(t0_0011001101110), .b(t0_0011001101111), .y(t0_001100110111));
wire t0_0011001101110, t0_0011001101111;
mixer mix_t0_001100111 (.a(t0_0011001110), .b(t0_0011001111), .y(t0_001100111));
wire t0_0011001110, t0_0011001111;
mixer mix_t0_0011001110 (.a(t0_00110011100), .b(t0_00110011101), .y(t0_0011001110));
wire t0_00110011100, t0_00110011101;
mixer mix_t0_00110011100 (.a(t0_001100111000), .b(t0_001100111001), .y(t0_00110011100));
wire t0_001100111000, t0_001100111001;
mixer mix_t0_001100111000 (.a(t0_0011001110000), .b(t0_0011001110001), .y(t0_001100111000));
wire t0_0011001110000, t0_0011001110001;
mixer mix_t0_001100111001 (.a(t0_0011001110010), .b(t0_0011001110011), .y(t0_001100111001));
wire t0_0011001110010, t0_0011001110011;
mixer mix_t0_00110011101 (.a(t0_001100111010), .b(t0_001100111011), .y(t0_00110011101));
wire t0_001100111010, t0_001100111011;
mixer mix_t0_001100111010 (.a(t0_0011001110100), .b(t0_0011001110101), .y(t0_001100111010));
wire t0_0011001110100, t0_0011001110101;
mixer mix_t0_001100111011 (.a(t0_0011001110110), .b(t0_0011001110111), .y(t0_001100111011));
wire t0_0011001110110, t0_0011001110111;
mixer mix_t0_0011001111 (.a(t0_00110011110), .b(t0_00110011111), .y(t0_0011001111));
wire t0_00110011110, t0_00110011111;
mixer mix_t0_00110011110 (.a(t0_001100111100), .b(t0_001100111101), .y(t0_00110011110));
wire t0_001100111100, t0_001100111101;
mixer mix_t0_001100111100 (.a(t0_0011001111000), .b(t0_0011001111001), .y(t0_001100111100));
wire t0_0011001111000, t0_0011001111001;
mixer mix_t0_001100111101 (.a(t0_0011001111010), .b(t0_0011001111011), .y(t0_001100111101));
wire t0_0011001111010, t0_0011001111011;
mixer mix_t0_00110011111 (.a(t0_001100111110), .b(t0_001100111111), .y(t0_00110011111));
wire t0_001100111110, t0_001100111111;
mixer mix_t0_001100111110 (.a(t0_0011001111100), .b(t0_0011001111101), .y(t0_001100111110));
wire t0_0011001111100, t0_0011001111101;
mixer mix_t0_001100111111 (.a(t0_0011001111110), .b(t0_0011001111111), .y(t0_001100111111));
wire t0_0011001111110, t0_0011001111111;
mixer mix_t0_001101 (.a(t0_0011010), .b(t0_0011011), .y(t0_001101));
wire t0_0011010, t0_0011011;
mixer mix_t0_0011010 (.a(t0_00110100), .b(t0_00110101), .y(t0_0011010));
wire t0_00110100, t0_00110101;
mixer mix_t0_00110100 (.a(t0_001101000), .b(t0_001101001), .y(t0_00110100));
wire t0_001101000, t0_001101001;
mixer mix_t0_001101000 (.a(t0_0011010000), .b(t0_0011010001), .y(t0_001101000));
wire t0_0011010000, t0_0011010001;
mixer mix_t0_0011010000 (.a(t0_00110100000), .b(t0_00110100001), .y(t0_0011010000));
wire t0_00110100000, t0_00110100001;
mixer mix_t0_00110100000 (.a(t0_001101000000), .b(t0_001101000001), .y(t0_00110100000));
wire t0_001101000000, t0_001101000001;
mixer mix_t0_001101000000 (.a(t0_0011010000000), .b(t0_0011010000001), .y(t0_001101000000));
wire t0_0011010000000, t0_0011010000001;
mixer mix_t0_001101000001 (.a(t0_0011010000010), .b(t0_0011010000011), .y(t0_001101000001));
wire t0_0011010000010, t0_0011010000011;
mixer mix_t0_00110100001 (.a(t0_001101000010), .b(t0_001101000011), .y(t0_00110100001));
wire t0_001101000010, t0_001101000011;
mixer mix_t0_001101000010 (.a(t0_0011010000100), .b(t0_0011010000101), .y(t0_001101000010));
wire t0_0011010000100, t0_0011010000101;
mixer mix_t0_001101000011 (.a(t0_0011010000110), .b(t0_0011010000111), .y(t0_001101000011));
wire t0_0011010000110, t0_0011010000111;
mixer mix_t0_0011010001 (.a(t0_00110100010), .b(t0_00110100011), .y(t0_0011010001));
wire t0_00110100010, t0_00110100011;
mixer mix_t0_00110100010 (.a(t0_001101000100), .b(t0_001101000101), .y(t0_00110100010));
wire t0_001101000100, t0_001101000101;
mixer mix_t0_001101000100 (.a(t0_0011010001000), .b(t0_0011010001001), .y(t0_001101000100));
wire t0_0011010001000, t0_0011010001001;
mixer mix_t0_001101000101 (.a(t0_0011010001010), .b(t0_0011010001011), .y(t0_001101000101));
wire t0_0011010001010, t0_0011010001011;
mixer mix_t0_00110100011 (.a(t0_001101000110), .b(t0_001101000111), .y(t0_00110100011));
wire t0_001101000110, t0_001101000111;
mixer mix_t0_001101000110 (.a(t0_0011010001100), .b(t0_0011010001101), .y(t0_001101000110));
wire t0_0011010001100, t0_0011010001101;
mixer mix_t0_001101000111 (.a(t0_0011010001110), .b(t0_0011010001111), .y(t0_001101000111));
wire t0_0011010001110, t0_0011010001111;
mixer mix_t0_001101001 (.a(t0_0011010010), .b(t0_0011010011), .y(t0_001101001));
wire t0_0011010010, t0_0011010011;
mixer mix_t0_0011010010 (.a(t0_00110100100), .b(t0_00110100101), .y(t0_0011010010));
wire t0_00110100100, t0_00110100101;
mixer mix_t0_00110100100 (.a(t0_001101001000), .b(t0_001101001001), .y(t0_00110100100));
wire t0_001101001000, t0_001101001001;
mixer mix_t0_001101001000 (.a(t0_0011010010000), .b(t0_0011010010001), .y(t0_001101001000));
wire t0_0011010010000, t0_0011010010001;
mixer mix_t0_001101001001 (.a(t0_0011010010010), .b(t0_0011010010011), .y(t0_001101001001));
wire t0_0011010010010, t0_0011010010011;
mixer mix_t0_00110100101 (.a(t0_001101001010), .b(t0_001101001011), .y(t0_00110100101));
wire t0_001101001010, t0_001101001011;
mixer mix_t0_001101001010 (.a(t0_0011010010100), .b(t0_0011010010101), .y(t0_001101001010));
wire t0_0011010010100, t0_0011010010101;
mixer mix_t0_001101001011 (.a(t0_0011010010110), .b(t0_0011010010111), .y(t0_001101001011));
wire t0_0011010010110, t0_0011010010111;
mixer mix_t0_0011010011 (.a(t0_00110100110), .b(t0_00110100111), .y(t0_0011010011));
wire t0_00110100110, t0_00110100111;
mixer mix_t0_00110100110 (.a(t0_001101001100), .b(t0_001101001101), .y(t0_00110100110));
wire t0_001101001100, t0_001101001101;
mixer mix_t0_001101001100 (.a(t0_0011010011000), .b(t0_0011010011001), .y(t0_001101001100));
wire t0_0011010011000, t0_0011010011001;
mixer mix_t0_001101001101 (.a(t0_0011010011010), .b(t0_0011010011011), .y(t0_001101001101));
wire t0_0011010011010, t0_0011010011011;
mixer mix_t0_00110100111 (.a(t0_001101001110), .b(t0_001101001111), .y(t0_00110100111));
wire t0_001101001110, t0_001101001111;
mixer mix_t0_001101001110 (.a(t0_0011010011100), .b(t0_0011010011101), .y(t0_001101001110));
wire t0_0011010011100, t0_0011010011101;
mixer mix_t0_001101001111 (.a(t0_0011010011110), .b(t0_0011010011111), .y(t0_001101001111));
wire t0_0011010011110, t0_0011010011111;
mixer mix_t0_00110101 (.a(t0_001101010), .b(t0_001101011), .y(t0_00110101));
wire t0_001101010, t0_001101011;
mixer mix_t0_001101010 (.a(t0_0011010100), .b(t0_0011010101), .y(t0_001101010));
wire t0_0011010100, t0_0011010101;
mixer mix_t0_0011010100 (.a(t0_00110101000), .b(t0_00110101001), .y(t0_0011010100));
wire t0_00110101000, t0_00110101001;
mixer mix_t0_00110101000 (.a(t0_001101010000), .b(t0_001101010001), .y(t0_00110101000));
wire t0_001101010000, t0_001101010001;
mixer mix_t0_001101010000 (.a(t0_0011010100000), .b(t0_0011010100001), .y(t0_001101010000));
wire t0_0011010100000, t0_0011010100001;
mixer mix_t0_001101010001 (.a(t0_0011010100010), .b(t0_0011010100011), .y(t0_001101010001));
wire t0_0011010100010, t0_0011010100011;
mixer mix_t0_00110101001 (.a(t0_001101010010), .b(t0_001101010011), .y(t0_00110101001));
wire t0_001101010010, t0_001101010011;
mixer mix_t0_001101010010 (.a(t0_0011010100100), .b(t0_0011010100101), .y(t0_001101010010));
wire t0_0011010100100, t0_0011010100101;
mixer mix_t0_001101010011 (.a(t0_0011010100110), .b(t0_0011010100111), .y(t0_001101010011));
wire t0_0011010100110, t0_0011010100111;
mixer mix_t0_0011010101 (.a(t0_00110101010), .b(t0_00110101011), .y(t0_0011010101));
wire t0_00110101010, t0_00110101011;
mixer mix_t0_00110101010 (.a(t0_001101010100), .b(t0_001101010101), .y(t0_00110101010));
wire t0_001101010100, t0_001101010101;
mixer mix_t0_001101010100 (.a(t0_0011010101000), .b(t0_0011010101001), .y(t0_001101010100));
wire t0_0011010101000, t0_0011010101001;
mixer mix_t0_001101010101 (.a(t0_0011010101010), .b(t0_0011010101011), .y(t0_001101010101));
wire t0_0011010101010, t0_0011010101011;
mixer mix_t0_00110101011 (.a(t0_001101010110), .b(t0_001101010111), .y(t0_00110101011));
wire t0_001101010110, t0_001101010111;
mixer mix_t0_001101010110 (.a(t0_0011010101100), .b(t0_0011010101101), .y(t0_001101010110));
wire t0_0011010101100, t0_0011010101101;
mixer mix_t0_001101010111 (.a(t0_0011010101110), .b(t0_0011010101111), .y(t0_001101010111));
wire t0_0011010101110, t0_0011010101111;
mixer mix_t0_001101011 (.a(t0_0011010110), .b(t0_0011010111), .y(t0_001101011));
wire t0_0011010110, t0_0011010111;
mixer mix_t0_0011010110 (.a(t0_00110101100), .b(t0_00110101101), .y(t0_0011010110));
wire t0_00110101100, t0_00110101101;
mixer mix_t0_00110101100 (.a(t0_001101011000), .b(t0_001101011001), .y(t0_00110101100));
wire t0_001101011000, t0_001101011001;
mixer mix_t0_001101011000 (.a(t0_0011010110000), .b(t0_0011010110001), .y(t0_001101011000));
wire t0_0011010110000, t0_0011010110001;
mixer mix_t0_001101011001 (.a(t0_0011010110010), .b(t0_0011010110011), .y(t0_001101011001));
wire t0_0011010110010, t0_0011010110011;
mixer mix_t0_00110101101 (.a(t0_001101011010), .b(t0_001101011011), .y(t0_00110101101));
wire t0_001101011010, t0_001101011011;
mixer mix_t0_001101011010 (.a(t0_0011010110100), .b(t0_0011010110101), .y(t0_001101011010));
wire t0_0011010110100, t0_0011010110101;
mixer mix_t0_001101011011 (.a(t0_0011010110110), .b(t0_0011010110111), .y(t0_001101011011));
wire t0_0011010110110, t0_0011010110111;
mixer mix_t0_0011010111 (.a(t0_00110101110), .b(t0_00110101111), .y(t0_0011010111));
wire t0_00110101110, t0_00110101111;
mixer mix_t0_00110101110 (.a(t0_001101011100), .b(t0_001101011101), .y(t0_00110101110));
wire t0_001101011100, t0_001101011101;
mixer mix_t0_001101011100 (.a(t0_0011010111000), .b(t0_0011010111001), .y(t0_001101011100));
wire t0_0011010111000, t0_0011010111001;
mixer mix_t0_001101011101 (.a(t0_0011010111010), .b(t0_0011010111011), .y(t0_001101011101));
wire t0_0011010111010, t0_0011010111011;
mixer mix_t0_00110101111 (.a(t0_001101011110), .b(t0_001101011111), .y(t0_00110101111));
wire t0_001101011110, t0_001101011111;
mixer mix_t0_001101011110 (.a(t0_0011010111100), .b(t0_0011010111101), .y(t0_001101011110));
wire t0_0011010111100, t0_0011010111101;
mixer mix_t0_001101011111 (.a(t0_0011010111110), .b(t0_0011010111111), .y(t0_001101011111));
wire t0_0011010111110, t0_0011010111111;
mixer mix_t0_0011011 (.a(t0_00110110), .b(t0_00110111), .y(t0_0011011));
wire t0_00110110, t0_00110111;
mixer mix_t0_00110110 (.a(t0_001101100), .b(t0_001101101), .y(t0_00110110));
wire t0_001101100, t0_001101101;
mixer mix_t0_001101100 (.a(t0_0011011000), .b(t0_0011011001), .y(t0_001101100));
wire t0_0011011000, t0_0011011001;
mixer mix_t0_0011011000 (.a(t0_00110110000), .b(t0_00110110001), .y(t0_0011011000));
wire t0_00110110000, t0_00110110001;
mixer mix_t0_00110110000 (.a(t0_001101100000), .b(t0_001101100001), .y(t0_00110110000));
wire t0_001101100000, t0_001101100001;
mixer mix_t0_001101100000 (.a(t0_0011011000000), .b(t0_0011011000001), .y(t0_001101100000));
wire t0_0011011000000, t0_0011011000001;
mixer mix_t0_001101100001 (.a(t0_0011011000010), .b(t0_0011011000011), .y(t0_001101100001));
wire t0_0011011000010, t0_0011011000011;
mixer mix_t0_00110110001 (.a(t0_001101100010), .b(t0_001101100011), .y(t0_00110110001));
wire t0_001101100010, t0_001101100011;
mixer mix_t0_001101100010 (.a(t0_0011011000100), .b(t0_0011011000101), .y(t0_001101100010));
wire t0_0011011000100, t0_0011011000101;
mixer mix_t0_001101100011 (.a(t0_0011011000110), .b(t0_0011011000111), .y(t0_001101100011));
wire t0_0011011000110, t0_0011011000111;
mixer mix_t0_0011011001 (.a(t0_00110110010), .b(t0_00110110011), .y(t0_0011011001));
wire t0_00110110010, t0_00110110011;
mixer mix_t0_00110110010 (.a(t0_001101100100), .b(t0_001101100101), .y(t0_00110110010));
wire t0_001101100100, t0_001101100101;
mixer mix_t0_001101100100 (.a(t0_0011011001000), .b(t0_0011011001001), .y(t0_001101100100));
wire t0_0011011001000, t0_0011011001001;
mixer mix_t0_001101100101 (.a(t0_0011011001010), .b(t0_0011011001011), .y(t0_001101100101));
wire t0_0011011001010, t0_0011011001011;
mixer mix_t0_00110110011 (.a(t0_001101100110), .b(t0_001101100111), .y(t0_00110110011));
wire t0_001101100110, t0_001101100111;
mixer mix_t0_001101100110 (.a(t0_0011011001100), .b(t0_0011011001101), .y(t0_001101100110));
wire t0_0011011001100, t0_0011011001101;
mixer mix_t0_001101100111 (.a(t0_0011011001110), .b(t0_0011011001111), .y(t0_001101100111));
wire t0_0011011001110, t0_0011011001111;
mixer mix_t0_001101101 (.a(t0_0011011010), .b(t0_0011011011), .y(t0_001101101));
wire t0_0011011010, t0_0011011011;
mixer mix_t0_0011011010 (.a(t0_00110110100), .b(t0_00110110101), .y(t0_0011011010));
wire t0_00110110100, t0_00110110101;
mixer mix_t0_00110110100 (.a(t0_001101101000), .b(t0_001101101001), .y(t0_00110110100));
wire t0_001101101000, t0_001101101001;
mixer mix_t0_001101101000 (.a(t0_0011011010000), .b(t0_0011011010001), .y(t0_001101101000));
wire t0_0011011010000, t0_0011011010001;
mixer mix_t0_001101101001 (.a(t0_0011011010010), .b(t0_0011011010011), .y(t0_001101101001));
wire t0_0011011010010, t0_0011011010011;
mixer mix_t0_00110110101 (.a(t0_001101101010), .b(t0_001101101011), .y(t0_00110110101));
wire t0_001101101010, t0_001101101011;
mixer mix_t0_001101101010 (.a(t0_0011011010100), .b(t0_0011011010101), .y(t0_001101101010));
wire t0_0011011010100, t0_0011011010101;
mixer mix_t0_001101101011 (.a(t0_0011011010110), .b(t0_0011011010111), .y(t0_001101101011));
wire t0_0011011010110, t0_0011011010111;
mixer mix_t0_0011011011 (.a(t0_00110110110), .b(t0_00110110111), .y(t0_0011011011));
wire t0_00110110110, t0_00110110111;
mixer mix_t0_00110110110 (.a(t0_001101101100), .b(t0_001101101101), .y(t0_00110110110));
wire t0_001101101100, t0_001101101101;
mixer mix_t0_001101101100 (.a(t0_0011011011000), .b(t0_0011011011001), .y(t0_001101101100));
wire t0_0011011011000, t0_0011011011001;
mixer mix_t0_001101101101 (.a(t0_0011011011010), .b(t0_0011011011011), .y(t0_001101101101));
wire t0_0011011011010, t0_0011011011011;
mixer mix_t0_00110110111 (.a(t0_001101101110), .b(t0_001101101111), .y(t0_00110110111));
wire t0_001101101110, t0_001101101111;
mixer mix_t0_001101101110 (.a(t0_0011011011100), .b(t0_0011011011101), .y(t0_001101101110));
wire t0_0011011011100, t0_0011011011101;
mixer mix_t0_001101101111 (.a(t0_0011011011110), .b(t0_0011011011111), .y(t0_001101101111));
wire t0_0011011011110, t0_0011011011111;
mixer mix_t0_00110111 (.a(t0_001101110), .b(t0_001101111), .y(t0_00110111));
wire t0_001101110, t0_001101111;
mixer mix_t0_001101110 (.a(t0_0011011100), .b(t0_0011011101), .y(t0_001101110));
wire t0_0011011100, t0_0011011101;
mixer mix_t0_0011011100 (.a(t0_00110111000), .b(t0_00110111001), .y(t0_0011011100));
wire t0_00110111000, t0_00110111001;
mixer mix_t0_00110111000 (.a(t0_001101110000), .b(t0_001101110001), .y(t0_00110111000));
wire t0_001101110000, t0_001101110001;
mixer mix_t0_001101110000 (.a(t0_0011011100000), .b(t0_0011011100001), .y(t0_001101110000));
wire t0_0011011100000, t0_0011011100001;
mixer mix_t0_001101110001 (.a(t0_0011011100010), .b(t0_0011011100011), .y(t0_001101110001));
wire t0_0011011100010, t0_0011011100011;
mixer mix_t0_00110111001 (.a(t0_001101110010), .b(t0_001101110011), .y(t0_00110111001));
wire t0_001101110010, t0_001101110011;
mixer mix_t0_001101110010 (.a(t0_0011011100100), .b(t0_0011011100101), .y(t0_001101110010));
wire t0_0011011100100, t0_0011011100101;
mixer mix_t0_001101110011 (.a(t0_0011011100110), .b(t0_0011011100111), .y(t0_001101110011));
wire t0_0011011100110, t0_0011011100111;
mixer mix_t0_0011011101 (.a(t0_00110111010), .b(t0_00110111011), .y(t0_0011011101));
wire t0_00110111010, t0_00110111011;
mixer mix_t0_00110111010 (.a(t0_001101110100), .b(t0_001101110101), .y(t0_00110111010));
wire t0_001101110100, t0_001101110101;
mixer mix_t0_001101110100 (.a(t0_0011011101000), .b(t0_0011011101001), .y(t0_001101110100));
wire t0_0011011101000, t0_0011011101001;
mixer mix_t0_001101110101 (.a(t0_0011011101010), .b(t0_0011011101011), .y(t0_001101110101));
wire t0_0011011101010, t0_0011011101011;
mixer mix_t0_00110111011 (.a(t0_001101110110), .b(t0_001101110111), .y(t0_00110111011));
wire t0_001101110110, t0_001101110111;
mixer mix_t0_001101110110 (.a(t0_0011011101100), .b(t0_0011011101101), .y(t0_001101110110));
wire t0_0011011101100, t0_0011011101101;
mixer mix_t0_001101110111 (.a(t0_0011011101110), .b(t0_0011011101111), .y(t0_001101110111));
wire t0_0011011101110, t0_0011011101111;
mixer mix_t0_001101111 (.a(t0_0011011110), .b(t0_0011011111), .y(t0_001101111));
wire t0_0011011110, t0_0011011111;
mixer mix_t0_0011011110 (.a(t0_00110111100), .b(t0_00110111101), .y(t0_0011011110));
wire t0_00110111100, t0_00110111101;
mixer mix_t0_00110111100 (.a(t0_001101111000), .b(t0_001101111001), .y(t0_00110111100));
wire t0_001101111000, t0_001101111001;
mixer mix_t0_001101111000 (.a(t0_0011011110000), .b(t0_0011011110001), .y(t0_001101111000));
wire t0_0011011110000, t0_0011011110001;
mixer mix_t0_001101111001 (.a(t0_0011011110010), .b(t0_0011011110011), .y(t0_001101111001));
wire t0_0011011110010, t0_0011011110011;
mixer mix_t0_00110111101 (.a(t0_001101111010), .b(t0_001101111011), .y(t0_00110111101));
wire t0_001101111010, t0_001101111011;
mixer mix_t0_001101111010 (.a(t0_0011011110100), .b(t0_0011011110101), .y(t0_001101111010));
wire t0_0011011110100, t0_0011011110101;
mixer mix_t0_001101111011 (.a(t0_0011011110110), .b(t0_0011011110111), .y(t0_001101111011));
wire t0_0011011110110, t0_0011011110111;
mixer mix_t0_0011011111 (.a(t0_00110111110), .b(t0_00110111111), .y(t0_0011011111));
wire t0_00110111110, t0_00110111111;
mixer mix_t0_00110111110 (.a(t0_001101111100), .b(t0_001101111101), .y(t0_00110111110));
wire t0_001101111100, t0_001101111101;
mixer mix_t0_001101111100 (.a(t0_0011011111000), .b(t0_0011011111001), .y(t0_001101111100));
wire t0_0011011111000, t0_0011011111001;
mixer mix_t0_001101111101 (.a(t0_0011011111010), .b(t0_0011011111011), .y(t0_001101111101));
wire t0_0011011111010, t0_0011011111011;
mixer mix_t0_00110111111 (.a(t0_001101111110), .b(t0_001101111111), .y(t0_00110111111));
wire t0_001101111110, t0_001101111111;
mixer mix_t0_001101111110 (.a(t0_0011011111100), .b(t0_0011011111101), .y(t0_001101111110));
wire t0_0011011111100, t0_0011011111101;
mixer mix_t0_001101111111 (.a(t0_0011011111110), .b(t0_0011011111111), .y(t0_001101111111));
wire t0_0011011111110, t0_0011011111111;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_001110 (.a(t0_0011100), .b(t0_0011101), .y(t0_001110));
wire t0_0011100, t0_0011101;
mixer mix_t0_0011100 (.a(t0_00111000), .b(t0_00111001), .y(t0_0011100));
wire t0_00111000, t0_00111001;
mixer mix_t0_00111000 (.a(t0_001110000), .b(t0_001110001), .y(t0_00111000));
wire t0_001110000, t0_001110001;
mixer mix_t0_001110000 (.a(t0_0011100000), .b(t0_0011100001), .y(t0_001110000));
wire t0_0011100000, t0_0011100001;
mixer mix_t0_0011100000 (.a(t0_00111000000), .b(t0_00111000001), .y(t0_0011100000));
wire t0_00111000000, t0_00111000001;
mixer mix_t0_00111000000 (.a(t0_001110000000), .b(t0_001110000001), .y(t0_00111000000));
wire t0_001110000000, t0_001110000001;
mixer mix_t0_001110000000 (.a(t0_0011100000000), .b(t0_0011100000001), .y(t0_001110000000));
wire t0_0011100000000, t0_0011100000001;
mixer mix_t0_001110000001 (.a(t0_0011100000010), .b(t0_0011100000011), .y(t0_001110000001));
wire t0_0011100000010, t0_0011100000011;
mixer mix_t0_00111000001 (.a(t0_001110000010), .b(t0_001110000011), .y(t0_00111000001));
wire t0_001110000010, t0_001110000011;
mixer mix_t0_001110000010 (.a(t0_0011100000100), .b(t0_0011100000101), .y(t0_001110000010));
wire t0_0011100000100, t0_0011100000101;
mixer mix_t0_001110000011 (.a(t0_0011100000110), .b(t0_0011100000111), .y(t0_001110000011));
wire t0_0011100000110, t0_0011100000111;
mixer mix_t0_0011100001 (.a(t0_00111000010), .b(t0_00111000011), .y(t0_0011100001));
wire t0_00111000010, t0_00111000011;
mixer mix_t0_00111000010 (.a(t0_001110000100), .b(t0_001110000101), .y(t0_00111000010));
wire t0_001110000100, t0_001110000101;
mixer mix_t0_001110000100 (.a(t0_0011100001000), .b(t0_0011100001001), .y(t0_001110000100));
wire t0_0011100001000, t0_0011100001001;
mixer mix_t0_001110000101 (.a(t0_0011100001010), .b(t0_0011100001011), .y(t0_001110000101));
wire t0_0011100001010, t0_0011100001011;
mixer mix_t0_00111000011 (.a(t0_001110000110), .b(t0_001110000111), .y(t0_00111000011));
wire t0_001110000110, t0_001110000111;
mixer mix_t0_001110000110 (.a(t0_0011100001100), .b(t0_0011100001101), .y(t0_001110000110));
wire t0_0011100001100, t0_0011100001101;
mixer mix_t0_001110000111 (.a(t0_0011100001110), .b(t0_0011100001111), .y(t0_001110000111));
wire t0_0011100001110, t0_0011100001111;
mixer mix_t0_001110001 (.a(t0_0011100010), .b(t0_0011100011), .y(t0_001110001));
wire t0_0011100010, t0_0011100011;
mixer mix_t0_0011100010 (.a(t0_00111000100), .b(t0_00111000101), .y(t0_0011100010));
wire t0_00111000100, t0_00111000101;
mixer mix_t0_00111000100 (.a(t0_001110001000), .b(t0_001110001001), .y(t0_00111000100));
wire t0_001110001000, t0_001110001001;
mixer mix_t0_001110001000 (.a(t0_0011100010000), .b(t0_0011100010001), .y(t0_001110001000));
wire t0_0011100010000, t0_0011100010001;
mixer mix_t0_001110001001 (.a(t0_0011100010010), .b(t0_0011100010011), .y(t0_001110001001));
wire t0_0011100010010, t0_0011100010011;
mixer mix_t0_00111000101 (.a(t0_001110001010), .b(t0_001110001011), .y(t0_00111000101));
wire t0_001110001010, t0_001110001011;
mixer mix_t0_001110001010 (.a(t0_0011100010100), .b(t0_0011100010101), .y(t0_001110001010));
wire t0_0011100010100, t0_0011100010101;
mixer mix_t0_001110001011 (.a(t0_0011100010110), .b(t0_0011100010111), .y(t0_001110001011));
wire t0_0011100010110, t0_0011100010111;
mixer mix_t0_0011100011 (.a(t0_00111000110), .b(t0_00111000111), .y(t0_0011100011));
wire t0_00111000110, t0_00111000111;
mixer mix_t0_00111000110 (.a(t0_001110001100), .b(t0_001110001101), .y(t0_00111000110));
wire t0_001110001100, t0_001110001101;
mixer mix_t0_001110001100 (.a(t0_0011100011000), .b(t0_0011100011001), .y(t0_001110001100));
wire t0_0011100011000, t0_0011100011001;
mixer mix_t0_001110001101 (.a(t0_0011100011010), .b(t0_0011100011011), .y(t0_001110001101));
wire t0_0011100011010, t0_0011100011011;
mixer mix_t0_00111000111 (.a(t0_001110001110), .b(t0_001110001111), .y(t0_00111000111));
wire t0_001110001110, t0_001110001111;
mixer mix_t0_001110001110 (.a(t0_0011100011100), .b(t0_0011100011101), .y(t0_001110001110));
wire t0_0011100011100, t0_0011100011101;
mixer mix_t0_001110001111 (.a(t0_0011100011110), .b(t0_0011100011111), .y(t0_001110001111));
wire t0_0011100011110, t0_0011100011111;
mixer mix_t0_00111001 (.a(t0_001110010), .b(t0_001110011), .y(t0_00111001));
wire t0_001110010, t0_001110011;
mixer mix_t0_001110010 (.a(t0_0011100100), .b(t0_0011100101), .y(t0_001110010));
wire t0_0011100100, t0_0011100101;
mixer mix_t0_0011100100 (.a(t0_00111001000), .b(t0_00111001001), .y(t0_0011100100));
wire t0_00111001000, t0_00111001001;
mixer mix_t0_00111001000 (.a(t0_001110010000), .b(t0_001110010001), .y(t0_00111001000));
wire t0_001110010000, t0_001110010001;
mixer mix_t0_001110010000 (.a(t0_0011100100000), .b(t0_0011100100001), .y(t0_001110010000));
wire t0_0011100100000, t0_0011100100001;
mixer mix_t0_001110010001 (.a(t0_0011100100010), .b(t0_0011100100011), .y(t0_001110010001));
wire t0_0011100100010, t0_0011100100011;
mixer mix_t0_00111001001 (.a(t0_001110010010), .b(t0_001110010011), .y(t0_00111001001));
wire t0_001110010010, t0_001110010011;
mixer mix_t0_001110010010 (.a(t0_0011100100100), .b(t0_0011100100101), .y(t0_001110010010));
wire t0_0011100100100, t0_0011100100101;
mixer mix_t0_001110010011 (.a(t0_0011100100110), .b(t0_0011100100111), .y(t0_001110010011));
wire t0_0011100100110, t0_0011100100111;
mixer mix_t0_0011100101 (.a(t0_00111001010), .b(t0_00111001011), .y(t0_0011100101));
wire t0_00111001010, t0_00111001011;
mixer mix_t0_00111001010 (.a(t0_001110010100), .b(t0_001110010101), .y(t0_00111001010));
wire t0_001110010100, t0_001110010101;
mixer mix_t0_001110010100 (.a(t0_0011100101000), .b(t0_0011100101001), .y(t0_001110010100));
wire t0_0011100101000, t0_0011100101001;
mixer mix_t0_001110010101 (.a(t0_0011100101010), .b(t0_0011100101011), .y(t0_001110010101));
wire t0_0011100101010, t0_0011100101011;
mixer mix_t0_00111001011 (.a(t0_001110010110), .b(t0_001110010111), .y(t0_00111001011));
wire t0_001110010110, t0_001110010111;
mixer mix_t0_001110010110 (.a(t0_0011100101100), .b(t0_0011100101101), .y(t0_001110010110));
wire t0_0011100101100, t0_0011100101101;
mixer mix_t0_001110010111 (.a(t0_0011100101110), .b(t0_0011100101111), .y(t0_001110010111));
wire t0_0011100101110, t0_0011100101111;
mixer mix_t0_001110011 (.a(t0_0011100110), .b(t0_0011100111), .y(t0_001110011));
wire t0_0011100110, t0_0011100111;
mixer mix_t0_0011100110 (.a(t0_00111001100), .b(t0_00111001101), .y(t0_0011100110));
wire t0_00111001100, t0_00111001101;
mixer mix_t0_00111001100 (.a(t0_001110011000), .b(t0_001110011001), .y(t0_00111001100));
wire t0_001110011000, t0_001110011001;
mixer mix_t0_001110011000 (.a(t0_0011100110000), .b(t0_0011100110001), .y(t0_001110011000));
wire t0_0011100110000, t0_0011100110001;
mixer mix_t0_001110011001 (.a(t0_0011100110010), .b(t0_0011100110011), .y(t0_001110011001));
wire t0_0011100110010, t0_0011100110011;
mixer mix_t0_00111001101 (.a(t0_001110011010), .b(t0_001110011011), .y(t0_00111001101));
wire t0_001110011010, t0_001110011011;
mixer mix_t0_001110011010 (.a(t0_0011100110100), .b(t0_0011100110101), .y(t0_001110011010));
wire t0_0011100110100, t0_0011100110101;
mixer mix_t0_001110011011 (.a(t0_0011100110110), .b(t0_0011100110111), .y(t0_001110011011));
wire t0_0011100110110, t0_0011100110111;
mixer mix_t0_0011100111 (.a(t0_00111001110), .b(t0_00111001111), .y(t0_0011100111));
wire t0_00111001110, t0_00111001111;
mixer mix_t0_00111001110 (.a(t0_001110011100), .b(t0_001110011101), .y(t0_00111001110));
wire t0_001110011100, t0_001110011101;
mixer mix_t0_001110011100 (.a(t0_0011100111000), .b(t0_0011100111001), .y(t0_001110011100));
wire t0_0011100111000, t0_0011100111001;
mixer mix_t0_001110011101 (.a(t0_0011100111010), .b(t0_0011100111011), .y(t0_001110011101));
wire t0_0011100111010, t0_0011100111011;
mixer mix_t0_00111001111 (.a(t0_001110011110), .b(t0_001110011111), .y(t0_00111001111));
wire t0_001110011110, t0_001110011111;
mixer mix_t0_001110011110 (.a(t0_0011100111100), .b(t0_0011100111101), .y(t0_001110011110));
wire t0_0011100111100, t0_0011100111101;
mixer mix_t0_001110011111 (.a(t0_0011100111110), .b(t0_0011100111111), .y(t0_001110011111));
wire t0_0011100111110, t0_0011100111111;
mixer mix_t0_0011101 (.a(t0_00111010), .b(t0_00111011), .y(t0_0011101));
wire t0_00111010, t0_00111011;
mixer mix_t0_00111010 (.a(t0_001110100), .b(t0_001110101), .y(t0_00111010));
wire t0_001110100, t0_001110101;
mixer mix_t0_001110100 (.a(t0_0011101000), .b(t0_0011101001), .y(t0_001110100));
wire t0_0011101000, t0_0011101001;
mixer mix_t0_0011101000 (.a(t0_00111010000), .b(t0_00111010001), .y(t0_0011101000));
wire t0_00111010000, t0_00111010001;
mixer mix_t0_00111010000 (.a(t0_001110100000), .b(t0_001110100001), .y(t0_00111010000));
wire t0_001110100000, t0_001110100001;
mixer mix_t0_001110100000 (.a(t0_0011101000000), .b(t0_0011101000001), .y(t0_001110100000));
wire t0_0011101000000, t0_0011101000001;
mixer mix_t0_001110100001 (.a(t0_0011101000010), .b(t0_0011101000011), .y(t0_001110100001));
wire t0_0011101000010, t0_0011101000011;
mixer mix_t0_00111010001 (.a(t0_001110100010), .b(t0_001110100011), .y(t0_00111010001));
wire t0_001110100010, t0_001110100011;
mixer mix_t0_001110100010 (.a(t0_0011101000100), .b(t0_0011101000101), .y(t0_001110100010));
wire t0_0011101000100, t0_0011101000101;
mixer mix_t0_001110100011 (.a(t0_0011101000110), .b(t0_0011101000111), .y(t0_001110100011));
wire t0_0011101000110, t0_0011101000111;
mixer mix_t0_0011101001 (.a(t0_00111010010), .b(t0_00111010011), .y(t0_0011101001));
wire t0_00111010010, t0_00111010011;
mixer mix_t0_00111010010 (.a(t0_001110100100), .b(t0_001110100101), .y(t0_00111010010));
wire t0_001110100100, t0_001110100101;
mixer mix_t0_001110100100 (.a(t0_0011101001000), .b(t0_0011101001001), .y(t0_001110100100));
wire t0_0011101001000, t0_0011101001001;
mixer mix_t0_001110100101 (.a(t0_0011101001010), .b(t0_0011101001011), .y(t0_001110100101));
wire t0_0011101001010, t0_0011101001011;
mixer mix_t0_00111010011 (.a(t0_001110100110), .b(t0_001110100111), .y(t0_00111010011));
wire t0_001110100110, t0_001110100111;
mixer mix_t0_001110100110 (.a(t0_0011101001100), .b(t0_0011101001101), .y(t0_001110100110));
wire t0_0011101001100, t0_0011101001101;
mixer mix_t0_001110100111 (.a(t0_0011101001110), .b(t0_0011101001111), .y(t0_001110100111));
wire t0_0011101001110, t0_0011101001111;
mixer mix_t0_001110101 (.a(t0_0011101010), .b(t0_0011101011), .y(t0_001110101));
wire t0_0011101010, t0_0011101011;
mixer mix_t0_0011101010 (.a(t0_00111010100), .b(t0_00111010101), .y(t0_0011101010));
wire t0_00111010100, t0_00111010101;
mixer mix_t0_00111010100 (.a(t0_001110101000), .b(t0_001110101001), .y(t0_00111010100));
wire t0_001110101000, t0_001110101001;
mixer mix_t0_001110101000 (.a(t0_0011101010000), .b(t0_0011101010001), .y(t0_001110101000));
wire t0_0011101010000, t0_0011101010001;
mixer mix_t0_001110101001 (.a(t0_0011101010010), .b(t0_0011101010011), .y(t0_001110101001));
wire t0_0011101010010, t0_0011101010011;
mixer mix_t0_00111010101 (.a(t0_001110101010), .b(t0_001110101011), .y(t0_00111010101));
wire t0_001110101010, t0_001110101011;
mixer mix_t0_001110101010 (.a(t0_0011101010100), .b(t0_0011101010101), .y(t0_001110101010));
wire t0_0011101010100, t0_0011101010101;
mixer mix_t0_001110101011 (.a(t0_0011101010110), .b(t0_0011101010111), .y(t0_001110101011));
wire t0_0011101010110, t0_0011101010111;
mixer mix_t0_0011101011 (.a(t0_00111010110), .b(t0_00111010111), .y(t0_0011101011));
wire t0_00111010110, t0_00111010111;
mixer mix_t0_00111010110 (.a(t0_001110101100), .b(t0_001110101101), .y(t0_00111010110));
wire t0_001110101100, t0_001110101101;
mixer mix_t0_001110101100 (.a(t0_0011101011000), .b(t0_0011101011001), .y(t0_001110101100));
wire t0_0011101011000, t0_0011101011001;
mixer mix_t0_001110101101 (.a(t0_0011101011010), .b(t0_0011101011011), .y(t0_001110101101));
wire t0_0011101011010, t0_0011101011011;
mixer mix_t0_00111010111 (.a(t0_001110101110), .b(t0_001110101111), .y(t0_00111010111));
wire t0_001110101110, t0_001110101111;
mixer mix_t0_001110101110 (.a(t0_0011101011100), .b(t0_0011101011101), .y(t0_001110101110));
wire t0_0011101011100, t0_0011101011101;
mixer mix_t0_001110101111 (.a(t0_0011101011110), .b(t0_0011101011111), .y(t0_001110101111));
wire t0_0011101011110, t0_0011101011111;
mixer mix_t0_00111011 (.a(t0_001110110), .b(t0_001110111), .y(t0_00111011));
wire t0_001110110, t0_001110111;
mixer mix_t0_001110110 (.a(t0_0011101100), .b(t0_0011101101), .y(t0_001110110));
wire t0_0011101100, t0_0011101101;
mixer mix_t0_0011101100 (.a(t0_00111011000), .b(t0_00111011001), .y(t0_0011101100));
wire t0_00111011000, t0_00111011001;
mixer mix_t0_00111011000 (.a(t0_001110110000), .b(t0_001110110001), .y(t0_00111011000));
wire t0_001110110000, t0_001110110001;
mixer mix_t0_001110110000 (.a(t0_0011101100000), .b(t0_0011101100001), .y(t0_001110110000));
wire t0_0011101100000, t0_0011101100001;
mixer mix_t0_001110110001 (.a(t0_0011101100010), .b(t0_0011101100011), .y(t0_001110110001));
wire t0_0011101100010, t0_0011101100011;
mixer mix_t0_00111011001 (.a(t0_001110110010), .b(t0_001110110011), .y(t0_00111011001));
wire t0_001110110010, t0_001110110011;
mixer mix_t0_001110110010 (.a(t0_0011101100100), .b(t0_0011101100101), .y(t0_001110110010));
wire t0_0011101100100, t0_0011101100101;
mixer mix_t0_001110110011 (.a(t0_0011101100110), .b(t0_0011101100111), .y(t0_001110110011));
wire t0_0011101100110, t0_0011101100111;
mixer mix_t0_0011101101 (.a(t0_00111011010), .b(t0_00111011011), .y(t0_0011101101));
wire t0_00111011010, t0_00111011011;
mixer mix_t0_00111011010 (.a(t0_001110110100), .b(t0_001110110101), .y(t0_00111011010));
wire t0_001110110100, t0_001110110101;
mixer mix_t0_001110110100 (.a(t0_0011101101000), .b(t0_0011101101001), .y(t0_001110110100));
wire t0_0011101101000, t0_0011101101001;
mixer mix_t0_001110110101 (.a(t0_0011101101010), .b(t0_0011101101011), .y(t0_001110110101));
wire t0_0011101101010, t0_0011101101011;
mixer mix_t0_00111011011 (.a(t0_001110110110), .b(t0_001110110111), .y(t0_00111011011));
wire t0_001110110110, t0_001110110111;
mixer mix_t0_001110110110 (.a(t0_0011101101100), .b(t0_0011101101101), .y(t0_001110110110));
wire t0_0011101101100, t0_0011101101101;
mixer mix_t0_001110110111 (.a(t0_0011101101110), .b(t0_0011101101111), .y(t0_001110110111));
wire t0_0011101101110, t0_0011101101111;
mixer mix_t0_001110111 (.a(t0_0011101110), .b(t0_0011101111), .y(t0_001110111));
wire t0_0011101110, t0_0011101111;
mixer mix_t0_0011101110 (.a(t0_00111011100), .b(t0_00111011101), .y(t0_0011101110));
wire t0_00111011100, t0_00111011101;
mixer mix_t0_00111011100 (.a(t0_001110111000), .b(t0_001110111001), .y(t0_00111011100));
wire t0_001110111000, t0_001110111001;
mixer mix_t0_001110111000 (.a(t0_0011101110000), .b(t0_0011101110001), .y(t0_001110111000));
wire t0_0011101110000, t0_0011101110001;
mixer mix_t0_001110111001 (.a(t0_0011101110010), .b(t0_0011101110011), .y(t0_001110111001));
wire t0_0011101110010, t0_0011101110011;
mixer mix_t0_00111011101 (.a(t0_001110111010), .b(t0_001110111011), .y(t0_00111011101));
wire t0_001110111010, t0_001110111011;
mixer mix_t0_001110111010 (.a(t0_0011101110100), .b(t0_0011101110101), .y(t0_001110111010));
wire t0_0011101110100, t0_0011101110101;
mixer mix_t0_001110111011 (.a(t0_0011101110110), .b(t0_0011101110111), .y(t0_001110111011));
wire t0_0011101110110, t0_0011101110111;
mixer mix_t0_0011101111 (.a(t0_00111011110), .b(t0_00111011111), .y(t0_0011101111));
wire t0_00111011110, t0_00111011111;
mixer mix_t0_00111011110 (.a(t0_001110111100), .b(t0_001110111101), .y(t0_00111011110));
wire t0_001110111100, t0_001110111101;
mixer mix_t0_001110111100 (.a(t0_0011101111000), .b(t0_0011101111001), .y(t0_001110111100));
wire t0_0011101111000, t0_0011101111001;
mixer mix_t0_001110111101 (.a(t0_0011101111010), .b(t0_0011101111011), .y(t0_001110111101));
wire t0_0011101111010, t0_0011101111011;
mixer mix_t0_00111011111 (.a(t0_001110111110), .b(t0_001110111111), .y(t0_00111011111));
wire t0_001110111110, t0_001110111111;
mixer mix_t0_001110111110 (.a(t0_0011101111100), .b(t0_0011101111101), .y(t0_001110111110));
wire t0_0011101111100, t0_0011101111101;
mixer mix_t0_001110111111 (.a(t0_0011101111110), .b(t0_0011101111111), .y(t0_001110111111));
wire t0_0011101111110, t0_0011101111111;
mixer mix_t0_001111 (.a(t0_0011110), .b(t0_0011111), .y(t0_001111));
wire t0_0011110, t0_0011111;
mixer mix_t0_0011110 (.a(t0_00111100), .b(t0_00111101), .y(t0_0011110));
wire t0_00111100, t0_00111101;
mixer mix_t0_00111100 (.a(t0_001111000), .b(t0_001111001), .y(t0_00111100));
wire t0_001111000, t0_001111001;
mixer mix_t0_001111000 (.a(t0_0011110000), .b(t0_0011110001), .y(t0_001111000));
wire t0_0011110000, t0_0011110001;
mixer mix_t0_0011110000 (.a(t0_00111100000), .b(t0_00111100001), .y(t0_0011110000));
wire t0_00111100000, t0_00111100001;
mixer mix_t0_00111100000 (.a(t0_001111000000), .b(t0_001111000001), .y(t0_00111100000));
wire t0_001111000000, t0_001111000001;
mixer mix_t0_001111000000 (.a(t0_0011110000000), .b(t0_0011110000001), .y(t0_001111000000));
wire t0_0011110000000, t0_0011110000001;
mixer mix_t0_001111000001 (.a(t0_0011110000010), .b(t0_0011110000011), .y(t0_001111000001));
wire t0_0011110000010, t0_0011110000011;
mixer mix_t0_00111100001 (.a(t0_001111000010), .b(t0_001111000011), .y(t0_00111100001));
wire t0_001111000010, t0_001111000011;
mixer mix_t0_001111000010 (.a(t0_0011110000100), .b(t0_0011110000101), .y(t0_001111000010));
wire t0_0011110000100, t0_0011110000101;
mixer mix_t0_001111000011 (.a(t0_0011110000110), .b(t0_0011110000111), .y(t0_001111000011));
wire t0_0011110000110, t0_0011110000111;
mixer mix_t0_0011110001 (.a(t0_00111100010), .b(t0_00111100011), .y(t0_0011110001));
wire t0_00111100010, t0_00111100011;
mixer mix_t0_00111100010 (.a(t0_001111000100), .b(t0_001111000101), .y(t0_00111100010));
wire t0_001111000100, t0_001111000101;
mixer mix_t0_001111000100 (.a(t0_0011110001000), .b(t0_0011110001001), .y(t0_001111000100));
wire t0_0011110001000, t0_0011110001001;
mixer mix_t0_001111000101 (.a(t0_0011110001010), .b(t0_0011110001011), .y(t0_001111000101));
wire t0_0011110001010, t0_0011110001011;
mixer mix_t0_00111100011 (.a(t0_001111000110), .b(t0_001111000111), .y(t0_00111100011));
wire t0_001111000110, t0_001111000111;
mixer mix_t0_001111000110 (.a(t0_0011110001100), .b(t0_0011110001101), .y(t0_001111000110));
wire t0_0011110001100, t0_0011110001101;
mixer mix_t0_001111000111 (.a(t0_0011110001110), .b(t0_0011110001111), .y(t0_001111000111));
wire t0_0011110001110, t0_0011110001111;
mixer mix_t0_001111001 (.a(t0_0011110010), .b(t0_0011110011), .y(t0_001111001));
wire t0_0011110010, t0_0011110011;
mixer mix_t0_0011110010 (.a(t0_00111100100), .b(t0_00111100101), .y(t0_0011110010));
wire t0_00111100100, t0_00111100101;
mixer mix_t0_00111100100 (.a(t0_001111001000), .b(t0_001111001001), .y(t0_00111100100));
wire t0_001111001000, t0_001111001001;
mixer mix_t0_001111001000 (.a(t0_0011110010000), .b(t0_0011110010001), .y(t0_001111001000));
wire t0_0011110010000, t0_0011110010001;
mixer mix_t0_001111001001 (.a(t0_0011110010010), .b(t0_0011110010011), .y(t0_001111001001));
wire t0_0011110010010, t0_0011110010011;
mixer mix_t0_00111100101 (.a(t0_001111001010), .b(t0_001111001011), .y(t0_00111100101));
wire t0_001111001010, t0_001111001011;
mixer mix_t0_001111001010 (.a(t0_0011110010100), .b(t0_0011110010101), .y(t0_001111001010));
wire t0_0011110010100, t0_0011110010101;
mixer mix_t0_001111001011 (.a(t0_0011110010110), .b(t0_0011110010111), .y(t0_001111001011));
wire t0_0011110010110, t0_0011110010111;
mixer mix_t0_0011110011 (.a(t0_00111100110), .b(t0_00111100111), .y(t0_0011110011));
wire t0_00111100110, t0_00111100111;
mixer mix_t0_00111100110 (.a(t0_001111001100), .b(t0_001111001101), .y(t0_00111100110));
wire t0_001111001100, t0_001111001101;
mixer mix_t0_001111001100 (.a(t0_0011110011000), .b(t0_0011110011001), .y(t0_001111001100));
wire t0_0011110011000, t0_0011110011001;
mixer mix_t0_001111001101 (.a(t0_0011110011010), .b(t0_0011110011011), .y(t0_001111001101));
wire t0_0011110011010, t0_0011110011011;
mixer mix_t0_00111100111 (.a(t0_001111001110), .b(t0_001111001111), .y(t0_00111100111));
wire t0_001111001110, t0_001111001111;
mixer mix_t0_001111001110 (.a(t0_0011110011100), .b(t0_0011110011101), .y(t0_001111001110));
wire t0_0011110011100, t0_0011110011101;
mixer mix_t0_001111001111 (.a(t0_0011110011110), .b(t0_0011110011111), .y(t0_001111001111));
wire t0_0011110011110, t0_0011110011111;
mixer mix_t0_00111101 (.a(t0_001111010), .b(t0_001111011), .y(t0_00111101));
wire t0_001111010, t0_001111011;
mixer mix_t0_001111010 (.a(t0_0011110100), .b(t0_0011110101), .y(t0_001111010));
wire t0_0011110100, t0_0011110101;
mixer mix_t0_0011110100 (.a(t0_00111101000), .b(t0_00111101001), .y(t0_0011110100));
wire t0_00111101000, t0_00111101001;
mixer mix_t0_00111101000 (.a(t0_001111010000), .b(t0_001111010001), .y(t0_00111101000));
wire t0_001111010000, t0_001111010001;
mixer mix_t0_001111010000 (.a(t0_0011110100000), .b(t0_0011110100001), .y(t0_001111010000));
wire t0_0011110100000, t0_0011110100001;
mixer mix_t0_001111010001 (.a(t0_0011110100010), .b(t0_0011110100011), .y(t0_001111010001));
wire t0_0011110100010, t0_0011110100011;
mixer mix_t0_00111101001 (.a(t0_001111010010), .b(t0_001111010011), .y(t0_00111101001));
wire t0_001111010010, t0_001111010011;
mixer mix_t0_001111010010 (.a(t0_0011110100100), .b(t0_0011110100101), .y(t0_001111010010));
wire t0_0011110100100, t0_0011110100101;
mixer mix_t0_001111010011 (.a(t0_0011110100110), .b(t0_0011110100111), .y(t0_001111010011));
wire t0_0011110100110, t0_0011110100111;
mixer mix_t0_0011110101 (.a(t0_00111101010), .b(t0_00111101011), .y(t0_0011110101));
wire t0_00111101010, t0_00111101011;
mixer mix_t0_00111101010 (.a(t0_001111010100), .b(t0_001111010101), .y(t0_00111101010));
wire t0_001111010100, t0_001111010101;
mixer mix_t0_001111010100 (.a(t0_0011110101000), .b(t0_0011110101001), .y(t0_001111010100));
wire t0_0011110101000, t0_0011110101001;
mixer mix_t0_001111010101 (.a(t0_0011110101010), .b(t0_0011110101011), .y(t0_001111010101));
wire t0_0011110101010, t0_0011110101011;
mixer mix_t0_00111101011 (.a(t0_001111010110), .b(t0_001111010111), .y(t0_00111101011));
wire t0_001111010110, t0_001111010111;
mixer mix_t0_001111010110 (.a(t0_0011110101100), .b(t0_0011110101101), .y(t0_001111010110));
wire t0_0011110101100, t0_0011110101101;
mixer mix_t0_001111010111 (.a(t0_0011110101110), .b(t0_0011110101111), .y(t0_001111010111));
wire t0_0011110101110, t0_0011110101111;
mixer mix_t0_001111011 (.a(t0_0011110110), .b(t0_0011110111), .y(t0_001111011));
wire t0_0011110110, t0_0011110111;
mixer mix_t0_0011110110 (.a(t0_00111101100), .b(t0_00111101101), .y(t0_0011110110));
wire t0_00111101100, t0_00111101101;
mixer mix_t0_00111101100 (.a(t0_001111011000), .b(t0_001111011001), .y(t0_00111101100));
wire t0_001111011000, t0_001111011001;
mixer mix_t0_001111011000 (.a(t0_0011110110000), .b(t0_0011110110001), .y(t0_001111011000));
wire t0_0011110110000, t0_0011110110001;
mixer mix_t0_001111011001 (.a(t0_0011110110010), .b(t0_0011110110011), .y(t0_001111011001));
wire t0_0011110110010, t0_0011110110011;
mixer mix_t0_00111101101 (.a(t0_001111011010), .b(t0_001111011011), .y(t0_00111101101));
wire t0_001111011010, t0_001111011011;
mixer mix_t0_001111011010 (.a(t0_0011110110100), .b(t0_0011110110101), .y(t0_001111011010));
wire t0_0011110110100, t0_0011110110101;
mixer mix_t0_001111011011 (.a(t0_0011110110110), .b(t0_0011110110111), .y(t0_001111011011));
wire t0_0011110110110, t0_0011110110111;
mixer mix_t0_0011110111 (.a(t0_00111101110), .b(t0_00111101111), .y(t0_0011110111));
wire t0_00111101110, t0_00111101111;
mixer mix_t0_00111101110 (.a(t0_001111011100), .b(t0_001111011101), .y(t0_00111101110));
wire t0_001111011100, t0_001111011101;
mixer mix_t0_001111011100 (.a(t0_0011110111000), .b(t0_0011110111001), .y(t0_001111011100));
wire t0_0011110111000, t0_0011110111001;
mixer mix_t0_001111011101 (.a(t0_0011110111010), .b(t0_0011110111011), .y(t0_001111011101));
wire t0_0011110111010, t0_0011110111011;
mixer mix_t0_00111101111 (.a(t0_001111011110), .b(t0_001111011111), .y(t0_00111101111));
wire t0_001111011110, t0_001111011111;
mixer mix_t0_001111011110 (.a(t0_0011110111100), .b(t0_0011110111101), .y(t0_001111011110));
wire t0_0011110111100, t0_0011110111101;
mixer mix_t0_001111011111 (.a(t0_0011110111110), .b(t0_0011110111111), .y(t0_001111011111));
wire t0_0011110111110, t0_0011110111111;
mixer mix_t0_0011111 (.a(t0_00111110), .b(t0_00111111), .y(t0_0011111));
wire t0_00111110, t0_00111111;
mixer mix_t0_00111110 (.a(t0_001111100), .b(t0_001111101), .y(t0_00111110));
wire t0_001111100, t0_001111101;
mixer mix_t0_001111100 (.a(t0_0011111000), .b(t0_0011111001), .y(t0_001111100));
wire t0_0011111000, t0_0011111001;
mixer mix_t0_0011111000 (.a(t0_00111110000), .b(t0_00111110001), .y(t0_0011111000));
wire t0_00111110000, t0_00111110001;
mixer mix_t0_00111110000 (.a(t0_001111100000), .b(t0_001111100001), .y(t0_00111110000));
wire t0_001111100000, t0_001111100001;
mixer mix_t0_001111100000 (.a(t0_0011111000000), .b(t0_0011111000001), .y(t0_001111100000));
wire t0_0011111000000, t0_0011111000001;
mixer mix_t0_001111100001 (.a(t0_0011111000010), .b(t0_0011111000011), .y(t0_001111100001));
wire t0_0011111000010, t0_0011111000011;
mixer mix_t0_00111110001 (.a(t0_001111100010), .b(t0_001111100011), .y(t0_00111110001));
wire t0_001111100010, t0_001111100011;
mixer mix_t0_001111100010 (.a(t0_0011111000100), .b(t0_0011111000101), .y(t0_001111100010));
wire t0_0011111000100, t0_0011111000101;
mixer mix_t0_001111100011 (.a(t0_0011111000110), .b(t0_0011111000111), .y(t0_001111100011));
wire t0_0011111000110, t0_0011111000111;
mixer mix_t0_0011111001 (.a(t0_00111110010), .b(t0_00111110011), .y(t0_0011111001));
wire t0_00111110010, t0_00111110011;
mixer mix_t0_00111110010 (.a(t0_001111100100), .b(t0_001111100101), .y(t0_00111110010));
wire t0_001111100100, t0_001111100101;
mixer mix_t0_001111100100 (.a(t0_0011111001000), .b(t0_0011111001001), .y(t0_001111100100));
wire t0_0011111001000, t0_0011111001001;
mixer mix_t0_001111100101 (.a(t0_0011111001010), .b(t0_0011111001011), .y(t0_001111100101));
wire t0_0011111001010, t0_0011111001011;
mixer mix_t0_00111110011 (.a(t0_001111100110), .b(t0_001111100111), .y(t0_00111110011));
wire t0_001111100110, t0_001111100111;
mixer mix_t0_001111100110 (.a(t0_0011111001100), .b(t0_0011111001101), .y(t0_001111100110));
wire t0_0011111001100, t0_0011111001101;
mixer mix_t0_001111100111 (.a(t0_0011111001110), .b(t0_0011111001111), .y(t0_001111100111));
wire t0_0011111001110, t0_0011111001111;
mixer mix_t0_001111101 (.a(t0_0011111010), .b(t0_0011111011), .y(t0_001111101));
wire t0_0011111010, t0_0011111011;
mixer mix_t0_0011111010 (.a(t0_00111110100), .b(t0_00111110101), .y(t0_0011111010));
wire t0_00111110100, t0_00111110101;
mixer mix_t0_00111110100 (.a(t0_001111101000), .b(t0_001111101001), .y(t0_00111110100));
wire t0_001111101000, t0_001111101001;
mixer mix_t0_001111101000 (.a(t0_0011111010000), .b(t0_0011111010001), .y(t0_001111101000));
wire t0_0011111010000, t0_0011111010001;
mixer mix_t0_001111101001 (.a(t0_0011111010010), .b(t0_0011111010011), .y(t0_001111101001));
wire t0_0011111010010, t0_0011111010011;
mixer mix_t0_00111110101 (.a(t0_001111101010), .b(t0_001111101011), .y(t0_00111110101));
wire t0_001111101010, t0_001111101011;
mixer mix_t0_001111101010 (.a(t0_0011111010100), .b(t0_0011111010101), .y(t0_001111101010));
wire t0_0011111010100, t0_0011111010101;
mixer mix_t0_001111101011 (.a(t0_0011111010110), .b(t0_0011111010111), .y(t0_001111101011));
wire t0_0011111010110, t0_0011111010111;
mixer mix_t0_0011111011 (.a(t0_00111110110), .b(t0_00111110111), .y(t0_0011111011));
wire t0_00111110110, t0_00111110111;
mixer mix_t0_00111110110 (.a(t0_001111101100), .b(t0_001111101101), .y(t0_00111110110));
wire t0_001111101100, t0_001111101101;
mixer mix_t0_001111101100 (.a(t0_0011111011000), .b(t0_0011111011001), .y(t0_001111101100));
wire t0_0011111011000, t0_0011111011001;
mixer mix_t0_001111101101 (.a(t0_0011111011010), .b(t0_0011111011011), .y(t0_001111101101));
wire t0_0011111011010, t0_0011111011011;
mixer mix_t0_00111110111 (.a(t0_001111101110), .b(t0_001111101111), .y(t0_00111110111));
wire t0_001111101110, t0_001111101111;
mixer mix_t0_001111101110 (.a(t0_0011111011100), .b(t0_0011111011101), .y(t0_001111101110));
wire t0_0011111011100, t0_0011111011101;
mixer mix_t0_001111101111 (.a(t0_0011111011110), .b(t0_0011111011111), .y(t0_001111101111));
wire t0_0011111011110, t0_0011111011111;
mixer mix_t0_00111111 (.a(t0_001111110), .b(t0_001111111), .y(t0_00111111));
wire t0_001111110, t0_001111111;
mixer mix_t0_001111110 (.a(t0_0011111100), .b(t0_0011111101), .y(t0_001111110));
wire t0_0011111100, t0_0011111101;
mixer mix_t0_0011111100 (.a(t0_00111111000), .b(t0_00111111001), .y(t0_0011111100));
wire t0_00111111000, t0_00111111001;
mixer mix_t0_00111111000 (.a(t0_001111110000), .b(t0_001111110001), .y(t0_00111111000));
wire t0_001111110000, t0_001111110001;
mixer mix_t0_001111110000 (.a(t0_0011111100000), .b(t0_0011111100001), .y(t0_001111110000));
wire t0_0011111100000, t0_0011111100001;
mixer mix_t0_001111110001 (.a(t0_0011111100010), .b(t0_0011111100011), .y(t0_001111110001));
wire t0_0011111100010, t0_0011111100011;
mixer mix_t0_00111111001 (.a(t0_001111110010), .b(t0_001111110011), .y(t0_00111111001));
wire t0_001111110010, t0_001111110011;
mixer mix_t0_001111110010 (.a(t0_0011111100100), .b(t0_0011111100101), .y(t0_001111110010));
wire t0_0011111100100, t0_0011111100101;
mixer mix_t0_001111110011 (.a(t0_0011111100110), .b(t0_0011111100111), .y(t0_001111110011));
wire t0_0011111100110, t0_0011111100111;
mixer mix_t0_0011111101 (.a(t0_00111111010), .b(t0_00111111011), .y(t0_0011111101));
wire t0_00111111010, t0_00111111011;
mixer mix_t0_00111111010 (.a(t0_001111110100), .b(t0_001111110101), .y(t0_00111111010));
wire t0_001111110100, t0_001111110101;
mixer mix_t0_001111110100 (.a(t0_0011111101000), .b(t0_0011111101001), .y(t0_001111110100));
wire t0_0011111101000, t0_0011111101001;
mixer mix_t0_001111110101 (.a(t0_0011111101010), .b(t0_0011111101011), .y(t0_001111110101));
wire t0_0011111101010, t0_0011111101011;
mixer mix_t0_00111111011 (.a(t0_001111110110), .b(t0_001111110111), .y(t0_00111111011));
wire t0_001111110110, t0_001111110111;
mixer mix_t0_001111110110 (.a(t0_0011111101100), .b(t0_0011111101101), .y(t0_001111110110));
wire t0_0011111101100, t0_0011111101101;
mixer mix_t0_001111110111 (.a(t0_0011111101110), .b(t0_0011111101111), .y(t0_001111110111));
wire t0_0011111101110, t0_0011111101111;
mixer mix_t0_001111111 (.a(t0_0011111110), .b(t0_0011111111), .y(t0_001111111));
wire t0_0011111110, t0_0011111111;
mixer mix_t0_0011111110 (.a(t0_00111111100), .b(t0_00111111101), .y(t0_0011111110));
wire t0_00111111100, t0_00111111101;
mixer mix_t0_00111111100 (.a(t0_001111111000), .b(t0_001111111001), .y(t0_00111111100));
wire t0_001111111000, t0_001111111001;
mixer mix_t0_001111111000 (.a(t0_0011111110000), .b(t0_0011111110001), .y(t0_001111111000));
wire t0_0011111110000, t0_0011111110001;
mixer mix_t0_001111111001 (.a(t0_0011111110010), .b(t0_0011111110011), .y(t0_001111111001));
wire t0_0011111110010, t0_0011111110011;
mixer mix_t0_00111111101 (.a(t0_001111111010), .b(t0_001111111011), .y(t0_00111111101));
wire t0_001111111010, t0_001111111011;
mixer mix_t0_001111111010 (.a(t0_0011111110100), .b(t0_0011111110101), .y(t0_001111111010));
wire t0_0011111110100, t0_0011111110101;
mixer mix_t0_001111111011 (.a(t0_0011111110110), .b(t0_0011111110111), .y(t0_001111111011));
wire t0_0011111110110, t0_0011111110111;
mixer mix_t0_0011111111 (.a(t0_00111111110), .b(t0_00111111111), .y(t0_0011111111));
wire t0_00111111110, t0_00111111111;
mixer mix_t0_00111111110 (.a(t0_001111111100), .b(t0_001111111101), .y(t0_00111111110));
wire t0_001111111100, t0_001111111101;
mixer mix_t0_001111111100 (.a(t0_0011111111000), .b(t0_0011111111001), .y(t0_001111111100));
wire t0_0011111111000, t0_0011111111001;
mixer mix_t0_001111111101 (.a(t0_0011111111010), .b(t0_0011111111011), .y(t0_001111111101));
wire t0_0011111111010, t0_0011111111011;
mixer mix_t0_00111111111 (.a(t0_001111111110), .b(t0_001111111111), .y(t0_00111111111));
wire t0_001111111110, t0_001111111111;
mixer mix_t0_001111111110 (.a(t0_0011111111100), .b(t0_0011111111101), .y(t0_001111111110));
wire t0_0011111111100, t0_0011111111101;
mixer mix_t0_001111111111 (.a(t0_0011111111110), .b(t0_0011111111111), .y(t0_001111111111));
wire t0_0011111111110, t0_0011111111111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_010000 (.a(t0_0100000), .b(t0_0100001), .y(t0_010000));
wire t0_0100000, t0_0100001;
mixer mix_t0_0100000 (.a(t0_01000000), .b(t0_01000001), .y(t0_0100000));
wire t0_01000000, t0_01000001;
mixer mix_t0_01000000 (.a(t0_010000000), .b(t0_010000001), .y(t0_01000000));
wire t0_010000000, t0_010000001;
mixer mix_t0_010000000 (.a(t0_0100000000), .b(t0_0100000001), .y(t0_010000000));
wire t0_0100000000, t0_0100000001;
mixer mix_t0_0100000000 (.a(t0_01000000000), .b(t0_01000000001), .y(t0_0100000000));
wire t0_01000000000, t0_01000000001;
mixer mix_t0_01000000000 (.a(t0_010000000000), .b(t0_010000000001), .y(t0_01000000000));
wire t0_010000000000, t0_010000000001;
mixer mix_t0_010000000000 (.a(t0_0100000000000), .b(t0_0100000000001), .y(t0_010000000000));
wire t0_0100000000000, t0_0100000000001;
mixer mix_t0_010000000001 (.a(t0_0100000000010), .b(t0_0100000000011), .y(t0_010000000001));
wire t0_0100000000010, t0_0100000000011;
mixer mix_t0_01000000001 (.a(t0_010000000010), .b(t0_010000000011), .y(t0_01000000001));
wire t0_010000000010, t0_010000000011;
mixer mix_t0_010000000010 (.a(t0_0100000000100), .b(t0_0100000000101), .y(t0_010000000010));
wire t0_0100000000100, t0_0100000000101;
mixer mix_t0_010000000011 (.a(t0_0100000000110), .b(t0_0100000000111), .y(t0_010000000011));
wire t0_0100000000110, t0_0100000000111;
mixer mix_t0_0100000001 (.a(t0_01000000010), .b(t0_01000000011), .y(t0_0100000001));
wire t0_01000000010, t0_01000000011;
mixer mix_t0_01000000010 (.a(t0_010000000100), .b(t0_010000000101), .y(t0_01000000010));
wire t0_010000000100, t0_010000000101;
mixer mix_t0_010000000100 (.a(t0_0100000001000), .b(t0_0100000001001), .y(t0_010000000100));
wire t0_0100000001000, t0_0100000001001;
mixer mix_t0_010000000101 (.a(t0_0100000001010), .b(t0_0100000001011), .y(t0_010000000101));
wire t0_0100000001010, t0_0100000001011;
mixer mix_t0_01000000011 (.a(t0_010000000110), .b(t0_010000000111), .y(t0_01000000011));
wire t0_010000000110, t0_010000000111;
mixer mix_t0_010000000110 (.a(t0_0100000001100), .b(t0_0100000001101), .y(t0_010000000110));
wire t0_0100000001100, t0_0100000001101;
mixer mix_t0_010000000111 (.a(t0_0100000001110), .b(t0_0100000001111), .y(t0_010000000111));
wire t0_0100000001110, t0_0100000001111;
mixer mix_t0_010000001 (.a(t0_0100000010), .b(t0_0100000011), .y(t0_010000001));
wire t0_0100000010, t0_0100000011;
mixer mix_t0_0100000010 (.a(t0_01000000100), .b(t0_01000000101), .y(t0_0100000010));
wire t0_01000000100, t0_01000000101;
mixer mix_t0_01000000100 (.a(t0_010000001000), .b(t0_010000001001), .y(t0_01000000100));
wire t0_010000001000, t0_010000001001;
mixer mix_t0_010000001000 (.a(t0_0100000010000), .b(t0_0100000010001), .y(t0_010000001000));
wire t0_0100000010000, t0_0100000010001;
mixer mix_t0_010000001001 (.a(t0_0100000010010), .b(t0_0100000010011), .y(t0_010000001001));
wire t0_0100000010010, t0_0100000010011;
mixer mix_t0_01000000101 (.a(t0_010000001010), .b(t0_010000001011), .y(t0_01000000101));
wire t0_010000001010, t0_010000001011;
mixer mix_t0_010000001010 (.a(t0_0100000010100), .b(t0_0100000010101), .y(t0_010000001010));
wire t0_0100000010100, t0_0100000010101;
mixer mix_t0_010000001011 (.a(t0_0100000010110), .b(t0_0100000010111), .y(t0_010000001011));
wire t0_0100000010110, t0_0100000010111;
mixer mix_t0_0100000011 (.a(t0_01000000110), .b(t0_01000000111), .y(t0_0100000011));
wire t0_01000000110, t0_01000000111;
mixer mix_t0_01000000110 (.a(t0_010000001100), .b(t0_010000001101), .y(t0_01000000110));
wire t0_010000001100, t0_010000001101;
mixer mix_t0_010000001100 (.a(t0_0100000011000), .b(t0_0100000011001), .y(t0_010000001100));
wire t0_0100000011000, t0_0100000011001;
mixer mix_t0_010000001101 (.a(t0_0100000011010), .b(t0_0100000011011), .y(t0_010000001101));
wire t0_0100000011010, t0_0100000011011;
mixer mix_t0_01000000111 (.a(t0_010000001110), .b(t0_010000001111), .y(t0_01000000111));
wire t0_010000001110, t0_010000001111;
mixer mix_t0_010000001110 (.a(t0_0100000011100), .b(t0_0100000011101), .y(t0_010000001110));
wire t0_0100000011100, t0_0100000011101;
mixer mix_t0_010000001111 (.a(t0_0100000011110), .b(t0_0100000011111), .y(t0_010000001111));
wire t0_0100000011110, t0_0100000011111;
mixer mix_t0_01000001 (.a(t0_010000010), .b(t0_010000011), .y(t0_01000001));
wire t0_010000010, t0_010000011;
mixer mix_t0_010000010 (.a(t0_0100000100), .b(t0_0100000101), .y(t0_010000010));
wire t0_0100000100, t0_0100000101;
mixer mix_t0_0100000100 (.a(t0_01000001000), .b(t0_01000001001), .y(t0_0100000100));
wire t0_01000001000, t0_01000001001;
mixer mix_t0_01000001000 (.a(t0_010000010000), .b(t0_010000010001), .y(t0_01000001000));
wire t0_010000010000, t0_010000010001;
mixer mix_t0_010000010000 (.a(t0_0100000100000), .b(t0_0100000100001), .y(t0_010000010000));
wire t0_0100000100000, t0_0100000100001;
mixer mix_t0_010000010001 (.a(t0_0100000100010), .b(t0_0100000100011), .y(t0_010000010001));
wire t0_0100000100010, t0_0100000100011;
mixer mix_t0_01000001001 (.a(t0_010000010010), .b(t0_010000010011), .y(t0_01000001001));
wire t0_010000010010, t0_010000010011;
mixer mix_t0_010000010010 (.a(t0_0100000100100), .b(t0_0100000100101), .y(t0_010000010010));
wire t0_0100000100100, t0_0100000100101;
mixer mix_t0_010000010011 (.a(t0_0100000100110), .b(t0_0100000100111), .y(t0_010000010011));
wire t0_0100000100110, t0_0100000100111;
mixer mix_t0_0100000101 (.a(t0_01000001010), .b(t0_01000001011), .y(t0_0100000101));
wire t0_01000001010, t0_01000001011;
mixer mix_t0_01000001010 (.a(t0_010000010100), .b(t0_010000010101), .y(t0_01000001010));
wire t0_010000010100, t0_010000010101;
mixer mix_t0_010000010100 (.a(t0_0100000101000), .b(t0_0100000101001), .y(t0_010000010100));
wire t0_0100000101000, t0_0100000101001;
mixer mix_t0_010000010101 (.a(t0_0100000101010), .b(t0_0100000101011), .y(t0_010000010101));
wire t0_0100000101010, t0_0100000101011;
mixer mix_t0_01000001011 (.a(t0_010000010110), .b(t0_010000010111), .y(t0_01000001011));
wire t0_010000010110, t0_010000010111;
mixer mix_t0_010000010110 (.a(t0_0100000101100), .b(t0_0100000101101), .y(t0_010000010110));
wire t0_0100000101100, t0_0100000101101;
mixer mix_t0_010000010111 (.a(t0_0100000101110), .b(t0_0100000101111), .y(t0_010000010111));
wire t0_0100000101110, t0_0100000101111;
mixer mix_t0_010000011 (.a(t0_0100000110), .b(t0_0100000111), .y(t0_010000011));
wire t0_0100000110, t0_0100000111;
mixer mix_t0_0100000110 (.a(t0_01000001100), .b(t0_01000001101), .y(t0_0100000110));
wire t0_01000001100, t0_01000001101;
mixer mix_t0_01000001100 (.a(t0_010000011000), .b(t0_010000011001), .y(t0_01000001100));
wire t0_010000011000, t0_010000011001;
mixer mix_t0_010000011000 (.a(t0_0100000110000), .b(t0_0100000110001), .y(t0_010000011000));
wire t0_0100000110000, t0_0100000110001;
mixer mix_t0_010000011001 (.a(t0_0100000110010), .b(t0_0100000110011), .y(t0_010000011001));
wire t0_0100000110010, t0_0100000110011;
mixer mix_t0_01000001101 (.a(t0_010000011010), .b(t0_010000011011), .y(t0_01000001101));
wire t0_010000011010, t0_010000011011;
mixer mix_t0_010000011010 (.a(t0_0100000110100), .b(t0_0100000110101), .y(t0_010000011010));
wire t0_0100000110100, t0_0100000110101;
mixer mix_t0_010000011011 (.a(t0_0100000110110), .b(t0_0100000110111), .y(t0_010000011011));
wire t0_0100000110110, t0_0100000110111;
mixer mix_t0_0100000111 (.a(t0_01000001110), .b(t0_01000001111), .y(t0_0100000111));
wire t0_01000001110, t0_01000001111;
mixer mix_t0_01000001110 (.a(t0_010000011100), .b(t0_010000011101), .y(t0_01000001110));
wire t0_010000011100, t0_010000011101;
mixer mix_t0_010000011100 (.a(t0_0100000111000), .b(t0_0100000111001), .y(t0_010000011100));
wire t0_0100000111000, t0_0100000111001;
mixer mix_t0_010000011101 (.a(t0_0100000111010), .b(t0_0100000111011), .y(t0_010000011101));
wire t0_0100000111010, t0_0100000111011;
mixer mix_t0_01000001111 (.a(t0_010000011110), .b(t0_010000011111), .y(t0_01000001111));
wire t0_010000011110, t0_010000011111;
mixer mix_t0_010000011110 (.a(t0_0100000111100), .b(t0_0100000111101), .y(t0_010000011110));
wire t0_0100000111100, t0_0100000111101;
mixer mix_t0_010000011111 (.a(t0_0100000111110), .b(t0_0100000111111), .y(t0_010000011111));
wire t0_0100000111110, t0_0100000111111;
mixer mix_t0_0100001 (.a(t0_01000010), .b(t0_01000011), .y(t0_0100001));
wire t0_01000010, t0_01000011;
mixer mix_t0_01000010 (.a(t0_010000100), .b(t0_010000101), .y(t0_01000010));
wire t0_010000100, t0_010000101;
mixer mix_t0_010000100 (.a(t0_0100001000), .b(t0_0100001001), .y(t0_010000100));
wire t0_0100001000, t0_0100001001;
mixer mix_t0_0100001000 (.a(t0_01000010000), .b(t0_01000010001), .y(t0_0100001000));
wire t0_01000010000, t0_01000010001;
mixer mix_t0_01000010000 (.a(t0_010000100000), .b(t0_010000100001), .y(t0_01000010000));
wire t0_010000100000, t0_010000100001;
mixer mix_t0_010000100000 (.a(t0_0100001000000), .b(t0_0100001000001), .y(t0_010000100000));
wire t0_0100001000000, t0_0100001000001;
mixer mix_t0_010000100001 (.a(t0_0100001000010), .b(t0_0100001000011), .y(t0_010000100001));
wire t0_0100001000010, t0_0100001000011;
mixer mix_t0_01000010001 (.a(t0_010000100010), .b(t0_010000100011), .y(t0_01000010001));
wire t0_010000100010, t0_010000100011;
mixer mix_t0_010000100010 (.a(t0_0100001000100), .b(t0_0100001000101), .y(t0_010000100010));
wire t0_0100001000100, t0_0100001000101;
mixer mix_t0_010000100011 (.a(t0_0100001000110), .b(t0_0100001000111), .y(t0_010000100011));
wire t0_0100001000110, t0_0100001000111;
mixer mix_t0_0100001001 (.a(t0_01000010010), .b(t0_01000010011), .y(t0_0100001001));
wire t0_01000010010, t0_01000010011;
mixer mix_t0_01000010010 (.a(t0_010000100100), .b(t0_010000100101), .y(t0_01000010010));
wire t0_010000100100, t0_010000100101;
mixer mix_t0_010000100100 (.a(t0_0100001001000), .b(t0_0100001001001), .y(t0_010000100100));
wire t0_0100001001000, t0_0100001001001;
mixer mix_t0_010000100101 (.a(t0_0100001001010), .b(t0_0100001001011), .y(t0_010000100101));
wire t0_0100001001010, t0_0100001001011;
mixer mix_t0_01000010011 (.a(t0_010000100110), .b(t0_010000100111), .y(t0_01000010011));
wire t0_010000100110, t0_010000100111;
mixer mix_t0_010000100110 (.a(t0_0100001001100), .b(t0_0100001001101), .y(t0_010000100110));
wire t0_0100001001100, t0_0100001001101;
mixer mix_t0_010000100111 (.a(t0_0100001001110), .b(t0_0100001001111), .y(t0_010000100111));
wire t0_0100001001110, t0_0100001001111;
mixer mix_t0_010000101 (.a(t0_0100001010), .b(t0_0100001011), .y(t0_010000101));
wire t0_0100001010, t0_0100001011;
mixer mix_t0_0100001010 (.a(t0_01000010100), .b(t0_01000010101), .y(t0_0100001010));
wire t0_01000010100, t0_01000010101;
mixer mix_t0_01000010100 (.a(t0_010000101000), .b(t0_010000101001), .y(t0_01000010100));
wire t0_010000101000, t0_010000101001;
mixer mix_t0_010000101000 (.a(t0_0100001010000), .b(t0_0100001010001), .y(t0_010000101000));
wire t0_0100001010000, t0_0100001010001;
mixer mix_t0_010000101001 (.a(t0_0100001010010), .b(t0_0100001010011), .y(t0_010000101001));
wire t0_0100001010010, t0_0100001010011;
mixer mix_t0_01000010101 (.a(t0_010000101010), .b(t0_010000101011), .y(t0_01000010101));
wire t0_010000101010, t0_010000101011;
mixer mix_t0_010000101010 (.a(t0_0100001010100), .b(t0_0100001010101), .y(t0_010000101010));
wire t0_0100001010100, t0_0100001010101;
mixer mix_t0_010000101011 (.a(t0_0100001010110), .b(t0_0100001010111), .y(t0_010000101011));
wire t0_0100001010110, t0_0100001010111;
mixer mix_t0_0100001011 (.a(t0_01000010110), .b(t0_01000010111), .y(t0_0100001011));
wire t0_01000010110, t0_01000010111;
mixer mix_t0_01000010110 (.a(t0_010000101100), .b(t0_010000101101), .y(t0_01000010110));
wire t0_010000101100, t0_010000101101;
mixer mix_t0_010000101100 (.a(t0_0100001011000), .b(t0_0100001011001), .y(t0_010000101100));
wire t0_0100001011000, t0_0100001011001;
mixer mix_t0_010000101101 (.a(t0_0100001011010), .b(t0_0100001011011), .y(t0_010000101101));
wire t0_0100001011010, t0_0100001011011;
mixer mix_t0_01000010111 (.a(t0_010000101110), .b(t0_010000101111), .y(t0_01000010111));
wire t0_010000101110, t0_010000101111;
mixer mix_t0_010000101110 (.a(t0_0100001011100), .b(t0_0100001011101), .y(t0_010000101110));
wire t0_0100001011100, t0_0100001011101;
mixer mix_t0_010000101111 (.a(t0_0100001011110), .b(t0_0100001011111), .y(t0_010000101111));
wire t0_0100001011110, t0_0100001011111;
mixer mix_t0_01000011 (.a(t0_010000110), .b(t0_010000111), .y(t0_01000011));
wire t0_010000110, t0_010000111;
mixer mix_t0_010000110 (.a(t0_0100001100), .b(t0_0100001101), .y(t0_010000110));
wire t0_0100001100, t0_0100001101;
mixer mix_t0_0100001100 (.a(t0_01000011000), .b(t0_01000011001), .y(t0_0100001100));
wire t0_01000011000, t0_01000011001;
mixer mix_t0_01000011000 (.a(t0_010000110000), .b(t0_010000110001), .y(t0_01000011000));
wire t0_010000110000, t0_010000110001;
mixer mix_t0_010000110000 (.a(t0_0100001100000), .b(t0_0100001100001), .y(t0_010000110000));
wire t0_0100001100000, t0_0100001100001;
mixer mix_t0_010000110001 (.a(t0_0100001100010), .b(t0_0100001100011), .y(t0_010000110001));
wire t0_0100001100010, t0_0100001100011;
mixer mix_t0_01000011001 (.a(t0_010000110010), .b(t0_010000110011), .y(t0_01000011001));
wire t0_010000110010, t0_010000110011;
mixer mix_t0_010000110010 (.a(t0_0100001100100), .b(t0_0100001100101), .y(t0_010000110010));
wire t0_0100001100100, t0_0100001100101;
mixer mix_t0_010000110011 (.a(t0_0100001100110), .b(t0_0100001100111), .y(t0_010000110011));
wire t0_0100001100110, t0_0100001100111;
mixer mix_t0_0100001101 (.a(t0_01000011010), .b(t0_01000011011), .y(t0_0100001101));
wire t0_01000011010, t0_01000011011;
mixer mix_t0_01000011010 (.a(t0_010000110100), .b(t0_010000110101), .y(t0_01000011010));
wire t0_010000110100, t0_010000110101;
mixer mix_t0_010000110100 (.a(t0_0100001101000), .b(t0_0100001101001), .y(t0_010000110100));
wire t0_0100001101000, t0_0100001101001;
mixer mix_t0_010000110101 (.a(t0_0100001101010), .b(t0_0100001101011), .y(t0_010000110101));
wire t0_0100001101010, t0_0100001101011;
mixer mix_t0_01000011011 (.a(t0_010000110110), .b(t0_010000110111), .y(t0_01000011011));
wire t0_010000110110, t0_010000110111;
mixer mix_t0_010000110110 (.a(t0_0100001101100), .b(t0_0100001101101), .y(t0_010000110110));
wire t0_0100001101100, t0_0100001101101;
mixer mix_t0_010000110111 (.a(t0_0100001101110), .b(t0_0100001101111), .y(t0_010000110111));
wire t0_0100001101110, t0_0100001101111;
mixer mix_t0_010000111 (.a(t0_0100001110), .b(t0_0100001111), .y(t0_010000111));
wire t0_0100001110, t0_0100001111;
mixer mix_t0_0100001110 (.a(t0_01000011100), .b(t0_01000011101), .y(t0_0100001110));
wire t0_01000011100, t0_01000011101;
mixer mix_t0_01000011100 (.a(t0_010000111000), .b(t0_010000111001), .y(t0_01000011100));
wire t0_010000111000, t0_010000111001;
mixer mix_t0_010000111000 (.a(t0_0100001110000), .b(t0_0100001110001), .y(t0_010000111000));
wire t0_0100001110000, t0_0100001110001;
mixer mix_t0_010000111001 (.a(t0_0100001110010), .b(t0_0100001110011), .y(t0_010000111001));
wire t0_0100001110010, t0_0100001110011;
mixer mix_t0_01000011101 (.a(t0_010000111010), .b(t0_010000111011), .y(t0_01000011101));
wire t0_010000111010, t0_010000111011;
mixer mix_t0_010000111010 (.a(t0_0100001110100), .b(t0_0100001110101), .y(t0_010000111010));
wire t0_0100001110100, t0_0100001110101;
mixer mix_t0_010000111011 (.a(t0_0100001110110), .b(t0_0100001110111), .y(t0_010000111011));
wire t0_0100001110110, t0_0100001110111;
mixer mix_t0_0100001111 (.a(t0_01000011110), .b(t0_01000011111), .y(t0_0100001111));
wire t0_01000011110, t0_01000011111;
mixer mix_t0_01000011110 (.a(t0_010000111100), .b(t0_010000111101), .y(t0_01000011110));
wire t0_010000111100, t0_010000111101;
mixer mix_t0_010000111100 (.a(t0_0100001111000), .b(t0_0100001111001), .y(t0_010000111100));
wire t0_0100001111000, t0_0100001111001;
mixer mix_t0_010000111101 (.a(t0_0100001111010), .b(t0_0100001111011), .y(t0_010000111101));
wire t0_0100001111010, t0_0100001111011;
mixer mix_t0_01000011111 (.a(t0_010000111110), .b(t0_010000111111), .y(t0_01000011111));
wire t0_010000111110, t0_010000111111;
mixer mix_t0_010000111110 (.a(t0_0100001111100), .b(t0_0100001111101), .y(t0_010000111110));
wire t0_0100001111100, t0_0100001111101;
mixer mix_t0_010000111111 (.a(t0_0100001111110), .b(t0_0100001111111), .y(t0_010000111111));
wire t0_0100001111110, t0_0100001111111;
mixer mix_t0_010001 (.a(t0_0100010), .b(t0_0100011), .y(t0_010001));
wire t0_0100010, t0_0100011;
mixer mix_t0_0100010 (.a(t0_01000100), .b(t0_01000101), .y(t0_0100010));
wire t0_01000100, t0_01000101;
mixer mix_t0_01000100 (.a(t0_010001000), .b(t0_010001001), .y(t0_01000100));
wire t0_010001000, t0_010001001;
mixer mix_t0_010001000 (.a(t0_0100010000), .b(t0_0100010001), .y(t0_010001000));
wire t0_0100010000, t0_0100010001;
mixer mix_t0_0100010000 (.a(t0_01000100000), .b(t0_01000100001), .y(t0_0100010000));
wire t0_01000100000, t0_01000100001;
mixer mix_t0_01000100000 (.a(t0_010001000000), .b(t0_010001000001), .y(t0_01000100000));
wire t0_010001000000, t0_010001000001;
mixer mix_t0_010001000000 (.a(t0_0100010000000), .b(t0_0100010000001), .y(t0_010001000000));
wire t0_0100010000000, t0_0100010000001;
mixer mix_t0_010001000001 (.a(t0_0100010000010), .b(t0_0100010000011), .y(t0_010001000001));
wire t0_0100010000010, t0_0100010000011;
mixer mix_t0_01000100001 (.a(t0_010001000010), .b(t0_010001000011), .y(t0_01000100001));
wire t0_010001000010, t0_010001000011;
mixer mix_t0_010001000010 (.a(t0_0100010000100), .b(t0_0100010000101), .y(t0_010001000010));
wire t0_0100010000100, t0_0100010000101;
mixer mix_t0_010001000011 (.a(t0_0100010000110), .b(t0_0100010000111), .y(t0_010001000011));
wire t0_0100010000110, t0_0100010000111;
mixer mix_t0_0100010001 (.a(t0_01000100010), .b(t0_01000100011), .y(t0_0100010001));
wire t0_01000100010, t0_01000100011;
mixer mix_t0_01000100010 (.a(t0_010001000100), .b(t0_010001000101), .y(t0_01000100010));
wire t0_010001000100, t0_010001000101;
mixer mix_t0_010001000100 (.a(t0_0100010001000), .b(t0_0100010001001), .y(t0_010001000100));
wire t0_0100010001000, t0_0100010001001;
mixer mix_t0_010001000101 (.a(t0_0100010001010), .b(t0_0100010001011), .y(t0_010001000101));
wire t0_0100010001010, t0_0100010001011;
mixer mix_t0_01000100011 (.a(t0_010001000110), .b(t0_010001000111), .y(t0_01000100011));
wire t0_010001000110, t0_010001000111;
mixer mix_t0_010001000110 (.a(t0_0100010001100), .b(t0_0100010001101), .y(t0_010001000110));
wire t0_0100010001100, t0_0100010001101;
mixer mix_t0_010001000111 (.a(t0_0100010001110), .b(t0_0100010001111), .y(t0_010001000111));
wire t0_0100010001110, t0_0100010001111;
mixer mix_t0_010001001 (.a(t0_0100010010), .b(t0_0100010011), .y(t0_010001001));
wire t0_0100010010, t0_0100010011;
mixer mix_t0_0100010010 (.a(t0_01000100100), .b(t0_01000100101), .y(t0_0100010010));
wire t0_01000100100, t0_01000100101;
mixer mix_t0_01000100100 (.a(t0_010001001000), .b(t0_010001001001), .y(t0_01000100100));
wire t0_010001001000, t0_010001001001;
mixer mix_t0_010001001000 (.a(t0_0100010010000), .b(t0_0100010010001), .y(t0_010001001000));
wire t0_0100010010000, t0_0100010010001;
mixer mix_t0_010001001001 (.a(t0_0100010010010), .b(t0_0100010010011), .y(t0_010001001001));
wire t0_0100010010010, t0_0100010010011;
mixer mix_t0_01000100101 (.a(t0_010001001010), .b(t0_010001001011), .y(t0_01000100101));
wire t0_010001001010, t0_010001001011;
mixer mix_t0_010001001010 (.a(t0_0100010010100), .b(t0_0100010010101), .y(t0_010001001010));
wire t0_0100010010100, t0_0100010010101;
mixer mix_t0_010001001011 (.a(t0_0100010010110), .b(t0_0100010010111), .y(t0_010001001011));
wire t0_0100010010110, t0_0100010010111;
mixer mix_t0_0100010011 (.a(t0_01000100110), .b(t0_01000100111), .y(t0_0100010011));
wire t0_01000100110, t0_01000100111;
mixer mix_t0_01000100110 (.a(t0_010001001100), .b(t0_010001001101), .y(t0_01000100110));
wire t0_010001001100, t0_010001001101;
mixer mix_t0_010001001100 (.a(t0_0100010011000), .b(t0_0100010011001), .y(t0_010001001100));
wire t0_0100010011000, t0_0100010011001;
mixer mix_t0_010001001101 (.a(t0_0100010011010), .b(t0_0100010011011), .y(t0_010001001101));
wire t0_0100010011010, t0_0100010011011;
mixer mix_t0_01000100111 (.a(t0_010001001110), .b(t0_010001001111), .y(t0_01000100111));
wire t0_010001001110, t0_010001001111;
mixer mix_t0_010001001110 (.a(t0_0100010011100), .b(t0_0100010011101), .y(t0_010001001110));
wire t0_0100010011100, t0_0100010011101;
mixer mix_t0_010001001111 (.a(t0_0100010011110), .b(t0_0100010011111), .y(t0_010001001111));
wire t0_0100010011110, t0_0100010011111;
mixer mix_t0_01000101 (.a(t0_010001010), .b(t0_010001011), .y(t0_01000101));
wire t0_010001010, t0_010001011;
mixer mix_t0_010001010 (.a(t0_0100010100), .b(t0_0100010101), .y(t0_010001010));
wire t0_0100010100, t0_0100010101;
mixer mix_t0_0100010100 (.a(t0_01000101000), .b(t0_01000101001), .y(t0_0100010100));
wire t0_01000101000, t0_01000101001;
mixer mix_t0_01000101000 (.a(t0_010001010000), .b(t0_010001010001), .y(t0_01000101000));
wire t0_010001010000, t0_010001010001;
mixer mix_t0_010001010000 (.a(t0_0100010100000), .b(t0_0100010100001), .y(t0_010001010000));
wire t0_0100010100000, t0_0100010100001;
mixer mix_t0_010001010001 (.a(t0_0100010100010), .b(t0_0100010100011), .y(t0_010001010001));
wire t0_0100010100010, t0_0100010100011;
mixer mix_t0_01000101001 (.a(t0_010001010010), .b(t0_010001010011), .y(t0_01000101001));
wire t0_010001010010, t0_010001010011;
mixer mix_t0_010001010010 (.a(t0_0100010100100), .b(t0_0100010100101), .y(t0_010001010010));
wire t0_0100010100100, t0_0100010100101;
mixer mix_t0_010001010011 (.a(t0_0100010100110), .b(t0_0100010100111), .y(t0_010001010011));
wire t0_0100010100110, t0_0100010100111;
mixer mix_t0_0100010101 (.a(t0_01000101010), .b(t0_01000101011), .y(t0_0100010101));
wire t0_01000101010, t0_01000101011;
mixer mix_t0_01000101010 (.a(t0_010001010100), .b(t0_010001010101), .y(t0_01000101010));
wire t0_010001010100, t0_010001010101;
mixer mix_t0_010001010100 (.a(t0_0100010101000), .b(t0_0100010101001), .y(t0_010001010100));
wire t0_0100010101000, t0_0100010101001;
mixer mix_t0_010001010101 (.a(t0_0100010101010), .b(t0_0100010101011), .y(t0_010001010101));
wire t0_0100010101010, t0_0100010101011;
mixer mix_t0_01000101011 (.a(t0_010001010110), .b(t0_010001010111), .y(t0_01000101011));
wire t0_010001010110, t0_010001010111;
mixer mix_t0_010001010110 (.a(t0_0100010101100), .b(t0_0100010101101), .y(t0_010001010110));
wire t0_0100010101100, t0_0100010101101;
mixer mix_t0_010001010111 (.a(t0_0100010101110), .b(t0_0100010101111), .y(t0_010001010111));
wire t0_0100010101110, t0_0100010101111;
mixer mix_t0_010001011 (.a(t0_0100010110), .b(t0_0100010111), .y(t0_010001011));
wire t0_0100010110, t0_0100010111;
mixer mix_t0_0100010110 (.a(t0_01000101100), .b(t0_01000101101), .y(t0_0100010110));
wire t0_01000101100, t0_01000101101;
mixer mix_t0_01000101100 (.a(t0_010001011000), .b(t0_010001011001), .y(t0_01000101100));
wire t0_010001011000, t0_010001011001;
mixer mix_t0_010001011000 (.a(t0_0100010110000), .b(t0_0100010110001), .y(t0_010001011000));
wire t0_0100010110000, t0_0100010110001;
mixer mix_t0_010001011001 (.a(t0_0100010110010), .b(t0_0100010110011), .y(t0_010001011001));
wire t0_0100010110010, t0_0100010110011;
mixer mix_t0_01000101101 (.a(t0_010001011010), .b(t0_010001011011), .y(t0_01000101101));
wire t0_010001011010, t0_010001011011;
mixer mix_t0_010001011010 (.a(t0_0100010110100), .b(t0_0100010110101), .y(t0_010001011010));
wire t0_0100010110100, t0_0100010110101;
mixer mix_t0_010001011011 (.a(t0_0100010110110), .b(t0_0100010110111), .y(t0_010001011011));
wire t0_0100010110110, t0_0100010110111;
mixer mix_t0_0100010111 (.a(t0_01000101110), .b(t0_01000101111), .y(t0_0100010111));
wire t0_01000101110, t0_01000101111;
mixer mix_t0_01000101110 (.a(t0_010001011100), .b(t0_010001011101), .y(t0_01000101110));
wire t0_010001011100, t0_010001011101;
mixer mix_t0_010001011100 (.a(t0_0100010111000), .b(t0_0100010111001), .y(t0_010001011100));
wire t0_0100010111000, t0_0100010111001;
mixer mix_t0_010001011101 (.a(t0_0100010111010), .b(t0_0100010111011), .y(t0_010001011101));
wire t0_0100010111010, t0_0100010111011;
mixer mix_t0_01000101111 (.a(t0_010001011110), .b(t0_010001011111), .y(t0_01000101111));
wire t0_010001011110, t0_010001011111;
mixer mix_t0_010001011110 (.a(t0_0100010111100), .b(t0_0100010111101), .y(t0_010001011110));
wire t0_0100010111100, t0_0100010111101;
mixer mix_t0_010001011111 (.a(t0_0100010111110), .b(t0_0100010111111), .y(t0_010001011111));
wire t0_0100010111110, t0_0100010111111;
mixer mix_t0_0100011 (.a(t0_01000110), .b(t0_01000111), .y(t0_0100011));
wire t0_01000110, t0_01000111;
mixer mix_t0_01000110 (.a(t0_010001100), .b(t0_010001101), .y(t0_01000110));
wire t0_010001100, t0_010001101;
mixer mix_t0_010001100 (.a(t0_0100011000), .b(t0_0100011001), .y(t0_010001100));
wire t0_0100011000, t0_0100011001;
mixer mix_t0_0100011000 (.a(t0_01000110000), .b(t0_01000110001), .y(t0_0100011000));
wire t0_01000110000, t0_01000110001;
mixer mix_t0_01000110000 (.a(t0_010001100000), .b(t0_010001100001), .y(t0_01000110000));
wire t0_010001100000, t0_010001100001;
mixer mix_t0_010001100000 (.a(t0_0100011000000), .b(t0_0100011000001), .y(t0_010001100000));
wire t0_0100011000000, t0_0100011000001;
mixer mix_t0_010001100001 (.a(t0_0100011000010), .b(t0_0100011000011), .y(t0_010001100001));
wire t0_0100011000010, t0_0100011000011;
mixer mix_t0_01000110001 (.a(t0_010001100010), .b(t0_010001100011), .y(t0_01000110001));
wire t0_010001100010, t0_010001100011;
mixer mix_t0_010001100010 (.a(t0_0100011000100), .b(t0_0100011000101), .y(t0_010001100010));
wire t0_0100011000100, t0_0100011000101;
mixer mix_t0_010001100011 (.a(t0_0100011000110), .b(t0_0100011000111), .y(t0_010001100011));
wire t0_0100011000110, t0_0100011000111;
mixer mix_t0_0100011001 (.a(t0_01000110010), .b(t0_01000110011), .y(t0_0100011001));
wire t0_01000110010, t0_01000110011;
mixer mix_t0_01000110010 (.a(t0_010001100100), .b(t0_010001100101), .y(t0_01000110010));
wire t0_010001100100, t0_010001100101;
mixer mix_t0_010001100100 (.a(t0_0100011001000), .b(t0_0100011001001), .y(t0_010001100100));
wire t0_0100011001000, t0_0100011001001;
mixer mix_t0_010001100101 (.a(t0_0100011001010), .b(t0_0100011001011), .y(t0_010001100101));
wire t0_0100011001010, t0_0100011001011;
mixer mix_t0_01000110011 (.a(t0_010001100110), .b(t0_010001100111), .y(t0_01000110011));
wire t0_010001100110, t0_010001100111;
mixer mix_t0_010001100110 (.a(t0_0100011001100), .b(t0_0100011001101), .y(t0_010001100110));
wire t0_0100011001100, t0_0100011001101;
mixer mix_t0_010001100111 (.a(t0_0100011001110), .b(t0_0100011001111), .y(t0_010001100111));
wire t0_0100011001110, t0_0100011001111;
mixer mix_t0_010001101 (.a(t0_0100011010), .b(t0_0100011011), .y(t0_010001101));
wire t0_0100011010, t0_0100011011;
mixer mix_t0_0100011010 (.a(t0_01000110100), .b(t0_01000110101), .y(t0_0100011010));
wire t0_01000110100, t0_01000110101;
mixer mix_t0_01000110100 (.a(t0_010001101000), .b(t0_010001101001), .y(t0_01000110100));
wire t0_010001101000, t0_010001101001;
mixer mix_t0_010001101000 (.a(t0_0100011010000), .b(t0_0100011010001), .y(t0_010001101000));
wire t0_0100011010000, t0_0100011010001;
mixer mix_t0_010001101001 (.a(t0_0100011010010), .b(t0_0100011010011), .y(t0_010001101001));
wire t0_0100011010010, t0_0100011010011;
mixer mix_t0_01000110101 (.a(t0_010001101010), .b(t0_010001101011), .y(t0_01000110101));
wire t0_010001101010, t0_010001101011;
mixer mix_t0_010001101010 (.a(t0_0100011010100), .b(t0_0100011010101), .y(t0_010001101010));
wire t0_0100011010100, t0_0100011010101;
mixer mix_t0_010001101011 (.a(t0_0100011010110), .b(t0_0100011010111), .y(t0_010001101011));
wire t0_0100011010110, t0_0100011010111;
mixer mix_t0_0100011011 (.a(t0_01000110110), .b(t0_01000110111), .y(t0_0100011011));
wire t0_01000110110, t0_01000110111;
mixer mix_t0_01000110110 (.a(t0_010001101100), .b(t0_010001101101), .y(t0_01000110110));
wire t0_010001101100, t0_010001101101;
mixer mix_t0_010001101100 (.a(t0_0100011011000), .b(t0_0100011011001), .y(t0_010001101100));
wire t0_0100011011000, t0_0100011011001;
mixer mix_t0_010001101101 (.a(t0_0100011011010), .b(t0_0100011011011), .y(t0_010001101101));
wire t0_0100011011010, t0_0100011011011;
mixer mix_t0_01000110111 (.a(t0_010001101110), .b(t0_010001101111), .y(t0_01000110111));
wire t0_010001101110, t0_010001101111;
mixer mix_t0_010001101110 (.a(t0_0100011011100), .b(t0_0100011011101), .y(t0_010001101110));
wire t0_0100011011100, t0_0100011011101;
mixer mix_t0_010001101111 (.a(t0_0100011011110), .b(t0_0100011011111), .y(t0_010001101111));
wire t0_0100011011110, t0_0100011011111;
mixer mix_t0_01000111 (.a(t0_010001110), .b(t0_010001111), .y(t0_01000111));
wire t0_010001110, t0_010001111;
mixer mix_t0_010001110 (.a(t0_0100011100), .b(t0_0100011101), .y(t0_010001110));
wire t0_0100011100, t0_0100011101;
mixer mix_t0_0100011100 (.a(t0_01000111000), .b(t0_01000111001), .y(t0_0100011100));
wire t0_01000111000, t0_01000111001;
mixer mix_t0_01000111000 (.a(t0_010001110000), .b(t0_010001110001), .y(t0_01000111000));
wire t0_010001110000, t0_010001110001;
mixer mix_t0_010001110000 (.a(t0_0100011100000), .b(t0_0100011100001), .y(t0_010001110000));
wire t0_0100011100000, t0_0100011100001;
mixer mix_t0_010001110001 (.a(t0_0100011100010), .b(t0_0100011100011), .y(t0_010001110001));
wire t0_0100011100010, t0_0100011100011;
mixer mix_t0_01000111001 (.a(t0_010001110010), .b(t0_010001110011), .y(t0_01000111001));
wire t0_010001110010, t0_010001110011;
mixer mix_t0_010001110010 (.a(t0_0100011100100), .b(t0_0100011100101), .y(t0_010001110010));
wire t0_0100011100100, t0_0100011100101;
mixer mix_t0_010001110011 (.a(t0_0100011100110), .b(t0_0100011100111), .y(t0_010001110011));
wire t0_0100011100110, t0_0100011100111;
mixer mix_t0_0100011101 (.a(t0_01000111010), .b(t0_01000111011), .y(t0_0100011101));
wire t0_01000111010, t0_01000111011;
mixer mix_t0_01000111010 (.a(t0_010001110100), .b(t0_010001110101), .y(t0_01000111010));
wire t0_010001110100, t0_010001110101;
mixer mix_t0_010001110100 (.a(t0_0100011101000), .b(t0_0100011101001), .y(t0_010001110100));
wire t0_0100011101000, t0_0100011101001;
mixer mix_t0_010001110101 (.a(t0_0100011101010), .b(t0_0100011101011), .y(t0_010001110101));
wire t0_0100011101010, t0_0100011101011;
mixer mix_t0_01000111011 (.a(t0_010001110110), .b(t0_010001110111), .y(t0_01000111011));
wire t0_010001110110, t0_010001110111;
mixer mix_t0_010001110110 (.a(t0_0100011101100), .b(t0_0100011101101), .y(t0_010001110110));
wire t0_0100011101100, t0_0100011101101;
mixer mix_t0_010001110111 (.a(t0_0100011101110), .b(t0_0100011101111), .y(t0_010001110111));
wire t0_0100011101110, t0_0100011101111;
mixer mix_t0_010001111 (.a(t0_0100011110), .b(t0_0100011111), .y(t0_010001111));
wire t0_0100011110, t0_0100011111;
mixer mix_t0_0100011110 (.a(t0_01000111100), .b(t0_01000111101), .y(t0_0100011110));
wire t0_01000111100, t0_01000111101;
mixer mix_t0_01000111100 (.a(t0_010001111000), .b(t0_010001111001), .y(t0_01000111100));
wire t0_010001111000, t0_010001111001;
mixer mix_t0_010001111000 (.a(t0_0100011110000), .b(t0_0100011110001), .y(t0_010001111000));
wire t0_0100011110000, t0_0100011110001;
mixer mix_t0_010001111001 (.a(t0_0100011110010), .b(t0_0100011110011), .y(t0_010001111001));
wire t0_0100011110010, t0_0100011110011;
mixer mix_t0_01000111101 (.a(t0_010001111010), .b(t0_010001111011), .y(t0_01000111101));
wire t0_010001111010, t0_010001111011;
mixer mix_t0_010001111010 (.a(t0_0100011110100), .b(t0_0100011110101), .y(t0_010001111010));
wire t0_0100011110100, t0_0100011110101;
mixer mix_t0_010001111011 (.a(t0_0100011110110), .b(t0_0100011110111), .y(t0_010001111011));
wire t0_0100011110110, t0_0100011110111;
mixer mix_t0_0100011111 (.a(t0_01000111110), .b(t0_01000111111), .y(t0_0100011111));
wire t0_01000111110, t0_01000111111;
mixer mix_t0_01000111110 (.a(t0_010001111100), .b(t0_010001111101), .y(t0_01000111110));
wire t0_010001111100, t0_010001111101;
mixer mix_t0_010001111100 (.a(t0_0100011111000), .b(t0_0100011111001), .y(t0_010001111100));
wire t0_0100011111000, t0_0100011111001;
mixer mix_t0_010001111101 (.a(t0_0100011111010), .b(t0_0100011111011), .y(t0_010001111101));
wire t0_0100011111010, t0_0100011111011;
mixer mix_t0_01000111111 (.a(t0_010001111110), .b(t0_010001111111), .y(t0_01000111111));
wire t0_010001111110, t0_010001111111;
mixer mix_t0_010001111110 (.a(t0_0100011111100), .b(t0_0100011111101), .y(t0_010001111110));
wire t0_0100011111100, t0_0100011111101;
mixer mix_t0_010001111111 (.a(t0_0100011111110), .b(t0_0100011111111), .y(t0_010001111111));
wire t0_0100011111110, t0_0100011111111;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_010010 (.a(t0_0100100), .b(t0_0100101), .y(t0_010010));
wire t0_0100100, t0_0100101;
mixer mix_t0_0100100 (.a(t0_01001000), .b(t0_01001001), .y(t0_0100100));
wire t0_01001000, t0_01001001;
mixer mix_t0_01001000 (.a(t0_010010000), .b(t0_010010001), .y(t0_01001000));
wire t0_010010000, t0_010010001;
mixer mix_t0_010010000 (.a(t0_0100100000), .b(t0_0100100001), .y(t0_010010000));
wire t0_0100100000, t0_0100100001;
mixer mix_t0_0100100000 (.a(t0_01001000000), .b(t0_01001000001), .y(t0_0100100000));
wire t0_01001000000, t0_01001000001;
mixer mix_t0_01001000000 (.a(t0_010010000000), .b(t0_010010000001), .y(t0_01001000000));
wire t0_010010000000, t0_010010000001;
mixer mix_t0_010010000000 (.a(t0_0100100000000), .b(t0_0100100000001), .y(t0_010010000000));
wire t0_0100100000000, t0_0100100000001;
mixer mix_t0_010010000001 (.a(t0_0100100000010), .b(t0_0100100000011), .y(t0_010010000001));
wire t0_0100100000010, t0_0100100000011;
mixer mix_t0_01001000001 (.a(t0_010010000010), .b(t0_010010000011), .y(t0_01001000001));
wire t0_010010000010, t0_010010000011;
mixer mix_t0_010010000010 (.a(t0_0100100000100), .b(t0_0100100000101), .y(t0_010010000010));
wire t0_0100100000100, t0_0100100000101;
mixer mix_t0_010010000011 (.a(t0_0100100000110), .b(t0_0100100000111), .y(t0_010010000011));
wire t0_0100100000110, t0_0100100000111;
mixer mix_t0_0100100001 (.a(t0_01001000010), .b(t0_01001000011), .y(t0_0100100001));
wire t0_01001000010, t0_01001000011;
mixer mix_t0_01001000010 (.a(t0_010010000100), .b(t0_010010000101), .y(t0_01001000010));
wire t0_010010000100, t0_010010000101;
mixer mix_t0_010010000100 (.a(t0_0100100001000), .b(t0_0100100001001), .y(t0_010010000100));
wire t0_0100100001000, t0_0100100001001;
mixer mix_t0_010010000101 (.a(t0_0100100001010), .b(t0_0100100001011), .y(t0_010010000101));
wire t0_0100100001010, t0_0100100001011;
mixer mix_t0_01001000011 (.a(t0_010010000110), .b(t0_010010000111), .y(t0_01001000011));
wire t0_010010000110, t0_010010000111;
mixer mix_t0_010010000110 (.a(t0_0100100001100), .b(t0_0100100001101), .y(t0_010010000110));
wire t0_0100100001100, t0_0100100001101;
mixer mix_t0_010010000111 (.a(t0_0100100001110), .b(t0_0100100001111), .y(t0_010010000111));
wire t0_0100100001110, t0_0100100001111;
mixer mix_t0_010010001 (.a(t0_0100100010), .b(t0_0100100011), .y(t0_010010001));
wire t0_0100100010, t0_0100100011;
mixer mix_t0_0100100010 (.a(t0_01001000100), .b(t0_01001000101), .y(t0_0100100010));
wire t0_01001000100, t0_01001000101;
mixer mix_t0_01001000100 (.a(t0_010010001000), .b(t0_010010001001), .y(t0_01001000100));
wire t0_010010001000, t0_010010001001;
mixer mix_t0_010010001000 (.a(t0_0100100010000), .b(t0_0100100010001), .y(t0_010010001000));
wire t0_0100100010000, t0_0100100010001;
mixer mix_t0_010010001001 (.a(t0_0100100010010), .b(t0_0100100010011), .y(t0_010010001001));
wire t0_0100100010010, t0_0100100010011;
mixer mix_t0_01001000101 (.a(t0_010010001010), .b(t0_010010001011), .y(t0_01001000101));
wire t0_010010001010, t0_010010001011;
mixer mix_t0_010010001010 (.a(t0_0100100010100), .b(t0_0100100010101), .y(t0_010010001010));
wire t0_0100100010100, t0_0100100010101;
mixer mix_t0_010010001011 (.a(t0_0100100010110), .b(t0_0100100010111), .y(t0_010010001011));
wire t0_0100100010110, t0_0100100010111;
mixer mix_t0_0100100011 (.a(t0_01001000110), .b(t0_01001000111), .y(t0_0100100011));
wire t0_01001000110, t0_01001000111;
mixer mix_t0_01001000110 (.a(t0_010010001100), .b(t0_010010001101), .y(t0_01001000110));
wire t0_010010001100, t0_010010001101;
mixer mix_t0_010010001100 (.a(t0_0100100011000), .b(t0_0100100011001), .y(t0_010010001100));
wire t0_0100100011000, t0_0100100011001;
mixer mix_t0_010010001101 (.a(t0_0100100011010), .b(t0_0100100011011), .y(t0_010010001101));
wire t0_0100100011010, t0_0100100011011;
mixer mix_t0_01001000111 (.a(t0_010010001110), .b(t0_010010001111), .y(t0_01001000111));
wire t0_010010001110, t0_010010001111;
mixer mix_t0_010010001110 (.a(t0_0100100011100), .b(t0_0100100011101), .y(t0_010010001110));
wire t0_0100100011100, t0_0100100011101;
mixer mix_t0_010010001111 (.a(t0_0100100011110), .b(t0_0100100011111), .y(t0_010010001111));
wire t0_0100100011110, t0_0100100011111;
mixer mix_t0_01001001 (.a(t0_010010010), .b(t0_010010011), .y(t0_01001001));
wire t0_010010010, t0_010010011;
mixer mix_t0_010010010 (.a(t0_0100100100), .b(t0_0100100101), .y(t0_010010010));
wire t0_0100100100, t0_0100100101;
mixer mix_t0_0100100100 (.a(t0_01001001000), .b(t0_01001001001), .y(t0_0100100100));
wire t0_01001001000, t0_01001001001;
mixer mix_t0_01001001000 (.a(t0_010010010000), .b(t0_010010010001), .y(t0_01001001000));
wire t0_010010010000, t0_010010010001;
mixer mix_t0_010010010000 (.a(t0_0100100100000), .b(t0_0100100100001), .y(t0_010010010000));
wire t0_0100100100000, t0_0100100100001;
mixer mix_t0_010010010001 (.a(t0_0100100100010), .b(t0_0100100100011), .y(t0_010010010001));
wire t0_0100100100010, t0_0100100100011;
mixer mix_t0_01001001001 (.a(t0_010010010010), .b(t0_010010010011), .y(t0_01001001001));
wire t0_010010010010, t0_010010010011;
mixer mix_t0_010010010010 (.a(t0_0100100100100), .b(t0_0100100100101), .y(t0_010010010010));
wire t0_0100100100100, t0_0100100100101;
mixer mix_t0_010010010011 (.a(t0_0100100100110), .b(t0_0100100100111), .y(t0_010010010011));
wire t0_0100100100110, t0_0100100100111;
mixer mix_t0_0100100101 (.a(t0_01001001010), .b(t0_01001001011), .y(t0_0100100101));
wire t0_01001001010, t0_01001001011;
mixer mix_t0_01001001010 (.a(t0_010010010100), .b(t0_010010010101), .y(t0_01001001010));
wire t0_010010010100, t0_010010010101;
mixer mix_t0_010010010100 (.a(t0_0100100101000), .b(t0_0100100101001), .y(t0_010010010100));
wire t0_0100100101000, t0_0100100101001;
mixer mix_t0_010010010101 (.a(t0_0100100101010), .b(t0_0100100101011), .y(t0_010010010101));
wire t0_0100100101010, t0_0100100101011;
mixer mix_t0_01001001011 (.a(t0_010010010110), .b(t0_010010010111), .y(t0_01001001011));
wire t0_010010010110, t0_010010010111;
mixer mix_t0_010010010110 (.a(t0_0100100101100), .b(t0_0100100101101), .y(t0_010010010110));
wire t0_0100100101100, t0_0100100101101;
mixer mix_t0_010010010111 (.a(t0_0100100101110), .b(t0_0100100101111), .y(t0_010010010111));
wire t0_0100100101110, t0_0100100101111;
mixer mix_t0_010010011 (.a(t0_0100100110), .b(t0_0100100111), .y(t0_010010011));
wire t0_0100100110, t0_0100100111;
mixer mix_t0_0100100110 (.a(t0_01001001100), .b(t0_01001001101), .y(t0_0100100110));
wire t0_01001001100, t0_01001001101;
mixer mix_t0_01001001100 (.a(t0_010010011000), .b(t0_010010011001), .y(t0_01001001100));
wire t0_010010011000, t0_010010011001;
mixer mix_t0_010010011000 (.a(t0_0100100110000), .b(t0_0100100110001), .y(t0_010010011000));
wire t0_0100100110000, t0_0100100110001;
mixer mix_t0_010010011001 (.a(t0_0100100110010), .b(t0_0100100110011), .y(t0_010010011001));
wire t0_0100100110010, t0_0100100110011;
mixer mix_t0_01001001101 (.a(t0_010010011010), .b(t0_010010011011), .y(t0_01001001101));
wire t0_010010011010, t0_010010011011;
mixer mix_t0_010010011010 (.a(t0_0100100110100), .b(t0_0100100110101), .y(t0_010010011010));
wire t0_0100100110100, t0_0100100110101;
mixer mix_t0_010010011011 (.a(t0_0100100110110), .b(t0_0100100110111), .y(t0_010010011011));
wire t0_0100100110110, t0_0100100110111;
mixer mix_t0_0100100111 (.a(t0_01001001110), .b(t0_01001001111), .y(t0_0100100111));
wire t0_01001001110, t0_01001001111;
mixer mix_t0_01001001110 (.a(t0_010010011100), .b(t0_010010011101), .y(t0_01001001110));
wire t0_010010011100, t0_010010011101;
mixer mix_t0_010010011100 (.a(t0_0100100111000), .b(t0_0100100111001), .y(t0_010010011100));
wire t0_0100100111000, t0_0100100111001;
mixer mix_t0_010010011101 (.a(t0_0100100111010), .b(t0_0100100111011), .y(t0_010010011101));
wire t0_0100100111010, t0_0100100111011;
mixer mix_t0_01001001111 (.a(t0_010010011110), .b(t0_010010011111), .y(t0_01001001111));
wire t0_010010011110, t0_010010011111;
mixer mix_t0_010010011110 (.a(t0_0100100111100), .b(t0_0100100111101), .y(t0_010010011110));
wire t0_0100100111100, t0_0100100111101;
mixer mix_t0_010010011111 (.a(t0_0100100111110), .b(t0_0100100111111), .y(t0_010010011111));
wire t0_0100100111110, t0_0100100111111;
mixer mix_t0_0100101 (.a(t0_01001010), .b(t0_01001011), .y(t0_0100101));
wire t0_01001010, t0_01001011;
mixer mix_t0_01001010 (.a(t0_010010100), .b(t0_010010101), .y(t0_01001010));
wire t0_010010100, t0_010010101;
mixer mix_t0_010010100 (.a(t0_0100101000), .b(t0_0100101001), .y(t0_010010100));
wire t0_0100101000, t0_0100101001;
mixer mix_t0_0100101000 (.a(t0_01001010000), .b(t0_01001010001), .y(t0_0100101000));
wire t0_01001010000, t0_01001010001;
mixer mix_t0_01001010000 (.a(t0_010010100000), .b(t0_010010100001), .y(t0_01001010000));
wire t0_010010100000, t0_010010100001;
mixer mix_t0_010010100000 (.a(t0_0100101000000), .b(t0_0100101000001), .y(t0_010010100000));
wire t0_0100101000000, t0_0100101000001;
mixer mix_t0_010010100001 (.a(t0_0100101000010), .b(t0_0100101000011), .y(t0_010010100001));
wire t0_0100101000010, t0_0100101000011;
mixer mix_t0_01001010001 (.a(t0_010010100010), .b(t0_010010100011), .y(t0_01001010001));
wire t0_010010100010, t0_010010100011;
mixer mix_t0_010010100010 (.a(t0_0100101000100), .b(t0_0100101000101), .y(t0_010010100010));
wire t0_0100101000100, t0_0100101000101;
mixer mix_t0_010010100011 (.a(t0_0100101000110), .b(t0_0100101000111), .y(t0_010010100011));
wire t0_0100101000110, t0_0100101000111;
mixer mix_t0_0100101001 (.a(t0_01001010010), .b(t0_01001010011), .y(t0_0100101001));
wire t0_01001010010, t0_01001010011;
mixer mix_t0_01001010010 (.a(t0_010010100100), .b(t0_010010100101), .y(t0_01001010010));
wire t0_010010100100, t0_010010100101;
mixer mix_t0_010010100100 (.a(t0_0100101001000), .b(t0_0100101001001), .y(t0_010010100100));
wire t0_0100101001000, t0_0100101001001;
mixer mix_t0_010010100101 (.a(t0_0100101001010), .b(t0_0100101001011), .y(t0_010010100101));
wire t0_0100101001010, t0_0100101001011;
mixer mix_t0_01001010011 (.a(t0_010010100110), .b(t0_010010100111), .y(t0_01001010011));
wire t0_010010100110, t0_010010100111;
mixer mix_t0_010010100110 (.a(t0_0100101001100), .b(t0_0100101001101), .y(t0_010010100110));
wire t0_0100101001100, t0_0100101001101;
mixer mix_t0_010010100111 (.a(t0_0100101001110), .b(t0_0100101001111), .y(t0_010010100111));
wire t0_0100101001110, t0_0100101001111;
mixer mix_t0_010010101 (.a(t0_0100101010), .b(t0_0100101011), .y(t0_010010101));
wire t0_0100101010, t0_0100101011;
mixer mix_t0_0100101010 (.a(t0_01001010100), .b(t0_01001010101), .y(t0_0100101010));
wire t0_01001010100, t0_01001010101;
mixer mix_t0_01001010100 (.a(t0_010010101000), .b(t0_010010101001), .y(t0_01001010100));
wire t0_010010101000, t0_010010101001;
mixer mix_t0_010010101000 (.a(t0_0100101010000), .b(t0_0100101010001), .y(t0_010010101000));
wire t0_0100101010000, t0_0100101010001;
mixer mix_t0_010010101001 (.a(t0_0100101010010), .b(t0_0100101010011), .y(t0_010010101001));
wire t0_0100101010010, t0_0100101010011;
mixer mix_t0_01001010101 (.a(t0_010010101010), .b(t0_010010101011), .y(t0_01001010101));
wire t0_010010101010, t0_010010101011;
mixer mix_t0_010010101010 (.a(t0_0100101010100), .b(t0_0100101010101), .y(t0_010010101010));
wire t0_0100101010100, t0_0100101010101;
mixer mix_t0_010010101011 (.a(t0_0100101010110), .b(t0_0100101010111), .y(t0_010010101011));
wire t0_0100101010110, t0_0100101010111;
mixer mix_t0_0100101011 (.a(t0_01001010110), .b(t0_01001010111), .y(t0_0100101011));
wire t0_01001010110, t0_01001010111;
mixer mix_t0_01001010110 (.a(t0_010010101100), .b(t0_010010101101), .y(t0_01001010110));
wire t0_010010101100, t0_010010101101;
mixer mix_t0_010010101100 (.a(t0_0100101011000), .b(t0_0100101011001), .y(t0_010010101100));
wire t0_0100101011000, t0_0100101011001;
mixer mix_t0_010010101101 (.a(t0_0100101011010), .b(t0_0100101011011), .y(t0_010010101101));
wire t0_0100101011010, t0_0100101011011;
mixer mix_t0_01001010111 (.a(t0_010010101110), .b(t0_010010101111), .y(t0_01001010111));
wire t0_010010101110, t0_010010101111;
mixer mix_t0_010010101110 (.a(t0_0100101011100), .b(t0_0100101011101), .y(t0_010010101110));
wire t0_0100101011100, t0_0100101011101;
mixer mix_t0_010010101111 (.a(t0_0100101011110), .b(t0_0100101011111), .y(t0_010010101111));
wire t0_0100101011110, t0_0100101011111;
mixer mix_t0_01001011 (.a(t0_010010110), .b(t0_010010111), .y(t0_01001011));
wire t0_010010110, t0_010010111;
mixer mix_t0_010010110 (.a(t0_0100101100), .b(t0_0100101101), .y(t0_010010110));
wire t0_0100101100, t0_0100101101;
mixer mix_t0_0100101100 (.a(t0_01001011000), .b(t0_01001011001), .y(t0_0100101100));
wire t0_01001011000, t0_01001011001;
mixer mix_t0_01001011000 (.a(t0_010010110000), .b(t0_010010110001), .y(t0_01001011000));
wire t0_010010110000, t0_010010110001;
mixer mix_t0_010010110000 (.a(t0_0100101100000), .b(t0_0100101100001), .y(t0_010010110000));
wire t0_0100101100000, t0_0100101100001;
mixer mix_t0_010010110001 (.a(t0_0100101100010), .b(t0_0100101100011), .y(t0_010010110001));
wire t0_0100101100010, t0_0100101100011;
mixer mix_t0_01001011001 (.a(t0_010010110010), .b(t0_010010110011), .y(t0_01001011001));
wire t0_010010110010, t0_010010110011;
mixer mix_t0_010010110010 (.a(t0_0100101100100), .b(t0_0100101100101), .y(t0_010010110010));
wire t0_0100101100100, t0_0100101100101;
mixer mix_t0_010010110011 (.a(t0_0100101100110), .b(t0_0100101100111), .y(t0_010010110011));
wire t0_0100101100110, t0_0100101100111;
mixer mix_t0_0100101101 (.a(t0_01001011010), .b(t0_01001011011), .y(t0_0100101101));
wire t0_01001011010, t0_01001011011;
mixer mix_t0_01001011010 (.a(t0_010010110100), .b(t0_010010110101), .y(t0_01001011010));
wire t0_010010110100, t0_010010110101;
mixer mix_t0_010010110100 (.a(t0_0100101101000), .b(t0_0100101101001), .y(t0_010010110100));
wire t0_0100101101000, t0_0100101101001;
mixer mix_t0_010010110101 (.a(t0_0100101101010), .b(t0_0100101101011), .y(t0_010010110101));
wire t0_0100101101010, t0_0100101101011;
mixer mix_t0_01001011011 (.a(t0_010010110110), .b(t0_010010110111), .y(t0_01001011011));
wire t0_010010110110, t0_010010110111;
mixer mix_t0_010010110110 (.a(t0_0100101101100), .b(t0_0100101101101), .y(t0_010010110110));
wire t0_0100101101100, t0_0100101101101;
mixer mix_t0_010010110111 (.a(t0_0100101101110), .b(t0_0100101101111), .y(t0_010010110111));
wire t0_0100101101110, t0_0100101101111;
mixer mix_t0_010010111 (.a(t0_0100101110), .b(t0_0100101111), .y(t0_010010111));
wire t0_0100101110, t0_0100101111;
mixer mix_t0_0100101110 (.a(t0_01001011100), .b(t0_01001011101), .y(t0_0100101110));
wire t0_01001011100, t0_01001011101;
mixer mix_t0_01001011100 (.a(t0_010010111000), .b(t0_010010111001), .y(t0_01001011100));
wire t0_010010111000, t0_010010111001;
mixer mix_t0_010010111000 (.a(t0_0100101110000), .b(t0_0100101110001), .y(t0_010010111000));
wire t0_0100101110000, t0_0100101110001;
mixer mix_t0_010010111001 (.a(t0_0100101110010), .b(t0_0100101110011), .y(t0_010010111001));
wire t0_0100101110010, t0_0100101110011;
mixer mix_t0_01001011101 (.a(t0_010010111010), .b(t0_010010111011), .y(t0_01001011101));
wire t0_010010111010, t0_010010111011;
mixer mix_t0_010010111010 (.a(t0_0100101110100), .b(t0_0100101110101), .y(t0_010010111010));
wire t0_0100101110100, t0_0100101110101;
mixer mix_t0_010010111011 (.a(t0_0100101110110), .b(t0_0100101110111), .y(t0_010010111011));
wire t0_0100101110110, t0_0100101110111;
mixer mix_t0_0100101111 (.a(t0_01001011110), .b(t0_01001011111), .y(t0_0100101111));
wire t0_01001011110, t0_01001011111;
mixer mix_t0_01001011110 (.a(t0_010010111100), .b(t0_010010111101), .y(t0_01001011110));
wire t0_010010111100, t0_010010111101;
mixer mix_t0_010010111100 (.a(t0_0100101111000), .b(t0_0100101111001), .y(t0_010010111100));
wire t0_0100101111000, t0_0100101111001;
mixer mix_t0_010010111101 (.a(t0_0100101111010), .b(t0_0100101111011), .y(t0_010010111101));
wire t0_0100101111010, t0_0100101111011;
mixer mix_t0_01001011111 (.a(t0_010010111110), .b(t0_010010111111), .y(t0_01001011111));
wire t0_010010111110, t0_010010111111;
mixer mix_t0_010010111110 (.a(t0_0100101111100), .b(t0_0100101111101), .y(t0_010010111110));
wire t0_0100101111100, t0_0100101111101;
mixer mix_t0_010010111111 (.a(t0_0100101111110), .b(t0_0100101111111), .y(t0_010010111111));
wire t0_0100101111110, t0_0100101111111;
mixer mix_t0_010011 (.a(t0_0100110), .b(t0_0100111), .y(t0_010011));
wire t0_0100110, t0_0100111;
mixer mix_t0_0100110 (.a(t0_01001100), .b(t0_01001101), .y(t0_0100110));
wire t0_01001100, t0_01001101;
mixer mix_t0_01001100 (.a(t0_010011000), .b(t0_010011001), .y(t0_01001100));
wire t0_010011000, t0_010011001;
mixer mix_t0_010011000 (.a(t0_0100110000), .b(t0_0100110001), .y(t0_010011000));
wire t0_0100110000, t0_0100110001;
mixer mix_t0_0100110000 (.a(t0_01001100000), .b(t0_01001100001), .y(t0_0100110000));
wire t0_01001100000, t0_01001100001;
mixer mix_t0_01001100000 (.a(t0_010011000000), .b(t0_010011000001), .y(t0_01001100000));
wire t0_010011000000, t0_010011000001;
mixer mix_t0_010011000000 (.a(t0_0100110000000), .b(t0_0100110000001), .y(t0_010011000000));
wire t0_0100110000000, t0_0100110000001;
mixer mix_t0_010011000001 (.a(t0_0100110000010), .b(t0_0100110000011), .y(t0_010011000001));
wire t0_0100110000010, t0_0100110000011;
mixer mix_t0_01001100001 (.a(t0_010011000010), .b(t0_010011000011), .y(t0_01001100001));
wire t0_010011000010, t0_010011000011;
mixer mix_t0_010011000010 (.a(t0_0100110000100), .b(t0_0100110000101), .y(t0_010011000010));
wire t0_0100110000100, t0_0100110000101;
mixer mix_t0_010011000011 (.a(t0_0100110000110), .b(t0_0100110000111), .y(t0_010011000011));
wire t0_0100110000110, t0_0100110000111;
mixer mix_t0_0100110001 (.a(t0_01001100010), .b(t0_01001100011), .y(t0_0100110001));
wire t0_01001100010, t0_01001100011;
mixer mix_t0_01001100010 (.a(t0_010011000100), .b(t0_010011000101), .y(t0_01001100010));
wire t0_010011000100, t0_010011000101;
mixer mix_t0_010011000100 (.a(t0_0100110001000), .b(t0_0100110001001), .y(t0_010011000100));
wire t0_0100110001000, t0_0100110001001;
mixer mix_t0_010011000101 (.a(t0_0100110001010), .b(t0_0100110001011), .y(t0_010011000101));
wire t0_0100110001010, t0_0100110001011;
mixer mix_t0_01001100011 (.a(t0_010011000110), .b(t0_010011000111), .y(t0_01001100011));
wire t0_010011000110, t0_010011000111;
mixer mix_t0_010011000110 (.a(t0_0100110001100), .b(t0_0100110001101), .y(t0_010011000110));
wire t0_0100110001100, t0_0100110001101;
mixer mix_t0_010011000111 (.a(t0_0100110001110), .b(t0_0100110001111), .y(t0_010011000111));
wire t0_0100110001110, t0_0100110001111;
mixer mix_t0_010011001 (.a(t0_0100110010), .b(t0_0100110011), .y(t0_010011001));
wire t0_0100110010, t0_0100110011;
mixer mix_t0_0100110010 (.a(t0_01001100100), .b(t0_01001100101), .y(t0_0100110010));
wire t0_01001100100, t0_01001100101;
mixer mix_t0_01001100100 (.a(t0_010011001000), .b(t0_010011001001), .y(t0_01001100100));
wire t0_010011001000, t0_010011001001;
mixer mix_t0_010011001000 (.a(t0_0100110010000), .b(t0_0100110010001), .y(t0_010011001000));
wire t0_0100110010000, t0_0100110010001;
mixer mix_t0_010011001001 (.a(t0_0100110010010), .b(t0_0100110010011), .y(t0_010011001001));
wire t0_0100110010010, t0_0100110010011;
mixer mix_t0_01001100101 (.a(t0_010011001010), .b(t0_010011001011), .y(t0_01001100101));
wire t0_010011001010, t0_010011001011;
mixer mix_t0_010011001010 (.a(t0_0100110010100), .b(t0_0100110010101), .y(t0_010011001010));
wire t0_0100110010100, t0_0100110010101;
mixer mix_t0_010011001011 (.a(t0_0100110010110), .b(t0_0100110010111), .y(t0_010011001011));
wire t0_0100110010110, t0_0100110010111;
mixer mix_t0_0100110011 (.a(t0_01001100110), .b(t0_01001100111), .y(t0_0100110011));
wire t0_01001100110, t0_01001100111;
mixer mix_t0_01001100110 (.a(t0_010011001100), .b(t0_010011001101), .y(t0_01001100110));
wire t0_010011001100, t0_010011001101;
mixer mix_t0_010011001100 (.a(t0_0100110011000), .b(t0_0100110011001), .y(t0_010011001100));
wire t0_0100110011000, t0_0100110011001;
mixer mix_t0_010011001101 (.a(t0_0100110011010), .b(t0_0100110011011), .y(t0_010011001101));
wire t0_0100110011010, t0_0100110011011;
mixer mix_t0_01001100111 (.a(t0_010011001110), .b(t0_010011001111), .y(t0_01001100111));
wire t0_010011001110, t0_010011001111;
mixer mix_t0_010011001110 (.a(t0_0100110011100), .b(t0_0100110011101), .y(t0_010011001110));
wire t0_0100110011100, t0_0100110011101;
mixer mix_t0_010011001111 (.a(t0_0100110011110), .b(t0_0100110011111), .y(t0_010011001111));
wire t0_0100110011110, t0_0100110011111;
mixer mix_t0_01001101 (.a(t0_010011010), .b(t0_010011011), .y(t0_01001101));
wire t0_010011010, t0_010011011;
mixer mix_t0_010011010 (.a(t0_0100110100), .b(t0_0100110101), .y(t0_010011010));
wire t0_0100110100, t0_0100110101;
mixer mix_t0_0100110100 (.a(t0_01001101000), .b(t0_01001101001), .y(t0_0100110100));
wire t0_01001101000, t0_01001101001;
mixer mix_t0_01001101000 (.a(t0_010011010000), .b(t0_010011010001), .y(t0_01001101000));
wire t0_010011010000, t0_010011010001;
mixer mix_t0_010011010000 (.a(t0_0100110100000), .b(t0_0100110100001), .y(t0_010011010000));
wire t0_0100110100000, t0_0100110100001;
mixer mix_t0_010011010001 (.a(t0_0100110100010), .b(t0_0100110100011), .y(t0_010011010001));
wire t0_0100110100010, t0_0100110100011;
mixer mix_t0_01001101001 (.a(t0_010011010010), .b(t0_010011010011), .y(t0_01001101001));
wire t0_010011010010, t0_010011010011;
mixer mix_t0_010011010010 (.a(t0_0100110100100), .b(t0_0100110100101), .y(t0_010011010010));
wire t0_0100110100100, t0_0100110100101;
mixer mix_t0_010011010011 (.a(t0_0100110100110), .b(t0_0100110100111), .y(t0_010011010011));
wire t0_0100110100110, t0_0100110100111;
mixer mix_t0_0100110101 (.a(t0_01001101010), .b(t0_01001101011), .y(t0_0100110101));
wire t0_01001101010, t0_01001101011;
mixer mix_t0_01001101010 (.a(t0_010011010100), .b(t0_010011010101), .y(t0_01001101010));
wire t0_010011010100, t0_010011010101;
mixer mix_t0_010011010100 (.a(t0_0100110101000), .b(t0_0100110101001), .y(t0_010011010100));
wire t0_0100110101000, t0_0100110101001;
mixer mix_t0_010011010101 (.a(t0_0100110101010), .b(t0_0100110101011), .y(t0_010011010101));
wire t0_0100110101010, t0_0100110101011;
mixer mix_t0_01001101011 (.a(t0_010011010110), .b(t0_010011010111), .y(t0_01001101011));
wire t0_010011010110, t0_010011010111;
mixer mix_t0_010011010110 (.a(t0_0100110101100), .b(t0_0100110101101), .y(t0_010011010110));
wire t0_0100110101100, t0_0100110101101;
mixer mix_t0_010011010111 (.a(t0_0100110101110), .b(t0_0100110101111), .y(t0_010011010111));
wire t0_0100110101110, t0_0100110101111;
mixer mix_t0_010011011 (.a(t0_0100110110), .b(t0_0100110111), .y(t0_010011011));
wire t0_0100110110, t0_0100110111;
mixer mix_t0_0100110110 (.a(t0_01001101100), .b(t0_01001101101), .y(t0_0100110110));
wire t0_01001101100, t0_01001101101;
mixer mix_t0_01001101100 (.a(t0_010011011000), .b(t0_010011011001), .y(t0_01001101100));
wire t0_010011011000, t0_010011011001;
mixer mix_t0_010011011000 (.a(t0_0100110110000), .b(t0_0100110110001), .y(t0_010011011000));
wire t0_0100110110000, t0_0100110110001;
mixer mix_t0_010011011001 (.a(t0_0100110110010), .b(t0_0100110110011), .y(t0_010011011001));
wire t0_0100110110010, t0_0100110110011;
mixer mix_t0_01001101101 (.a(t0_010011011010), .b(t0_010011011011), .y(t0_01001101101));
wire t0_010011011010, t0_010011011011;
mixer mix_t0_010011011010 (.a(t0_0100110110100), .b(t0_0100110110101), .y(t0_010011011010));
wire t0_0100110110100, t0_0100110110101;
mixer mix_t0_010011011011 (.a(t0_0100110110110), .b(t0_0100110110111), .y(t0_010011011011));
wire t0_0100110110110, t0_0100110110111;
mixer mix_t0_0100110111 (.a(t0_01001101110), .b(t0_01001101111), .y(t0_0100110111));
wire t0_01001101110, t0_01001101111;
mixer mix_t0_01001101110 (.a(t0_010011011100), .b(t0_010011011101), .y(t0_01001101110));
wire t0_010011011100, t0_010011011101;
mixer mix_t0_010011011100 (.a(t0_0100110111000), .b(t0_0100110111001), .y(t0_010011011100));
wire t0_0100110111000, t0_0100110111001;
mixer mix_t0_010011011101 (.a(t0_0100110111010), .b(t0_0100110111011), .y(t0_010011011101));
wire t0_0100110111010, t0_0100110111011;
mixer mix_t0_01001101111 (.a(t0_010011011110), .b(t0_010011011111), .y(t0_01001101111));
wire t0_010011011110, t0_010011011111;
mixer mix_t0_010011011110 (.a(t0_0100110111100), .b(t0_0100110111101), .y(t0_010011011110));
wire t0_0100110111100, t0_0100110111101;
mixer mix_t0_010011011111 (.a(t0_0100110111110), .b(t0_0100110111111), .y(t0_010011011111));
wire t0_0100110111110, t0_0100110111111;
mixer mix_t0_0100111 (.a(t0_01001110), .b(t0_01001111), .y(t0_0100111));
wire t0_01001110, t0_01001111;
mixer mix_t0_01001110 (.a(t0_010011100), .b(t0_010011101), .y(t0_01001110));
wire t0_010011100, t0_010011101;
mixer mix_t0_010011100 (.a(t0_0100111000), .b(t0_0100111001), .y(t0_010011100));
wire t0_0100111000, t0_0100111001;
mixer mix_t0_0100111000 (.a(t0_01001110000), .b(t0_01001110001), .y(t0_0100111000));
wire t0_01001110000, t0_01001110001;
mixer mix_t0_01001110000 (.a(t0_010011100000), .b(t0_010011100001), .y(t0_01001110000));
wire t0_010011100000, t0_010011100001;
mixer mix_t0_010011100000 (.a(t0_0100111000000), .b(t0_0100111000001), .y(t0_010011100000));
wire t0_0100111000000, t0_0100111000001;
mixer mix_t0_010011100001 (.a(t0_0100111000010), .b(t0_0100111000011), .y(t0_010011100001));
wire t0_0100111000010, t0_0100111000011;
mixer mix_t0_01001110001 (.a(t0_010011100010), .b(t0_010011100011), .y(t0_01001110001));
wire t0_010011100010, t0_010011100011;
mixer mix_t0_010011100010 (.a(t0_0100111000100), .b(t0_0100111000101), .y(t0_010011100010));
wire t0_0100111000100, t0_0100111000101;
mixer mix_t0_010011100011 (.a(t0_0100111000110), .b(t0_0100111000111), .y(t0_010011100011));
wire t0_0100111000110, t0_0100111000111;
mixer mix_t0_0100111001 (.a(t0_01001110010), .b(t0_01001110011), .y(t0_0100111001));
wire t0_01001110010, t0_01001110011;
mixer mix_t0_01001110010 (.a(t0_010011100100), .b(t0_010011100101), .y(t0_01001110010));
wire t0_010011100100, t0_010011100101;
mixer mix_t0_010011100100 (.a(t0_0100111001000), .b(t0_0100111001001), .y(t0_010011100100));
wire t0_0100111001000, t0_0100111001001;
mixer mix_t0_010011100101 (.a(t0_0100111001010), .b(t0_0100111001011), .y(t0_010011100101));
wire t0_0100111001010, t0_0100111001011;
mixer mix_t0_01001110011 (.a(t0_010011100110), .b(t0_010011100111), .y(t0_01001110011));
wire t0_010011100110, t0_010011100111;
mixer mix_t0_010011100110 (.a(t0_0100111001100), .b(t0_0100111001101), .y(t0_010011100110));
wire t0_0100111001100, t0_0100111001101;
mixer mix_t0_010011100111 (.a(t0_0100111001110), .b(t0_0100111001111), .y(t0_010011100111));
wire t0_0100111001110, t0_0100111001111;
mixer mix_t0_010011101 (.a(t0_0100111010), .b(t0_0100111011), .y(t0_010011101));
wire t0_0100111010, t0_0100111011;
mixer mix_t0_0100111010 (.a(t0_01001110100), .b(t0_01001110101), .y(t0_0100111010));
wire t0_01001110100, t0_01001110101;
mixer mix_t0_01001110100 (.a(t0_010011101000), .b(t0_010011101001), .y(t0_01001110100));
wire t0_010011101000, t0_010011101001;
mixer mix_t0_010011101000 (.a(t0_0100111010000), .b(t0_0100111010001), .y(t0_010011101000));
wire t0_0100111010000, t0_0100111010001;
mixer mix_t0_010011101001 (.a(t0_0100111010010), .b(t0_0100111010011), .y(t0_010011101001));
wire t0_0100111010010, t0_0100111010011;
mixer mix_t0_01001110101 (.a(t0_010011101010), .b(t0_010011101011), .y(t0_01001110101));
wire t0_010011101010, t0_010011101011;
mixer mix_t0_010011101010 (.a(t0_0100111010100), .b(t0_0100111010101), .y(t0_010011101010));
wire t0_0100111010100, t0_0100111010101;
mixer mix_t0_010011101011 (.a(t0_0100111010110), .b(t0_0100111010111), .y(t0_010011101011));
wire t0_0100111010110, t0_0100111010111;
mixer mix_t0_0100111011 (.a(t0_01001110110), .b(t0_01001110111), .y(t0_0100111011));
wire t0_01001110110, t0_01001110111;
mixer mix_t0_01001110110 (.a(t0_010011101100), .b(t0_010011101101), .y(t0_01001110110));
wire t0_010011101100, t0_010011101101;
mixer mix_t0_010011101100 (.a(t0_0100111011000), .b(t0_0100111011001), .y(t0_010011101100));
wire t0_0100111011000, t0_0100111011001;
mixer mix_t0_010011101101 (.a(t0_0100111011010), .b(t0_0100111011011), .y(t0_010011101101));
wire t0_0100111011010, t0_0100111011011;
mixer mix_t0_01001110111 (.a(t0_010011101110), .b(t0_010011101111), .y(t0_01001110111));
wire t0_010011101110, t0_010011101111;
mixer mix_t0_010011101110 (.a(t0_0100111011100), .b(t0_0100111011101), .y(t0_010011101110));
wire t0_0100111011100, t0_0100111011101;
mixer mix_t0_010011101111 (.a(t0_0100111011110), .b(t0_0100111011111), .y(t0_010011101111));
wire t0_0100111011110, t0_0100111011111;
mixer mix_t0_01001111 (.a(t0_010011110), .b(t0_010011111), .y(t0_01001111));
wire t0_010011110, t0_010011111;
mixer mix_t0_010011110 (.a(t0_0100111100), .b(t0_0100111101), .y(t0_010011110));
wire t0_0100111100, t0_0100111101;
mixer mix_t0_0100111100 (.a(t0_01001111000), .b(t0_01001111001), .y(t0_0100111100));
wire t0_01001111000, t0_01001111001;
mixer mix_t0_01001111000 (.a(t0_010011110000), .b(t0_010011110001), .y(t0_01001111000));
wire t0_010011110000, t0_010011110001;
mixer mix_t0_010011110000 (.a(t0_0100111100000), .b(t0_0100111100001), .y(t0_010011110000));
wire t0_0100111100000, t0_0100111100001;
mixer mix_t0_010011110001 (.a(t0_0100111100010), .b(t0_0100111100011), .y(t0_010011110001));
wire t0_0100111100010, t0_0100111100011;
mixer mix_t0_01001111001 (.a(t0_010011110010), .b(t0_010011110011), .y(t0_01001111001));
wire t0_010011110010, t0_010011110011;
mixer mix_t0_010011110010 (.a(t0_0100111100100), .b(t0_0100111100101), .y(t0_010011110010));
wire t0_0100111100100, t0_0100111100101;
mixer mix_t0_010011110011 (.a(t0_0100111100110), .b(t0_0100111100111), .y(t0_010011110011));
wire t0_0100111100110, t0_0100111100111;
mixer mix_t0_0100111101 (.a(t0_01001111010), .b(t0_01001111011), .y(t0_0100111101));
wire t0_01001111010, t0_01001111011;
mixer mix_t0_01001111010 (.a(t0_010011110100), .b(t0_010011110101), .y(t0_01001111010));
wire t0_010011110100, t0_010011110101;
mixer mix_t0_010011110100 (.a(t0_0100111101000), .b(t0_0100111101001), .y(t0_010011110100));
wire t0_0100111101000, t0_0100111101001;
mixer mix_t0_010011110101 (.a(t0_0100111101010), .b(t0_0100111101011), .y(t0_010011110101));
wire t0_0100111101010, t0_0100111101011;
mixer mix_t0_01001111011 (.a(t0_010011110110), .b(t0_010011110111), .y(t0_01001111011));
wire t0_010011110110, t0_010011110111;
mixer mix_t0_010011110110 (.a(t0_0100111101100), .b(t0_0100111101101), .y(t0_010011110110));
wire t0_0100111101100, t0_0100111101101;
mixer mix_t0_010011110111 (.a(t0_0100111101110), .b(t0_0100111101111), .y(t0_010011110111));
wire t0_0100111101110, t0_0100111101111;
mixer mix_t0_010011111 (.a(t0_0100111110), .b(t0_0100111111), .y(t0_010011111));
wire t0_0100111110, t0_0100111111;
mixer mix_t0_0100111110 (.a(t0_01001111100), .b(t0_01001111101), .y(t0_0100111110));
wire t0_01001111100, t0_01001111101;
mixer mix_t0_01001111100 (.a(t0_010011111000), .b(t0_010011111001), .y(t0_01001111100));
wire t0_010011111000, t0_010011111001;
mixer mix_t0_010011111000 (.a(t0_0100111110000), .b(t0_0100111110001), .y(t0_010011111000));
wire t0_0100111110000, t0_0100111110001;
mixer mix_t0_010011111001 (.a(t0_0100111110010), .b(t0_0100111110011), .y(t0_010011111001));
wire t0_0100111110010, t0_0100111110011;
mixer mix_t0_01001111101 (.a(t0_010011111010), .b(t0_010011111011), .y(t0_01001111101));
wire t0_010011111010, t0_010011111011;
mixer mix_t0_010011111010 (.a(t0_0100111110100), .b(t0_0100111110101), .y(t0_010011111010));
wire t0_0100111110100, t0_0100111110101;
mixer mix_t0_010011111011 (.a(t0_0100111110110), .b(t0_0100111110111), .y(t0_010011111011));
wire t0_0100111110110, t0_0100111110111;
mixer mix_t0_0100111111 (.a(t0_01001111110), .b(t0_01001111111), .y(t0_0100111111));
wire t0_01001111110, t0_01001111111;
mixer mix_t0_01001111110 (.a(t0_010011111100), .b(t0_010011111101), .y(t0_01001111110));
wire t0_010011111100, t0_010011111101;
mixer mix_t0_010011111100 (.a(t0_0100111111000), .b(t0_0100111111001), .y(t0_010011111100));
wire t0_0100111111000, t0_0100111111001;
mixer mix_t0_010011111101 (.a(t0_0100111111010), .b(t0_0100111111011), .y(t0_010011111101));
wire t0_0100111111010, t0_0100111111011;
mixer mix_t0_01001111111 (.a(t0_010011111110), .b(t0_010011111111), .y(t0_01001111111));
wire t0_010011111110, t0_010011111111;
mixer mix_t0_010011111110 (.a(t0_0100111111100), .b(t0_0100111111101), .y(t0_010011111110));
wire t0_0100111111100, t0_0100111111101;
mixer mix_t0_010011111111 (.a(t0_0100111111110), .b(t0_0100111111111), .y(t0_010011111111));
wire t0_0100111111110, t0_0100111111111;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_010100 (.a(t0_0101000), .b(t0_0101001), .y(t0_010100));
wire t0_0101000, t0_0101001;
mixer mix_t0_0101000 (.a(t0_01010000), .b(t0_01010001), .y(t0_0101000));
wire t0_01010000, t0_01010001;
mixer mix_t0_01010000 (.a(t0_010100000), .b(t0_010100001), .y(t0_01010000));
wire t0_010100000, t0_010100001;
mixer mix_t0_010100000 (.a(t0_0101000000), .b(t0_0101000001), .y(t0_010100000));
wire t0_0101000000, t0_0101000001;
mixer mix_t0_0101000000 (.a(t0_01010000000), .b(t0_01010000001), .y(t0_0101000000));
wire t0_01010000000, t0_01010000001;
mixer mix_t0_01010000000 (.a(t0_010100000000), .b(t0_010100000001), .y(t0_01010000000));
wire t0_010100000000, t0_010100000001;
mixer mix_t0_010100000000 (.a(t0_0101000000000), .b(t0_0101000000001), .y(t0_010100000000));
wire t0_0101000000000, t0_0101000000001;
mixer mix_t0_010100000001 (.a(t0_0101000000010), .b(t0_0101000000011), .y(t0_010100000001));
wire t0_0101000000010, t0_0101000000011;
mixer mix_t0_01010000001 (.a(t0_010100000010), .b(t0_010100000011), .y(t0_01010000001));
wire t0_010100000010, t0_010100000011;
mixer mix_t0_010100000010 (.a(t0_0101000000100), .b(t0_0101000000101), .y(t0_010100000010));
wire t0_0101000000100, t0_0101000000101;
mixer mix_t0_010100000011 (.a(t0_0101000000110), .b(t0_0101000000111), .y(t0_010100000011));
wire t0_0101000000110, t0_0101000000111;
mixer mix_t0_0101000001 (.a(t0_01010000010), .b(t0_01010000011), .y(t0_0101000001));
wire t0_01010000010, t0_01010000011;
mixer mix_t0_01010000010 (.a(t0_010100000100), .b(t0_010100000101), .y(t0_01010000010));
wire t0_010100000100, t0_010100000101;
mixer mix_t0_010100000100 (.a(t0_0101000001000), .b(t0_0101000001001), .y(t0_010100000100));
wire t0_0101000001000, t0_0101000001001;
mixer mix_t0_010100000101 (.a(t0_0101000001010), .b(t0_0101000001011), .y(t0_010100000101));
wire t0_0101000001010, t0_0101000001011;
mixer mix_t0_01010000011 (.a(t0_010100000110), .b(t0_010100000111), .y(t0_01010000011));
wire t0_010100000110, t0_010100000111;
mixer mix_t0_010100000110 (.a(t0_0101000001100), .b(t0_0101000001101), .y(t0_010100000110));
wire t0_0101000001100, t0_0101000001101;
mixer mix_t0_010100000111 (.a(t0_0101000001110), .b(t0_0101000001111), .y(t0_010100000111));
wire t0_0101000001110, t0_0101000001111;
mixer mix_t0_010100001 (.a(t0_0101000010), .b(t0_0101000011), .y(t0_010100001));
wire t0_0101000010, t0_0101000011;
mixer mix_t0_0101000010 (.a(t0_01010000100), .b(t0_01010000101), .y(t0_0101000010));
wire t0_01010000100, t0_01010000101;
mixer mix_t0_01010000100 (.a(t0_010100001000), .b(t0_010100001001), .y(t0_01010000100));
wire t0_010100001000, t0_010100001001;
mixer mix_t0_010100001000 (.a(t0_0101000010000), .b(t0_0101000010001), .y(t0_010100001000));
wire t0_0101000010000, t0_0101000010001;
mixer mix_t0_010100001001 (.a(t0_0101000010010), .b(t0_0101000010011), .y(t0_010100001001));
wire t0_0101000010010, t0_0101000010011;
mixer mix_t0_01010000101 (.a(t0_010100001010), .b(t0_010100001011), .y(t0_01010000101));
wire t0_010100001010, t0_010100001011;
mixer mix_t0_010100001010 (.a(t0_0101000010100), .b(t0_0101000010101), .y(t0_010100001010));
wire t0_0101000010100, t0_0101000010101;
mixer mix_t0_010100001011 (.a(t0_0101000010110), .b(t0_0101000010111), .y(t0_010100001011));
wire t0_0101000010110, t0_0101000010111;
mixer mix_t0_0101000011 (.a(t0_01010000110), .b(t0_01010000111), .y(t0_0101000011));
wire t0_01010000110, t0_01010000111;
mixer mix_t0_01010000110 (.a(t0_010100001100), .b(t0_010100001101), .y(t0_01010000110));
wire t0_010100001100, t0_010100001101;
mixer mix_t0_010100001100 (.a(t0_0101000011000), .b(t0_0101000011001), .y(t0_010100001100));
wire t0_0101000011000, t0_0101000011001;
mixer mix_t0_010100001101 (.a(t0_0101000011010), .b(t0_0101000011011), .y(t0_010100001101));
wire t0_0101000011010, t0_0101000011011;
mixer mix_t0_01010000111 (.a(t0_010100001110), .b(t0_010100001111), .y(t0_01010000111));
wire t0_010100001110, t0_010100001111;
mixer mix_t0_010100001110 (.a(t0_0101000011100), .b(t0_0101000011101), .y(t0_010100001110));
wire t0_0101000011100, t0_0101000011101;
mixer mix_t0_010100001111 (.a(t0_0101000011110), .b(t0_0101000011111), .y(t0_010100001111));
wire t0_0101000011110, t0_0101000011111;
mixer mix_t0_01010001 (.a(t0_010100010), .b(t0_010100011), .y(t0_01010001));
wire t0_010100010, t0_010100011;
mixer mix_t0_010100010 (.a(t0_0101000100), .b(t0_0101000101), .y(t0_010100010));
wire t0_0101000100, t0_0101000101;
mixer mix_t0_0101000100 (.a(t0_01010001000), .b(t0_01010001001), .y(t0_0101000100));
wire t0_01010001000, t0_01010001001;
mixer mix_t0_01010001000 (.a(t0_010100010000), .b(t0_010100010001), .y(t0_01010001000));
wire t0_010100010000, t0_010100010001;
mixer mix_t0_010100010000 (.a(t0_0101000100000), .b(t0_0101000100001), .y(t0_010100010000));
wire t0_0101000100000, t0_0101000100001;
mixer mix_t0_010100010001 (.a(t0_0101000100010), .b(t0_0101000100011), .y(t0_010100010001));
wire t0_0101000100010, t0_0101000100011;
mixer mix_t0_01010001001 (.a(t0_010100010010), .b(t0_010100010011), .y(t0_01010001001));
wire t0_010100010010, t0_010100010011;
mixer mix_t0_010100010010 (.a(t0_0101000100100), .b(t0_0101000100101), .y(t0_010100010010));
wire t0_0101000100100, t0_0101000100101;
mixer mix_t0_010100010011 (.a(t0_0101000100110), .b(t0_0101000100111), .y(t0_010100010011));
wire t0_0101000100110, t0_0101000100111;
mixer mix_t0_0101000101 (.a(t0_01010001010), .b(t0_01010001011), .y(t0_0101000101));
wire t0_01010001010, t0_01010001011;
mixer mix_t0_01010001010 (.a(t0_010100010100), .b(t0_010100010101), .y(t0_01010001010));
wire t0_010100010100, t0_010100010101;
mixer mix_t0_010100010100 (.a(t0_0101000101000), .b(t0_0101000101001), .y(t0_010100010100));
wire t0_0101000101000, t0_0101000101001;
mixer mix_t0_010100010101 (.a(t0_0101000101010), .b(t0_0101000101011), .y(t0_010100010101));
wire t0_0101000101010, t0_0101000101011;
mixer mix_t0_01010001011 (.a(t0_010100010110), .b(t0_010100010111), .y(t0_01010001011));
wire t0_010100010110, t0_010100010111;
mixer mix_t0_010100010110 (.a(t0_0101000101100), .b(t0_0101000101101), .y(t0_010100010110));
wire t0_0101000101100, t0_0101000101101;
mixer mix_t0_010100010111 (.a(t0_0101000101110), .b(t0_0101000101111), .y(t0_010100010111));
wire t0_0101000101110, t0_0101000101111;
mixer mix_t0_010100011 (.a(t0_0101000110), .b(t0_0101000111), .y(t0_010100011));
wire t0_0101000110, t0_0101000111;
mixer mix_t0_0101000110 (.a(t0_01010001100), .b(t0_01010001101), .y(t0_0101000110));
wire t0_01010001100, t0_01010001101;
mixer mix_t0_01010001100 (.a(t0_010100011000), .b(t0_010100011001), .y(t0_01010001100));
wire t0_010100011000, t0_010100011001;
mixer mix_t0_010100011000 (.a(t0_0101000110000), .b(t0_0101000110001), .y(t0_010100011000));
wire t0_0101000110000, t0_0101000110001;
mixer mix_t0_010100011001 (.a(t0_0101000110010), .b(t0_0101000110011), .y(t0_010100011001));
wire t0_0101000110010, t0_0101000110011;
mixer mix_t0_01010001101 (.a(t0_010100011010), .b(t0_010100011011), .y(t0_01010001101));
wire t0_010100011010, t0_010100011011;
mixer mix_t0_010100011010 (.a(t0_0101000110100), .b(t0_0101000110101), .y(t0_010100011010));
wire t0_0101000110100, t0_0101000110101;
mixer mix_t0_010100011011 (.a(t0_0101000110110), .b(t0_0101000110111), .y(t0_010100011011));
wire t0_0101000110110, t0_0101000110111;
mixer mix_t0_0101000111 (.a(t0_01010001110), .b(t0_01010001111), .y(t0_0101000111));
wire t0_01010001110, t0_01010001111;
mixer mix_t0_01010001110 (.a(t0_010100011100), .b(t0_010100011101), .y(t0_01010001110));
wire t0_010100011100, t0_010100011101;
mixer mix_t0_010100011100 (.a(t0_0101000111000), .b(t0_0101000111001), .y(t0_010100011100));
wire t0_0101000111000, t0_0101000111001;
mixer mix_t0_010100011101 (.a(t0_0101000111010), .b(t0_0101000111011), .y(t0_010100011101));
wire t0_0101000111010, t0_0101000111011;
mixer mix_t0_01010001111 (.a(t0_010100011110), .b(t0_010100011111), .y(t0_01010001111));
wire t0_010100011110, t0_010100011111;
mixer mix_t0_010100011110 (.a(t0_0101000111100), .b(t0_0101000111101), .y(t0_010100011110));
wire t0_0101000111100, t0_0101000111101;
mixer mix_t0_010100011111 (.a(t0_0101000111110), .b(t0_0101000111111), .y(t0_010100011111));
wire t0_0101000111110, t0_0101000111111;
mixer mix_t0_0101001 (.a(t0_01010010), .b(t0_01010011), .y(t0_0101001));
wire t0_01010010, t0_01010011;
mixer mix_t0_01010010 (.a(t0_010100100), .b(t0_010100101), .y(t0_01010010));
wire t0_010100100, t0_010100101;
mixer mix_t0_010100100 (.a(t0_0101001000), .b(t0_0101001001), .y(t0_010100100));
wire t0_0101001000, t0_0101001001;
mixer mix_t0_0101001000 (.a(t0_01010010000), .b(t0_01010010001), .y(t0_0101001000));
wire t0_01010010000, t0_01010010001;
mixer mix_t0_01010010000 (.a(t0_010100100000), .b(t0_010100100001), .y(t0_01010010000));
wire t0_010100100000, t0_010100100001;
mixer mix_t0_010100100000 (.a(t0_0101001000000), .b(t0_0101001000001), .y(t0_010100100000));
wire t0_0101001000000, t0_0101001000001;
mixer mix_t0_010100100001 (.a(t0_0101001000010), .b(t0_0101001000011), .y(t0_010100100001));
wire t0_0101001000010, t0_0101001000011;
mixer mix_t0_01010010001 (.a(t0_010100100010), .b(t0_010100100011), .y(t0_01010010001));
wire t0_010100100010, t0_010100100011;
mixer mix_t0_010100100010 (.a(t0_0101001000100), .b(t0_0101001000101), .y(t0_010100100010));
wire t0_0101001000100, t0_0101001000101;
mixer mix_t0_010100100011 (.a(t0_0101001000110), .b(t0_0101001000111), .y(t0_010100100011));
wire t0_0101001000110, t0_0101001000111;
mixer mix_t0_0101001001 (.a(t0_01010010010), .b(t0_01010010011), .y(t0_0101001001));
wire t0_01010010010, t0_01010010011;
mixer mix_t0_01010010010 (.a(t0_010100100100), .b(t0_010100100101), .y(t0_01010010010));
wire t0_010100100100, t0_010100100101;
mixer mix_t0_010100100100 (.a(t0_0101001001000), .b(t0_0101001001001), .y(t0_010100100100));
wire t0_0101001001000, t0_0101001001001;
mixer mix_t0_010100100101 (.a(t0_0101001001010), .b(t0_0101001001011), .y(t0_010100100101));
wire t0_0101001001010, t0_0101001001011;
mixer mix_t0_01010010011 (.a(t0_010100100110), .b(t0_010100100111), .y(t0_01010010011));
wire t0_010100100110, t0_010100100111;
mixer mix_t0_010100100110 (.a(t0_0101001001100), .b(t0_0101001001101), .y(t0_010100100110));
wire t0_0101001001100, t0_0101001001101;
mixer mix_t0_010100100111 (.a(t0_0101001001110), .b(t0_0101001001111), .y(t0_010100100111));
wire t0_0101001001110, t0_0101001001111;
mixer mix_t0_010100101 (.a(t0_0101001010), .b(t0_0101001011), .y(t0_010100101));
wire t0_0101001010, t0_0101001011;
mixer mix_t0_0101001010 (.a(t0_01010010100), .b(t0_01010010101), .y(t0_0101001010));
wire t0_01010010100, t0_01010010101;
mixer mix_t0_01010010100 (.a(t0_010100101000), .b(t0_010100101001), .y(t0_01010010100));
wire t0_010100101000, t0_010100101001;
mixer mix_t0_010100101000 (.a(t0_0101001010000), .b(t0_0101001010001), .y(t0_010100101000));
wire t0_0101001010000, t0_0101001010001;
mixer mix_t0_010100101001 (.a(t0_0101001010010), .b(t0_0101001010011), .y(t0_010100101001));
wire t0_0101001010010, t0_0101001010011;
mixer mix_t0_01010010101 (.a(t0_010100101010), .b(t0_010100101011), .y(t0_01010010101));
wire t0_010100101010, t0_010100101011;
mixer mix_t0_010100101010 (.a(t0_0101001010100), .b(t0_0101001010101), .y(t0_010100101010));
wire t0_0101001010100, t0_0101001010101;
mixer mix_t0_010100101011 (.a(t0_0101001010110), .b(t0_0101001010111), .y(t0_010100101011));
wire t0_0101001010110, t0_0101001010111;
mixer mix_t0_0101001011 (.a(t0_01010010110), .b(t0_01010010111), .y(t0_0101001011));
wire t0_01010010110, t0_01010010111;
mixer mix_t0_01010010110 (.a(t0_010100101100), .b(t0_010100101101), .y(t0_01010010110));
wire t0_010100101100, t0_010100101101;
mixer mix_t0_010100101100 (.a(t0_0101001011000), .b(t0_0101001011001), .y(t0_010100101100));
wire t0_0101001011000, t0_0101001011001;
mixer mix_t0_010100101101 (.a(t0_0101001011010), .b(t0_0101001011011), .y(t0_010100101101));
wire t0_0101001011010, t0_0101001011011;
mixer mix_t0_01010010111 (.a(t0_010100101110), .b(t0_010100101111), .y(t0_01010010111));
wire t0_010100101110, t0_010100101111;
mixer mix_t0_010100101110 (.a(t0_0101001011100), .b(t0_0101001011101), .y(t0_010100101110));
wire t0_0101001011100, t0_0101001011101;
mixer mix_t0_010100101111 (.a(t0_0101001011110), .b(t0_0101001011111), .y(t0_010100101111));
wire t0_0101001011110, t0_0101001011111;
mixer mix_t0_01010011 (.a(t0_010100110), .b(t0_010100111), .y(t0_01010011));
wire t0_010100110, t0_010100111;
mixer mix_t0_010100110 (.a(t0_0101001100), .b(t0_0101001101), .y(t0_010100110));
wire t0_0101001100, t0_0101001101;
mixer mix_t0_0101001100 (.a(t0_01010011000), .b(t0_01010011001), .y(t0_0101001100));
wire t0_01010011000, t0_01010011001;
mixer mix_t0_01010011000 (.a(t0_010100110000), .b(t0_010100110001), .y(t0_01010011000));
wire t0_010100110000, t0_010100110001;
mixer mix_t0_010100110000 (.a(t0_0101001100000), .b(t0_0101001100001), .y(t0_010100110000));
wire t0_0101001100000, t0_0101001100001;
mixer mix_t0_010100110001 (.a(t0_0101001100010), .b(t0_0101001100011), .y(t0_010100110001));
wire t0_0101001100010, t0_0101001100011;
mixer mix_t0_01010011001 (.a(t0_010100110010), .b(t0_010100110011), .y(t0_01010011001));
wire t0_010100110010, t0_010100110011;
mixer mix_t0_010100110010 (.a(t0_0101001100100), .b(t0_0101001100101), .y(t0_010100110010));
wire t0_0101001100100, t0_0101001100101;
mixer mix_t0_010100110011 (.a(t0_0101001100110), .b(t0_0101001100111), .y(t0_010100110011));
wire t0_0101001100110, t0_0101001100111;
mixer mix_t0_0101001101 (.a(t0_01010011010), .b(t0_01010011011), .y(t0_0101001101));
wire t0_01010011010, t0_01010011011;
mixer mix_t0_01010011010 (.a(t0_010100110100), .b(t0_010100110101), .y(t0_01010011010));
wire t0_010100110100, t0_010100110101;
mixer mix_t0_010100110100 (.a(t0_0101001101000), .b(t0_0101001101001), .y(t0_010100110100));
wire t0_0101001101000, t0_0101001101001;
mixer mix_t0_010100110101 (.a(t0_0101001101010), .b(t0_0101001101011), .y(t0_010100110101));
wire t0_0101001101010, t0_0101001101011;
mixer mix_t0_01010011011 (.a(t0_010100110110), .b(t0_010100110111), .y(t0_01010011011));
wire t0_010100110110, t0_010100110111;
mixer mix_t0_010100110110 (.a(t0_0101001101100), .b(t0_0101001101101), .y(t0_010100110110));
wire t0_0101001101100, t0_0101001101101;
mixer mix_t0_010100110111 (.a(t0_0101001101110), .b(t0_0101001101111), .y(t0_010100110111));
wire t0_0101001101110, t0_0101001101111;
mixer mix_t0_010100111 (.a(t0_0101001110), .b(t0_0101001111), .y(t0_010100111));
wire t0_0101001110, t0_0101001111;
mixer mix_t0_0101001110 (.a(t0_01010011100), .b(t0_01010011101), .y(t0_0101001110));
wire t0_01010011100, t0_01010011101;
mixer mix_t0_01010011100 (.a(t0_010100111000), .b(t0_010100111001), .y(t0_01010011100));
wire t0_010100111000, t0_010100111001;
mixer mix_t0_010100111000 (.a(t0_0101001110000), .b(t0_0101001110001), .y(t0_010100111000));
wire t0_0101001110000, t0_0101001110001;
mixer mix_t0_010100111001 (.a(t0_0101001110010), .b(t0_0101001110011), .y(t0_010100111001));
wire t0_0101001110010, t0_0101001110011;
mixer mix_t0_01010011101 (.a(t0_010100111010), .b(t0_010100111011), .y(t0_01010011101));
wire t0_010100111010, t0_010100111011;
mixer mix_t0_010100111010 (.a(t0_0101001110100), .b(t0_0101001110101), .y(t0_010100111010));
wire t0_0101001110100, t0_0101001110101;
mixer mix_t0_010100111011 (.a(t0_0101001110110), .b(t0_0101001110111), .y(t0_010100111011));
wire t0_0101001110110, t0_0101001110111;
mixer mix_t0_0101001111 (.a(t0_01010011110), .b(t0_01010011111), .y(t0_0101001111));
wire t0_01010011110, t0_01010011111;
mixer mix_t0_01010011110 (.a(t0_010100111100), .b(t0_010100111101), .y(t0_01010011110));
wire t0_010100111100, t0_010100111101;
mixer mix_t0_010100111100 (.a(t0_0101001111000), .b(t0_0101001111001), .y(t0_010100111100));
wire t0_0101001111000, t0_0101001111001;
mixer mix_t0_010100111101 (.a(t0_0101001111010), .b(t0_0101001111011), .y(t0_010100111101));
wire t0_0101001111010, t0_0101001111011;
mixer mix_t0_01010011111 (.a(t0_010100111110), .b(t0_010100111111), .y(t0_01010011111));
wire t0_010100111110, t0_010100111111;
mixer mix_t0_010100111110 (.a(t0_0101001111100), .b(t0_0101001111101), .y(t0_010100111110));
wire t0_0101001111100, t0_0101001111101;
mixer mix_t0_010100111111 (.a(t0_0101001111110), .b(t0_0101001111111), .y(t0_010100111111));
wire t0_0101001111110, t0_0101001111111;
mixer mix_t0_010101 (.a(t0_0101010), .b(t0_0101011), .y(t0_010101));
wire t0_0101010, t0_0101011;
mixer mix_t0_0101010 (.a(t0_01010100), .b(t0_01010101), .y(t0_0101010));
wire t0_01010100, t0_01010101;
mixer mix_t0_01010100 (.a(t0_010101000), .b(t0_010101001), .y(t0_01010100));
wire t0_010101000, t0_010101001;
mixer mix_t0_010101000 (.a(t0_0101010000), .b(t0_0101010001), .y(t0_010101000));
wire t0_0101010000, t0_0101010001;
mixer mix_t0_0101010000 (.a(t0_01010100000), .b(t0_01010100001), .y(t0_0101010000));
wire t0_01010100000, t0_01010100001;
mixer mix_t0_01010100000 (.a(t0_010101000000), .b(t0_010101000001), .y(t0_01010100000));
wire t0_010101000000, t0_010101000001;
mixer mix_t0_010101000000 (.a(t0_0101010000000), .b(t0_0101010000001), .y(t0_010101000000));
wire t0_0101010000000, t0_0101010000001;
mixer mix_t0_010101000001 (.a(t0_0101010000010), .b(t0_0101010000011), .y(t0_010101000001));
wire t0_0101010000010, t0_0101010000011;
mixer mix_t0_01010100001 (.a(t0_010101000010), .b(t0_010101000011), .y(t0_01010100001));
wire t0_010101000010, t0_010101000011;
mixer mix_t0_010101000010 (.a(t0_0101010000100), .b(t0_0101010000101), .y(t0_010101000010));
wire t0_0101010000100, t0_0101010000101;
mixer mix_t0_010101000011 (.a(t0_0101010000110), .b(t0_0101010000111), .y(t0_010101000011));
wire t0_0101010000110, t0_0101010000111;
mixer mix_t0_0101010001 (.a(t0_01010100010), .b(t0_01010100011), .y(t0_0101010001));
wire t0_01010100010, t0_01010100011;
mixer mix_t0_01010100010 (.a(t0_010101000100), .b(t0_010101000101), .y(t0_01010100010));
wire t0_010101000100, t0_010101000101;
mixer mix_t0_010101000100 (.a(t0_0101010001000), .b(t0_0101010001001), .y(t0_010101000100));
wire t0_0101010001000, t0_0101010001001;
mixer mix_t0_010101000101 (.a(t0_0101010001010), .b(t0_0101010001011), .y(t0_010101000101));
wire t0_0101010001010, t0_0101010001011;
mixer mix_t0_01010100011 (.a(t0_010101000110), .b(t0_010101000111), .y(t0_01010100011));
wire t0_010101000110, t0_010101000111;
mixer mix_t0_010101000110 (.a(t0_0101010001100), .b(t0_0101010001101), .y(t0_010101000110));
wire t0_0101010001100, t0_0101010001101;
mixer mix_t0_010101000111 (.a(t0_0101010001110), .b(t0_0101010001111), .y(t0_010101000111));
wire t0_0101010001110, t0_0101010001111;
mixer mix_t0_010101001 (.a(t0_0101010010), .b(t0_0101010011), .y(t0_010101001));
wire t0_0101010010, t0_0101010011;
mixer mix_t0_0101010010 (.a(t0_01010100100), .b(t0_01010100101), .y(t0_0101010010));
wire t0_01010100100, t0_01010100101;
mixer mix_t0_01010100100 (.a(t0_010101001000), .b(t0_010101001001), .y(t0_01010100100));
wire t0_010101001000, t0_010101001001;
mixer mix_t0_010101001000 (.a(t0_0101010010000), .b(t0_0101010010001), .y(t0_010101001000));
wire t0_0101010010000, t0_0101010010001;
mixer mix_t0_010101001001 (.a(t0_0101010010010), .b(t0_0101010010011), .y(t0_010101001001));
wire t0_0101010010010, t0_0101010010011;
mixer mix_t0_01010100101 (.a(t0_010101001010), .b(t0_010101001011), .y(t0_01010100101));
wire t0_010101001010, t0_010101001011;
mixer mix_t0_010101001010 (.a(t0_0101010010100), .b(t0_0101010010101), .y(t0_010101001010));
wire t0_0101010010100, t0_0101010010101;
mixer mix_t0_010101001011 (.a(t0_0101010010110), .b(t0_0101010010111), .y(t0_010101001011));
wire t0_0101010010110, t0_0101010010111;
mixer mix_t0_0101010011 (.a(t0_01010100110), .b(t0_01010100111), .y(t0_0101010011));
wire t0_01010100110, t0_01010100111;
mixer mix_t0_01010100110 (.a(t0_010101001100), .b(t0_010101001101), .y(t0_01010100110));
wire t0_010101001100, t0_010101001101;
mixer mix_t0_010101001100 (.a(t0_0101010011000), .b(t0_0101010011001), .y(t0_010101001100));
wire t0_0101010011000, t0_0101010011001;
mixer mix_t0_010101001101 (.a(t0_0101010011010), .b(t0_0101010011011), .y(t0_010101001101));
wire t0_0101010011010, t0_0101010011011;
mixer mix_t0_01010100111 (.a(t0_010101001110), .b(t0_010101001111), .y(t0_01010100111));
wire t0_010101001110, t0_010101001111;
mixer mix_t0_010101001110 (.a(t0_0101010011100), .b(t0_0101010011101), .y(t0_010101001110));
wire t0_0101010011100, t0_0101010011101;
mixer mix_t0_010101001111 (.a(t0_0101010011110), .b(t0_0101010011111), .y(t0_010101001111));
wire t0_0101010011110, t0_0101010011111;
mixer mix_t0_01010101 (.a(t0_010101010), .b(t0_010101011), .y(t0_01010101));
wire t0_010101010, t0_010101011;
mixer mix_t0_010101010 (.a(t0_0101010100), .b(t0_0101010101), .y(t0_010101010));
wire t0_0101010100, t0_0101010101;
mixer mix_t0_0101010100 (.a(t0_01010101000), .b(t0_01010101001), .y(t0_0101010100));
wire t0_01010101000, t0_01010101001;
mixer mix_t0_01010101000 (.a(t0_010101010000), .b(t0_010101010001), .y(t0_01010101000));
wire t0_010101010000, t0_010101010001;
mixer mix_t0_010101010000 (.a(t0_0101010100000), .b(t0_0101010100001), .y(t0_010101010000));
wire t0_0101010100000, t0_0101010100001;
mixer mix_t0_010101010001 (.a(t0_0101010100010), .b(t0_0101010100011), .y(t0_010101010001));
wire t0_0101010100010, t0_0101010100011;
mixer mix_t0_01010101001 (.a(t0_010101010010), .b(t0_010101010011), .y(t0_01010101001));
wire t0_010101010010, t0_010101010011;
mixer mix_t0_010101010010 (.a(t0_0101010100100), .b(t0_0101010100101), .y(t0_010101010010));
wire t0_0101010100100, t0_0101010100101;
mixer mix_t0_010101010011 (.a(t0_0101010100110), .b(t0_0101010100111), .y(t0_010101010011));
wire t0_0101010100110, t0_0101010100111;
mixer mix_t0_0101010101 (.a(t0_01010101010), .b(t0_01010101011), .y(t0_0101010101));
wire t0_01010101010, t0_01010101011;
mixer mix_t0_01010101010 (.a(t0_010101010100), .b(t0_010101010101), .y(t0_01010101010));
wire t0_010101010100, t0_010101010101;
mixer mix_t0_010101010100 (.a(t0_0101010101000), .b(t0_0101010101001), .y(t0_010101010100));
wire t0_0101010101000, t0_0101010101001;
mixer mix_t0_010101010101 (.a(t0_0101010101010), .b(t0_0101010101011), .y(t0_010101010101));
wire t0_0101010101010, t0_0101010101011;
mixer mix_t0_01010101011 (.a(t0_010101010110), .b(t0_010101010111), .y(t0_01010101011));
wire t0_010101010110, t0_010101010111;
mixer mix_t0_010101010110 (.a(t0_0101010101100), .b(t0_0101010101101), .y(t0_010101010110));
wire t0_0101010101100, t0_0101010101101;
mixer mix_t0_010101010111 (.a(t0_0101010101110), .b(t0_0101010101111), .y(t0_010101010111));
wire t0_0101010101110, t0_0101010101111;
mixer mix_t0_010101011 (.a(t0_0101010110), .b(t0_0101010111), .y(t0_010101011));
wire t0_0101010110, t0_0101010111;
mixer mix_t0_0101010110 (.a(t0_01010101100), .b(t0_01010101101), .y(t0_0101010110));
wire t0_01010101100, t0_01010101101;
mixer mix_t0_01010101100 (.a(t0_010101011000), .b(t0_010101011001), .y(t0_01010101100));
wire t0_010101011000, t0_010101011001;
mixer mix_t0_010101011000 (.a(t0_0101010110000), .b(t0_0101010110001), .y(t0_010101011000));
wire t0_0101010110000, t0_0101010110001;
mixer mix_t0_010101011001 (.a(t0_0101010110010), .b(t0_0101010110011), .y(t0_010101011001));
wire t0_0101010110010, t0_0101010110011;
mixer mix_t0_01010101101 (.a(t0_010101011010), .b(t0_010101011011), .y(t0_01010101101));
wire t0_010101011010, t0_010101011011;
mixer mix_t0_010101011010 (.a(t0_0101010110100), .b(t0_0101010110101), .y(t0_010101011010));
wire t0_0101010110100, t0_0101010110101;
mixer mix_t0_010101011011 (.a(t0_0101010110110), .b(t0_0101010110111), .y(t0_010101011011));
wire t0_0101010110110, t0_0101010110111;
mixer mix_t0_0101010111 (.a(t0_01010101110), .b(t0_01010101111), .y(t0_0101010111));
wire t0_01010101110, t0_01010101111;
mixer mix_t0_01010101110 (.a(t0_010101011100), .b(t0_010101011101), .y(t0_01010101110));
wire t0_010101011100, t0_010101011101;
mixer mix_t0_010101011100 (.a(t0_0101010111000), .b(t0_0101010111001), .y(t0_010101011100));
wire t0_0101010111000, t0_0101010111001;
mixer mix_t0_010101011101 (.a(t0_0101010111010), .b(t0_0101010111011), .y(t0_010101011101));
wire t0_0101010111010, t0_0101010111011;
mixer mix_t0_01010101111 (.a(t0_010101011110), .b(t0_010101011111), .y(t0_01010101111));
wire t0_010101011110, t0_010101011111;
mixer mix_t0_010101011110 (.a(t0_0101010111100), .b(t0_0101010111101), .y(t0_010101011110));
wire t0_0101010111100, t0_0101010111101;
mixer mix_t0_010101011111 (.a(t0_0101010111110), .b(t0_0101010111111), .y(t0_010101011111));
wire t0_0101010111110, t0_0101010111111;
mixer mix_t0_0101011 (.a(t0_01010110), .b(t0_01010111), .y(t0_0101011));
wire t0_01010110, t0_01010111;
mixer mix_t0_01010110 (.a(t0_010101100), .b(t0_010101101), .y(t0_01010110));
wire t0_010101100, t0_010101101;
mixer mix_t0_010101100 (.a(t0_0101011000), .b(t0_0101011001), .y(t0_010101100));
wire t0_0101011000, t0_0101011001;
mixer mix_t0_0101011000 (.a(t0_01010110000), .b(t0_01010110001), .y(t0_0101011000));
wire t0_01010110000, t0_01010110001;
mixer mix_t0_01010110000 (.a(t0_010101100000), .b(t0_010101100001), .y(t0_01010110000));
wire t0_010101100000, t0_010101100001;
mixer mix_t0_010101100000 (.a(t0_0101011000000), .b(t0_0101011000001), .y(t0_010101100000));
wire t0_0101011000000, t0_0101011000001;
mixer mix_t0_010101100001 (.a(t0_0101011000010), .b(t0_0101011000011), .y(t0_010101100001));
wire t0_0101011000010, t0_0101011000011;
mixer mix_t0_01010110001 (.a(t0_010101100010), .b(t0_010101100011), .y(t0_01010110001));
wire t0_010101100010, t0_010101100011;
mixer mix_t0_010101100010 (.a(t0_0101011000100), .b(t0_0101011000101), .y(t0_010101100010));
wire t0_0101011000100, t0_0101011000101;
mixer mix_t0_010101100011 (.a(t0_0101011000110), .b(t0_0101011000111), .y(t0_010101100011));
wire t0_0101011000110, t0_0101011000111;
mixer mix_t0_0101011001 (.a(t0_01010110010), .b(t0_01010110011), .y(t0_0101011001));
wire t0_01010110010, t0_01010110011;
mixer mix_t0_01010110010 (.a(t0_010101100100), .b(t0_010101100101), .y(t0_01010110010));
wire t0_010101100100, t0_010101100101;
mixer mix_t0_010101100100 (.a(t0_0101011001000), .b(t0_0101011001001), .y(t0_010101100100));
wire t0_0101011001000, t0_0101011001001;
mixer mix_t0_010101100101 (.a(t0_0101011001010), .b(t0_0101011001011), .y(t0_010101100101));
wire t0_0101011001010, t0_0101011001011;
mixer mix_t0_01010110011 (.a(t0_010101100110), .b(t0_010101100111), .y(t0_01010110011));
wire t0_010101100110, t0_010101100111;
mixer mix_t0_010101100110 (.a(t0_0101011001100), .b(t0_0101011001101), .y(t0_010101100110));
wire t0_0101011001100, t0_0101011001101;
mixer mix_t0_010101100111 (.a(t0_0101011001110), .b(t0_0101011001111), .y(t0_010101100111));
wire t0_0101011001110, t0_0101011001111;
mixer mix_t0_010101101 (.a(t0_0101011010), .b(t0_0101011011), .y(t0_010101101));
wire t0_0101011010, t0_0101011011;
mixer mix_t0_0101011010 (.a(t0_01010110100), .b(t0_01010110101), .y(t0_0101011010));
wire t0_01010110100, t0_01010110101;
mixer mix_t0_01010110100 (.a(t0_010101101000), .b(t0_010101101001), .y(t0_01010110100));
wire t0_010101101000, t0_010101101001;
mixer mix_t0_010101101000 (.a(t0_0101011010000), .b(t0_0101011010001), .y(t0_010101101000));
wire t0_0101011010000, t0_0101011010001;
mixer mix_t0_010101101001 (.a(t0_0101011010010), .b(t0_0101011010011), .y(t0_010101101001));
wire t0_0101011010010, t0_0101011010011;
mixer mix_t0_01010110101 (.a(t0_010101101010), .b(t0_010101101011), .y(t0_01010110101));
wire t0_010101101010, t0_010101101011;
mixer mix_t0_010101101010 (.a(t0_0101011010100), .b(t0_0101011010101), .y(t0_010101101010));
wire t0_0101011010100, t0_0101011010101;
mixer mix_t0_010101101011 (.a(t0_0101011010110), .b(t0_0101011010111), .y(t0_010101101011));
wire t0_0101011010110, t0_0101011010111;
mixer mix_t0_0101011011 (.a(t0_01010110110), .b(t0_01010110111), .y(t0_0101011011));
wire t0_01010110110, t0_01010110111;
mixer mix_t0_01010110110 (.a(t0_010101101100), .b(t0_010101101101), .y(t0_01010110110));
wire t0_010101101100, t0_010101101101;
mixer mix_t0_010101101100 (.a(t0_0101011011000), .b(t0_0101011011001), .y(t0_010101101100));
wire t0_0101011011000, t0_0101011011001;
mixer mix_t0_010101101101 (.a(t0_0101011011010), .b(t0_0101011011011), .y(t0_010101101101));
wire t0_0101011011010, t0_0101011011011;
mixer mix_t0_01010110111 (.a(t0_010101101110), .b(t0_010101101111), .y(t0_01010110111));
wire t0_010101101110, t0_010101101111;
mixer mix_t0_010101101110 (.a(t0_0101011011100), .b(t0_0101011011101), .y(t0_010101101110));
wire t0_0101011011100, t0_0101011011101;
mixer mix_t0_010101101111 (.a(t0_0101011011110), .b(t0_0101011011111), .y(t0_010101101111));
wire t0_0101011011110, t0_0101011011111;
mixer mix_t0_01010111 (.a(t0_010101110), .b(t0_010101111), .y(t0_01010111));
wire t0_010101110, t0_010101111;
mixer mix_t0_010101110 (.a(t0_0101011100), .b(t0_0101011101), .y(t0_010101110));
wire t0_0101011100, t0_0101011101;
mixer mix_t0_0101011100 (.a(t0_01010111000), .b(t0_01010111001), .y(t0_0101011100));
wire t0_01010111000, t0_01010111001;
mixer mix_t0_01010111000 (.a(t0_010101110000), .b(t0_010101110001), .y(t0_01010111000));
wire t0_010101110000, t0_010101110001;
mixer mix_t0_010101110000 (.a(t0_0101011100000), .b(t0_0101011100001), .y(t0_010101110000));
wire t0_0101011100000, t0_0101011100001;
mixer mix_t0_010101110001 (.a(t0_0101011100010), .b(t0_0101011100011), .y(t0_010101110001));
wire t0_0101011100010, t0_0101011100011;
mixer mix_t0_01010111001 (.a(t0_010101110010), .b(t0_010101110011), .y(t0_01010111001));
wire t0_010101110010, t0_010101110011;
mixer mix_t0_010101110010 (.a(t0_0101011100100), .b(t0_0101011100101), .y(t0_010101110010));
wire t0_0101011100100, t0_0101011100101;
mixer mix_t0_010101110011 (.a(t0_0101011100110), .b(t0_0101011100111), .y(t0_010101110011));
wire t0_0101011100110, t0_0101011100111;
mixer mix_t0_0101011101 (.a(t0_01010111010), .b(t0_01010111011), .y(t0_0101011101));
wire t0_01010111010, t0_01010111011;
mixer mix_t0_01010111010 (.a(t0_010101110100), .b(t0_010101110101), .y(t0_01010111010));
wire t0_010101110100, t0_010101110101;
mixer mix_t0_010101110100 (.a(t0_0101011101000), .b(t0_0101011101001), .y(t0_010101110100));
wire t0_0101011101000, t0_0101011101001;
mixer mix_t0_010101110101 (.a(t0_0101011101010), .b(t0_0101011101011), .y(t0_010101110101));
wire t0_0101011101010, t0_0101011101011;
mixer mix_t0_01010111011 (.a(t0_010101110110), .b(t0_010101110111), .y(t0_01010111011));
wire t0_010101110110, t0_010101110111;
mixer mix_t0_010101110110 (.a(t0_0101011101100), .b(t0_0101011101101), .y(t0_010101110110));
wire t0_0101011101100, t0_0101011101101;
mixer mix_t0_010101110111 (.a(t0_0101011101110), .b(t0_0101011101111), .y(t0_010101110111));
wire t0_0101011101110, t0_0101011101111;
mixer mix_t0_010101111 (.a(t0_0101011110), .b(t0_0101011111), .y(t0_010101111));
wire t0_0101011110, t0_0101011111;
mixer mix_t0_0101011110 (.a(t0_01010111100), .b(t0_01010111101), .y(t0_0101011110));
wire t0_01010111100, t0_01010111101;
mixer mix_t0_01010111100 (.a(t0_010101111000), .b(t0_010101111001), .y(t0_01010111100));
wire t0_010101111000, t0_010101111001;
mixer mix_t0_010101111000 (.a(t0_0101011110000), .b(t0_0101011110001), .y(t0_010101111000));
wire t0_0101011110000, t0_0101011110001;
mixer mix_t0_010101111001 (.a(t0_0101011110010), .b(t0_0101011110011), .y(t0_010101111001));
wire t0_0101011110010, t0_0101011110011;
mixer mix_t0_01010111101 (.a(t0_010101111010), .b(t0_010101111011), .y(t0_01010111101));
wire t0_010101111010, t0_010101111011;
mixer mix_t0_010101111010 (.a(t0_0101011110100), .b(t0_0101011110101), .y(t0_010101111010));
wire t0_0101011110100, t0_0101011110101;
mixer mix_t0_010101111011 (.a(t0_0101011110110), .b(t0_0101011110111), .y(t0_010101111011));
wire t0_0101011110110, t0_0101011110111;
mixer mix_t0_0101011111 (.a(t0_01010111110), .b(t0_01010111111), .y(t0_0101011111));
wire t0_01010111110, t0_01010111111;
mixer mix_t0_01010111110 (.a(t0_010101111100), .b(t0_010101111101), .y(t0_01010111110));
wire t0_010101111100, t0_010101111101;
mixer mix_t0_010101111100 (.a(t0_0101011111000), .b(t0_0101011111001), .y(t0_010101111100));
wire t0_0101011111000, t0_0101011111001;
mixer mix_t0_010101111101 (.a(t0_0101011111010), .b(t0_0101011111011), .y(t0_010101111101));
wire t0_0101011111010, t0_0101011111011;
mixer mix_t0_01010111111 (.a(t0_010101111110), .b(t0_010101111111), .y(t0_01010111111));
wire t0_010101111110, t0_010101111111;
mixer mix_t0_010101111110 (.a(t0_0101011111100), .b(t0_0101011111101), .y(t0_010101111110));
wire t0_0101011111100, t0_0101011111101;
mixer mix_t0_010101111111 (.a(t0_0101011111110), .b(t0_0101011111111), .y(t0_010101111111));
wire t0_0101011111110, t0_0101011111111;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_010110 (.a(t0_0101100), .b(t0_0101101), .y(t0_010110));
wire t0_0101100, t0_0101101;
mixer mix_t0_0101100 (.a(t0_01011000), .b(t0_01011001), .y(t0_0101100));
wire t0_01011000, t0_01011001;
mixer mix_t0_01011000 (.a(t0_010110000), .b(t0_010110001), .y(t0_01011000));
wire t0_010110000, t0_010110001;
mixer mix_t0_010110000 (.a(t0_0101100000), .b(t0_0101100001), .y(t0_010110000));
wire t0_0101100000, t0_0101100001;
mixer mix_t0_0101100000 (.a(t0_01011000000), .b(t0_01011000001), .y(t0_0101100000));
wire t0_01011000000, t0_01011000001;
mixer mix_t0_01011000000 (.a(t0_010110000000), .b(t0_010110000001), .y(t0_01011000000));
wire t0_010110000000, t0_010110000001;
mixer mix_t0_010110000000 (.a(t0_0101100000000), .b(t0_0101100000001), .y(t0_010110000000));
wire t0_0101100000000, t0_0101100000001;
mixer mix_t0_010110000001 (.a(t0_0101100000010), .b(t0_0101100000011), .y(t0_010110000001));
wire t0_0101100000010, t0_0101100000011;
mixer mix_t0_01011000001 (.a(t0_010110000010), .b(t0_010110000011), .y(t0_01011000001));
wire t0_010110000010, t0_010110000011;
mixer mix_t0_010110000010 (.a(t0_0101100000100), .b(t0_0101100000101), .y(t0_010110000010));
wire t0_0101100000100, t0_0101100000101;
mixer mix_t0_010110000011 (.a(t0_0101100000110), .b(t0_0101100000111), .y(t0_010110000011));
wire t0_0101100000110, t0_0101100000111;
mixer mix_t0_0101100001 (.a(t0_01011000010), .b(t0_01011000011), .y(t0_0101100001));
wire t0_01011000010, t0_01011000011;
mixer mix_t0_01011000010 (.a(t0_010110000100), .b(t0_010110000101), .y(t0_01011000010));
wire t0_010110000100, t0_010110000101;
mixer mix_t0_010110000100 (.a(t0_0101100001000), .b(t0_0101100001001), .y(t0_010110000100));
wire t0_0101100001000, t0_0101100001001;
mixer mix_t0_010110000101 (.a(t0_0101100001010), .b(t0_0101100001011), .y(t0_010110000101));
wire t0_0101100001010, t0_0101100001011;
mixer mix_t0_01011000011 (.a(t0_010110000110), .b(t0_010110000111), .y(t0_01011000011));
wire t0_010110000110, t0_010110000111;
mixer mix_t0_010110000110 (.a(t0_0101100001100), .b(t0_0101100001101), .y(t0_010110000110));
wire t0_0101100001100, t0_0101100001101;
mixer mix_t0_010110000111 (.a(t0_0101100001110), .b(t0_0101100001111), .y(t0_010110000111));
wire t0_0101100001110, t0_0101100001111;
mixer mix_t0_010110001 (.a(t0_0101100010), .b(t0_0101100011), .y(t0_010110001));
wire t0_0101100010, t0_0101100011;
mixer mix_t0_0101100010 (.a(t0_01011000100), .b(t0_01011000101), .y(t0_0101100010));
wire t0_01011000100, t0_01011000101;
mixer mix_t0_01011000100 (.a(t0_010110001000), .b(t0_010110001001), .y(t0_01011000100));
wire t0_010110001000, t0_010110001001;
mixer mix_t0_010110001000 (.a(t0_0101100010000), .b(t0_0101100010001), .y(t0_010110001000));
wire t0_0101100010000, t0_0101100010001;
mixer mix_t0_010110001001 (.a(t0_0101100010010), .b(t0_0101100010011), .y(t0_010110001001));
wire t0_0101100010010, t0_0101100010011;
mixer mix_t0_01011000101 (.a(t0_010110001010), .b(t0_010110001011), .y(t0_01011000101));
wire t0_010110001010, t0_010110001011;
mixer mix_t0_010110001010 (.a(t0_0101100010100), .b(t0_0101100010101), .y(t0_010110001010));
wire t0_0101100010100, t0_0101100010101;
mixer mix_t0_010110001011 (.a(t0_0101100010110), .b(t0_0101100010111), .y(t0_010110001011));
wire t0_0101100010110, t0_0101100010111;
mixer mix_t0_0101100011 (.a(t0_01011000110), .b(t0_01011000111), .y(t0_0101100011));
wire t0_01011000110, t0_01011000111;
mixer mix_t0_01011000110 (.a(t0_010110001100), .b(t0_010110001101), .y(t0_01011000110));
wire t0_010110001100, t0_010110001101;
mixer mix_t0_010110001100 (.a(t0_0101100011000), .b(t0_0101100011001), .y(t0_010110001100));
wire t0_0101100011000, t0_0101100011001;
mixer mix_t0_010110001101 (.a(t0_0101100011010), .b(t0_0101100011011), .y(t0_010110001101));
wire t0_0101100011010, t0_0101100011011;
mixer mix_t0_01011000111 (.a(t0_010110001110), .b(t0_010110001111), .y(t0_01011000111));
wire t0_010110001110, t0_010110001111;
mixer mix_t0_010110001110 (.a(t0_0101100011100), .b(t0_0101100011101), .y(t0_010110001110));
wire t0_0101100011100, t0_0101100011101;
mixer mix_t0_010110001111 (.a(t0_0101100011110), .b(t0_0101100011111), .y(t0_010110001111));
wire t0_0101100011110, t0_0101100011111;
mixer mix_t0_01011001 (.a(t0_010110010), .b(t0_010110011), .y(t0_01011001));
wire t0_010110010, t0_010110011;
mixer mix_t0_010110010 (.a(t0_0101100100), .b(t0_0101100101), .y(t0_010110010));
wire t0_0101100100, t0_0101100101;
mixer mix_t0_0101100100 (.a(t0_01011001000), .b(t0_01011001001), .y(t0_0101100100));
wire t0_01011001000, t0_01011001001;
mixer mix_t0_01011001000 (.a(t0_010110010000), .b(t0_010110010001), .y(t0_01011001000));
wire t0_010110010000, t0_010110010001;
mixer mix_t0_010110010000 (.a(t0_0101100100000), .b(t0_0101100100001), .y(t0_010110010000));
wire t0_0101100100000, t0_0101100100001;
mixer mix_t0_010110010001 (.a(t0_0101100100010), .b(t0_0101100100011), .y(t0_010110010001));
wire t0_0101100100010, t0_0101100100011;
mixer mix_t0_01011001001 (.a(t0_010110010010), .b(t0_010110010011), .y(t0_01011001001));
wire t0_010110010010, t0_010110010011;
mixer mix_t0_010110010010 (.a(t0_0101100100100), .b(t0_0101100100101), .y(t0_010110010010));
wire t0_0101100100100, t0_0101100100101;
mixer mix_t0_010110010011 (.a(t0_0101100100110), .b(t0_0101100100111), .y(t0_010110010011));
wire t0_0101100100110, t0_0101100100111;
mixer mix_t0_0101100101 (.a(t0_01011001010), .b(t0_01011001011), .y(t0_0101100101));
wire t0_01011001010, t0_01011001011;
mixer mix_t0_01011001010 (.a(t0_010110010100), .b(t0_010110010101), .y(t0_01011001010));
wire t0_010110010100, t0_010110010101;
mixer mix_t0_010110010100 (.a(t0_0101100101000), .b(t0_0101100101001), .y(t0_010110010100));
wire t0_0101100101000, t0_0101100101001;
mixer mix_t0_010110010101 (.a(t0_0101100101010), .b(t0_0101100101011), .y(t0_010110010101));
wire t0_0101100101010, t0_0101100101011;
mixer mix_t0_01011001011 (.a(t0_010110010110), .b(t0_010110010111), .y(t0_01011001011));
wire t0_010110010110, t0_010110010111;
mixer mix_t0_010110010110 (.a(t0_0101100101100), .b(t0_0101100101101), .y(t0_010110010110));
wire t0_0101100101100, t0_0101100101101;
mixer mix_t0_010110010111 (.a(t0_0101100101110), .b(t0_0101100101111), .y(t0_010110010111));
wire t0_0101100101110, t0_0101100101111;
mixer mix_t0_010110011 (.a(t0_0101100110), .b(t0_0101100111), .y(t0_010110011));
wire t0_0101100110, t0_0101100111;
mixer mix_t0_0101100110 (.a(t0_01011001100), .b(t0_01011001101), .y(t0_0101100110));
wire t0_01011001100, t0_01011001101;
mixer mix_t0_01011001100 (.a(t0_010110011000), .b(t0_010110011001), .y(t0_01011001100));
wire t0_010110011000, t0_010110011001;
mixer mix_t0_010110011000 (.a(t0_0101100110000), .b(t0_0101100110001), .y(t0_010110011000));
wire t0_0101100110000, t0_0101100110001;
mixer mix_t0_010110011001 (.a(t0_0101100110010), .b(t0_0101100110011), .y(t0_010110011001));
wire t0_0101100110010, t0_0101100110011;
mixer mix_t0_01011001101 (.a(t0_010110011010), .b(t0_010110011011), .y(t0_01011001101));
wire t0_010110011010, t0_010110011011;
mixer mix_t0_010110011010 (.a(t0_0101100110100), .b(t0_0101100110101), .y(t0_010110011010));
wire t0_0101100110100, t0_0101100110101;
mixer mix_t0_010110011011 (.a(t0_0101100110110), .b(t0_0101100110111), .y(t0_010110011011));
wire t0_0101100110110, t0_0101100110111;
mixer mix_t0_0101100111 (.a(t0_01011001110), .b(t0_01011001111), .y(t0_0101100111));
wire t0_01011001110, t0_01011001111;
mixer mix_t0_01011001110 (.a(t0_010110011100), .b(t0_010110011101), .y(t0_01011001110));
wire t0_010110011100, t0_010110011101;
mixer mix_t0_010110011100 (.a(t0_0101100111000), .b(t0_0101100111001), .y(t0_010110011100));
wire t0_0101100111000, t0_0101100111001;
mixer mix_t0_010110011101 (.a(t0_0101100111010), .b(t0_0101100111011), .y(t0_010110011101));
wire t0_0101100111010, t0_0101100111011;
mixer mix_t0_01011001111 (.a(t0_010110011110), .b(t0_010110011111), .y(t0_01011001111));
wire t0_010110011110, t0_010110011111;
mixer mix_t0_010110011110 (.a(t0_0101100111100), .b(t0_0101100111101), .y(t0_010110011110));
wire t0_0101100111100, t0_0101100111101;
mixer mix_t0_010110011111 (.a(t0_0101100111110), .b(t0_0101100111111), .y(t0_010110011111));
wire t0_0101100111110, t0_0101100111111;
mixer mix_t0_0101101 (.a(t0_01011010), .b(t0_01011011), .y(t0_0101101));
wire t0_01011010, t0_01011011;
mixer mix_t0_01011010 (.a(t0_010110100), .b(t0_010110101), .y(t0_01011010));
wire t0_010110100, t0_010110101;
mixer mix_t0_010110100 (.a(t0_0101101000), .b(t0_0101101001), .y(t0_010110100));
wire t0_0101101000, t0_0101101001;
mixer mix_t0_0101101000 (.a(t0_01011010000), .b(t0_01011010001), .y(t0_0101101000));
wire t0_01011010000, t0_01011010001;
mixer mix_t0_01011010000 (.a(t0_010110100000), .b(t0_010110100001), .y(t0_01011010000));
wire t0_010110100000, t0_010110100001;
mixer mix_t0_010110100000 (.a(t0_0101101000000), .b(t0_0101101000001), .y(t0_010110100000));
wire t0_0101101000000, t0_0101101000001;
mixer mix_t0_010110100001 (.a(t0_0101101000010), .b(t0_0101101000011), .y(t0_010110100001));
wire t0_0101101000010, t0_0101101000011;
mixer mix_t0_01011010001 (.a(t0_010110100010), .b(t0_010110100011), .y(t0_01011010001));
wire t0_010110100010, t0_010110100011;
mixer mix_t0_010110100010 (.a(t0_0101101000100), .b(t0_0101101000101), .y(t0_010110100010));
wire t0_0101101000100, t0_0101101000101;
mixer mix_t0_010110100011 (.a(t0_0101101000110), .b(t0_0101101000111), .y(t0_010110100011));
wire t0_0101101000110, t0_0101101000111;
mixer mix_t0_0101101001 (.a(t0_01011010010), .b(t0_01011010011), .y(t0_0101101001));
wire t0_01011010010, t0_01011010011;
mixer mix_t0_01011010010 (.a(t0_010110100100), .b(t0_010110100101), .y(t0_01011010010));
wire t0_010110100100, t0_010110100101;
mixer mix_t0_010110100100 (.a(t0_0101101001000), .b(t0_0101101001001), .y(t0_010110100100));
wire t0_0101101001000, t0_0101101001001;
mixer mix_t0_010110100101 (.a(t0_0101101001010), .b(t0_0101101001011), .y(t0_010110100101));
wire t0_0101101001010, t0_0101101001011;
mixer mix_t0_01011010011 (.a(t0_010110100110), .b(t0_010110100111), .y(t0_01011010011));
wire t0_010110100110, t0_010110100111;
mixer mix_t0_010110100110 (.a(t0_0101101001100), .b(t0_0101101001101), .y(t0_010110100110));
wire t0_0101101001100, t0_0101101001101;
mixer mix_t0_010110100111 (.a(t0_0101101001110), .b(t0_0101101001111), .y(t0_010110100111));
wire t0_0101101001110, t0_0101101001111;
mixer mix_t0_010110101 (.a(t0_0101101010), .b(t0_0101101011), .y(t0_010110101));
wire t0_0101101010, t0_0101101011;
mixer mix_t0_0101101010 (.a(t0_01011010100), .b(t0_01011010101), .y(t0_0101101010));
wire t0_01011010100, t0_01011010101;
mixer mix_t0_01011010100 (.a(t0_010110101000), .b(t0_010110101001), .y(t0_01011010100));
wire t0_010110101000, t0_010110101001;
mixer mix_t0_010110101000 (.a(t0_0101101010000), .b(t0_0101101010001), .y(t0_010110101000));
wire t0_0101101010000, t0_0101101010001;
mixer mix_t0_010110101001 (.a(t0_0101101010010), .b(t0_0101101010011), .y(t0_010110101001));
wire t0_0101101010010, t0_0101101010011;
mixer mix_t0_01011010101 (.a(t0_010110101010), .b(t0_010110101011), .y(t0_01011010101));
wire t0_010110101010, t0_010110101011;
mixer mix_t0_010110101010 (.a(t0_0101101010100), .b(t0_0101101010101), .y(t0_010110101010));
wire t0_0101101010100, t0_0101101010101;
mixer mix_t0_010110101011 (.a(t0_0101101010110), .b(t0_0101101010111), .y(t0_010110101011));
wire t0_0101101010110, t0_0101101010111;
mixer mix_t0_0101101011 (.a(t0_01011010110), .b(t0_01011010111), .y(t0_0101101011));
wire t0_01011010110, t0_01011010111;
mixer mix_t0_01011010110 (.a(t0_010110101100), .b(t0_010110101101), .y(t0_01011010110));
wire t0_010110101100, t0_010110101101;
mixer mix_t0_010110101100 (.a(t0_0101101011000), .b(t0_0101101011001), .y(t0_010110101100));
wire t0_0101101011000, t0_0101101011001;
mixer mix_t0_010110101101 (.a(t0_0101101011010), .b(t0_0101101011011), .y(t0_010110101101));
wire t0_0101101011010, t0_0101101011011;
mixer mix_t0_01011010111 (.a(t0_010110101110), .b(t0_010110101111), .y(t0_01011010111));
wire t0_010110101110, t0_010110101111;
mixer mix_t0_010110101110 (.a(t0_0101101011100), .b(t0_0101101011101), .y(t0_010110101110));
wire t0_0101101011100, t0_0101101011101;
mixer mix_t0_010110101111 (.a(t0_0101101011110), .b(t0_0101101011111), .y(t0_010110101111));
wire t0_0101101011110, t0_0101101011111;
mixer mix_t0_01011011 (.a(t0_010110110), .b(t0_010110111), .y(t0_01011011));
wire t0_010110110, t0_010110111;
mixer mix_t0_010110110 (.a(t0_0101101100), .b(t0_0101101101), .y(t0_010110110));
wire t0_0101101100, t0_0101101101;
mixer mix_t0_0101101100 (.a(t0_01011011000), .b(t0_01011011001), .y(t0_0101101100));
wire t0_01011011000, t0_01011011001;
mixer mix_t0_01011011000 (.a(t0_010110110000), .b(t0_010110110001), .y(t0_01011011000));
wire t0_010110110000, t0_010110110001;
mixer mix_t0_010110110000 (.a(t0_0101101100000), .b(t0_0101101100001), .y(t0_010110110000));
wire t0_0101101100000, t0_0101101100001;
mixer mix_t0_010110110001 (.a(t0_0101101100010), .b(t0_0101101100011), .y(t0_010110110001));
wire t0_0101101100010, t0_0101101100011;
mixer mix_t0_01011011001 (.a(t0_010110110010), .b(t0_010110110011), .y(t0_01011011001));
wire t0_010110110010, t0_010110110011;
mixer mix_t0_010110110010 (.a(t0_0101101100100), .b(t0_0101101100101), .y(t0_010110110010));
wire t0_0101101100100, t0_0101101100101;
mixer mix_t0_010110110011 (.a(t0_0101101100110), .b(t0_0101101100111), .y(t0_010110110011));
wire t0_0101101100110, t0_0101101100111;
mixer mix_t0_0101101101 (.a(t0_01011011010), .b(t0_01011011011), .y(t0_0101101101));
wire t0_01011011010, t0_01011011011;
mixer mix_t0_01011011010 (.a(t0_010110110100), .b(t0_010110110101), .y(t0_01011011010));
wire t0_010110110100, t0_010110110101;
mixer mix_t0_010110110100 (.a(t0_0101101101000), .b(t0_0101101101001), .y(t0_010110110100));
wire t0_0101101101000, t0_0101101101001;
mixer mix_t0_010110110101 (.a(t0_0101101101010), .b(t0_0101101101011), .y(t0_010110110101));
wire t0_0101101101010, t0_0101101101011;
mixer mix_t0_01011011011 (.a(t0_010110110110), .b(t0_010110110111), .y(t0_01011011011));
wire t0_010110110110, t0_010110110111;
mixer mix_t0_010110110110 (.a(t0_0101101101100), .b(t0_0101101101101), .y(t0_010110110110));
wire t0_0101101101100, t0_0101101101101;
mixer mix_t0_010110110111 (.a(t0_0101101101110), .b(t0_0101101101111), .y(t0_010110110111));
wire t0_0101101101110, t0_0101101101111;
mixer mix_t0_010110111 (.a(t0_0101101110), .b(t0_0101101111), .y(t0_010110111));
wire t0_0101101110, t0_0101101111;
mixer mix_t0_0101101110 (.a(t0_01011011100), .b(t0_01011011101), .y(t0_0101101110));
wire t0_01011011100, t0_01011011101;
mixer mix_t0_01011011100 (.a(t0_010110111000), .b(t0_010110111001), .y(t0_01011011100));
wire t0_010110111000, t0_010110111001;
mixer mix_t0_010110111000 (.a(t0_0101101110000), .b(t0_0101101110001), .y(t0_010110111000));
wire t0_0101101110000, t0_0101101110001;
mixer mix_t0_010110111001 (.a(t0_0101101110010), .b(t0_0101101110011), .y(t0_010110111001));
wire t0_0101101110010, t0_0101101110011;
mixer mix_t0_01011011101 (.a(t0_010110111010), .b(t0_010110111011), .y(t0_01011011101));
wire t0_010110111010, t0_010110111011;
mixer mix_t0_010110111010 (.a(t0_0101101110100), .b(t0_0101101110101), .y(t0_010110111010));
wire t0_0101101110100, t0_0101101110101;
mixer mix_t0_010110111011 (.a(t0_0101101110110), .b(t0_0101101110111), .y(t0_010110111011));
wire t0_0101101110110, t0_0101101110111;
mixer mix_t0_0101101111 (.a(t0_01011011110), .b(t0_01011011111), .y(t0_0101101111));
wire t0_01011011110, t0_01011011111;
mixer mix_t0_01011011110 (.a(t0_010110111100), .b(t0_010110111101), .y(t0_01011011110));
wire t0_010110111100, t0_010110111101;
mixer mix_t0_010110111100 (.a(t0_0101101111000), .b(t0_0101101111001), .y(t0_010110111100));
wire t0_0101101111000, t0_0101101111001;
mixer mix_t0_010110111101 (.a(t0_0101101111010), .b(t0_0101101111011), .y(t0_010110111101));
wire t0_0101101111010, t0_0101101111011;
mixer mix_t0_01011011111 (.a(t0_010110111110), .b(t0_010110111111), .y(t0_01011011111));
wire t0_010110111110, t0_010110111111;
mixer mix_t0_010110111110 (.a(t0_0101101111100), .b(t0_0101101111101), .y(t0_010110111110));
wire t0_0101101111100, t0_0101101111101;
mixer mix_t0_010110111111 (.a(t0_0101101111110), .b(t0_0101101111111), .y(t0_010110111111));
wire t0_0101101111110, t0_0101101111111;
mixer mix_t0_010111 (.a(t0_0101110), .b(t0_0101111), .y(t0_010111));
wire t0_0101110, t0_0101111;
mixer mix_t0_0101110 (.a(t0_01011100), .b(t0_01011101), .y(t0_0101110));
wire t0_01011100, t0_01011101;
mixer mix_t0_01011100 (.a(t0_010111000), .b(t0_010111001), .y(t0_01011100));
wire t0_010111000, t0_010111001;
mixer mix_t0_010111000 (.a(t0_0101110000), .b(t0_0101110001), .y(t0_010111000));
wire t0_0101110000, t0_0101110001;
mixer mix_t0_0101110000 (.a(t0_01011100000), .b(t0_01011100001), .y(t0_0101110000));
wire t0_01011100000, t0_01011100001;
mixer mix_t0_01011100000 (.a(t0_010111000000), .b(t0_010111000001), .y(t0_01011100000));
wire t0_010111000000, t0_010111000001;
mixer mix_t0_010111000000 (.a(t0_0101110000000), .b(t0_0101110000001), .y(t0_010111000000));
wire t0_0101110000000, t0_0101110000001;
mixer mix_t0_010111000001 (.a(t0_0101110000010), .b(t0_0101110000011), .y(t0_010111000001));
wire t0_0101110000010, t0_0101110000011;
mixer mix_t0_01011100001 (.a(t0_010111000010), .b(t0_010111000011), .y(t0_01011100001));
wire t0_010111000010, t0_010111000011;
mixer mix_t0_010111000010 (.a(t0_0101110000100), .b(t0_0101110000101), .y(t0_010111000010));
wire t0_0101110000100, t0_0101110000101;
mixer mix_t0_010111000011 (.a(t0_0101110000110), .b(t0_0101110000111), .y(t0_010111000011));
wire t0_0101110000110, t0_0101110000111;
mixer mix_t0_0101110001 (.a(t0_01011100010), .b(t0_01011100011), .y(t0_0101110001));
wire t0_01011100010, t0_01011100011;
mixer mix_t0_01011100010 (.a(t0_010111000100), .b(t0_010111000101), .y(t0_01011100010));
wire t0_010111000100, t0_010111000101;
mixer mix_t0_010111000100 (.a(t0_0101110001000), .b(t0_0101110001001), .y(t0_010111000100));
wire t0_0101110001000, t0_0101110001001;
mixer mix_t0_010111000101 (.a(t0_0101110001010), .b(t0_0101110001011), .y(t0_010111000101));
wire t0_0101110001010, t0_0101110001011;
mixer mix_t0_01011100011 (.a(t0_010111000110), .b(t0_010111000111), .y(t0_01011100011));
wire t0_010111000110, t0_010111000111;
mixer mix_t0_010111000110 (.a(t0_0101110001100), .b(t0_0101110001101), .y(t0_010111000110));
wire t0_0101110001100, t0_0101110001101;
mixer mix_t0_010111000111 (.a(t0_0101110001110), .b(t0_0101110001111), .y(t0_010111000111));
wire t0_0101110001110, t0_0101110001111;
mixer mix_t0_010111001 (.a(t0_0101110010), .b(t0_0101110011), .y(t0_010111001));
wire t0_0101110010, t0_0101110011;
mixer mix_t0_0101110010 (.a(t0_01011100100), .b(t0_01011100101), .y(t0_0101110010));
wire t0_01011100100, t0_01011100101;
mixer mix_t0_01011100100 (.a(t0_010111001000), .b(t0_010111001001), .y(t0_01011100100));
wire t0_010111001000, t0_010111001001;
mixer mix_t0_010111001000 (.a(t0_0101110010000), .b(t0_0101110010001), .y(t0_010111001000));
wire t0_0101110010000, t0_0101110010001;
mixer mix_t0_010111001001 (.a(t0_0101110010010), .b(t0_0101110010011), .y(t0_010111001001));
wire t0_0101110010010, t0_0101110010011;
mixer mix_t0_01011100101 (.a(t0_010111001010), .b(t0_010111001011), .y(t0_01011100101));
wire t0_010111001010, t0_010111001011;
mixer mix_t0_010111001010 (.a(t0_0101110010100), .b(t0_0101110010101), .y(t0_010111001010));
wire t0_0101110010100, t0_0101110010101;
mixer mix_t0_010111001011 (.a(t0_0101110010110), .b(t0_0101110010111), .y(t0_010111001011));
wire t0_0101110010110, t0_0101110010111;
mixer mix_t0_0101110011 (.a(t0_01011100110), .b(t0_01011100111), .y(t0_0101110011));
wire t0_01011100110, t0_01011100111;
mixer mix_t0_01011100110 (.a(t0_010111001100), .b(t0_010111001101), .y(t0_01011100110));
wire t0_010111001100, t0_010111001101;
mixer mix_t0_010111001100 (.a(t0_0101110011000), .b(t0_0101110011001), .y(t0_010111001100));
wire t0_0101110011000, t0_0101110011001;
mixer mix_t0_010111001101 (.a(t0_0101110011010), .b(t0_0101110011011), .y(t0_010111001101));
wire t0_0101110011010, t0_0101110011011;
mixer mix_t0_01011100111 (.a(t0_010111001110), .b(t0_010111001111), .y(t0_01011100111));
wire t0_010111001110, t0_010111001111;
mixer mix_t0_010111001110 (.a(t0_0101110011100), .b(t0_0101110011101), .y(t0_010111001110));
wire t0_0101110011100, t0_0101110011101;
mixer mix_t0_010111001111 (.a(t0_0101110011110), .b(t0_0101110011111), .y(t0_010111001111));
wire t0_0101110011110, t0_0101110011111;
mixer mix_t0_01011101 (.a(t0_010111010), .b(t0_010111011), .y(t0_01011101));
wire t0_010111010, t0_010111011;
mixer mix_t0_010111010 (.a(t0_0101110100), .b(t0_0101110101), .y(t0_010111010));
wire t0_0101110100, t0_0101110101;
mixer mix_t0_0101110100 (.a(t0_01011101000), .b(t0_01011101001), .y(t0_0101110100));
wire t0_01011101000, t0_01011101001;
mixer mix_t0_01011101000 (.a(t0_010111010000), .b(t0_010111010001), .y(t0_01011101000));
wire t0_010111010000, t0_010111010001;
mixer mix_t0_010111010000 (.a(t0_0101110100000), .b(t0_0101110100001), .y(t0_010111010000));
wire t0_0101110100000, t0_0101110100001;
mixer mix_t0_010111010001 (.a(t0_0101110100010), .b(t0_0101110100011), .y(t0_010111010001));
wire t0_0101110100010, t0_0101110100011;
mixer mix_t0_01011101001 (.a(t0_010111010010), .b(t0_010111010011), .y(t0_01011101001));
wire t0_010111010010, t0_010111010011;
mixer mix_t0_010111010010 (.a(t0_0101110100100), .b(t0_0101110100101), .y(t0_010111010010));
wire t0_0101110100100, t0_0101110100101;
mixer mix_t0_010111010011 (.a(t0_0101110100110), .b(t0_0101110100111), .y(t0_010111010011));
wire t0_0101110100110, t0_0101110100111;
mixer mix_t0_0101110101 (.a(t0_01011101010), .b(t0_01011101011), .y(t0_0101110101));
wire t0_01011101010, t0_01011101011;
mixer mix_t0_01011101010 (.a(t0_010111010100), .b(t0_010111010101), .y(t0_01011101010));
wire t0_010111010100, t0_010111010101;
mixer mix_t0_010111010100 (.a(t0_0101110101000), .b(t0_0101110101001), .y(t0_010111010100));
wire t0_0101110101000, t0_0101110101001;
mixer mix_t0_010111010101 (.a(t0_0101110101010), .b(t0_0101110101011), .y(t0_010111010101));
wire t0_0101110101010, t0_0101110101011;
mixer mix_t0_01011101011 (.a(t0_010111010110), .b(t0_010111010111), .y(t0_01011101011));
wire t0_010111010110, t0_010111010111;
mixer mix_t0_010111010110 (.a(t0_0101110101100), .b(t0_0101110101101), .y(t0_010111010110));
wire t0_0101110101100, t0_0101110101101;
mixer mix_t0_010111010111 (.a(t0_0101110101110), .b(t0_0101110101111), .y(t0_010111010111));
wire t0_0101110101110, t0_0101110101111;
mixer mix_t0_010111011 (.a(t0_0101110110), .b(t0_0101110111), .y(t0_010111011));
wire t0_0101110110, t0_0101110111;
mixer mix_t0_0101110110 (.a(t0_01011101100), .b(t0_01011101101), .y(t0_0101110110));
wire t0_01011101100, t0_01011101101;
mixer mix_t0_01011101100 (.a(t0_010111011000), .b(t0_010111011001), .y(t0_01011101100));
wire t0_010111011000, t0_010111011001;
mixer mix_t0_010111011000 (.a(t0_0101110110000), .b(t0_0101110110001), .y(t0_010111011000));
wire t0_0101110110000, t0_0101110110001;
mixer mix_t0_010111011001 (.a(t0_0101110110010), .b(t0_0101110110011), .y(t0_010111011001));
wire t0_0101110110010, t0_0101110110011;
mixer mix_t0_01011101101 (.a(t0_010111011010), .b(t0_010111011011), .y(t0_01011101101));
wire t0_010111011010, t0_010111011011;
mixer mix_t0_010111011010 (.a(t0_0101110110100), .b(t0_0101110110101), .y(t0_010111011010));
wire t0_0101110110100, t0_0101110110101;
mixer mix_t0_010111011011 (.a(t0_0101110110110), .b(t0_0101110110111), .y(t0_010111011011));
wire t0_0101110110110, t0_0101110110111;
mixer mix_t0_0101110111 (.a(t0_01011101110), .b(t0_01011101111), .y(t0_0101110111));
wire t0_01011101110, t0_01011101111;
mixer mix_t0_01011101110 (.a(t0_010111011100), .b(t0_010111011101), .y(t0_01011101110));
wire t0_010111011100, t0_010111011101;
mixer mix_t0_010111011100 (.a(t0_0101110111000), .b(t0_0101110111001), .y(t0_010111011100));
wire t0_0101110111000, t0_0101110111001;
mixer mix_t0_010111011101 (.a(t0_0101110111010), .b(t0_0101110111011), .y(t0_010111011101));
wire t0_0101110111010, t0_0101110111011;
mixer mix_t0_01011101111 (.a(t0_010111011110), .b(t0_010111011111), .y(t0_01011101111));
wire t0_010111011110, t0_010111011111;
mixer mix_t0_010111011110 (.a(t0_0101110111100), .b(t0_0101110111101), .y(t0_010111011110));
wire t0_0101110111100, t0_0101110111101;
mixer mix_t0_010111011111 (.a(t0_0101110111110), .b(t0_0101110111111), .y(t0_010111011111));
wire t0_0101110111110, t0_0101110111111;
mixer mix_t0_0101111 (.a(t0_01011110), .b(t0_01011111), .y(t0_0101111));
wire t0_01011110, t0_01011111;
mixer mix_t0_01011110 (.a(t0_010111100), .b(t0_010111101), .y(t0_01011110));
wire t0_010111100, t0_010111101;
mixer mix_t0_010111100 (.a(t0_0101111000), .b(t0_0101111001), .y(t0_010111100));
wire t0_0101111000, t0_0101111001;
mixer mix_t0_0101111000 (.a(t0_01011110000), .b(t0_01011110001), .y(t0_0101111000));
wire t0_01011110000, t0_01011110001;
mixer mix_t0_01011110000 (.a(t0_010111100000), .b(t0_010111100001), .y(t0_01011110000));
wire t0_010111100000, t0_010111100001;
mixer mix_t0_010111100000 (.a(t0_0101111000000), .b(t0_0101111000001), .y(t0_010111100000));
wire t0_0101111000000, t0_0101111000001;
mixer mix_t0_010111100001 (.a(t0_0101111000010), .b(t0_0101111000011), .y(t0_010111100001));
wire t0_0101111000010, t0_0101111000011;
mixer mix_t0_01011110001 (.a(t0_010111100010), .b(t0_010111100011), .y(t0_01011110001));
wire t0_010111100010, t0_010111100011;
mixer mix_t0_010111100010 (.a(t0_0101111000100), .b(t0_0101111000101), .y(t0_010111100010));
wire t0_0101111000100, t0_0101111000101;
mixer mix_t0_010111100011 (.a(t0_0101111000110), .b(t0_0101111000111), .y(t0_010111100011));
wire t0_0101111000110, t0_0101111000111;
mixer mix_t0_0101111001 (.a(t0_01011110010), .b(t0_01011110011), .y(t0_0101111001));
wire t0_01011110010, t0_01011110011;
mixer mix_t0_01011110010 (.a(t0_010111100100), .b(t0_010111100101), .y(t0_01011110010));
wire t0_010111100100, t0_010111100101;
mixer mix_t0_010111100100 (.a(t0_0101111001000), .b(t0_0101111001001), .y(t0_010111100100));
wire t0_0101111001000, t0_0101111001001;
mixer mix_t0_010111100101 (.a(t0_0101111001010), .b(t0_0101111001011), .y(t0_010111100101));
wire t0_0101111001010, t0_0101111001011;
mixer mix_t0_01011110011 (.a(t0_010111100110), .b(t0_010111100111), .y(t0_01011110011));
wire t0_010111100110, t0_010111100111;
mixer mix_t0_010111100110 (.a(t0_0101111001100), .b(t0_0101111001101), .y(t0_010111100110));
wire t0_0101111001100, t0_0101111001101;
mixer mix_t0_010111100111 (.a(t0_0101111001110), .b(t0_0101111001111), .y(t0_010111100111));
wire t0_0101111001110, t0_0101111001111;
mixer mix_t0_010111101 (.a(t0_0101111010), .b(t0_0101111011), .y(t0_010111101));
wire t0_0101111010, t0_0101111011;
mixer mix_t0_0101111010 (.a(t0_01011110100), .b(t0_01011110101), .y(t0_0101111010));
wire t0_01011110100, t0_01011110101;
mixer mix_t0_01011110100 (.a(t0_010111101000), .b(t0_010111101001), .y(t0_01011110100));
wire t0_010111101000, t0_010111101001;
mixer mix_t0_010111101000 (.a(t0_0101111010000), .b(t0_0101111010001), .y(t0_010111101000));
wire t0_0101111010000, t0_0101111010001;
mixer mix_t0_010111101001 (.a(t0_0101111010010), .b(t0_0101111010011), .y(t0_010111101001));
wire t0_0101111010010, t0_0101111010011;
mixer mix_t0_01011110101 (.a(t0_010111101010), .b(t0_010111101011), .y(t0_01011110101));
wire t0_010111101010, t0_010111101011;
mixer mix_t0_010111101010 (.a(t0_0101111010100), .b(t0_0101111010101), .y(t0_010111101010));
wire t0_0101111010100, t0_0101111010101;
mixer mix_t0_010111101011 (.a(t0_0101111010110), .b(t0_0101111010111), .y(t0_010111101011));
wire t0_0101111010110, t0_0101111010111;
mixer mix_t0_0101111011 (.a(t0_01011110110), .b(t0_01011110111), .y(t0_0101111011));
wire t0_01011110110, t0_01011110111;
mixer mix_t0_01011110110 (.a(t0_010111101100), .b(t0_010111101101), .y(t0_01011110110));
wire t0_010111101100, t0_010111101101;
mixer mix_t0_010111101100 (.a(t0_0101111011000), .b(t0_0101111011001), .y(t0_010111101100));
wire t0_0101111011000, t0_0101111011001;
mixer mix_t0_010111101101 (.a(t0_0101111011010), .b(t0_0101111011011), .y(t0_010111101101));
wire t0_0101111011010, t0_0101111011011;
mixer mix_t0_01011110111 (.a(t0_010111101110), .b(t0_010111101111), .y(t0_01011110111));
wire t0_010111101110, t0_010111101111;
mixer mix_t0_010111101110 (.a(t0_0101111011100), .b(t0_0101111011101), .y(t0_010111101110));
wire t0_0101111011100, t0_0101111011101;
mixer mix_t0_010111101111 (.a(t0_0101111011110), .b(t0_0101111011111), .y(t0_010111101111));
wire t0_0101111011110, t0_0101111011111;
mixer mix_t0_01011111 (.a(t0_010111110), .b(t0_010111111), .y(t0_01011111));
wire t0_010111110, t0_010111111;
mixer mix_t0_010111110 (.a(t0_0101111100), .b(t0_0101111101), .y(t0_010111110));
wire t0_0101111100, t0_0101111101;
mixer mix_t0_0101111100 (.a(t0_01011111000), .b(t0_01011111001), .y(t0_0101111100));
wire t0_01011111000, t0_01011111001;
mixer mix_t0_01011111000 (.a(t0_010111110000), .b(t0_010111110001), .y(t0_01011111000));
wire t0_010111110000, t0_010111110001;
mixer mix_t0_010111110000 (.a(t0_0101111100000), .b(t0_0101111100001), .y(t0_010111110000));
wire t0_0101111100000, t0_0101111100001;
mixer mix_t0_010111110001 (.a(t0_0101111100010), .b(t0_0101111100011), .y(t0_010111110001));
wire t0_0101111100010, t0_0101111100011;
mixer mix_t0_01011111001 (.a(t0_010111110010), .b(t0_010111110011), .y(t0_01011111001));
wire t0_010111110010, t0_010111110011;
mixer mix_t0_010111110010 (.a(t0_0101111100100), .b(t0_0101111100101), .y(t0_010111110010));
wire t0_0101111100100, t0_0101111100101;
mixer mix_t0_010111110011 (.a(t0_0101111100110), .b(t0_0101111100111), .y(t0_010111110011));
wire t0_0101111100110, t0_0101111100111;
mixer mix_t0_0101111101 (.a(t0_01011111010), .b(t0_01011111011), .y(t0_0101111101));
wire t0_01011111010, t0_01011111011;
mixer mix_t0_01011111010 (.a(t0_010111110100), .b(t0_010111110101), .y(t0_01011111010));
wire t0_010111110100, t0_010111110101;
mixer mix_t0_010111110100 (.a(t0_0101111101000), .b(t0_0101111101001), .y(t0_010111110100));
wire t0_0101111101000, t0_0101111101001;
mixer mix_t0_010111110101 (.a(t0_0101111101010), .b(t0_0101111101011), .y(t0_010111110101));
wire t0_0101111101010, t0_0101111101011;
mixer mix_t0_01011111011 (.a(t0_010111110110), .b(t0_010111110111), .y(t0_01011111011));
wire t0_010111110110, t0_010111110111;
mixer mix_t0_010111110110 (.a(t0_0101111101100), .b(t0_0101111101101), .y(t0_010111110110));
wire t0_0101111101100, t0_0101111101101;
mixer mix_t0_010111110111 (.a(t0_0101111101110), .b(t0_0101111101111), .y(t0_010111110111));
wire t0_0101111101110, t0_0101111101111;
mixer mix_t0_010111111 (.a(t0_0101111110), .b(t0_0101111111), .y(t0_010111111));
wire t0_0101111110, t0_0101111111;
mixer mix_t0_0101111110 (.a(t0_01011111100), .b(t0_01011111101), .y(t0_0101111110));
wire t0_01011111100, t0_01011111101;
mixer mix_t0_01011111100 (.a(t0_010111111000), .b(t0_010111111001), .y(t0_01011111100));
wire t0_010111111000, t0_010111111001;
mixer mix_t0_010111111000 (.a(t0_0101111110000), .b(t0_0101111110001), .y(t0_010111111000));
wire t0_0101111110000, t0_0101111110001;
mixer mix_t0_010111111001 (.a(t0_0101111110010), .b(t0_0101111110011), .y(t0_010111111001));
wire t0_0101111110010, t0_0101111110011;
mixer mix_t0_01011111101 (.a(t0_010111111010), .b(t0_010111111011), .y(t0_01011111101));
wire t0_010111111010, t0_010111111011;
mixer mix_t0_010111111010 (.a(t0_0101111110100), .b(t0_0101111110101), .y(t0_010111111010));
wire t0_0101111110100, t0_0101111110101;
mixer mix_t0_010111111011 (.a(t0_0101111110110), .b(t0_0101111110111), .y(t0_010111111011));
wire t0_0101111110110, t0_0101111110111;
mixer mix_t0_0101111111 (.a(t0_01011111110), .b(t0_01011111111), .y(t0_0101111111));
wire t0_01011111110, t0_01011111111;
mixer mix_t0_01011111110 (.a(t0_010111111100), .b(t0_010111111101), .y(t0_01011111110));
wire t0_010111111100, t0_010111111101;
mixer mix_t0_010111111100 (.a(t0_0101111111000), .b(t0_0101111111001), .y(t0_010111111100));
wire t0_0101111111000, t0_0101111111001;
mixer mix_t0_010111111101 (.a(t0_0101111111010), .b(t0_0101111111011), .y(t0_010111111101));
wire t0_0101111111010, t0_0101111111011;
mixer mix_t0_01011111111 (.a(t0_010111111110), .b(t0_010111111111), .y(t0_01011111111));
wire t0_010111111110, t0_010111111111;
mixer mix_t0_010111111110 (.a(t0_0101111111100), .b(t0_0101111111101), .y(t0_010111111110));
wire t0_0101111111100, t0_0101111111101;
mixer mix_t0_010111111111 (.a(t0_0101111111110), .b(t0_0101111111111), .y(t0_010111111111));
wire t0_0101111111110, t0_0101111111111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_011000 (.a(t0_0110000), .b(t0_0110001), .y(t0_011000));
wire t0_0110000, t0_0110001;
mixer mix_t0_0110000 (.a(t0_01100000), .b(t0_01100001), .y(t0_0110000));
wire t0_01100000, t0_01100001;
mixer mix_t0_01100000 (.a(t0_011000000), .b(t0_011000001), .y(t0_01100000));
wire t0_011000000, t0_011000001;
mixer mix_t0_011000000 (.a(t0_0110000000), .b(t0_0110000001), .y(t0_011000000));
wire t0_0110000000, t0_0110000001;
mixer mix_t0_0110000000 (.a(t0_01100000000), .b(t0_01100000001), .y(t0_0110000000));
wire t0_01100000000, t0_01100000001;
mixer mix_t0_01100000000 (.a(t0_011000000000), .b(t0_011000000001), .y(t0_01100000000));
wire t0_011000000000, t0_011000000001;
mixer mix_t0_011000000000 (.a(t0_0110000000000), .b(t0_0110000000001), .y(t0_011000000000));
wire t0_0110000000000, t0_0110000000001;
mixer mix_t0_011000000001 (.a(t0_0110000000010), .b(t0_0110000000011), .y(t0_011000000001));
wire t0_0110000000010, t0_0110000000011;
mixer mix_t0_01100000001 (.a(t0_011000000010), .b(t0_011000000011), .y(t0_01100000001));
wire t0_011000000010, t0_011000000011;
mixer mix_t0_011000000010 (.a(t0_0110000000100), .b(t0_0110000000101), .y(t0_011000000010));
wire t0_0110000000100, t0_0110000000101;
mixer mix_t0_011000000011 (.a(t0_0110000000110), .b(t0_0110000000111), .y(t0_011000000011));
wire t0_0110000000110, t0_0110000000111;
mixer mix_t0_0110000001 (.a(t0_01100000010), .b(t0_01100000011), .y(t0_0110000001));
wire t0_01100000010, t0_01100000011;
mixer mix_t0_01100000010 (.a(t0_011000000100), .b(t0_011000000101), .y(t0_01100000010));
wire t0_011000000100, t0_011000000101;
mixer mix_t0_011000000100 (.a(t0_0110000001000), .b(t0_0110000001001), .y(t0_011000000100));
wire t0_0110000001000, t0_0110000001001;
mixer mix_t0_011000000101 (.a(t0_0110000001010), .b(t0_0110000001011), .y(t0_011000000101));
wire t0_0110000001010, t0_0110000001011;
mixer mix_t0_01100000011 (.a(t0_011000000110), .b(t0_011000000111), .y(t0_01100000011));
wire t0_011000000110, t0_011000000111;
mixer mix_t0_011000000110 (.a(t0_0110000001100), .b(t0_0110000001101), .y(t0_011000000110));
wire t0_0110000001100, t0_0110000001101;
mixer mix_t0_011000000111 (.a(t0_0110000001110), .b(t0_0110000001111), .y(t0_011000000111));
wire t0_0110000001110, t0_0110000001111;
mixer mix_t0_011000001 (.a(t0_0110000010), .b(t0_0110000011), .y(t0_011000001));
wire t0_0110000010, t0_0110000011;
mixer mix_t0_0110000010 (.a(t0_01100000100), .b(t0_01100000101), .y(t0_0110000010));
wire t0_01100000100, t0_01100000101;
mixer mix_t0_01100000100 (.a(t0_011000001000), .b(t0_011000001001), .y(t0_01100000100));
wire t0_011000001000, t0_011000001001;
mixer mix_t0_011000001000 (.a(t0_0110000010000), .b(t0_0110000010001), .y(t0_011000001000));
wire t0_0110000010000, t0_0110000010001;
mixer mix_t0_011000001001 (.a(t0_0110000010010), .b(t0_0110000010011), .y(t0_011000001001));
wire t0_0110000010010, t0_0110000010011;
mixer mix_t0_01100000101 (.a(t0_011000001010), .b(t0_011000001011), .y(t0_01100000101));
wire t0_011000001010, t0_011000001011;
mixer mix_t0_011000001010 (.a(t0_0110000010100), .b(t0_0110000010101), .y(t0_011000001010));
wire t0_0110000010100, t0_0110000010101;
mixer mix_t0_011000001011 (.a(t0_0110000010110), .b(t0_0110000010111), .y(t0_011000001011));
wire t0_0110000010110, t0_0110000010111;
mixer mix_t0_0110000011 (.a(t0_01100000110), .b(t0_01100000111), .y(t0_0110000011));
wire t0_01100000110, t0_01100000111;
mixer mix_t0_01100000110 (.a(t0_011000001100), .b(t0_011000001101), .y(t0_01100000110));
wire t0_011000001100, t0_011000001101;
mixer mix_t0_011000001100 (.a(t0_0110000011000), .b(t0_0110000011001), .y(t0_011000001100));
wire t0_0110000011000, t0_0110000011001;
mixer mix_t0_011000001101 (.a(t0_0110000011010), .b(t0_0110000011011), .y(t0_011000001101));
wire t0_0110000011010, t0_0110000011011;
mixer mix_t0_01100000111 (.a(t0_011000001110), .b(t0_011000001111), .y(t0_01100000111));
wire t0_011000001110, t0_011000001111;
mixer mix_t0_011000001110 (.a(t0_0110000011100), .b(t0_0110000011101), .y(t0_011000001110));
wire t0_0110000011100, t0_0110000011101;
mixer mix_t0_011000001111 (.a(t0_0110000011110), .b(t0_0110000011111), .y(t0_011000001111));
wire t0_0110000011110, t0_0110000011111;
mixer mix_t0_01100001 (.a(t0_011000010), .b(t0_011000011), .y(t0_01100001));
wire t0_011000010, t0_011000011;
mixer mix_t0_011000010 (.a(t0_0110000100), .b(t0_0110000101), .y(t0_011000010));
wire t0_0110000100, t0_0110000101;
mixer mix_t0_0110000100 (.a(t0_01100001000), .b(t0_01100001001), .y(t0_0110000100));
wire t0_01100001000, t0_01100001001;
mixer mix_t0_01100001000 (.a(t0_011000010000), .b(t0_011000010001), .y(t0_01100001000));
wire t0_011000010000, t0_011000010001;
mixer mix_t0_011000010000 (.a(t0_0110000100000), .b(t0_0110000100001), .y(t0_011000010000));
wire t0_0110000100000, t0_0110000100001;
mixer mix_t0_011000010001 (.a(t0_0110000100010), .b(t0_0110000100011), .y(t0_011000010001));
wire t0_0110000100010, t0_0110000100011;
mixer mix_t0_01100001001 (.a(t0_011000010010), .b(t0_011000010011), .y(t0_01100001001));
wire t0_011000010010, t0_011000010011;
mixer mix_t0_011000010010 (.a(t0_0110000100100), .b(t0_0110000100101), .y(t0_011000010010));
wire t0_0110000100100, t0_0110000100101;
mixer mix_t0_011000010011 (.a(t0_0110000100110), .b(t0_0110000100111), .y(t0_011000010011));
wire t0_0110000100110, t0_0110000100111;
mixer mix_t0_0110000101 (.a(t0_01100001010), .b(t0_01100001011), .y(t0_0110000101));
wire t0_01100001010, t0_01100001011;
mixer mix_t0_01100001010 (.a(t0_011000010100), .b(t0_011000010101), .y(t0_01100001010));
wire t0_011000010100, t0_011000010101;
mixer mix_t0_011000010100 (.a(t0_0110000101000), .b(t0_0110000101001), .y(t0_011000010100));
wire t0_0110000101000, t0_0110000101001;
mixer mix_t0_011000010101 (.a(t0_0110000101010), .b(t0_0110000101011), .y(t0_011000010101));
wire t0_0110000101010, t0_0110000101011;
mixer mix_t0_01100001011 (.a(t0_011000010110), .b(t0_011000010111), .y(t0_01100001011));
wire t0_011000010110, t0_011000010111;
mixer mix_t0_011000010110 (.a(t0_0110000101100), .b(t0_0110000101101), .y(t0_011000010110));
wire t0_0110000101100, t0_0110000101101;
mixer mix_t0_011000010111 (.a(t0_0110000101110), .b(t0_0110000101111), .y(t0_011000010111));
wire t0_0110000101110, t0_0110000101111;
mixer mix_t0_011000011 (.a(t0_0110000110), .b(t0_0110000111), .y(t0_011000011));
wire t0_0110000110, t0_0110000111;
mixer mix_t0_0110000110 (.a(t0_01100001100), .b(t0_01100001101), .y(t0_0110000110));
wire t0_01100001100, t0_01100001101;
mixer mix_t0_01100001100 (.a(t0_011000011000), .b(t0_011000011001), .y(t0_01100001100));
wire t0_011000011000, t0_011000011001;
mixer mix_t0_011000011000 (.a(t0_0110000110000), .b(t0_0110000110001), .y(t0_011000011000));
wire t0_0110000110000, t0_0110000110001;
mixer mix_t0_011000011001 (.a(t0_0110000110010), .b(t0_0110000110011), .y(t0_011000011001));
wire t0_0110000110010, t0_0110000110011;
mixer mix_t0_01100001101 (.a(t0_011000011010), .b(t0_011000011011), .y(t0_01100001101));
wire t0_011000011010, t0_011000011011;
mixer mix_t0_011000011010 (.a(t0_0110000110100), .b(t0_0110000110101), .y(t0_011000011010));
wire t0_0110000110100, t0_0110000110101;
mixer mix_t0_011000011011 (.a(t0_0110000110110), .b(t0_0110000110111), .y(t0_011000011011));
wire t0_0110000110110, t0_0110000110111;
mixer mix_t0_0110000111 (.a(t0_01100001110), .b(t0_01100001111), .y(t0_0110000111));
wire t0_01100001110, t0_01100001111;
mixer mix_t0_01100001110 (.a(t0_011000011100), .b(t0_011000011101), .y(t0_01100001110));
wire t0_011000011100, t0_011000011101;
mixer mix_t0_011000011100 (.a(t0_0110000111000), .b(t0_0110000111001), .y(t0_011000011100));
wire t0_0110000111000, t0_0110000111001;
mixer mix_t0_011000011101 (.a(t0_0110000111010), .b(t0_0110000111011), .y(t0_011000011101));
wire t0_0110000111010, t0_0110000111011;
mixer mix_t0_01100001111 (.a(t0_011000011110), .b(t0_011000011111), .y(t0_01100001111));
wire t0_011000011110, t0_011000011111;
mixer mix_t0_011000011110 (.a(t0_0110000111100), .b(t0_0110000111101), .y(t0_011000011110));
wire t0_0110000111100, t0_0110000111101;
mixer mix_t0_011000011111 (.a(t0_0110000111110), .b(t0_0110000111111), .y(t0_011000011111));
wire t0_0110000111110, t0_0110000111111;
mixer mix_t0_0110001 (.a(t0_01100010), .b(t0_01100011), .y(t0_0110001));
wire t0_01100010, t0_01100011;
mixer mix_t0_01100010 (.a(t0_011000100), .b(t0_011000101), .y(t0_01100010));
wire t0_011000100, t0_011000101;
mixer mix_t0_011000100 (.a(t0_0110001000), .b(t0_0110001001), .y(t0_011000100));
wire t0_0110001000, t0_0110001001;
mixer mix_t0_0110001000 (.a(t0_01100010000), .b(t0_01100010001), .y(t0_0110001000));
wire t0_01100010000, t0_01100010001;
mixer mix_t0_01100010000 (.a(t0_011000100000), .b(t0_011000100001), .y(t0_01100010000));
wire t0_011000100000, t0_011000100001;
mixer mix_t0_011000100000 (.a(t0_0110001000000), .b(t0_0110001000001), .y(t0_011000100000));
wire t0_0110001000000, t0_0110001000001;
mixer mix_t0_011000100001 (.a(t0_0110001000010), .b(t0_0110001000011), .y(t0_011000100001));
wire t0_0110001000010, t0_0110001000011;
mixer mix_t0_01100010001 (.a(t0_011000100010), .b(t0_011000100011), .y(t0_01100010001));
wire t0_011000100010, t0_011000100011;
mixer mix_t0_011000100010 (.a(t0_0110001000100), .b(t0_0110001000101), .y(t0_011000100010));
wire t0_0110001000100, t0_0110001000101;
mixer mix_t0_011000100011 (.a(t0_0110001000110), .b(t0_0110001000111), .y(t0_011000100011));
wire t0_0110001000110, t0_0110001000111;
mixer mix_t0_0110001001 (.a(t0_01100010010), .b(t0_01100010011), .y(t0_0110001001));
wire t0_01100010010, t0_01100010011;
mixer mix_t0_01100010010 (.a(t0_011000100100), .b(t0_011000100101), .y(t0_01100010010));
wire t0_011000100100, t0_011000100101;
mixer mix_t0_011000100100 (.a(t0_0110001001000), .b(t0_0110001001001), .y(t0_011000100100));
wire t0_0110001001000, t0_0110001001001;
mixer mix_t0_011000100101 (.a(t0_0110001001010), .b(t0_0110001001011), .y(t0_011000100101));
wire t0_0110001001010, t0_0110001001011;
mixer mix_t0_01100010011 (.a(t0_011000100110), .b(t0_011000100111), .y(t0_01100010011));
wire t0_011000100110, t0_011000100111;
mixer mix_t0_011000100110 (.a(t0_0110001001100), .b(t0_0110001001101), .y(t0_011000100110));
wire t0_0110001001100, t0_0110001001101;
mixer mix_t0_011000100111 (.a(t0_0110001001110), .b(t0_0110001001111), .y(t0_011000100111));
wire t0_0110001001110, t0_0110001001111;
mixer mix_t0_011000101 (.a(t0_0110001010), .b(t0_0110001011), .y(t0_011000101));
wire t0_0110001010, t0_0110001011;
mixer mix_t0_0110001010 (.a(t0_01100010100), .b(t0_01100010101), .y(t0_0110001010));
wire t0_01100010100, t0_01100010101;
mixer mix_t0_01100010100 (.a(t0_011000101000), .b(t0_011000101001), .y(t0_01100010100));
wire t0_011000101000, t0_011000101001;
mixer mix_t0_011000101000 (.a(t0_0110001010000), .b(t0_0110001010001), .y(t0_011000101000));
wire t0_0110001010000, t0_0110001010001;
mixer mix_t0_011000101001 (.a(t0_0110001010010), .b(t0_0110001010011), .y(t0_011000101001));
wire t0_0110001010010, t0_0110001010011;
mixer mix_t0_01100010101 (.a(t0_011000101010), .b(t0_011000101011), .y(t0_01100010101));
wire t0_011000101010, t0_011000101011;
mixer mix_t0_011000101010 (.a(t0_0110001010100), .b(t0_0110001010101), .y(t0_011000101010));
wire t0_0110001010100, t0_0110001010101;
mixer mix_t0_011000101011 (.a(t0_0110001010110), .b(t0_0110001010111), .y(t0_011000101011));
wire t0_0110001010110, t0_0110001010111;
mixer mix_t0_0110001011 (.a(t0_01100010110), .b(t0_01100010111), .y(t0_0110001011));
wire t0_01100010110, t0_01100010111;
mixer mix_t0_01100010110 (.a(t0_011000101100), .b(t0_011000101101), .y(t0_01100010110));
wire t0_011000101100, t0_011000101101;
mixer mix_t0_011000101100 (.a(t0_0110001011000), .b(t0_0110001011001), .y(t0_011000101100));
wire t0_0110001011000, t0_0110001011001;
mixer mix_t0_011000101101 (.a(t0_0110001011010), .b(t0_0110001011011), .y(t0_011000101101));
wire t0_0110001011010, t0_0110001011011;
mixer mix_t0_01100010111 (.a(t0_011000101110), .b(t0_011000101111), .y(t0_01100010111));
wire t0_011000101110, t0_011000101111;
mixer mix_t0_011000101110 (.a(t0_0110001011100), .b(t0_0110001011101), .y(t0_011000101110));
wire t0_0110001011100, t0_0110001011101;
mixer mix_t0_011000101111 (.a(t0_0110001011110), .b(t0_0110001011111), .y(t0_011000101111));
wire t0_0110001011110, t0_0110001011111;
mixer mix_t0_01100011 (.a(t0_011000110), .b(t0_011000111), .y(t0_01100011));
wire t0_011000110, t0_011000111;
mixer mix_t0_011000110 (.a(t0_0110001100), .b(t0_0110001101), .y(t0_011000110));
wire t0_0110001100, t0_0110001101;
mixer mix_t0_0110001100 (.a(t0_01100011000), .b(t0_01100011001), .y(t0_0110001100));
wire t0_01100011000, t0_01100011001;
mixer mix_t0_01100011000 (.a(t0_011000110000), .b(t0_011000110001), .y(t0_01100011000));
wire t0_011000110000, t0_011000110001;
mixer mix_t0_011000110000 (.a(t0_0110001100000), .b(t0_0110001100001), .y(t0_011000110000));
wire t0_0110001100000, t0_0110001100001;
mixer mix_t0_011000110001 (.a(t0_0110001100010), .b(t0_0110001100011), .y(t0_011000110001));
wire t0_0110001100010, t0_0110001100011;
mixer mix_t0_01100011001 (.a(t0_011000110010), .b(t0_011000110011), .y(t0_01100011001));
wire t0_011000110010, t0_011000110011;
mixer mix_t0_011000110010 (.a(t0_0110001100100), .b(t0_0110001100101), .y(t0_011000110010));
wire t0_0110001100100, t0_0110001100101;
mixer mix_t0_011000110011 (.a(t0_0110001100110), .b(t0_0110001100111), .y(t0_011000110011));
wire t0_0110001100110, t0_0110001100111;
mixer mix_t0_0110001101 (.a(t0_01100011010), .b(t0_01100011011), .y(t0_0110001101));
wire t0_01100011010, t0_01100011011;
mixer mix_t0_01100011010 (.a(t0_011000110100), .b(t0_011000110101), .y(t0_01100011010));
wire t0_011000110100, t0_011000110101;
mixer mix_t0_011000110100 (.a(t0_0110001101000), .b(t0_0110001101001), .y(t0_011000110100));
wire t0_0110001101000, t0_0110001101001;
mixer mix_t0_011000110101 (.a(t0_0110001101010), .b(t0_0110001101011), .y(t0_011000110101));
wire t0_0110001101010, t0_0110001101011;
mixer mix_t0_01100011011 (.a(t0_011000110110), .b(t0_011000110111), .y(t0_01100011011));
wire t0_011000110110, t0_011000110111;
mixer mix_t0_011000110110 (.a(t0_0110001101100), .b(t0_0110001101101), .y(t0_011000110110));
wire t0_0110001101100, t0_0110001101101;
mixer mix_t0_011000110111 (.a(t0_0110001101110), .b(t0_0110001101111), .y(t0_011000110111));
wire t0_0110001101110, t0_0110001101111;
mixer mix_t0_011000111 (.a(t0_0110001110), .b(t0_0110001111), .y(t0_011000111));
wire t0_0110001110, t0_0110001111;
mixer mix_t0_0110001110 (.a(t0_01100011100), .b(t0_01100011101), .y(t0_0110001110));
wire t0_01100011100, t0_01100011101;
mixer mix_t0_01100011100 (.a(t0_011000111000), .b(t0_011000111001), .y(t0_01100011100));
wire t0_011000111000, t0_011000111001;
mixer mix_t0_011000111000 (.a(t0_0110001110000), .b(t0_0110001110001), .y(t0_011000111000));
wire t0_0110001110000, t0_0110001110001;
mixer mix_t0_011000111001 (.a(t0_0110001110010), .b(t0_0110001110011), .y(t0_011000111001));
wire t0_0110001110010, t0_0110001110011;
mixer mix_t0_01100011101 (.a(t0_011000111010), .b(t0_011000111011), .y(t0_01100011101));
wire t0_011000111010, t0_011000111011;
mixer mix_t0_011000111010 (.a(t0_0110001110100), .b(t0_0110001110101), .y(t0_011000111010));
wire t0_0110001110100, t0_0110001110101;
mixer mix_t0_011000111011 (.a(t0_0110001110110), .b(t0_0110001110111), .y(t0_011000111011));
wire t0_0110001110110, t0_0110001110111;
mixer mix_t0_0110001111 (.a(t0_01100011110), .b(t0_01100011111), .y(t0_0110001111));
wire t0_01100011110, t0_01100011111;
mixer mix_t0_01100011110 (.a(t0_011000111100), .b(t0_011000111101), .y(t0_01100011110));
wire t0_011000111100, t0_011000111101;
mixer mix_t0_011000111100 (.a(t0_0110001111000), .b(t0_0110001111001), .y(t0_011000111100));
wire t0_0110001111000, t0_0110001111001;
mixer mix_t0_011000111101 (.a(t0_0110001111010), .b(t0_0110001111011), .y(t0_011000111101));
wire t0_0110001111010, t0_0110001111011;
mixer mix_t0_01100011111 (.a(t0_011000111110), .b(t0_011000111111), .y(t0_01100011111));
wire t0_011000111110, t0_011000111111;
mixer mix_t0_011000111110 (.a(t0_0110001111100), .b(t0_0110001111101), .y(t0_011000111110));
wire t0_0110001111100, t0_0110001111101;
mixer mix_t0_011000111111 (.a(t0_0110001111110), .b(t0_0110001111111), .y(t0_011000111111));
wire t0_0110001111110, t0_0110001111111;
mixer mix_t0_011001 (.a(t0_0110010), .b(t0_0110011), .y(t0_011001));
wire t0_0110010, t0_0110011;
mixer mix_t0_0110010 (.a(t0_01100100), .b(t0_01100101), .y(t0_0110010));
wire t0_01100100, t0_01100101;
mixer mix_t0_01100100 (.a(t0_011001000), .b(t0_011001001), .y(t0_01100100));
wire t0_011001000, t0_011001001;
mixer mix_t0_011001000 (.a(t0_0110010000), .b(t0_0110010001), .y(t0_011001000));
wire t0_0110010000, t0_0110010001;
mixer mix_t0_0110010000 (.a(t0_01100100000), .b(t0_01100100001), .y(t0_0110010000));
wire t0_01100100000, t0_01100100001;
mixer mix_t0_01100100000 (.a(t0_011001000000), .b(t0_011001000001), .y(t0_01100100000));
wire t0_011001000000, t0_011001000001;
mixer mix_t0_011001000000 (.a(t0_0110010000000), .b(t0_0110010000001), .y(t0_011001000000));
wire t0_0110010000000, t0_0110010000001;
mixer mix_t0_011001000001 (.a(t0_0110010000010), .b(t0_0110010000011), .y(t0_011001000001));
wire t0_0110010000010, t0_0110010000011;
mixer mix_t0_01100100001 (.a(t0_011001000010), .b(t0_011001000011), .y(t0_01100100001));
wire t0_011001000010, t0_011001000011;
mixer mix_t0_011001000010 (.a(t0_0110010000100), .b(t0_0110010000101), .y(t0_011001000010));
wire t0_0110010000100, t0_0110010000101;
mixer mix_t0_011001000011 (.a(t0_0110010000110), .b(t0_0110010000111), .y(t0_011001000011));
wire t0_0110010000110, t0_0110010000111;
mixer mix_t0_0110010001 (.a(t0_01100100010), .b(t0_01100100011), .y(t0_0110010001));
wire t0_01100100010, t0_01100100011;
mixer mix_t0_01100100010 (.a(t0_011001000100), .b(t0_011001000101), .y(t0_01100100010));
wire t0_011001000100, t0_011001000101;
mixer mix_t0_011001000100 (.a(t0_0110010001000), .b(t0_0110010001001), .y(t0_011001000100));
wire t0_0110010001000, t0_0110010001001;
mixer mix_t0_011001000101 (.a(t0_0110010001010), .b(t0_0110010001011), .y(t0_011001000101));
wire t0_0110010001010, t0_0110010001011;
mixer mix_t0_01100100011 (.a(t0_011001000110), .b(t0_011001000111), .y(t0_01100100011));
wire t0_011001000110, t0_011001000111;
mixer mix_t0_011001000110 (.a(t0_0110010001100), .b(t0_0110010001101), .y(t0_011001000110));
wire t0_0110010001100, t0_0110010001101;
mixer mix_t0_011001000111 (.a(t0_0110010001110), .b(t0_0110010001111), .y(t0_011001000111));
wire t0_0110010001110, t0_0110010001111;
mixer mix_t0_011001001 (.a(t0_0110010010), .b(t0_0110010011), .y(t0_011001001));
wire t0_0110010010, t0_0110010011;
mixer mix_t0_0110010010 (.a(t0_01100100100), .b(t0_01100100101), .y(t0_0110010010));
wire t0_01100100100, t0_01100100101;
mixer mix_t0_01100100100 (.a(t0_011001001000), .b(t0_011001001001), .y(t0_01100100100));
wire t0_011001001000, t0_011001001001;
mixer mix_t0_011001001000 (.a(t0_0110010010000), .b(t0_0110010010001), .y(t0_011001001000));
wire t0_0110010010000, t0_0110010010001;
mixer mix_t0_011001001001 (.a(t0_0110010010010), .b(t0_0110010010011), .y(t0_011001001001));
wire t0_0110010010010, t0_0110010010011;
mixer mix_t0_01100100101 (.a(t0_011001001010), .b(t0_011001001011), .y(t0_01100100101));
wire t0_011001001010, t0_011001001011;
mixer mix_t0_011001001010 (.a(t0_0110010010100), .b(t0_0110010010101), .y(t0_011001001010));
wire t0_0110010010100, t0_0110010010101;
mixer mix_t0_011001001011 (.a(t0_0110010010110), .b(t0_0110010010111), .y(t0_011001001011));
wire t0_0110010010110, t0_0110010010111;
mixer mix_t0_0110010011 (.a(t0_01100100110), .b(t0_01100100111), .y(t0_0110010011));
wire t0_01100100110, t0_01100100111;
mixer mix_t0_01100100110 (.a(t0_011001001100), .b(t0_011001001101), .y(t0_01100100110));
wire t0_011001001100, t0_011001001101;
mixer mix_t0_011001001100 (.a(t0_0110010011000), .b(t0_0110010011001), .y(t0_011001001100));
wire t0_0110010011000, t0_0110010011001;
mixer mix_t0_011001001101 (.a(t0_0110010011010), .b(t0_0110010011011), .y(t0_011001001101));
wire t0_0110010011010, t0_0110010011011;
mixer mix_t0_01100100111 (.a(t0_011001001110), .b(t0_011001001111), .y(t0_01100100111));
wire t0_011001001110, t0_011001001111;
mixer mix_t0_011001001110 (.a(t0_0110010011100), .b(t0_0110010011101), .y(t0_011001001110));
wire t0_0110010011100, t0_0110010011101;
mixer mix_t0_011001001111 (.a(t0_0110010011110), .b(t0_0110010011111), .y(t0_011001001111));
wire t0_0110010011110, t0_0110010011111;
mixer mix_t0_01100101 (.a(t0_011001010), .b(t0_011001011), .y(t0_01100101));
wire t0_011001010, t0_011001011;
mixer mix_t0_011001010 (.a(t0_0110010100), .b(t0_0110010101), .y(t0_011001010));
wire t0_0110010100, t0_0110010101;
mixer mix_t0_0110010100 (.a(t0_01100101000), .b(t0_01100101001), .y(t0_0110010100));
wire t0_01100101000, t0_01100101001;
mixer mix_t0_01100101000 (.a(t0_011001010000), .b(t0_011001010001), .y(t0_01100101000));
wire t0_011001010000, t0_011001010001;
mixer mix_t0_011001010000 (.a(t0_0110010100000), .b(t0_0110010100001), .y(t0_011001010000));
wire t0_0110010100000, t0_0110010100001;
mixer mix_t0_011001010001 (.a(t0_0110010100010), .b(t0_0110010100011), .y(t0_011001010001));
wire t0_0110010100010, t0_0110010100011;
mixer mix_t0_01100101001 (.a(t0_011001010010), .b(t0_011001010011), .y(t0_01100101001));
wire t0_011001010010, t0_011001010011;
mixer mix_t0_011001010010 (.a(t0_0110010100100), .b(t0_0110010100101), .y(t0_011001010010));
wire t0_0110010100100, t0_0110010100101;
mixer mix_t0_011001010011 (.a(t0_0110010100110), .b(t0_0110010100111), .y(t0_011001010011));
wire t0_0110010100110, t0_0110010100111;
mixer mix_t0_0110010101 (.a(t0_01100101010), .b(t0_01100101011), .y(t0_0110010101));
wire t0_01100101010, t0_01100101011;
mixer mix_t0_01100101010 (.a(t0_011001010100), .b(t0_011001010101), .y(t0_01100101010));
wire t0_011001010100, t0_011001010101;
mixer mix_t0_011001010100 (.a(t0_0110010101000), .b(t0_0110010101001), .y(t0_011001010100));
wire t0_0110010101000, t0_0110010101001;
mixer mix_t0_011001010101 (.a(t0_0110010101010), .b(t0_0110010101011), .y(t0_011001010101));
wire t0_0110010101010, t0_0110010101011;
mixer mix_t0_01100101011 (.a(t0_011001010110), .b(t0_011001010111), .y(t0_01100101011));
wire t0_011001010110, t0_011001010111;
mixer mix_t0_011001010110 (.a(t0_0110010101100), .b(t0_0110010101101), .y(t0_011001010110));
wire t0_0110010101100, t0_0110010101101;
mixer mix_t0_011001010111 (.a(t0_0110010101110), .b(t0_0110010101111), .y(t0_011001010111));
wire t0_0110010101110, t0_0110010101111;
mixer mix_t0_011001011 (.a(t0_0110010110), .b(t0_0110010111), .y(t0_011001011));
wire t0_0110010110, t0_0110010111;
mixer mix_t0_0110010110 (.a(t0_01100101100), .b(t0_01100101101), .y(t0_0110010110));
wire t0_01100101100, t0_01100101101;
mixer mix_t0_01100101100 (.a(t0_011001011000), .b(t0_011001011001), .y(t0_01100101100));
wire t0_011001011000, t0_011001011001;
mixer mix_t0_011001011000 (.a(t0_0110010110000), .b(t0_0110010110001), .y(t0_011001011000));
wire t0_0110010110000, t0_0110010110001;
mixer mix_t0_011001011001 (.a(t0_0110010110010), .b(t0_0110010110011), .y(t0_011001011001));
wire t0_0110010110010, t0_0110010110011;
mixer mix_t0_01100101101 (.a(t0_011001011010), .b(t0_011001011011), .y(t0_01100101101));
wire t0_011001011010, t0_011001011011;
mixer mix_t0_011001011010 (.a(t0_0110010110100), .b(t0_0110010110101), .y(t0_011001011010));
wire t0_0110010110100, t0_0110010110101;
mixer mix_t0_011001011011 (.a(t0_0110010110110), .b(t0_0110010110111), .y(t0_011001011011));
wire t0_0110010110110, t0_0110010110111;
mixer mix_t0_0110010111 (.a(t0_01100101110), .b(t0_01100101111), .y(t0_0110010111));
wire t0_01100101110, t0_01100101111;
mixer mix_t0_01100101110 (.a(t0_011001011100), .b(t0_011001011101), .y(t0_01100101110));
wire t0_011001011100, t0_011001011101;
mixer mix_t0_011001011100 (.a(t0_0110010111000), .b(t0_0110010111001), .y(t0_011001011100));
wire t0_0110010111000, t0_0110010111001;
mixer mix_t0_011001011101 (.a(t0_0110010111010), .b(t0_0110010111011), .y(t0_011001011101));
wire t0_0110010111010, t0_0110010111011;
mixer mix_t0_01100101111 (.a(t0_011001011110), .b(t0_011001011111), .y(t0_01100101111));
wire t0_011001011110, t0_011001011111;
mixer mix_t0_011001011110 (.a(t0_0110010111100), .b(t0_0110010111101), .y(t0_011001011110));
wire t0_0110010111100, t0_0110010111101;
mixer mix_t0_011001011111 (.a(t0_0110010111110), .b(t0_0110010111111), .y(t0_011001011111));
wire t0_0110010111110, t0_0110010111111;
mixer mix_t0_0110011 (.a(t0_01100110), .b(t0_01100111), .y(t0_0110011));
wire t0_01100110, t0_01100111;
mixer mix_t0_01100110 (.a(t0_011001100), .b(t0_011001101), .y(t0_01100110));
wire t0_011001100, t0_011001101;
mixer mix_t0_011001100 (.a(t0_0110011000), .b(t0_0110011001), .y(t0_011001100));
wire t0_0110011000, t0_0110011001;
mixer mix_t0_0110011000 (.a(t0_01100110000), .b(t0_01100110001), .y(t0_0110011000));
wire t0_01100110000, t0_01100110001;
mixer mix_t0_01100110000 (.a(t0_011001100000), .b(t0_011001100001), .y(t0_01100110000));
wire t0_011001100000, t0_011001100001;
mixer mix_t0_011001100000 (.a(t0_0110011000000), .b(t0_0110011000001), .y(t0_011001100000));
wire t0_0110011000000, t0_0110011000001;
mixer mix_t0_011001100001 (.a(t0_0110011000010), .b(t0_0110011000011), .y(t0_011001100001));
wire t0_0110011000010, t0_0110011000011;
mixer mix_t0_01100110001 (.a(t0_011001100010), .b(t0_011001100011), .y(t0_01100110001));
wire t0_011001100010, t0_011001100011;
mixer mix_t0_011001100010 (.a(t0_0110011000100), .b(t0_0110011000101), .y(t0_011001100010));
wire t0_0110011000100, t0_0110011000101;
mixer mix_t0_011001100011 (.a(t0_0110011000110), .b(t0_0110011000111), .y(t0_011001100011));
wire t0_0110011000110, t0_0110011000111;
mixer mix_t0_0110011001 (.a(t0_01100110010), .b(t0_01100110011), .y(t0_0110011001));
wire t0_01100110010, t0_01100110011;
mixer mix_t0_01100110010 (.a(t0_011001100100), .b(t0_011001100101), .y(t0_01100110010));
wire t0_011001100100, t0_011001100101;
mixer mix_t0_011001100100 (.a(t0_0110011001000), .b(t0_0110011001001), .y(t0_011001100100));
wire t0_0110011001000, t0_0110011001001;
mixer mix_t0_011001100101 (.a(t0_0110011001010), .b(t0_0110011001011), .y(t0_011001100101));
wire t0_0110011001010, t0_0110011001011;
mixer mix_t0_01100110011 (.a(t0_011001100110), .b(t0_011001100111), .y(t0_01100110011));
wire t0_011001100110, t0_011001100111;
mixer mix_t0_011001100110 (.a(t0_0110011001100), .b(t0_0110011001101), .y(t0_011001100110));
wire t0_0110011001100, t0_0110011001101;
mixer mix_t0_011001100111 (.a(t0_0110011001110), .b(t0_0110011001111), .y(t0_011001100111));
wire t0_0110011001110, t0_0110011001111;
mixer mix_t0_011001101 (.a(t0_0110011010), .b(t0_0110011011), .y(t0_011001101));
wire t0_0110011010, t0_0110011011;
mixer mix_t0_0110011010 (.a(t0_01100110100), .b(t0_01100110101), .y(t0_0110011010));
wire t0_01100110100, t0_01100110101;
mixer mix_t0_01100110100 (.a(t0_011001101000), .b(t0_011001101001), .y(t0_01100110100));
wire t0_011001101000, t0_011001101001;
mixer mix_t0_011001101000 (.a(t0_0110011010000), .b(t0_0110011010001), .y(t0_011001101000));
wire t0_0110011010000, t0_0110011010001;
mixer mix_t0_011001101001 (.a(t0_0110011010010), .b(t0_0110011010011), .y(t0_011001101001));
wire t0_0110011010010, t0_0110011010011;
mixer mix_t0_01100110101 (.a(t0_011001101010), .b(t0_011001101011), .y(t0_01100110101));
wire t0_011001101010, t0_011001101011;
mixer mix_t0_011001101010 (.a(t0_0110011010100), .b(t0_0110011010101), .y(t0_011001101010));
wire t0_0110011010100, t0_0110011010101;
mixer mix_t0_011001101011 (.a(t0_0110011010110), .b(t0_0110011010111), .y(t0_011001101011));
wire t0_0110011010110, t0_0110011010111;
mixer mix_t0_0110011011 (.a(t0_01100110110), .b(t0_01100110111), .y(t0_0110011011));
wire t0_01100110110, t0_01100110111;
mixer mix_t0_01100110110 (.a(t0_011001101100), .b(t0_011001101101), .y(t0_01100110110));
wire t0_011001101100, t0_011001101101;
mixer mix_t0_011001101100 (.a(t0_0110011011000), .b(t0_0110011011001), .y(t0_011001101100));
wire t0_0110011011000, t0_0110011011001;
mixer mix_t0_011001101101 (.a(t0_0110011011010), .b(t0_0110011011011), .y(t0_011001101101));
wire t0_0110011011010, t0_0110011011011;
mixer mix_t0_01100110111 (.a(t0_011001101110), .b(t0_011001101111), .y(t0_01100110111));
wire t0_011001101110, t0_011001101111;
mixer mix_t0_011001101110 (.a(t0_0110011011100), .b(t0_0110011011101), .y(t0_011001101110));
wire t0_0110011011100, t0_0110011011101;
mixer mix_t0_011001101111 (.a(t0_0110011011110), .b(t0_0110011011111), .y(t0_011001101111));
wire t0_0110011011110, t0_0110011011111;
mixer mix_t0_01100111 (.a(t0_011001110), .b(t0_011001111), .y(t0_01100111));
wire t0_011001110, t0_011001111;
mixer mix_t0_011001110 (.a(t0_0110011100), .b(t0_0110011101), .y(t0_011001110));
wire t0_0110011100, t0_0110011101;
mixer mix_t0_0110011100 (.a(t0_01100111000), .b(t0_01100111001), .y(t0_0110011100));
wire t0_01100111000, t0_01100111001;
mixer mix_t0_01100111000 (.a(t0_011001110000), .b(t0_011001110001), .y(t0_01100111000));
wire t0_011001110000, t0_011001110001;
mixer mix_t0_011001110000 (.a(t0_0110011100000), .b(t0_0110011100001), .y(t0_011001110000));
wire t0_0110011100000, t0_0110011100001;
mixer mix_t0_011001110001 (.a(t0_0110011100010), .b(t0_0110011100011), .y(t0_011001110001));
wire t0_0110011100010, t0_0110011100011;
mixer mix_t0_01100111001 (.a(t0_011001110010), .b(t0_011001110011), .y(t0_01100111001));
wire t0_011001110010, t0_011001110011;
mixer mix_t0_011001110010 (.a(t0_0110011100100), .b(t0_0110011100101), .y(t0_011001110010));
wire t0_0110011100100, t0_0110011100101;
mixer mix_t0_011001110011 (.a(t0_0110011100110), .b(t0_0110011100111), .y(t0_011001110011));
wire t0_0110011100110, t0_0110011100111;
mixer mix_t0_0110011101 (.a(t0_01100111010), .b(t0_01100111011), .y(t0_0110011101));
wire t0_01100111010, t0_01100111011;
mixer mix_t0_01100111010 (.a(t0_011001110100), .b(t0_011001110101), .y(t0_01100111010));
wire t0_011001110100, t0_011001110101;
mixer mix_t0_011001110100 (.a(t0_0110011101000), .b(t0_0110011101001), .y(t0_011001110100));
wire t0_0110011101000, t0_0110011101001;
mixer mix_t0_011001110101 (.a(t0_0110011101010), .b(t0_0110011101011), .y(t0_011001110101));
wire t0_0110011101010, t0_0110011101011;
mixer mix_t0_01100111011 (.a(t0_011001110110), .b(t0_011001110111), .y(t0_01100111011));
wire t0_011001110110, t0_011001110111;
mixer mix_t0_011001110110 (.a(t0_0110011101100), .b(t0_0110011101101), .y(t0_011001110110));
wire t0_0110011101100, t0_0110011101101;
mixer mix_t0_011001110111 (.a(t0_0110011101110), .b(t0_0110011101111), .y(t0_011001110111));
wire t0_0110011101110, t0_0110011101111;
mixer mix_t0_011001111 (.a(t0_0110011110), .b(t0_0110011111), .y(t0_011001111));
wire t0_0110011110, t0_0110011111;
mixer mix_t0_0110011110 (.a(t0_01100111100), .b(t0_01100111101), .y(t0_0110011110));
wire t0_01100111100, t0_01100111101;
mixer mix_t0_01100111100 (.a(t0_011001111000), .b(t0_011001111001), .y(t0_01100111100));
wire t0_011001111000, t0_011001111001;
mixer mix_t0_011001111000 (.a(t0_0110011110000), .b(t0_0110011110001), .y(t0_011001111000));
wire t0_0110011110000, t0_0110011110001;
mixer mix_t0_011001111001 (.a(t0_0110011110010), .b(t0_0110011110011), .y(t0_011001111001));
wire t0_0110011110010, t0_0110011110011;
mixer mix_t0_01100111101 (.a(t0_011001111010), .b(t0_011001111011), .y(t0_01100111101));
wire t0_011001111010, t0_011001111011;
mixer mix_t0_011001111010 (.a(t0_0110011110100), .b(t0_0110011110101), .y(t0_011001111010));
wire t0_0110011110100, t0_0110011110101;
mixer mix_t0_011001111011 (.a(t0_0110011110110), .b(t0_0110011110111), .y(t0_011001111011));
wire t0_0110011110110, t0_0110011110111;
mixer mix_t0_0110011111 (.a(t0_01100111110), .b(t0_01100111111), .y(t0_0110011111));
wire t0_01100111110, t0_01100111111;
mixer mix_t0_01100111110 (.a(t0_011001111100), .b(t0_011001111101), .y(t0_01100111110));
wire t0_011001111100, t0_011001111101;
mixer mix_t0_011001111100 (.a(t0_0110011111000), .b(t0_0110011111001), .y(t0_011001111100));
wire t0_0110011111000, t0_0110011111001;
mixer mix_t0_011001111101 (.a(t0_0110011111010), .b(t0_0110011111011), .y(t0_011001111101));
wire t0_0110011111010, t0_0110011111011;
mixer mix_t0_01100111111 (.a(t0_011001111110), .b(t0_011001111111), .y(t0_01100111111));
wire t0_011001111110, t0_011001111111;
mixer mix_t0_011001111110 (.a(t0_0110011111100), .b(t0_0110011111101), .y(t0_011001111110));
wire t0_0110011111100, t0_0110011111101;
mixer mix_t0_011001111111 (.a(t0_0110011111110), .b(t0_0110011111111), .y(t0_011001111111));
wire t0_0110011111110, t0_0110011111111;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_011010 (.a(t0_0110100), .b(t0_0110101), .y(t0_011010));
wire t0_0110100, t0_0110101;
mixer mix_t0_0110100 (.a(t0_01101000), .b(t0_01101001), .y(t0_0110100));
wire t0_01101000, t0_01101001;
mixer mix_t0_01101000 (.a(t0_011010000), .b(t0_011010001), .y(t0_01101000));
wire t0_011010000, t0_011010001;
mixer mix_t0_011010000 (.a(t0_0110100000), .b(t0_0110100001), .y(t0_011010000));
wire t0_0110100000, t0_0110100001;
mixer mix_t0_0110100000 (.a(t0_01101000000), .b(t0_01101000001), .y(t0_0110100000));
wire t0_01101000000, t0_01101000001;
mixer mix_t0_01101000000 (.a(t0_011010000000), .b(t0_011010000001), .y(t0_01101000000));
wire t0_011010000000, t0_011010000001;
mixer mix_t0_011010000000 (.a(t0_0110100000000), .b(t0_0110100000001), .y(t0_011010000000));
wire t0_0110100000000, t0_0110100000001;
mixer mix_t0_011010000001 (.a(t0_0110100000010), .b(t0_0110100000011), .y(t0_011010000001));
wire t0_0110100000010, t0_0110100000011;
mixer mix_t0_01101000001 (.a(t0_011010000010), .b(t0_011010000011), .y(t0_01101000001));
wire t0_011010000010, t0_011010000011;
mixer mix_t0_011010000010 (.a(t0_0110100000100), .b(t0_0110100000101), .y(t0_011010000010));
wire t0_0110100000100, t0_0110100000101;
mixer mix_t0_011010000011 (.a(t0_0110100000110), .b(t0_0110100000111), .y(t0_011010000011));
wire t0_0110100000110, t0_0110100000111;
mixer mix_t0_0110100001 (.a(t0_01101000010), .b(t0_01101000011), .y(t0_0110100001));
wire t0_01101000010, t0_01101000011;
mixer mix_t0_01101000010 (.a(t0_011010000100), .b(t0_011010000101), .y(t0_01101000010));
wire t0_011010000100, t0_011010000101;
mixer mix_t0_011010000100 (.a(t0_0110100001000), .b(t0_0110100001001), .y(t0_011010000100));
wire t0_0110100001000, t0_0110100001001;
mixer mix_t0_011010000101 (.a(t0_0110100001010), .b(t0_0110100001011), .y(t0_011010000101));
wire t0_0110100001010, t0_0110100001011;
mixer mix_t0_01101000011 (.a(t0_011010000110), .b(t0_011010000111), .y(t0_01101000011));
wire t0_011010000110, t0_011010000111;
mixer mix_t0_011010000110 (.a(t0_0110100001100), .b(t0_0110100001101), .y(t0_011010000110));
wire t0_0110100001100, t0_0110100001101;
mixer mix_t0_011010000111 (.a(t0_0110100001110), .b(t0_0110100001111), .y(t0_011010000111));
wire t0_0110100001110, t0_0110100001111;
mixer mix_t0_011010001 (.a(t0_0110100010), .b(t0_0110100011), .y(t0_011010001));
wire t0_0110100010, t0_0110100011;
mixer mix_t0_0110100010 (.a(t0_01101000100), .b(t0_01101000101), .y(t0_0110100010));
wire t0_01101000100, t0_01101000101;
mixer mix_t0_01101000100 (.a(t0_011010001000), .b(t0_011010001001), .y(t0_01101000100));
wire t0_011010001000, t0_011010001001;
mixer mix_t0_011010001000 (.a(t0_0110100010000), .b(t0_0110100010001), .y(t0_011010001000));
wire t0_0110100010000, t0_0110100010001;
mixer mix_t0_011010001001 (.a(t0_0110100010010), .b(t0_0110100010011), .y(t0_011010001001));
wire t0_0110100010010, t0_0110100010011;
mixer mix_t0_01101000101 (.a(t0_011010001010), .b(t0_011010001011), .y(t0_01101000101));
wire t0_011010001010, t0_011010001011;
mixer mix_t0_011010001010 (.a(t0_0110100010100), .b(t0_0110100010101), .y(t0_011010001010));
wire t0_0110100010100, t0_0110100010101;
mixer mix_t0_011010001011 (.a(t0_0110100010110), .b(t0_0110100010111), .y(t0_011010001011));
wire t0_0110100010110, t0_0110100010111;
mixer mix_t0_0110100011 (.a(t0_01101000110), .b(t0_01101000111), .y(t0_0110100011));
wire t0_01101000110, t0_01101000111;
mixer mix_t0_01101000110 (.a(t0_011010001100), .b(t0_011010001101), .y(t0_01101000110));
wire t0_011010001100, t0_011010001101;
mixer mix_t0_011010001100 (.a(t0_0110100011000), .b(t0_0110100011001), .y(t0_011010001100));
wire t0_0110100011000, t0_0110100011001;
mixer mix_t0_011010001101 (.a(t0_0110100011010), .b(t0_0110100011011), .y(t0_011010001101));
wire t0_0110100011010, t0_0110100011011;
mixer mix_t0_01101000111 (.a(t0_011010001110), .b(t0_011010001111), .y(t0_01101000111));
wire t0_011010001110, t0_011010001111;
mixer mix_t0_011010001110 (.a(t0_0110100011100), .b(t0_0110100011101), .y(t0_011010001110));
wire t0_0110100011100, t0_0110100011101;
mixer mix_t0_011010001111 (.a(t0_0110100011110), .b(t0_0110100011111), .y(t0_011010001111));
wire t0_0110100011110, t0_0110100011111;
mixer mix_t0_01101001 (.a(t0_011010010), .b(t0_011010011), .y(t0_01101001));
wire t0_011010010, t0_011010011;
mixer mix_t0_011010010 (.a(t0_0110100100), .b(t0_0110100101), .y(t0_011010010));
wire t0_0110100100, t0_0110100101;
mixer mix_t0_0110100100 (.a(t0_01101001000), .b(t0_01101001001), .y(t0_0110100100));
wire t0_01101001000, t0_01101001001;
mixer mix_t0_01101001000 (.a(t0_011010010000), .b(t0_011010010001), .y(t0_01101001000));
wire t0_011010010000, t0_011010010001;
mixer mix_t0_011010010000 (.a(t0_0110100100000), .b(t0_0110100100001), .y(t0_011010010000));
wire t0_0110100100000, t0_0110100100001;
mixer mix_t0_011010010001 (.a(t0_0110100100010), .b(t0_0110100100011), .y(t0_011010010001));
wire t0_0110100100010, t0_0110100100011;
mixer mix_t0_01101001001 (.a(t0_011010010010), .b(t0_011010010011), .y(t0_01101001001));
wire t0_011010010010, t0_011010010011;
mixer mix_t0_011010010010 (.a(t0_0110100100100), .b(t0_0110100100101), .y(t0_011010010010));
wire t0_0110100100100, t0_0110100100101;
mixer mix_t0_011010010011 (.a(t0_0110100100110), .b(t0_0110100100111), .y(t0_011010010011));
wire t0_0110100100110, t0_0110100100111;
mixer mix_t0_0110100101 (.a(t0_01101001010), .b(t0_01101001011), .y(t0_0110100101));
wire t0_01101001010, t0_01101001011;
mixer mix_t0_01101001010 (.a(t0_011010010100), .b(t0_011010010101), .y(t0_01101001010));
wire t0_011010010100, t0_011010010101;
mixer mix_t0_011010010100 (.a(t0_0110100101000), .b(t0_0110100101001), .y(t0_011010010100));
wire t0_0110100101000, t0_0110100101001;
mixer mix_t0_011010010101 (.a(t0_0110100101010), .b(t0_0110100101011), .y(t0_011010010101));
wire t0_0110100101010, t0_0110100101011;
mixer mix_t0_01101001011 (.a(t0_011010010110), .b(t0_011010010111), .y(t0_01101001011));
wire t0_011010010110, t0_011010010111;
mixer mix_t0_011010010110 (.a(t0_0110100101100), .b(t0_0110100101101), .y(t0_011010010110));
wire t0_0110100101100, t0_0110100101101;
mixer mix_t0_011010010111 (.a(t0_0110100101110), .b(t0_0110100101111), .y(t0_011010010111));
wire t0_0110100101110, t0_0110100101111;
mixer mix_t0_011010011 (.a(t0_0110100110), .b(t0_0110100111), .y(t0_011010011));
wire t0_0110100110, t0_0110100111;
mixer mix_t0_0110100110 (.a(t0_01101001100), .b(t0_01101001101), .y(t0_0110100110));
wire t0_01101001100, t0_01101001101;
mixer mix_t0_01101001100 (.a(t0_011010011000), .b(t0_011010011001), .y(t0_01101001100));
wire t0_011010011000, t0_011010011001;
mixer mix_t0_011010011000 (.a(t0_0110100110000), .b(t0_0110100110001), .y(t0_011010011000));
wire t0_0110100110000, t0_0110100110001;
mixer mix_t0_011010011001 (.a(t0_0110100110010), .b(t0_0110100110011), .y(t0_011010011001));
wire t0_0110100110010, t0_0110100110011;
mixer mix_t0_01101001101 (.a(t0_011010011010), .b(t0_011010011011), .y(t0_01101001101));
wire t0_011010011010, t0_011010011011;
mixer mix_t0_011010011010 (.a(t0_0110100110100), .b(t0_0110100110101), .y(t0_011010011010));
wire t0_0110100110100, t0_0110100110101;
mixer mix_t0_011010011011 (.a(t0_0110100110110), .b(t0_0110100110111), .y(t0_011010011011));
wire t0_0110100110110, t0_0110100110111;
mixer mix_t0_0110100111 (.a(t0_01101001110), .b(t0_01101001111), .y(t0_0110100111));
wire t0_01101001110, t0_01101001111;
mixer mix_t0_01101001110 (.a(t0_011010011100), .b(t0_011010011101), .y(t0_01101001110));
wire t0_011010011100, t0_011010011101;
mixer mix_t0_011010011100 (.a(t0_0110100111000), .b(t0_0110100111001), .y(t0_011010011100));
wire t0_0110100111000, t0_0110100111001;
mixer mix_t0_011010011101 (.a(t0_0110100111010), .b(t0_0110100111011), .y(t0_011010011101));
wire t0_0110100111010, t0_0110100111011;
mixer mix_t0_01101001111 (.a(t0_011010011110), .b(t0_011010011111), .y(t0_01101001111));
wire t0_011010011110, t0_011010011111;
mixer mix_t0_011010011110 (.a(t0_0110100111100), .b(t0_0110100111101), .y(t0_011010011110));
wire t0_0110100111100, t0_0110100111101;
mixer mix_t0_011010011111 (.a(t0_0110100111110), .b(t0_0110100111111), .y(t0_011010011111));
wire t0_0110100111110, t0_0110100111111;
mixer mix_t0_0110101 (.a(t0_01101010), .b(t0_01101011), .y(t0_0110101));
wire t0_01101010, t0_01101011;
mixer mix_t0_01101010 (.a(t0_011010100), .b(t0_011010101), .y(t0_01101010));
wire t0_011010100, t0_011010101;
mixer mix_t0_011010100 (.a(t0_0110101000), .b(t0_0110101001), .y(t0_011010100));
wire t0_0110101000, t0_0110101001;
mixer mix_t0_0110101000 (.a(t0_01101010000), .b(t0_01101010001), .y(t0_0110101000));
wire t0_01101010000, t0_01101010001;
mixer mix_t0_01101010000 (.a(t0_011010100000), .b(t0_011010100001), .y(t0_01101010000));
wire t0_011010100000, t0_011010100001;
mixer mix_t0_011010100000 (.a(t0_0110101000000), .b(t0_0110101000001), .y(t0_011010100000));
wire t0_0110101000000, t0_0110101000001;
mixer mix_t0_011010100001 (.a(t0_0110101000010), .b(t0_0110101000011), .y(t0_011010100001));
wire t0_0110101000010, t0_0110101000011;
mixer mix_t0_01101010001 (.a(t0_011010100010), .b(t0_011010100011), .y(t0_01101010001));
wire t0_011010100010, t0_011010100011;
mixer mix_t0_011010100010 (.a(t0_0110101000100), .b(t0_0110101000101), .y(t0_011010100010));
wire t0_0110101000100, t0_0110101000101;
mixer mix_t0_011010100011 (.a(t0_0110101000110), .b(t0_0110101000111), .y(t0_011010100011));
wire t0_0110101000110, t0_0110101000111;
mixer mix_t0_0110101001 (.a(t0_01101010010), .b(t0_01101010011), .y(t0_0110101001));
wire t0_01101010010, t0_01101010011;
mixer mix_t0_01101010010 (.a(t0_011010100100), .b(t0_011010100101), .y(t0_01101010010));
wire t0_011010100100, t0_011010100101;
mixer mix_t0_011010100100 (.a(t0_0110101001000), .b(t0_0110101001001), .y(t0_011010100100));
wire t0_0110101001000, t0_0110101001001;
mixer mix_t0_011010100101 (.a(t0_0110101001010), .b(t0_0110101001011), .y(t0_011010100101));
wire t0_0110101001010, t0_0110101001011;
mixer mix_t0_01101010011 (.a(t0_011010100110), .b(t0_011010100111), .y(t0_01101010011));
wire t0_011010100110, t0_011010100111;
mixer mix_t0_011010100110 (.a(t0_0110101001100), .b(t0_0110101001101), .y(t0_011010100110));
wire t0_0110101001100, t0_0110101001101;
mixer mix_t0_011010100111 (.a(t0_0110101001110), .b(t0_0110101001111), .y(t0_011010100111));
wire t0_0110101001110, t0_0110101001111;
mixer mix_t0_011010101 (.a(t0_0110101010), .b(t0_0110101011), .y(t0_011010101));
wire t0_0110101010, t0_0110101011;
mixer mix_t0_0110101010 (.a(t0_01101010100), .b(t0_01101010101), .y(t0_0110101010));
wire t0_01101010100, t0_01101010101;
mixer mix_t0_01101010100 (.a(t0_011010101000), .b(t0_011010101001), .y(t0_01101010100));
wire t0_011010101000, t0_011010101001;
mixer mix_t0_011010101000 (.a(t0_0110101010000), .b(t0_0110101010001), .y(t0_011010101000));
wire t0_0110101010000, t0_0110101010001;
mixer mix_t0_011010101001 (.a(t0_0110101010010), .b(t0_0110101010011), .y(t0_011010101001));
wire t0_0110101010010, t0_0110101010011;
mixer mix_t0_01101010101 (.a(t0_011010101010), .b(t0_011010101011), .y(t0_01101010101));
wire t0_011010101010, t0_011010101011;
mixer mix_t0_011010101010 (.a(t0_0110101010100), .b(t0_0110101010101), .y(t0_011010101010));
wire t0_0110101010100, t0_0110101010101;
mixer mix_t0_011010101011 (.a(t0_0110101010110), .b(t0_0110101010111), .y(t0_011010101011));
wire t0_0110101010110, t0_0110101010111;
mixer mix_t0_0110101011 (.a(t0_01101010110), .b(t0_01101010111), .y(t0_0110101011));
wire t0_01101010110, t0_01101010111;
mixer mix_t0_01101010110 (.a(t0_011010101100), .b(t0_011010101101), .y(t0_01101010110));
wire t0_011010101100, t0_011010101101;
mixer mix_t0_011010101100 (.a(t0_0110101011000), .b(t0_0110101011001), .y(t0_011010101100));
wire t0_0110101011000, t0_0110101011001;
mixer mix_t0_011010101101 (.a(t0_0110101011010), .b(t0_0110101011011), .y(t0_011010101101));
wire t0_0110101011010, t0_0110101011011;
mixer mix_t0_01101010111 (.a(t0_011010101110), .b(t0_011010101111), .y(t0_01101010111));
wire t0_011010101110, t0_011010101111;
mixer mix_t0_011010101110 (.a(t0_0110101011100), .b(t0_0110101011101), .y(t0_011010101110));
wire t0_0110101011100, t0_0110101011101;
mixer mix_t0_011010101111 (.a(t0_0110101011110), .b(t0_0110101011111), .y(t0_011010101111));
wire t0_0110101011110, t0_0110101011111;
mixer mix_t0_01101011 (.a(t0_011010110), .b(t0_011010111), .y(t0_01101011));
wire t0_011010110, t0_011010111;
mixer mix_t0_011010110 (.a(t0_0110101100), .b(t0_0110101101), .y(t0_011010110));
wire t0_0110101100, t0_0110101101;
mixer mix_t0_0110101100 (.a(t0_01101011000), .b(t0_01101011001), .y(t0_0110101100));
wire t0_01101011000, t0_01101011001;
mixer mix_t0_01101011000 (.a(t0_011010110000), .b(t0_011010110001), .y(t0_01101011000));
wire t0_011010110000, t0_011010110001;
mixer mix_t0_011010110000 (.a(t0_0110101100000), .b(t0_0110101100001), .y(t0_011010110000));
wire t0_0110101100000, t0_0110101100001;
mixer mix_t0_011010110001 (.a(t0_0110101100010), .b(t0_0110101100011), .y(t0_011010110001));
wire t0_0110101100010, t0_0110101100011;
mixer mix_t0_01101011001 (.a(t0_011010110010), .b(t0_011010110011), .y(t0_01101011001));
wire t0_011010110010, t0_011010110011;
mixer mix_t0_011010110010 (.a(t0_0110101100100), .b(t0_0110101100101), .y(t0_011010110010));
wire t0_0110101100100, t0_0110101100101;
mixer mix_t0_011010110011 (.a(t0_0110101100110), .b(t0_0110101100111), .y(t0_011010110011));
wire t0_0110101100110, t0_0110101100111;
mixer mix_t0_0110101101 (.a(t0_01101011010), .b(t0_01101011011), .y(t0_0110101101));
wire t0_01101011010, t0_01101011011;
mixer mix_t0_01101011010 (.a(t0_011010110100), .b(t0_011010110101), .y(t0_01101011010));
wire t0_011010110100, t0_011010110101;
mixer mix_t0_011010110100 (.a(t0_0110101101000), .b(t0_0110101101001), .y(t0_011010110100));
wire t0_0110101101000, t0_0110101101001;
mixer mix_t0_011010110101 (.a(t0_0110101101010), .b(t0_0110101101011), .y(t0_011010110101));
wire t0_0110101101010, t0_0110101101011;
mixer mix_t0_01101011011 (.a(t0_011010110110), .b(t0_011010110111), .y(t0_01101011011));
wire t0_011010110110, t0_011010110111;
mixer mix_t0_011010110110 (.a(t0_0110101101100), .b(t0_0110101101101), .y(t0_011010110110));
wire t0_0110101101100, t0_0110101101101;
mixer mix_t0_011010110111 (.a(t0_0110101101110), .b(t0_0110101101111), .y(t0_011010110111));
wire t0_0110101101110, t0_0110101101111;
mixer mix_t0_011010111 (.a(t0_0110101110), .b(t0_0110101111), .y(t0_011010111));
wire t0_0110101110, t0_0110101111;
mixer mix_t0_0110101110 (.a(t0_01101011100), .b(t0_01101011101), .y(t0_0110101110));
wire t0_01101011100, t0_01101011101;
mixer mix_t0_01101011100 (.a(t0_011010111000), .b(t0_011010111001), .y(t0_01101011100));
wire t0_011010111000, t0_011010111001;
mixer mix_t0_011010111000 (.a(t0_0110101110000), .b(t0_0110101110001), .y(t0_011010111000));
wire t0_0110101110000, t0_0110101110001;
mixer mix_t0_011010111001 (.a(t0_0110101110010), .b(t0_0110101110011), .y(t0_011010111001));
wire t0_0110101110010, t0_0110101110011;
mixer mix_t0_01101011101 (.a(t0_011010111010), .b(t0_011010111011), .y(t0_01101011101));
wire t0_011010111010, t0_011010111011;
mixer mix_t0_011010111010 (.a(t0_0110101110100), .b(t0_0110101110101), .y(t0_011010111010));
wire t0_0110101110100, t0_0110101110101;
mixer mix_t0_011010111011 (.a(t0_0110101110110), .b(t0_0110101110111), .y(t0_011010111011));
wire t0_0110101110110, t0_0110101110111;
mixer mix_t0_0110101111 (.a(t0_01101011110), .b(t0_01101011111), .y(t0_0110101111));
wire t0_01101011110, t0_01101011111;
mixer mix_t0_01101011110 (.a(t0_011010111100), .b(t0_011010111101), .y(t0_01101011110));
wire t0_011010111100, t0_011010111101;
mixer mix_t0_011010111100 (.a(t0_0110101111000), .b(t0_0110101111001), .y(t0_011010111100));
wire t0_0110101111000, t0_0110101111001;
mixer mix_t0_011010111101 (.a(t0_0110101111010), .b(t0_0110101111011), .y(t0_011010111101));
wire t0_0110101111010, t0_0110101111011;
mixer mix_t0_01101011111 (.a(t0_011010111110), .b(t0_011010111111), .y(t0_01101011111));
wire t0_011010111110, t0_011010111111;
mixer mix_t0_011010111110 (.a(t0_0110101111100), .b(t0_0110101111101), .y(t0_011010111110));
wire t0_0110101111100, t0_0110101111101;
mixer mix_t0_011010111111 (.a(t0_0110101111110), .b(t0_0110101111111), .y(t0_011010111111));
wire t0_0110101111110, t0_0110101111111;
mixer mix_t0_011011 (.a(t0_0110110), .b(t0_0110111), .y(t0_011011));
wire t0_0110110, t0_0110111;
mixer mix_t0_0110110 (.a(t0_01101100), .b(t0_01101101), .y(t0_0110110));
wire t0_01101100, t0_01101101;
mixer mix_t0_01101100 (.a(t0_011011000), .b(t0_011011001), .y(t0_01101100));
wire t0_011011000, t0_011011001;
mixer mix_t0_011011000 (.a(t0_0110110000), .b(t0_0110110001), .y(t0_011011000));
wire t0_0110110000, t0_0110110001;
mixer mix_t0_0110110000 (.a(t0_01101100000), .b(t0_01101100001), .y(t0_0110110000));
wire t0_01101100000, t0_01101100001;
mixer mix_t0_01101100000 (.a(t0_011011000000), .b(t0_011011000001), .y(t0_01101100000));
wire t0_011011000000, t0_011011000001;
mixer mix_t0_011011000000 (.a(t0_0110110000000), .b(t0_0110110000001), .y(t0_011011000000));
wire t0_0110110000000, t0_0110110000001;
mixer mix_t0_011011000001 (.a(t0_0110110000010), .b(t0_0110110000011), .y(t0_011011000001));
wire t0_0110110000010, t0_0110110000011;
mixer mix_t0_01101100001 (.a(t0_011011000010), .b(t0_011011000011), .y(t0_01101100001));
wire t0_011011000010, t0_011011000011;
mixer mix_t0_011011000010 (.a(t0_0110110000100), .b(t0_0110110000101), .y(t0_011011000010));
wire t0_0110110000100, t0_0110110000101;
mixer mix_t0_011011000011 (.a(t0_0110110000110), .b(t0_0110110000111), .y(t0_011011000011));
wire t0_0110110000110, t0_0110110000111;
mixer mix_t0_0110110001 (.a(t0_01101100010), .b(t0_01101100011), .y(t0_0110110001));
wire t0_01101100010, t0_01101100011;
mixer mix_t0_01101100010 (.a(t0_011011000100), .b(t0_011011000101), .y(t0_01101100010));
wire t0_011011000100, t0_011011000101;
mixer mix_t0_011011000100 (.a(t0_0110110001000), .b(t0_0110110001001), .y(t0_011011000100));
wire t0_0110110001000, t0_0110110001001;
mixer mix_t0_011011000101 (.a(t0_0110110001010), .b(t0_0110110001011), .y(t0_011011000101));
wire t0_0110110001010, t0_0110110001011;
mixer mix_t0_01101100011 (.a(t0_011011000110), .b(t0_011011000111), .y(t0_01101100011));
wire t0_011011000110, t0_011011000111;
mixer mix_t0_011011000110 (.a(t0_0110110001100), .b(t0_0110110001101), .y(t0_011011000110));
wire t0_0110110001100, t0_0110110001101;
mixer mix_t0_011011000111 (.a(t0_0110110001110), .b(t0_0110110001111), .y(t0_011011000111));
wire t0_0110110001110, t0_0110110001111;
mixer mix_t0_011011001 (.a(t0_0110110010), .b(t0_0110110011), .y(t0_011011001));
wire t0_0110110010, t0_0110110011;
mixer mix_t0_0110110010 (.a(t0_01101100100), .b(t0_01101100101), .y(t0_0110110010));
wire t0_01101100100, t0_01101100101;
mixer mix_t0_01101100100 (.a(t0_011011001000), .b(t0_011011001001), .y(t0_01101100100));
wire t0_011011001000, t0_011011001001;
mixer mix_t0_011011001000 (.a(t0_0110110010000), .b(t0_0110110010001), .y(t0_011011001000));
wire t0_0110110010000, t0_0110110010001;
mixer mix_t0_011011001001 (.a(t0_0110110010010), .b(t0_0110110010011), .y(t0_011011001001));
wire t0_0110110010010, t0_0110110010011;
mixer mix_t0_01101100101 (.a(t0_011011001010), .b(t0_011011001011), .y(t0_01101100101));
wire t0_011011001010, t0_011011001011;
mixer mix_t0_011011001010 (.a(t0_0110110010100), .b(t0_0110110010101), .y(t0_011011001010));
wire t0_0110110010100, t0_0110110010101;
mixer mix_t0_011011001011 (.a(t0_0110110010110), .b(t0_0110110010111), .y(t0_011011001011));
wire t0_0110110010110, t0_0110110010111;
mixer mix_t0_0110110011 (.a(t0_01101100110), .b(t0_01101100111), .y(t0_0110110011));
wire t0_01101100110, t0_01101100111;
mixer mix_t0_01101100110 (.a(t0_011011001100), .b(t0_011011001101), .y(t0_01101100110));
wire t0_011011001100, t0_011011001101;
mixer mix_t0_011011001100 (.a(t0_0110110011000), .b(t0_0110110011001), .y(t0_011011001100));
wire t0_0110110011000, t0_0110110011001;
mixer mix_t0_011011001101 (.a(t0_0110110011010), .b(t0_0110110011011), .y(t0_011011001101));
wire t0_0110110011010, t0_0110110011011;
mixer mix_t0_01101100111 (.a(t0_011011001110), .b(t0_011011001111), .y(t0_01101100111));
wire t0_011011001110, t0_011011001111;
mixer mix_t0_011011001110 (.a(t0_0110110011100), .b(t0_0110110011101), .y(t0_011011001110));
wire t0_0110110011100, t0_0110110011101;
mixer mix_t0_011011001111 (.a(t0_0110110011110), .b(t0_0110110011111), .y(t0_011011001111));
wire t0_0110110011110, t0_0110110011111;
mixer mix_t0_01101101 (.a(t0_011011010), .b(t0_011011011), .y(t0_01101101));
wire t0_011011010, t0_011011011;
mixer mix_t0_011011010 (.a(t0_0110110100), .b(t0_0110110101), .y(t0_011011010));
wire t0_0110110100, t0_0110110101;
mixer mix_t0_0110110100 (.a(t0_01101101000), .b(t0_01101101001), .y(t0_0110110100));
wire t0_01101101000, t0_01101101001;
mixer mix_t0_01101101000 (.a(t0_011011010000), .b(t0_011011010001), .y(t0_01101101000));
wire t0_011011010000, t0_011011010001;
mixer mix_t0_011011010000 (.a(t0_0110110100000), .b(t0_0110110100001), .y(t0_011011010000));
wire t0_0110110100000, t0_0110110100001;
mixer mix_t0_011011010001 (.a(t0_0110110100010), .b(t0_0110110100011), .y(t0_011011010001));
wire t0_0110110100010, t0_0110110100011;
mixer mix_t0_01101101001 (.a(t0_011011010010), .b(t0_011011010011), .y(t0_01101101001));
wire t0_011011010010, t0_011011010011;
mixer mix_t0_011011010010 (.a(t0_0110110100100), .b(t0_0110110100101), .y(t0_011011010010));
wire t0_0110110100100, t0_0110110100101;
mixer mix_t0_011011010011 (.a(t0_0110110100110), .b(t0_0110110100111), .y(t0_011011010011));
wire t0_0110110100110, t0_0110110100111;
mixer mix_t0_0110110101 (.a(t0_01101101010), .b(t0_01101101011), .y(t0_0110110101));
wire t0_01101101010, t0_01101101011;
mixer mix_t0_01101101010 (.a(t0_011011010100), .b(t0_011011010101), .y(t0_01101101010));
wire t0_011011010100, t0_011011010101;
mixer mix_t0_011011010100 (.a(t0_0110110101000), .b(t0_0110110101001), .y(t0_011011010100));
wire t0_0110110101000, t0_0110110101001;
mixer mix_t0_011011010101 (.a(t0_0110110101010), .b(t0_0110110101011), .y(t0_011011010101));
wire t0_0110110101010, t0_0110110101011;
mixer mix_t0_01101101011 (.a(t0_011011010110), .b(t0_011011010111), .y(t0_01101101011));
wire t0_011011010110, t0_011011010111;
mixer mix_t0_011011010110 (.a(t0_0110110101100), .b(t0_0110110101101), .y(t0_011011010110));
wire t0_0110110101100, t0_0110110101101;
mixer mix_t0_011011010111 (.a(t0_0110110101110), .b(t0_0110110101111), .y(t0_011011010111));
wire t0_0110110101110, t0_0110110101111;
mixer mix_t0_011011011 (.a(t0_0110110110), .b(t0_0110110111), .y(t0_011011011));
wire t0_0110110110, t0_0110110111;
mixer mix_t0_0110110110 (.a(t0_01101101100), .b(t0_01101101101), .y(t0_0110110110));
wire t0_01101101100, t0_01101101101;
mixer mix_t0_01101101100 (.a(t0_011011011000), .b(t0_011011011001), .y(t0_01101101100));
wire t0_011011011000, t0_011011011001;
mixer mix_t0_011011011000 (.a(t0_0110110110000), .b(t0_0110110110001), .y(t0_011011011000));
wire t0_0110110110000, t0_0110110110001;
mixer mix_t0_011011011001 (.a(t0_0110110110010), .b(t0_0110110110011), .y(t0_011011011001));
wire t0_0110110110010, t0_0110110110011;
mixer mix_t0_01101101101 (.a(t0_011011011010), .b(t0_011011011011), .y(t0_01101101101));
wire t0_011011011010, t0_011011011011;
mixer mix_t0_011011011010 (.a(t0_0110110110100), .b(t0_0110110110101), .y(t0_011011011010));
wire t0_0110110110100, t0_0110110110101;
mixer mix_t0_011011011011 (.a(t0_0110110110110), .b(t0_0110110110111), .y(t0_011011011011));
wire t0_0110110110110, t0_0110110110111;
mixer mix_t0_0110110111 (.a(t0_01101101110), .b(t0_01101101111), .y(t0_0110110111));
wire t0_01101101110, t0_01101101111;
mixer mix_t0_01101101110 (.a(t0_011011011100), .b(t0_011011011101), .y(t0_01101101110));
wire t0_011011011100, t0_011011011101;
mixer mix_t0_011011011100 (.a(t0_0110110111000), .b(t0_0110110111001), .y(t0_011011011100));
wire t0_0110110111000, t0_0110110111001;
mixer mix_t0_011011011101 (.a(t0_0110110111010), .b(t0_0110110111011), .y(t0_011011011101));
wire t0_0110110111010, t0_0110110111011;
mixer mix_t0_01101101111 (.a(t0_011011011110), .b(t0_011011011111), .y(t0_01101101111));
wire t0_011011011110, t0_011011011111;
mixer mix_t0_011011011110 (.a(t0_0110110111100), .b(t0_0110110111101), .y(t0_011011011110));
wire t0_0110110111100, t0_0110110111101;
mixer mix_t0_011011011111 (.a(t0_0110110111110), .b(t0_0110110111111), .y(t0_011011011111));
wire t0_0110110111110, t0_0110110111111;
mixer mix_t0_0110111 (.a(t0_01101110), .b(t0_01101111), .y(t0_0110111));
wire t0_01101110, t0_01101111;
mixer mix_t0_01101110 (.a(t0_011011100), .b(t0_011011101), .y(t0_01101110));
wire t0_011011100, t0_011011101;
mixer mix_t0_011011100 (.a(t0_0110111000), .b(t0_0110111001), .y(t0_011011100));
wire t0_0110111000, t0_0110111001;
mixer mix_t0_0110111000 (.a(t0_01101110000), .b(t0_01101110001), .y(t0_0110111000));
wire t0_01101110000, t0_01101110001;
mixer mix_t0_01101110000 (.a(t0_011011100000), .b(t0_011011100001), .y(t0_01101110000));
wire t0_011011100000, t0_011011100001;
mixer mix_t0_011011100000 (.a(t0_0110111000000), .b(t0_0110111000001), .y(t0_011011100000));
wire t0_0110111000000, t0_0110111000001;
mixer mix_t0_011011100001 (.a(t0_0110111000010), .b(t0_0110111000011), .y(t0_011011100001));
wire t0_0110111000010, t0_0110111000011;
mixer mix_t0_01101110001 (.a(t0_011011100010), .b(t0_011011100011), .y(t0_01101110001));
wire t0_011011100010, t0_011011100011;
mixer mix_t0_011011100010 (.a(t0_0110111000100), .b(t0_0110111000101), .y(t0_011011100010));
wire t0_0110111000100, t0_0110111000101;
mixer mix_t0_011011100011 (.a(t0_0110111000110), .b(t0_0110111000111), .y(t0_011011100011));
wire t0_0110111000110, t0_0110111000111;
mixer mix_t0_0110111001 (.a(t0_01101110010), .b(t0_01101110011), .y(t0_0110111001));
wire t0_01101110010, t0_01101110011;
mixer mix_t0_01101110010 (.a(t0_011011100100), .b(t0_011011100101), .y(t0_01101110010));
wire t0_011011100100, t0_011011100101;
mixer mix_t0_011011100100 (.a(t0_0110111001000), .b(t0_0110111001001), .y(t0_011011100100));
wire t0_0110111001000, t0_0110111001001;
mixer mix_t0_011011100101 (.a(t0_0110111001010), .b(t0_0110111001011), .y(t0_011011100101));
wire t0_0110111001010, t0_0110111001011;
mixer mix_t0_01101110011 (.a(t0_011011100110), .b(t0_011011100111), .y(t0_01101110011));
wire t0_011011100110, t0_011011100111;
mixer mix_t0_011011100110 (.a(t0_0110111001100), .b(t0_0110111001101), .y(t0_011011100110));
wire t0_0110111001100, t0_0110111001101;
mixer mix_t0_011011100111 (.a(t0_0110111001110), .b(t0_0110111001111), .y(t0_011011100111));
wire t0_0110111001110, t0_0110111001111;
mixer mix_t0_011011101 (.a(t0_0110111010), .b(t0_0110111011), .y(t0_011011101));
wire t0_0110111010, t0_0110111011;
mixer mix_t0_0110111010 (.a(t0_01101110100), .b(t0_01101110101), .y(t0_0110111010));
wire t0_01101110100, t0_01101110101;
mixer mix_t0_01101110100 (.a(t0_011011101000), .b(t0_011011101001), .y(t0_01101110100));
wire t0_011011101000, t0_011011101001;
mixer mix_t0_011011101000 (.a(t0_0110111010000), .b(t0_0110111010001), .y(t0_011011101000));
wire t0_0110111010000, t0_0110111010001;
mixer mix_t0_011011101001 (.a(t0_0110111010010), .b(t0_0110111010011), .y(t0_011011101001));
wire t0_0110111010010, t0_0110111010011;
mixer mix_t0_01101110101 (.a(t0_011011101010), .b(t0_011011101011), .y(t0_01101110101));
wire t0_011011101010, t0_011011101011;
mixer mix_t0_011011101010 (.a(t0_0110111010100), .b(t0_0110111010101), .y(t0_011011101010));
wire t0_0110111010100, t0_0110111010101;
mixer mix_t0_011011101011 (.a(t0_0110111010110), .b(t0_0110111010111), .y(t0_011011101011));
wire t0_0110111010110, t0_0110111010111;
mixer mix_t0_0110111011 (.a(t0_01101110110), .b(t0_01101110111), .y(t0_0110111011));
wire t0_01101110110, t0_01101110111;
mixer mix_t0_01101110110 (.a(t0_011011101100), .b(t0_011011101101), .y(t0_01101110110));
wire t0_011011101100, t0_011011101101;
mixer mix_t0_011011101100 (.a(t0_0110111011000), .b(t0_0110111011001), .y(t0_011011101100));
wire t0_0110111011000, t0_0110111011001;
mixer mix_t0_011011101101 (.a(t0_0110111011010), .b(t0_0110111011011), .y(t0_011011101101));
wire t0_0110111011010, t0_0110111011011;
mixer mix_t0_01101110111 (.a(t0_011011101110), .b(t0_011011101111), .y(t0_01101110111));
wire t0_011011101110, t0_011011101111;
mixer mix_t0_011011101110 (.a(t0_0110111011100), .b(t0_0110111011101), .y(t0_011011101110));
wire t0_0110111011100, t0_0110111011101;
mixer mix_t0_011011101111 (.a(t0_0110111011110), .b(t0_0110111011111), .y(t0_011011101111));
wire t0_0110111011110, t0_0110111011111;
mixer mix_t0_01101111 (.a(t0_011011110), .b(t0_011011111), .y(t0_01101111));
wire t0_011011110, t0_011011111;
mixer mix_t0_011011110 (.a(t0_0110111100), .b(t0_0110111101), .y(t0_011011110));
wire t0_0110111100, t0_0110111101;
mixer mix_t0_0110111100 (.a(t0_01101111000), .b(t0_01101111001), .y(t0_0110111100));
wire t0_01101111000, t0_01101111001;
mixer mix_t0_01101111000 (.a(t0_011011110000), .b(t0_011011110001), .y(t0_01101111000));
wire t0_011011110000, t0_011011110001;
mixer mix_t0_011011110000 (.a(t0_0110111100000), .b(t0_0110111100001), .y(t0_011011110000));
wire t0_0110111100000, t0_0110111100001;
mixer mix_t0_011011110001 (.a(t0_0110111100010), .b(t0_0110111100011), .y(t0_011011110001));
wire t0_0110111100010, t0_0110111100011;
mixer mix_t0_01101111001 (.a(t0_011011110010), .b(t0_011011110011), .y(t0_01101111001));
wire t0_011011110010, t0_011011110011;
mixer mix_t0_011011110010 (.a(t0_0110111100100), .b(t0_0110111100101), .y(t0_011011110010));
wire t0_0110111100100, t0_0110111100101;
mixer mix_t0_011011110011 (.a(t0_0110111100110), .b(t0_0110111100111), .y(t0_011011110011));
wire t0_0110111100110, t0_0110111100111;
mixer mix_t0_0110111101 (.a(t0_01101111010), .b(t0_01101111011), .y(t0_0110111101));
wire t0_01101111010, t0_01101111011;
mixer mix_t0_01101111010 (.a(t0_011011110100), .b(t0_011011110101), .y(t0_01101111010));
wire t0_011011110100, t0_011011110101;
mixer mix_t0_011011110100 (.a(t0_0110111101000), .b(t0_0110111101001), .y(t0_011011110100));
wire t0_0110111101000, t0_0110111101001;
mixer mix_t0_011011110101 (.a(t0_0110111101010), .b(t0_0110111101011), .y(t0_011011110101));
wire t0_0110111101010, t0_0110111101011;
mixer mix_t0_01101111011 (.a(t0_011011110110), .b(t0_011011110111), .y(t0_01101111011));
wire t0_011011110110, t0_011011110111;
mixer mix_t0_011011110110 (.a(t0_0110111101100), .b(t0_0110111101101), .y(t0_011011110110));
wire t0_0110111101100, t0_0110111101101;
mixer mix_t0_011011110111 (.a(t0_0110111101110), .b(t0_0110111101111), .y(t0_011011110111));
wire t0_0110111101110, t0_0110111101111;
mixer mix_t0_011011111 (.a(t0_0110111110), .b(t0_0110111111), .y(t0_011011111));
wire t0_0110111110, t0_0110111111;
mixer mix_t0_0110111110 (.a(t0_01101111100), .b(t0_01101111101), .y(t0_0110111110));
wire t0_01101111100, t0_01101111101;
mixer mix_t0_01101111100 (.a(t0_011011111000), .b(t0_011011111001), .y(t0_01101111100));
wire t0_011011111000, t0_011011111001;
mixer mix_t0_011011111000 (.a(t0_0110111110000), .b(t0_0110111110001), .y(t0_011011111000));
wire t0_0110111110000, t0_0110111110001;
mixer mix_t0_011011111001 (.a(t0_0110111110010), .b(t0_0110111110011), .y(t0_011011111001));
wire t0_0110111110010, t0_0110111110011;
mixer mix_t0_01101111101 (.a(t0_011011111010), .b(t0_011011111011), .y(t0_01101111101));
wire t0_011011111010, t0_011011111011;
mixer mix_t0_011011111010 (.a(t0_0110111110100), .b(t0_0110111110101), .y(t0_011011111010));
wire t0_0110111110100, t0_0110111110101;
mixer mix_t0_011011111011 (.a(t0_0110111110110), .b(t0_0110111110111), .y(t0_011011111011));
wire t0_0110111110110, t0_0110111110111;
mixer mix_t0_0110111111 (.a(t0_01101111110), .b(t0_01101111111), .y(t0_0110111111));
wire t0_01101111110, t0_01101111111;
mixer mix_t0_01101111110 (.a(t0_011011111100), .b(t0_011011111101), .y(t0_01101111110));
wire t0_011011111100, t0_011011111101;
mixer mix_t0_011011111100 (.a(t0_0110111111000), .b(t0_0110111111001), .y(t0_011011111100));
wire t0_0110111111000, t0_0110111111001;
mixer mix_t0_011011111101 (.a(t0_0110111111010), .b(t0_0110111111011), .y(t0_011011111101));
wire t0_0110111111010, t0_0110111111011;
mixer mix_t0_01101111111 (.a(t0_011011111110), .b(t0_011011111111), .y(t0_01101111111));
wire t0_011011111110, t0_011011111111;
mixer mix_t0_011011111110 (.a(t0_0110111111100), .b(t0_0110111111101), .y(t0_011011111110));
wire t0_0110111111100, t0_0110111111101;
mixer mix_t0_011011111111 (.a(t0_0110111111110), .b(t0_0110111111111), .y(t0_011011111111));
wire t0_0110111111110, t0_0110111111111;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_011100 (.a(t0_0111000), .b(t0_0111001), .y(t0_011100));
wire t0_0111000, t0_0111001;
mixer mix_t0_0111000 (.a(t0_01110000), .b(t0_01110001), .y(t0_0111000));
wire t0_01110000, t0_01110001;
mixer mix_t0_01110000 (.a(t0_011100000), .b(t0_011100001), .y(t0_01110000));
wire t0_011100000, t0_011100001;
mixer mix_t0_011100000 (.a(t0_0111000000), .b(t0_0111000001), .y(t0_011100000));
wire t0_0111000000, t0_0111000001;
mixer mix_t0_0111000000 (.a(t0_01110000000), .b(t0_01110000001), .y(t0_0111000000));
wire t0_01110000000, t0_01110000001;
mixer mix_t0_01110000000 (.a(t0_011100000000), .b(t0_011100000001), .y(t0_01110000000));
wire t0_011100000000, t0_011100000001;
mixer mix_t0_011100000000 (.a(t0_0111000000000), .b(t0_0111000000001), .y(t0_011100000000));
wire t0_0111000000000, t0_0111000000001;
mixer mix_t0_011100000001 (.a(t0_0111000000010), .b(t0_0111000000011), .y(t0_011100000001));
wire t0_0111000000010, t0_0111000000011;
mixer mix_t0_01110000001 (.a(t0_011100000010), .b(t0_011100000011), .y(t0_01110000001));
wire t0_011100000010, t0_011100000011;
mixer mix_t0_011100000010 (.a(t0_0111000000100), .b(t0_0111000000101), .y(t0_011100000010));
wire t0_0111000000100, t0_0111000000101;
mixer mix_t0_011100000011 (.a(t0_0111000000110), .b(t0_0111000000111), .y(t0_011100000011));
wire t0_0111000000110, t0_0111000000111;
mixer mix_t0_0111000001 (.a(t0_01110000010), .b(t0_01110000011), .y(t0_0111000001));
wire t0_01110000010, t0_01110000011;
mixer mix_t0_01110000010 (.a(t0_011100000100), .b(t0_011100000101), .y(t0_01110000010));
wire t0_011100000100, t0_011100000101;
mixer mix_t0_011100000100 (.a(t0_0111000001000), .b(t0_0111000001001), .y(t0_011100000100));
wire t0_0111000001000, t0_0111000001001;
mixer mix_t0_011100000101 (.a(t0_0111000001010), .b(t0_0111000001011), .y(t0_011100000101));
wire t0_0111000001010, t0_0111000001011;
mixer mix_t0_01110000011 (.a(t0_011100000110), .b(t0_011100000111), .y(t0_01110000011));
wire t0_011100000110, t0_011100000111;
mixer mix_t0_011100000110 (.a(t0_0111000001100), .b(t0_0111000001101), .y(t0_011100000110));
wire t0_0111000001100, t0_0111000001101;
mixer mix_t0_011100000111 (.a(t0_0111000001110), .b(t0_0111000001111), .y(t0_011100000111));
wire t0_0111000001110, t0_0111000001111;
mixer mix_t0_011100001 (.a(t0_0111000010), .b(t0_0111000011), .y(t0_011100001));
wire t0_0111000010, t0_0111000011;
mixer mix_t0_0111000010 (.a(t0_01110000100), .b(t0_01110000101), .y(t0_0111000010));
wire t0_01110000100, t0_01110000101;
mixer mix_t0_01110000100 (.a(t0_011100001000), .b(t0_011100001001), .y(t0_01110000100));
wire t0_011100001000, t0_011100001001;
mixer mix_t0_011100001000 (.a(t0_0111000010000), .b(t0_0111000010001), .y(t0_011100001000));
wire t0_0111000010000, t0_0111000010001;
mixer mix_t0_011100001001 (.a(t0_0111000010010), .b(t0_0111000010011), .y(t0_011100001001));
wire t0_0111000010010, t0_0111000010011;
mixer mix_t0_01110000101 (.a(t0_011100001010), .b(t0_011100001011), .y(t0_01110000101));
wire t0_011100001010, t0_011100001011;
mixer mix_t0_011100001010 (.a(t0_0111000010100), .b(t0_0111000010101), .y(t0_011100001010));
wire t0_0111000010100, t0_0111000010101;
mixer mix_t0_011100001011 (.a(t0_0111000010110), .b(t0_0111000010111), .y(t0_011100001011));
wire t0_0111000010110, t0_0111000010111;
mixer mix_t0_0111000011 (.a(t0_01110000110), .b(t0_01110000111), .y(t0_0111000011));
wire t0_01110000110, t0_01110000111;
mixer mix_t0_01110000110 (.a(t0_011100001100), .b(t0_011100001101), .y(t0_01110000110));
wire t0_011100001100, t0_011100001101;
mixer mix_t0_011100001100 (.a(t0_0111000011000), .b(t0_0111000011001), .y(t0_011100001100));
wire t0_0111000011000, t0_0111000011001;
mixer mix_t0_011100001101 (.a(t0_0111000011010), .b(t0_0111000011011), .y(t0_011100001101));
wire t0_0111000011010, t0_0111000011011;
mixer mix_t0_01110000111 (.a(t0_011100001110), .b(t0_011100001111), .y(t0_01110000111));
wire t0_011100001110, t0_011100001111;
mixer mix_t0_011100001110 (.a(t0_0111000011100), .b(t0_0111000011101), .y(t0_011100001110));
wire t0_0111000011100, t0_0111000011101;
mixer mix_t0_011100001111 (.a(t0_0111000011110), .b(t0_0111000011111), .y(t0_011100001111));
wire t0_0111000011110, t0_0111000011111;
mixer mix_t0_01110001 (.a(t0_011100010), .b(t0_011100011), .y(t0_01110001));
wire t0_011100010, t0_011100011;
mixer mix_t0_011100010 (.a(t0_0111000100), .b(t0_0111000101), .y(t0_011100010));
wire t0_0111000100, t0_0111000101;
mixer mix_t0_0111000100 (.a(t0_01110001000), .b(t0_01110001001), .y(t0_0111000100));
wire t0_01110001000, t0_01110001001;
mixer mix_t0_01110001000 (.a(t0_011100010000), .b(t0_011100010001), .y(t0_01110001000));
wire t0_011100010000, t0_011100010001;
mixer mix_t0_011100010000 (.a(t0_0111000100000), .b(t0_0111000100001), .y(t0_011100010000));
wire t0_0111000100000, t0_0111000100001;
mixer mix_t0_011100010001 (.a(t0_0111000100010), .b(t0_0111000100011), .y(t0_011100010001));
wire t0_0111000100010, t0_0111000100011;
mixer mix_t0_01110001001 (.a(t0_011100010010), .b(t0_011100010011), .y(t0_01110001001));
wire t0_011100010010, t0_011100010011;
mixer mix_t0_011100010010 (.a(t0_0111000100100), .b(t0_0111000100101), .y(t0_011100010010));
wire t0_0111000100100, t0_0111000100101;
mixer mix_t0_011100010011 (.a(t0_0111000100110), .b(t0_0111000100111), .y(t0_011100010011));
wire t0_0111000100110, t0_0111000100111;
mixer mix_t0_0111000101 (.a(t0_01110001010), .b(t0_01110001011), .y(t0_0111000101));
wire t0_01110001010, t0_01110001011;
mixer mix_t0_01110001010 (.a(t0_011100010100), .b(t0_011100010101), .y(t0_01110001010));
wire t0_011100010100, t0_011100010101;
mixer mix_t0_011100010100 (.a(t0_0111000101000), .b(t0_0111000101001), .y(t0_011100010100));
wire t0_0111000101000, t0_0111000101001;
mixer mix_t0_011100010101 (.a(t0_0111000101010), .b(t0_0111000101011), .y(t0_011100010101));
wire t0_0111000101010, t0_0111000101011;
mixer mix_t0_01110001011 (.a(t0_011100010110), .b(t0_011100010111), .y(t0_01110001011));
wire t0_011100010110, t0_011100010111;
mixer mix_t0_011100010110 (.a(t0_0111000101100), .b(t0_0111000101101), .y(t0_011100010110));
wire t0_0111000101100, t0_0111000101101;
mixer mix_t0_011100010111 (.a(t0_0111000101110), .b(t0_0111000101111), .y(t0_011100010111));
wire t0_0111000101110, t0_0111000101111;
mixer mix_t0_011100011 (.a(t0_0111000110), .b(t0_0111000111), .y(t0_011100011));
wire t0_0111000110, t0_0111000111;
mixer mix_t0_0111000110 (.a(t0_01110001100), .b(t0_01110001101), .y(t0_0111000110));
wire t0_01110001100, t0_01110001101;
mixer mix_t0_01110001100 (.a(t0_011100011000), .b(t0_011100011001), .y(t0_01110001100));
wire t0_011100011000, t0_011100011001;
mixer mix_t0_011100011000 (.a(t0_0111000110000), .b(t0_0111000110001), .y(t0_011100011000));
wire t0_0111000110000, t0_0111000110001;
mixer mix_t0_011100011001 (.a(t0_0111000110010), .b(t0_0111000110011), .y(t0_011100011001));
wire t0_0111000110010, t0_0111000110011;
mixer mix_t0_01110001101 (.a(t0_011100011010), .b(t0_011100011011), .y(t0_01110001101));
wire t0_011100011010, t0_011100011011;
mixer mix_t0_011100011010 (.a(t0_0111000110100), .b(t0_0111000110101), .y(t0_011100011010));
wire t0_0111000110100, t0_0111000110101;
mixer mix_t0_011100011011 (.a(t0_0111000110110), .b(t0_0111000110111), .y(t0_011100011011));
wire t0_0111000110110, t0_0111000110111;
mixer mix_t0_0111000111 (.a(t0_01110001110), .b(t0_01110001111), .y(t0_0111000111));
wire t0_01110001110, t0_01110001111;
mixer mix_t0_01110001110 (.a(t0_011100011100), .b(t0_011100011101), .y(t0_01110001110));
wire t0_011100011100, t0_011100011101;
mixer mix_t0_011100011100 (.a(t0_0111000111000), .b(t0_0111000111001), .y(t0_011100011100));
wire t0_0111000111000, t0_0111000111001;
mixer mix_t0_011100011101 (.a(t0_0111000111010), .b(t0_0111000111011), .y(t0_011100011101));
wire t0_0111000111010, t0_0111000111011;
mixer mix_t0_01110001111 (.a(t0_011100011110), .b(t0_011100011111), .y(t0_01110001111));
wire t0_011100011110, t0_011100011111;
mixer mix_t0_011100011110 (.a(t0_0111000111100), .b(t0_0111000111101), .y(t0_011100011110));
wire t0_0111000111100, t0_0111000111101;
mixer mix_t0_011100011111 (.a(t0_0111000111110), .b(t0_0111000111111), .y(t0_011100011111));
wire t0_0111000111110, t0_0111000111111;
mixer mix_t0_0111001 (.a(t0_01110010), .b(t0_01110011), .y(t0_0111001));
wire t0_01110010, t0_01110011;
mixer mix_t0_01110010 (.a(t0_011100100), .b(t0_011100101), .y(t0_01110010));
wire t0_011100100, t0_011100101;
mixer mix_t0_011100100 (.a(t0_0111001000), .b(t0_0111001001), .y(t0_011100100));
wire t0_0111001000, t0_0111001001;
mixer mix_t0_0111001000 (.a(t0_01110010000), .b(t0_01110010001), .y(t0_0111001000));
wire t0_01110010000, t0_01110010001;
mixer mix_t0_01110010000 (.a(t0_011100100000), .b(t0_011100100001), .y(t0_01110010000));
wire t0_011100100000, t0_011100100001;
mixer mix_t0_011100100000 (.a(t0_0111001000000), .b(t0_0111001000001), .y(t0_011100100000));
wire t0_0111001000000, t0_0111001000001;
mixer mix_t0_011100100001 (.a(t0_0111001000010), .b(t0_0111001000011), .y(t0_011100100001));
wire t0_0111001000010, t0_0111001000011;
mixer mix_t0_01110010001 (.a(t0_011100100010), .b(t0_011100100011), .y(t0_01110010001));
wire t0_011100100010, t0_011100100011;
mixer mix_t0_011100100010 (.a(t0_0111001000100), .b(t0_0111001000101), .y(t0_011100100010));
wire t0_0111001000100, t0_0111001000101;
mixer mix_t0_011100100011 (.a(t0_0111001000110), .b(t0_0111001000111), .y(t0_011100100011));
wire t0_0111001000110, t0_0111001000111;
mixer mix_t0_0111001001 (.a(t0_01110010010), .b(t0_01110010011), .y(t0_0111001001));
wire t0_01110010010, t0_01110010011;
mixer mix_t0_01110010010 (.a(t0_011100100100), .b(t0_011100100101), .y(t0_01110010010));
wire t0_011100100100, t0_011100100101;
mixer mix_t0_011100100100 (.a(t0_0111001001000), .b(t0_0111001001001), .y(t0_011100100100));
wire t0_0111001001000, t0_0111001001001;
mixer mix_t0_011100100101 (.a(t0_0111001001010), .b(t0_0111001001011), .y(t0_011100100101));
wire t0_0111001001010, t0_0111001001011;
mixer mix_t0_01110010011 (.a(t0_011100100110), .b(t0_011100100111), .y(t0_01110010011));
wire t0_011100100110, t0_011100100111;
mixer mix_t0_011100100110 (.a(t0_0111001001100), .b(t0_0111001001101), .y(t0_011100100110));
wire t0_0111001001100, t0_0111001001101;
mixer mix_t0_011100100111 (.a(t0_0111001001110), .b(t0_0111001001111), .y(t0_011100100111));
wire t0_0111001001110, t0_0111001001111;
mixer mix_t0_011100101 (.a(t0_0111001010), .b(t0_0111001011), .y(t0_011100101));
wire t0_0111001010, t0_0111001011;
mixer mix_t0_0111001010 (.a(t0_01110010100), .b(t0_01110010101), .y(t0_0111001010));
wire t0_01110010100, t0_01110010101;
mixer mix_t0_01110010100 (.a(t0_011100101000), .b(t0_011100101001), .y(t0_01110010100));
wire t0_011100101000, t0_011100101001;
mixer mix_t0_011100101000 (.a(t0_0111001010000), .b(t0_0111001010001), .y(t0_011100101000));
wire t0_0111001010000, t0_0111001010001;
mixer mix_t0_011100101001 (.a(t0_0111001010010), .b(t0_0111001010011), .y(t0_011100101001));
wire t0_0111001010010, t0_0111001010011;
mixer mix_t0_01110010101 (.a(t0_011100101010), .b(t0_011100101011), .y(t0_01110010101));
wire t0_011100101010, t0_011100101011;
mixer mix_t0_011100101010 (.a(t0_0111001010100), .b(t0_0111001010101), .y(t0_011100101010));
wire t0_0111001010100, t0_0111001010101;
mixer mix_t0_011100101011 (.a(t0_0111001010110), .b(t0_0111001010111), .y(t0_011100101011));
wire t0_0111001010110, t0_0111001010111;
mixer mix_t0_0111001011 (.a(t0_01110010110), .b(t0_01110010111), .y(t0_0111001011));
wire t0_01110010110, t0_01110010111;
mixer mix_t0_01110010110 (.a(t0_011100101100), .b(t0_011100101101), .y(t0_01110010110));
wire t0_011100101100, t0_011100101101;
mixer mix_t0_011100101100 (.a(t0_0111001011000), .b(t0_0111001011001), .y(t0_011100101100));
wire t0_0111001011000, t0_0111001011001;
mixer mix_t0_011100101101 (.a(t0_0111001011010), .b(t0_0111001011011), .y(t0_011100101101));
wire t0_0111001011010, t0_0111001011011;
mixer mix_t0_01110010111 (.a(t0_011100101110), .b(t0_011100101111), .y(t0_01110010111));
wire t0_011100101110, t0_011100101111;
mixer mix_t0_011100101110 (.a(t0_0111001011100), .b(t0_0111001011101), .y(t0_011100101110));
wire t0_0111001011100, t0_0111001011101;
mixer mix_t0_011100101111 (.a(t0_0111001011110), .b(t0_0111001011111), .y(t0_011100101111));
wire t0_0111001011110, t0_0111001011111;
mixer mix_t0_01110011 (.a(t0_011100110), .b(t0_011100111), .y(t0_01110011));
wire t0_011100110, t0_011100111;
mixer mix_t0_011100110 (.a(t0_0111001100), .b(t0_0111001101), .y(t0_011100110));
wire t0_0111001100, t0_0111001101;
mixer mix_t0_0111001100 (.a(t0_01110011000), .b(t0_01110011001), .y(t0_0111001100));
wire t0_01110011000, t0_01110011001;
mixer mix_t0_01110011000 (.a(t0_011100110000), .b(t0_011100110001), .y(t0_01110011000));
wire t0_011100110000, t0_011100110001;
mixer mix_t0_011100110000 (.a(t0_0111001100000), .b(t0_0111001100001), .y(t0_011100110000));
wire t0_0111001100000, t0_0111001100001;
mixer mix_t0_011100110001 (.a(t0_0111001100010), .b(t0_0111001100011), .y(t0_011100110001));
wire t0_0111001100010, t0_0111001100011;
mixer mix_t0_01110011001 (.a(t0_011100110010), .b(t0_011100110011), .y(t0_01110011001));
wire t0_011100110010, t0_011100110011;
mixer mix_t0_011100110010 (.a(t0_0111001100100), .b(t0_0111001100101), .y(t0_011100110010));
wire t0_0111001100100, t0_0111001100101;
mixer mix_t0_011100110011 (.a(t0_0111001100110), .b(t0_0111001100111), .y(t0_011100110011));
wire t0_0111001100110, t0_0111001100111;
mixer mix_t0_0111001101 (.a(t0_01110011010), .b(t0_01110011011), .y(t0_0111001101));
wire t0_01110011010, t0_01110011011;
mixer mix_t0_01110011010 (.a(t0_011100110100), .b(t0_011100110101), .y(t0_01110011010));
wire t0_011100110100, t0_011100110101;
mixer mix_t0_011100110100 (.a(t0_0111001101000), .b(t0_0111001101001), .y(t0_011100110100));
wire t0_0111001101000, t0_0111001101001;
mixer mix_t0_011100110101 (.a(t0_0111001101010), .b(t0_0111001101011), .y(t0_011100110101));
wire t0_0111001101010, t0_0111001101011;
mixer mix_t0_01110011011 (.a(t0_011100110110), .b(t0_011100110111), .y(t0_01110011011));
wire t0_011100110110, t0_011100110111;
mixer mix_t0_011100110110 (.a(t0_0111001101100), .b(t0_0111001101101), .y(t0_011100110110));
wire t0_0111001101100, t0_0111001101101;
mixer mix_t0_011100110111 (.a(t0_0111001101110), .b(t0_0111001101111), .y(t0_011100110111));
wire t0_0111001101110, t0_0111001101111;
mixer mix_t0_011100111 (.a(t0_0111001110), .b(t0_0111001111), .y(t0_011100111));
wire t0_0111001110, t0_0111001111;
mixer mix_t0_0111001110 (.a(t0_01110011100), .b(t0_01110011101), .y(t0_0111001110));
wire t0_01110011100, t0_01110011101;
mixer mix_t0_01110011100 (.a(t0_011100111000), .b(t0_011100111001), .y(t0_01110011100));
wire t0_011100111000, t0_011100111001;
mixer mix_t0_011100111000 (.a(t0_0111001110000), .b(t0_0111001110001), .y(t0_011100111000));
wire t0_0111001110000, t0_0111001110001;
mixer mix_t0_011100111001 (.a(t0_0111001110010), .b(t0_0111001110011), .y(t0_011100111001));
wire t0_0111001110010, t0_0111001110011;
mixer mix_t0_01110011101 (.a(t0_011100111010), .b(t0_011100111011), .y(t0_01110011101));
wire t0_011100111010, t0_011100111011;
mixer mix_t0_011100111010 (.a(t0_0111001110100), .b(t0_0111001110101), .y(t0_011100111010));
wire t0_0111001110100, t0_0111001110101;
mixer mix_t0_011100111011 (.a(t0_0111001110110), .b(t0_0111001110111), .y(t0_011100111011));
wire t0_0111001110110, t0_0111001110111;
mixer mix_t0_0111001111 (.a(t0_01110011110), .b(t0_01110011111), .y(t0_0111001111));
wire t0_01110011110, t0_01110011111;
mixer mix_t0_01110011110 (.a(t0_011100111100), .b(t0_011100111101), .y(t0_01110011110));
wire t0_011100111100, t0_011100111101;
mixer mix_t0_011100111100 (.a(t0_0111001111000), .b(t0_0111001111001), .y(t0_011100111100));
wire t0_0111001111000, t0_0111001111001;
mixer mix_t0_011100111101 (.a(t0_0111001111010), .b(t0_0111001111011), .y(t0_011100111101));
wire t0_0111001111010, t0_0111001111011;
mixer mix_t0_01110011111 (.a(t0_011100111110), .b(t0_011100111111), .y(t0_01110011111));
wire t0_011100111110, t0_011100111111;
mixer mix_t0_011100111110 (.a(t0_0111001111100), .b(t0_0111001111101), .y(t0_011100111110));
wire t0_0111001111100, t0_0111001111101;
mixer mix_t0_011100111111 (.a(t0_0111001111110), .b(t0_0111001111111), .y(t0_011100111111));
wire t0_0111001111110, t0_0111001111111;
mixer mix_t0_011101 (.a(t0_0111010), .b(t0_0111011), .y(t0_011101));
wire t0_0111010, t0_0111011;
mixer mix_t0_0111010 (.a(t0_01110100), .b(t0_01110101), .y(t0_0111010));
wire t0_01110100, t0_01110101;
mixer mix_t0_01110100 (.a(t0_011101000), .b(t0_011101001), .y(t0_01110100));
wire t0_011101000, t0_011101001;
mixer mix_t0_011101000 (.a(t0_0111010000), .b(t0_0111010001), .y(t0_011101000));
wire t0_0111010000, t0_0111010001;
mixer mix_t0_0111010000 (.a(t0_01110100000), .b(t0_01110100001), .y(t0_0111010000));
wire t0_01110100000, t0_01110100001;
mixer mix_t0_01110100000 (.a(t0_011101000000), .b(t0_011101000001), .y(t0_01110100000));
wire t0_011101000000, t0_011101000001;
mixer mix_t0_011101000000 (.a(t0_0111010000000), .b(t0_0111010000001), .y(t0_011101000000));
wire t0_0111010000000, t0_0111010000001;
mixer mix_t0_011101000001 (.a(t0_0111010000010), .b(t0_0111010000011), .y(t0_011101000001));
wire t0_0111010000010, t0_0111010000011;
mixer mix_t0_01110100001 (.a(t0_011101000010), .b(t0_011101000011), .y(t0_01110100001));
wire t0_011101000010, t0_011101000011;
mixer mix_t0_011101000010 (.a(t0_0111010000100), .b(t0_0111010000101), .y(t0_011101000010));
wire t0_0111010000100, t0_0111010000101;
mixer mix_t0_011101000011 (.a(t0_0111010000110), .b(t0_0111010000111), .y(t0_011101000011));
wire t0_0111010000110, t0_0111010000111;
mixer mix_t0_0111010001 (.a(t0_01110100010), .b(t0_01110100011), .y(t0_0111010001));
wire t0_01110100010, t0_01110100011;
mixer mix_t0_01110100010 (.a(t0_011101000100), .b(t0_011101000101), .y(t0_01110100010));
wire t0_011101000100, t0_011101000101;
mixer mix_t0_011101000100 (.a(t0_0111010001000), .b(t0_0111010001001), .y(t0_011101000100));
wire t0_0111010001000, t0_0111010001001;
mixer mix_t0_011101000101 (.a(t0_0111010001010), .b(t0_0111010001011), .y(t0_011101000101));
wire t0_0111010001010, t0_0111010001011;
mixer mix_t0_01110100011 (.a(t0_011101000110), .b(t0_011101000111), .y(t0_01110100011));
wire t0_011101000110, t0_011101000111;
mixer mix_t0_011101000110 (.a(t0_0111010001100), .b(t0_0111010001101), .y(t0_011101000110));
wire t0_0111010001100, t0_0111010001101;
mixer mix_t0_011101000111 (.a(t0_0111010001110), .b(t0_0111010001111), .y(t0_011101000111));
wire t0_0111010001110, t0_0111010001111;
mixer mix_t0_011101001 (.a(t0_0111010010), .b(t0_0111010011), .y(t0_011101001));
wire t0_0111010010, t0_0111010011;
mixer mix_t0_0111010010 (.a(t0_01110100100), .b(t0_01110100101), .y(t0_0111010010));
wire t0_01110100100, t0_01110100101;
mixer mix_t0_01110100100 (.a(t0_011101001000), .b(t0_011101001001), .y(t0_01110100100));
wire t0_011101001000, t0_011101001001;
mixer mix_t0_011101001000 (.a(t0_0111010010000), .b(t0_0111010010001), .y(t0_011101001000));
wire t0_0111010010000, t0_0111010010001;
mixer mix_t0_011101001001 (.a(t0_0111010010010), .b(t0_0111010010011), .y(t0_011101001001));
wire t0_0111010010010, t0_0111010010011;
mixer mix_t0_01110100101 (.a(t0_011101001010), .b(t0_011101001011), .y(t0_01110100101));
wire t0_011101001010, t0_011101001011;
mixer mix_t0_011101001010 (.a(t0_0111010010100), .b(t0_0111010010101), .y(t0_011101001010));
wire t0_0111010010100, t0_0111010010101;
mixer mix_t0_011101001011 (.a(t0_0111010010110), .b(t0_0111010010111), .y(t0_011101001011));
wire t0_0111010010110, t0_0111010010111;
mixer mix_t0_0111010011 (.a(t0_01110100110), .b(t0_01110100111), .y(t0_0111010011));
wire t0_01110100110, t0_01110100111;
mixer mix_t0_01110100110 (.a(t0_011101001100), .b(t0_011101001101), .y(t0_01110100110));
wire t0_011101001100, t0_011101001101;
mixer mix_t0_011101001100 (.a(t0_0111010011000), .b(t0_0111010011001), .y(t0_011101001100));
wire t0_0111010011000, t0_0111010011001;
mixer mix_t0_011101001101 (.a(t0_0111010011010), .b(t0_0111010011011), .y(t0_011101001101));
wire t0_0111010011010, t0_0111010011011;
mixer mix_t0_01110100111 (.a(t0_011101001110), .b(t0_011101001111), .y(t0_01110100111));
wire t0_011101001110, t0_011101001111;
mixer mix_t0_011101001110 (.a(t0_0111010011100), .b(t0_0111010011101), .y(t0_011101001110));
wire t0_0111010011100, t0_0111010011101;
mixer mix_t0_011101001111 (.a(t0_0111010011110), .b(t0_0111010011111), .y(t0_011101001111));
wire t0_0111010011110, t0_0111010011111;
mixer mix_t0_01110101 (.a(t0_011101010), .b(t0_011101011), .y(t0_01110101));
wire t0_011101010, t0_011101011;
mixer mix_t0_011101010 (.a(t0_0111010100), .b(t0_0111010101), .y(t0_011101010));
wire t0_0111010100, t0_0111010101;
mixer mix_t0_0111010100 (.a(t0_01110101000), .b(t0_01110101001), .y(t0_0111010100));
wire t0_01110101000, t0_01110101001;
mixer mix_t0_01110101000 (.a(t0_011101010000), .b(t0_011101010001), .y(t0_01110101000));
wire t0_011101010000, t0_011101010001;
mixer mix_t0_011101010000 (.a(t0_0111010100000), .b(t0_0111010100001), .y(t0_011101010000));
wire t0_0111010100000, t0_0111010100001;
mixer mix_t0_011101010001 (.a(t0_0111010100010), .b(t0_0111010100011), .y(t0_011101010001));
wire t0_0111010100010, t0_0111010100011;
mixer mix_t0_01110101001 (.a(t0_011101010010), .b(t0_011101010011), .y(t0_01110101001));
wire t0_011101010010, t0_011101010011;
mixer mix_t0_011101010010 (.a(t0_0111010100100), .b(t0_0111010100101), .y(t0_011101010010));
wire t0_0111010100100, t0_0111010100101;
mixer mix_t0_011101010011 (.a(t0_0111010100110), .b(t0_0111010100111), .y(t0_011101010011));
wire t0_0111010100110, t0_0111010100111;
mixer mix_t0_0111010101 (.a(t0_01110101010), .b(t0_01110101011), .y(t0_0111010101));
wire t0_01110101010, t0_01110101011;
mixer mix_t0_01110101010 (.a(t0_011101010100), .b(t0_011101010101), .y(t0_01110101010));
wire t0_011101010100, t0_011101010101;
mixer mix_t0_011101010100 (.a(t0_0111010101000), .b(t0_0111010101001), .y(t0_011101010100));
wire t0_0111010101000, t0_0111010101001;
mixer mix_t0_011101010101 (.a(t0_0111010101010), .b(t0_0111010101011), .y(t0_011101010101));
wire t0_0111010101010, t0_0111010101011;
mixer mix_t0_01110101011 (.a(t0_011101010110), .b(t0_011101010111), .y(t0_01110101011));
wire t0_011101010110, t0_011101010111;
mixer mix_t0_011101010110 (.a(t0_0111010101100), .b(t0_0111010101101), .y(t0_011101010110));
wire t0_0111010101100, t0_0111010101101;
mixer mix_t0_011101010111 (.a(t0_0111010101110), .b(t0_0111010101111), .y(t0_011101010111));
wire t0_0111010101110, t0_0111010101111;
mixer mix_t0_011101011 (.a(t0_0111010110), .b(t0_0111010111), .y(t0_011101011));
wire t0_0111010110, t0_0111010111;
mixer mix_t0_0111010110 (.a(t0_01110101100), .b(t0_01110101101), .y(t0_0111010110));
wire t0_01110101100, t0_01110101101;
mixer mix_t0_01110101100 (.a(t0_011101011000), .b(t0_011101011001), .y(t0_01110101100));
wire t0_011101011000, t0_011101011001;
mixer mix_t0_011101011000 (.a(t0_0111010110000), .b(t0_0111010110001), .y(t0_011101011000));
wire t0_0111010110000, t0_0111010110001;
mixer mix_t0_011101011001 (.a(t0_0111010110010), .b(t0_0111010110011), .y(t0_011101011001));
wire t0_0111010110010, t0_0111010110011;
mixer mix_t0_01110101101 (.a(t0_011101011010), .b(t0_011101011011), .y(t0_01110101101));
wire t0_011101011010, t0_011101011011;
mixer mix_t0_011101011010 (.a(t0_0111010110100), .b(t0_0111010110101), .y(t0_011101011010));
wire t0_0111010110100, t0_0111010110101;
mixer mix_t0_011101011011 (.a(t0_0111010110110), .b(t0_0111010110111), .y(t0_011101011011));
wire t0_0111010110110, t0_0111010110111;
mixer mix_t0_0111010111 (.a(t0_01110101110), .b(t0_01110101111), .y(t0_0111010111));
wire t0_01110101110, t0_01110101111;
mixer mix_t0_01110101110 (.a(t0_011101011100), .b(t0_011101011101), .y(t0_01110101110));
wire t0_011101011100, t0_011101011101;
mixer mix_t0_011101011100 (.a(t0_0111010111000), .b(t0_0111010111001), .y(t0_011101011100));
wire t0_0111010111000, t0_0111010111001;
mixer mix_t0_011101011101 (.a(t0_0111010111010), .b(t0_0111010111011), .y(t0_011101011101));
wire t0_0111010111010, t0_0111010111011;
mixer mix_t0_01110101111 (.a(t0_011101011110), .b(t0_011101011111), .y(t0_01110101111));
wire t0_011101011110, t0_011101011111;
mixer mix_t0_011101011110 (.a(t0_0111010111100), .b(t0_0111010111101), .y(t0_011101011110));
wire t0_0111010111100, t0_0111010111101;
mixer mix_t0_011101011111 (.a(t0_0111010111110), .b(t0_0111010111111), .y(t0_011101011111));
wire t0_0111010111110, t0_0111010111111;
mixer mix_t0_0111011 (.a(t0_01110110), .b(t0_01110111), .y(t0_0111011));
wire t0_01110110, t0_01110111;
mixer mix_t0_01110110 (.a(t0_011101100), .b(t0_011101101), .y(t0_01110110));
wire t0_011101100, t0_011101101;
mixer mix_t0_011101100 (.a(t0_0111011000), .b(t0_0111011001), .y(t0_011101100));
wire t0_0111011000, t0_0111011001;
mixer mix_t0_0111011000 (.a(t0_01110110000), .b(t0_01110110001), .y(t0_0111011000));
wire t0_01110110000, t0_01110110001;
mixer mix_t0_01110110000 (.a(t0_011101100000), .b(t0_011101100001), .y(t0_01110110000));
wire t0_011101100000, t0_011101100001;
mixer mix_t0_011101100000 (.a(t0_0111011000000), .b(t0_0111011000001), .y(t0_011101100000));
wire t0_0111011000000, t0_0111011000001;
mixer mix_t0_011101100001 (.a(t0_0111011000010), .b(t0_0111011000011), .y(t0_011101100001));
wire t0_0111011000010, t0_0111011000011;
mixer mix_t0_01110110001 (.a(t0_011101100010), .b(t0_011101100011), .y(t0_01110110001));
wire t0_011101100010, t0_011101100011;
mixer mix_t0_011101100010 (.a(t0_0111011000100), .b(t0_0111011000101), .y(t0_011101100010));
wire t0_0111011000100, t0_0111011000101;
mixer mix_t0_011101100011 (.a(t0_0111011000110), .b(t0_0111011000111), .y(t0_011101100011));
wire t0_0111011000110, t0_0111011000111;
mixer mix_t0_0111011001 (.a(t0_01110110010), .b(t0_01110110011), .y(t0_0111011001));
wire t0_01110110010, t0_01110110011;
mixer mix_t0_01110110010 (.a(t0_011101100100), .b(t0_011101100101), .y(t0_01110110010));
wire t0_011101100100, t0_011101100101;
mixer mix_t0_011101100100 (.a(t0_0111011001000), .b(t0_0111011001001), .y(t0_011101100100));
wire t0_0111011001000, t0_0111011001001;
mixer mix_t0_011101100101 (.a(t0_0111011001010), .b(t0_0111011001011), .y(t0_011101100101));
wire t0_0111011001010, t0_0111011001011;
mixer mix_t0_01110110011 (.a(t0_011101100110), .b(t0_011101100111), .y(t0_01110110011));
wire t0_011101100110, t0_011101100111;
mixer mix_t0_011101100110 (.a(t0_0111011001100), .b(t0_0111011001101), .y(t0_011101100110));
wire t0_0111011001100, t0_0111011001101;
mixer mix_t0_011101100111 (.a(t0_0111011001110), .b(t0_0111011001111), .y(t0_011101100111));
wire t0_0111011001110, t0_0111011001111;
mixer mix_t0_011101101 (.a(t0_0111011010), .b(t0_0111011011), .y(t0_011101101));
wire t0_0111011010, t0_0111011011;
mixer mix_t0_0111011010 (.a(t0_01110110100), .b(t0_01110110101), .y(t0_0111011010));
wire t0_01110110100, t0_01110110101;
mixer mix_t0_01110110100 (.a(t0_011101101000), .b(t0_011101101001), .y(t0_01110110100));
wire t0_011101101000, t0_011101101001;
mixer mix_t0_011101101000 (.a(t0_0111011010000), .b(t0_0111011010001), .y(t0_011101101000));
wire t0_0111011010000, t0_0111011010001;
mixer mix_t0_011101101001 (.a(t0_0111011010010), .b(t0_0111011010011), .y(t0_011101101001));
wire t0_0111011010010, t0_0111011010011;
mixer mix_t0_01110110101 (.a(t0_011101101010), .b(t0_011101101011), .y(t0_01110110101));
wire t0_011101101010, t0_011101101011;
mixer mix_t0_011101101010 (.a(t0_0111011010100), .b(t0_0111011010101), .y(t0_011101101010));
wire t0_0111011010100, t0_0111011010101;
mixer mix_t0_011101101011 (.a(t0_0111011010110), .b(t0_0111011010111), .y(t0_011101101011));
wire t0_0111011010110, t0_0111011010111;
mixer mix_t0_0111011011 (.a(t0_01110110110), .b(t0_01110110111), .y(t0_0111011011));
wire t0_01110110110, t0_01110110111;
mixer mix_t0_01110110110 (.a(t0_011101101100), .b(t0_011101101101), .y(t0_01110110110));
wire t0_011101101100, t0_011101101101;
mixer mix_t0_011101101100 (.a(t0_0111011011000), .b(t0_0111011011001), .y(t0_011101101100));
wire t0_0111011011000, t0_0111011011001;
mixer mix_t0_011101101101 (.a(t0_0111011011010), .b(t0_0111011011011), .y(t0_011101101101));
wire t0_0111011011010, t0_0111011011011;
mixer mix_t0_01110110111 (.a(t0_011101101110), .b(t0_011101101111), .y(t0_01110110111));
wire t0_011101101110, t0_011101101111;
mixer mix_t0_011101101110 (.a(t0_0111011011100), .b(t0_0111011011101), .y(t0_011101101110));
wire t0_0111011011100, t0_0111011011101;
mixer mix_t0_011101101111 (.a(t0_0111011011110), .b(t0_0111011011111), .y(t0_011101101111));
wire t0_0111011011110, t0_0111011011111;
mixer mix_t0_01110111 (.a(t0_011101110), .b(t0_011101111), .y(t0_01110111));
wire t0_011101110, t0_011101111;
mixer mix_t0_011101110 (.a(t0_0111011100), .b(t0_0111011101), .y(t0_011101110));
wire t0_0111011100, t0_0111011101;
mixer mix_t0_0111011100 (.a(t0_01110111000), .b(t0_01110111001), .y(t0_0111011100));
wire t0_01110111000, t0_01110111001;
mixer mix_t0_01110111000 (.a(t0_011101110000), .b(t0_011101110001), .y(t0_01110111000));
wire t0_011101110000, t0_011101110001;
mixer mix_t0_011101110000 (.a(t0_0111011100000), .b(t0_0111011100001), .y(t0_011101110000));
wire t0_0111011100000, t0_0111011100001;
mixer mix_t0_011101110001 (.a(t0_0111011100010), .b(t0_0111011100011), .y(t0_011101110001));
wire t0_0111011100010, t0_0111011100011;
mixer mix_t0_01110111001 (.a(t0_011101110010), .b(t0_011101110011), .y(t0_01110111001));
wire t0_011101110010, t0_011101110011;
mixer mix_t0_011101110010 (.a(t0_0111011100100), .b(t0_0111011100101), .y(t0_011101110010));
wire t0_0111011100100, t0_0111011100101;
mixer mix_t0_011101110011 (.a(t0_0111011100110), .b(t0_0111011100111), .y(t0_011101110011));
wire t0_0111011100110, t0_0111011100111;
mixer mix_t0_0111011101 (.a(t0_01110111010), .b(t0_01110111011), .y(t0_0111011101));
wire t0_01110111010, t0_01110111011;
mixer mix_t0_01110111010 (.a(t0_011101110100), .b(t0_011101110101), .y(t0_01110111010));
wire t0_011101110100, t0_011101110101;
mixer mix_t0_011101110100 (.a(t0_0111011101000), .b(t0_0111011101001), .y(t0_011101110100));
wire t0_0111011101000, t0_0111011101001;
mixer mix_t0_011101110101 (.a(t0_0111011101010), .b(t0_0111011101011), .y(t0_011101110101));
wire t0_0111011101010, t0_0111011101011;
mixer mix_t0_01110111011 (.a(t0_011101110110), .b(t0_011101110111), .y(t0_01110111011));
wire t0_011101110110, t0_011101110111;
mixer mix_t0_011101110110 (.a(t0_0111011101100), .b(t0_0111011101101), .y(t0_011101110110));
wire t0_0111011101100, t0_0111011101101;
mixer mix_t0_011101110111 (.a(t0_0111011101110), .b(t0_0111011101111), .y(t0_011101110111));
wire t0_0111011101110, t0_0111011101111;
mixer mix_t0_011101111 (.a(t0_0111011110), .b(t0_0111011111), .y(t0_011101111));
wire t0_0111011110, t0_0111011111;
mixer mix_t0_0111011110 (.a(t0_01110111100), .b(t0_01110111101), .y(t0_0111011110));
wire t0_01110111100, t0_01110111101;
mixer mix_t0_01110111100 (.a(t0_011101111000), .b(t0_011101111001), .y(t0_01110111100));
wire t0_011101111000, t0_011101111001;
mixer mix_t0_011101111000 (.a(t0_0111011110000), .b(t0_0111011110001), .y(t0_011101111000));
wire t0_0111011110000, t0_0111011110001;
mixer mix_t0_011101111001 (.a(t0_0111011110010), .b(t0_0111011110011), .y(t0_011101111001));
wire t0_0111011110010, t0_0111011110011;
mixer mix_t0_01110111101 (.a(t0_011101111010), .b(t0_011101111011), .y(t0_01110111101));
wire t0_011101111010, t0_011101111011;
mixer mix_t0_011101111010 (.a(t0_0111011110100), .b(t0_0111011110101), .y(t0_011101111010));
wire t0_0111011110100, t0_0111011110101;
mixer mix_t0_011101111011 (.a(t0_0111011110110), .b(t0_0111011110111), .y(t0_011101111011));
wire t0_0111011110110, t0_0111011110111;
mixer mix_t0_0111011111 (.a(t0_01110111110), .b(t0_01110111111), .y(t0_0111011111));
wire t0_01110111110, t0_01110111111;
mixer mix_t0_01110111110 (.a(t0_011101111100), .b(t0_011101111101), .y(t0_01110111110));
wire t0_011101111100, t0_011101111101;
mixer mix_t0_011101111100 (.a(t0_0111011111000), .b(t0_0111011111001), .y(t0_011101111100));
wire t0_0111011111000, t0_0111011111001;
mixer mix_t0_011101111101 (.a(t0_0111011111010), .b(t0_0111011111011), .y(t0_011101111101));
wire t0_0111011111010, t0_0111011111011;
mixer mix_t0_01110111111 (.a(t0_011101111110), .b(t0_011101111111), .y(t0_01110111111));
wire t0_011101111110, t0_011101111111;
mixer mix_t0_011101111110 (.a(t0_0111011111100), .b(t0_0111011111101), .y(t0_011101111110));
wire t0_0111011111100, t0_0111011111101;
mixer mix_t0_011101111111 (.a(t0_0111011111110), .b(t0_0111011111111), .y(t0_011101111111));
wire t0_0111011111110, t0_0111011111111;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
mixer mix_t0_011110 (.a(t0_0111100), .b(t0_0111101), .y(t0_011110));
wire t0_0111100, t0_0111101;
mixer mix_t0_0111100 (.a(t0_01111000), .b(t0_01111001), .y(t0_0111100));
wire t0_01111000, t0_01111001;
mixer mix_t0_01111000 (.a(t0_011110000), .b(t0_011110001), .y(t0_01111000));
wire t0_011110000, t0_011110001;
mixer mix_t0_011110000 (.a(t0_0111100000), .b(t0_0111100001), .y(t0_011110000));
wire t0_0111100000, t0_0111100001;
mixer mix_t0_0111100000 (.a(t0_01111000000), .b(t0_01111000001), .y(t0_0111100000));
wire t0_01111000000, t0_01111000001;
mixer mix_t0_01111000000 (.a(t0_011110000000), .b(t0_011110000001), .y(t0_01111000000));
wire t0_011110000000, t0_011110000001;
mixer mix_t0_011110000000 (.a(t0_0111100000000), .b(t0_0111100000001), .y(t0_011110000000));
wire t0_0111100000000, t0_0111100000001;
mixer mix_t0_011110000001 (.a(t0_0111100000010), .b(t0_0111100000011), .y(t0_011110000001));
wire t0_0111100000010, t0_0111100000011;
mixer mix_t0_01111000001 (.a(t0_011110000010), .b(t0_011110000011), .y(t0_01111000001));
wire t0_011110000010, t0_011110000011;
mixer mix_t0_011110000010 (.a(t0_0111100000100), .b(t0_0111100000101), .y(t0_011110000010));
wire t0_0111100000100, t0_0111100000101;
mixer mix_t0_011110000011 (.a(t0_0111100000110), .b(t0_0111100000111), .y(t0_011110000011));
wire t0_0111100000110, t0_0111100000111;
mixer mix_t0_0111100001 (.a(t0_01111000010), .b(t0_01111000011), .y(t0_0111100001));
wire t0_01111000010, t0_01111000011;
mixer mix_t0_01111000010 (.a(t0_011110000100), .b(t0_011110000101), .y(t0_01111000010));
wire t0_011110000100, t0_011110000101;
mixer mix_t0_011110000100 (.a(t0_0111100001000), .b(t0_0111100001001), .y(t0_011110000100));
wire t0_0111100001000, t0_0111100001001;
mixer mix_t0_011110000101 (.a(t0_0111100001010), .b(t0_0111100001011), .y(t0_011110000101));
wire t0_0111100001010, t0_0111100001011;
mixer mix_t0_01111000011 (.a(t0_011110000110), .b(t0_011110000111), .y(t0_01111000011));
wire t0_011110000110, t0_011110000111;
mixer mix_t0_011110000110 (.a(t0_0111100001100), .b(t0_0111100001101), .y(t0_011110000110));
wire t0_0111100001100, t0_0111100001101;
mixer mix_t0_011110000111 (.a(t0_0111100001110), .b(t0_0111100001111), .y(t0_011110000111));
wire t0_0111100001110, t0_0111100001111;
mixer mix_t0_011110001 (.a(t0_0111100010), .b(t0_0111100011), .y(t0_011110001));
wire t0_0111100010, t0_0111100011;
mixer mix_t0_0111100010 (.a(t0_01111000100), .b(t0_01111000101), .y(t0_0111100010));
wire t0_01111000100, t0_01111000101;
mixer mix_t0_01111000100 (.a(t0_011110001000), .b(t0_011110001001), .y(t0_01111000100));
wire t0_011110001000, t0_011110001001;
mixer mix_t0_011110001000 (.a(t0_0111100010000), .b(t0_0111100010001), .y(t0_011110001000));
wire t0_0111100010000, t0_0111100010001;
mixer mix_t0_011110001001 (.a(t0_0111100010010), .b(t0_0111100010011), .y(t0_011110001001));
wire t0_0111100010010, t0_0111100010011;
mixer mix_t0_01111000101 (.a(t0_011110001010), .b(t0_011110001011), .y(t0_01111000101));
wire t0_011110001010, t0_011110001011;
mixer mix_t0_011110001010 (.a(t0_0111100010100), .b(t0_0111100010101), .y(t0_011110001010));
wire t0_0111100010100, t0_0111100010101;
mixer mix_t0_011110001011 (.a(t0_0111100010110), .b(t0_0111100010111), .y(t0_011110001011));
wire t0_0111100010110, t0_0111100010111;
mixer mix_t0_0111100011 (.a(t0_01111000110), .b(t0_01111000111), .y(t0_0111100011));
wire t0_01111000110, t0_01111000111;
mixer mix_t0_01111000110 (.a(t0_011110001100), .b(t0_011110001101), .y(t0_01111000110));
wire t0_011110001100, t0_011110001101;
mixer mix_t0_011110001100 (.a(t0_0111100011000), .b(t0_0111100011001), .y(t0_011110001100));
wire t0_0111100011000, t0_0111100011001;
mixer mix_t0_011110001101 (.a(t0_0111100011010), .b(t0_0111100011011), .y(t0_011110001101));
wire t0_0111100011010, t0_0111100011011;
mixer mix_t0_01111000111 (.a(t0_011110001110), .b(t0_011110001111), .y(t0_01111000111));
wire t0_011110001110, t0_011110001111;
mixer mix_t0_011110001110 (.a(t0_0111100011100), .b(t0_0111100011101), .y(t0_011110001110));
wire t0_0111100011100, t0_0111100011101;
mixer mix_t0_011110001111 (.a(t0_0111100011110), .b(t0_0111100011111), .y(t0_011110001111));
wire t0_0111100011110, t0_0111100011111;
mixer mix_t0_01111001 (.a(t0_011110010), .b(t0_011110011), .y(t0_01111001));
wire t0_011110010, t0_011110011;
mixer mix_t0_011110010 (.a(t0_0111100100), .b(t0_0111100101), .y(t0_011110010));
wire t0_0111100100, t0_0111100101;
mixer mix_t0_0111100100 (.a(t0_01111001000), .b(t0_01111001001), .y(t0_0111100100));
wire t0_01111001000, t0_01111001001;
mixer mix_t0_01111001000 (.a(t0_011110010000), .b(t0_011110010001), .y(t0_01111001000));
wire t0_011110010000, t0_011110010001;
mixer mix_t0_011110010000 (.a(t0_0111100100000), .b(t0_0111100100001), .y(t0_011110010000));
wire t0_0111100100000, t0_0111100100001;
mixer mix_t0_011110010001 (.a(t0_0111100100010), .b(t0_0111100100011), .y(t0_011110010001));
wire t0_0111100100010, t0_0111100100011;
mixer mix_t0_01111001001 (.a(t0_011110010010), .b(t0_011110010011), .y(t0_01111001001));
wire t0_011110010010, t0_011110010011;
mixer mix_t0_011110010010 (.a(t0_0111100100100), .b(t0_0111100100101), .y(t0_011110010010));
wire t0_0111100100100, t0_0111100100101;
mixer mix_t0_011110010011 (.a(t0_0111100100110), .b(t0_0111100100111), .y(t0_011110010011));
wire t0_0111100100110, t0_0111100100111;
mixer mix_t0_0111100101 (.a(t0_01111001010), .b(t0_01111001011), .y(t0_0111100101));
wire t0_01111001010, t0_01111001011;
mixer mix_t0_01111001010 (.a(t0_011110010100), .b(t0_011110010101), .y(t0_01111001010));
wire t0_011110010100, t0_011110010101;
mixer mix_t0_011110010100 (.a(t0_0111100101000), .b(t0_0111100101001), .y(t0_011110010100));
wire t0_0111100101000, t0_0111100101001;
mixer mix_t0_011110010101 (.a(t0_0111100101010), .b(t0_0111100101011), .y(t0_011110010101));
wire t0_0111100101010, t0_0111100101011;
mixer mix_t0_01111001011 (.a(t0_011110010110), .b(t0_011110010111), .y(t0_01111001011));
wire t0_011110010110, t0_011110010111;
mixer mix_t0_011110010110 (.a(t0_0111100101100), .b(t0_0111100101101), .y(t0_011110010110));
wire t0_0111100101100, t0_0111100101101;
mixer mix_t0_011110010111 (.a(t0_0111100101110), .b(t0_0111100101111), .y(t0_011110010111));
wire t0_0111100101110, t0_0111100101111;
mixer mix_t0_011110011 (.a(t0_0111100110), .b(t0_0111100111), .y(t0_011110011));
wire t0_0111100110, t0_0111100111;
mixer mix_t0_0111100110 (.a(t0_01111001100), .b(t0_01111001101), .y(t0_0111100110));
wire t0_01111001100, t0_01111001101;
mixer mix_t0_01111001100 (.a(t0_011110011000), .b(t0_011110011001), .y(t0_01111001100));
wire t0_011110011000, t0_011110011001;
mixer mix_t0_011110011000 (.a(t0_0111100110000), .b(t0_0111100110001), .y(t0_011110011000));
wire t0_0111100110000, t0_0111100110001;
mixer mix_t0_011110011001 (.a(t0_0111100110010), .b(t0_0111100110011), .y(t0_011110011001));
wire t0_0111100110010, t0_0111100110011;
mixer mix_t0_01111001101 (.a(t0_011110011010), .b(t0_011110011011), .y(t0_01111001101));
wire t0_011110011010, t0_011110011011;
mixer mix_t0_011110011010 (.a(t0_0111100110100), .b(t0_0111100110101), .y(t0_011110011010));
wire t0_0111100110100, t0_0111100110101;
mixer mix_t0_011110011011 (.a(t0_0111100110110), .b(t0_0111100110111), .y(t0_011110011011));
wire t0_0111100110110, t0_0111100110111;
mixer mix_t0_0111100111 (.a(t0_01111001110), .b(t0_01111001111), .y(t0_0111100111));
wire t0_01111001110, t0_01111001111;
mixer mix_t0_01111001110 (.a(t0_011110011100), .b(t0_011110011101), .y(t0_01111001110));
wire t0_011110011100, t0_011110011101;
mixer mix_t0_011110011100 (.a(t0_0111100111000), .b(t0_0111100111001), .y(t0_011110011100));
wire t0_0111100111000, t0_0111100111001;
mixer mix_t0_011110011101 (.a(t0_0111100111010), .b(t0_0111100111011), .y(t0_011110011101));
wire t0_0111100111010, t0_0111100111011;
mixer mix_t0_01111001111 (.a(t0_011110011110), .b(t0_011110011111), .y(t0_01111001111));
wire t0_011110011110, t0_011110011111;
mixer mix_t0_011110011110 (.a(t0_0111100111100), .b(t0_0111100111101), .y(t0_011110011110));
wire t0_0111100111100, t0_0111100111101;
mixer mix_t0_011110011111 (.a(t0_0111100111110), .b(t0_0111100111111), .y(t0_011110011111));
wire t0_0111100111110, t0_0111100111111;
mixer mix_t0_0111101 (.a(t0_01111010), .b(t0_01111011), .y(t0_0111101));
wire t0_01111010, t0_01111011;
mixer mix_t0_01111010 (.a(t0_011110100), .b(t0_011110101), .y(t0_01111010));
wire t0_011110100, t0_011110101;
mixer mix_t0_011110100 (.a(t0_0111101000), .b(t0_0111101001), .y(t0_011110100));
wire t0_0111101000, t0_0111101001;
mixer mix_t0_0111101000 (.a(t0_01111010000), .b(t0_01111010001), .y(t0_0111101000));
wire t0_01111010000, t0_01111010001;
mixer mix_t0_01111010000 (.a(t0_011110100000), .b(t0_011110100001), .y(t0_01111010000));
wire t0_011110100000, t0_011110100001;
mixer mix_t0_011110100000 (.a(t0_0111101000000), .b(t0_0111101000001), .y(t0_011110100000));
wire t0_0111101000000, t0_0111101000001;
mixer mix_t0_011110100001 (.a(t0_0111101000010), .b(t0_0111101000011), .y(t0_011110100001));
wire t0_0111101000010, t0_0111101000011;
mixer mix_t0_01111010001 (.a(t0_011110100010), .b(t0_011110100011), .y(t0_01111010001));
wire t0_011110100010, t0_011110100011;
mixer mix_t0_011110100010 (.a(t0_0111101000100), .b(t0_0111101000101), .y(t0_011110100010));
wire t0_0111101000100, t0_0111101000101;
mixer mix_t0_011110100011 (.a(t0_0111101000110), .b(t0_0111101000111), .y(t0_011110100011));
wire t0_0111101000110, t0_0111101000111;
mixer mix_t0_0111101001 (.a(t0_01111010010), .b(t0_01111010011), .y(t0_0111101001));
wire t0_01111010010, t0_01111010011;
mixer mix_t0_01111010010 (.a(t0_011110100100), .b(t0_011110100101), .y(t0_01111010010));
wire t0_011110100100, t0_011110100101;
mixer mix_t0_011110100100 (.a(t0_0111101001000), .b(t0_0111101001001), .y(t0_011110100100));
wire t0_0111101001000, t0_0111101001001;
mixer mix_t0_011110100101 (.a(t0_0111101001010), .b(t0_0111101001011), .y(t0_011110100101));
wire t0_0111101001010, t0_0111101001011;
mixer mix_t0_01111010011 (.a(t0_011110100110), .b(t0_011110100111), .y(t0_01111010011));
wire t0_011110100110, t0_011110100111;
mixer mix_t0_011110100110 (.a(t0_0111101001100), .b(t0_0111101001101), .y(t0_011110100110));
wire t0_0111101001100, t0_0111101001101;
mixer mix_t0_011110100111 (.a(t0_0111101001110), .b(t0_0111101001111), .y(t0_011110100111));
wire t0_0111101001110, t0_0111101001111;
mixer mix_t0_011110101 (.a(t0_0111101010), .b(t0_0111101011), .y(t0_011110101));
wire t0_0111101010, t0_0111101011;
mixer mix_t0_0111101010 (.a(t0_01111010100), .b(t0_01111010101), .y(t0_0111101010));
wire t0_01111010100, t0_01111010101;
mixer mix_t0_01111010100 (.a(t0_011110101000), .b(t0_011110101001), .y(t0_01111010100));
wire t0_011110101000, t0_011110101001;
mixer mix_t0_011110101000 (.a(t0_0111101010000), .b(t0_0111101010001), .y(t0_011110101000));
wire t0_0111101010000, t0_0111101010001;
mixer mix_t0_011110101001 (.a(t0_0111101010010), .b(t0_0111101010011), .y(t0_011110101001));
wire t0_0111101010010, t0_0111101010011;
mixer mix_t0_01111010101 (.a(t0_011110101010), .b(t0_011110101011), .y(t0_01111010101));
wire t0_011110101010, t0_011110101011;
mixer mix_t0_011110101010 (.a(t0_0111101010100), .b(t0_0111101010101), .y(t0_011110101010));
wire t0_0111101010100, t0_0111101010101;
mixer mix_t0_011110101011 (.a(t0_0111101010110), .b(t0_0111101010111), .y(t0_011110101011));
wire t0_0111101010110, t0_0111101010111;
mixer mix_t0_0111101011 (.a(t0_01111010110), .b(t0_01111010111), .y(t0_0111101011));
wire t0_01111010110, t0_01111010111;
mixer mix_t0_01111010110 (.a(t0_011110101100), .b(t0_011110101101), .y(t0_01111010110));
wire t0_011110101100, t0_011110101101;
mixer mix_t0_011110101100 (.a(t0_0111101011000), .b(t0_0111101011001), .y(t0_011110101100));
wire t0_0111101011000, t0_0111101011001;
mixer mix_t0_011110101101 (.a(t0_0111101011010), .b(t0_0111101011011), .y(t0_011110101101));
wire t0_0111101011010, t0_0111101011011;
mixer mix_t0_01111010111 (.a(t0_011110101110), .b(t0_011110101111), .y(t0_01111010111));
wire t0_011110101110, t0_011110101111;
mixer mix_t0_011110101110 (.a(t0_0111101011100), .b(t0_0111101011101), .y(t0_011110101110));
wire t0_0111101011100, t0_0111101011101;
mixer mix_t0_011110101111 (.a(t0_0111101011110), .b(t0_0111101011111), .y(t0_011110101111));
wire t0_0111101011110, t0_0111101011111;
mixer mix_t0_01111011 (.a(t0_011110110), .b(t0_011110111), .y(t0_01111011));
wire t0_011110110, t0_011110111;
mixer mix_t0_011110110 (.a(t0_0111101100), .b(t0_0111101101), .y(t0_011110110));
wire t0_0111101100, t0_0111101101;
mixer mix_t0_0111101100 (.a(t0_01111011000), .b(t0_01111011001), .y(t0_0111101100));
wire t0_01111011000, t0_01111011001;
mixer mix_t0_01111011000 (.a(t0_011110110000), .b(t0_011110110001), .y(t0_01111011000));
wire t0_011110110000, t0_011110110001;
mixer mix_t0_011110110000 (.a(t0_0111101100000), .b(t0_0111101100001), .y(t0_011110110000));
wire t0_0111101100000, t0_0111101100001;
mixer mix_t0_011110110001 (.a(t0_0111101100010), .b(t0_0111101100011), .y(t0_011110110001));
wire t0_0111101100010, t0_0111101100011;
mixer mix_t0_01111011001 (.a(t0_011110110010), .b(t0_011110110011), .y(t0_01111011001));
wire t0_011110110010, t0_011110110011;
mixer mix_t0_011110110010 (.a(t0_0111101100100), .b(t0_0111101100101), .y(t0_011110110010));
wire t0_0111101100100, t0_0111101100101;
mixer mix_t0_011110110011 (.a(t0_0111101100110), .b(t0_0111101100111), .y(t0_011110110011));
wire t0_0111101100110, t0_0111101100111;
mixer mix_t0_0111101101 (.a(t0_01111011010), .b(t0_01111011011), .y(t0_0111101101));
wire t0_01111011010, t0_01111011011;
mixer mix_t0_01111011010 (.a(t0_011110110100), .b(t0_011110110101), .y(t0_01111011010));
wire t0_011110110100, t0_011110110101;
mixer mix_t0_011110110100 (.a(t0_0111101101000), .b(t0_0111101101001), .y(t0_011110110100));
wire t0_0111101101000, t0_0111101101001;
mixer mix_t0_011110110101 (.a(t0_0111101101010), .b(t0_0111101101011), .y(t0_011110110101));
wire t0_0111101101010, t0_0111101101011;
mixer mix_t0_01111011011 (.a(t0_011110110110), .b(t0_011110110111), .y(t0_01111011011));
wire t0_011110110110, t0_011110110111;
mixer mix_t0_011110110110 (.a(t0_0111101101100), .b(t0_0111101101101), .y(t0_011110110110));
wire t0_0111101101100, t0_0111101101101;
mixer mix_t0_011110110111 (.a(t0_0111101101110), .b(t0_0111101101111), .y(t0_011110110111));
wire t0_0111101101110, t0_0111101101111;
mixer mix_t0_011110111 (.a(t0_0111101110), .b(t0_0111101111), .y(t0_011110111));
wire t0_0111101110, t0_0111101111;
mixer mix_t0_0111101110 (.a(t0_01111011100), .b(t0_01111011101), .y(t0_0111101110));
wire t0_01111011100, t0_01111011101;
mixer mix_t0_01111011100 (.a(t0_011110111000), .b(t0_011110111001), .y(t0_01111011100));
wire t0_011110111000, t0_011110111001;
mixer mix_t0_011110111000 (.a(t0_0111101110000), .b(t0_0111101110001), .y(t0_011110111000));
wire t0_0111101110000, t0_0111101110001;
mixer mix_t0_011110111001 (.a(t0_0111101110010), .b(t0_0111101110011), .y(t0_011110111001));
wire t0_0111101110010, t0_0111101110011;
mixer mix_t0_01111011101 (.a(t0_011110111010), .b(t0_011110111011), .y(t0_01111011101));
wire t0_011110111010, t0_011110111011;
mixer mix_t0_011110111010 (.a(t0_0111101110100), .b(t0_0111101110101), .y(t0_011110111010));
wire t0_0111101110100, t0_0111101110101;
mixer mix_t0_011110111011 (.a(t0_0111101110110), .b(t0_0111101110111), .y(t0_011110111011));
wire t0_0111101110110, t0_0111101110111;
mixer mix_t0_0111101111 (.a(t0_01111011110), .b(t0_01111011111), .y(t0_0111101111));
wire t0_01111011110, t0_01111011111;
mixer mix_t0_01111011110 (.a(t0_011110111100), .b(t0_011110111101), .y(t0_01111011110));
wire t0_011110111100, t0_011110111101;
mixer mix_t0_011110111100 (.a(t0_0111101111000), .b(t0_0111101111001), .y(t0_011110111100));
wire t0_0111101111000, t0_0111101111001;
mixer mix_t0_011110111101 (.a(t0_0111101111010), .b(t0_0111101111011), .y(t0_011110111101));
wire t0_0111101111010, t0_0111101111011;
mixer mix_t0_01111011111 (.a(t0_011110111110), .b(t0_011110111111), .y(t0_01111011111));
wire t0_011110111110, t0_011110111111;
mixer mix_t0_011110111110 (.a(t0_0111101111100), .b(t0_0111101111101), .y(t0_011110111110));
wire t0_0111101111100, t0_0111101111101;
mixer mix_t0_011110111111 (.a(t0_0111101111110), .b(t0_0111101111111), .y(t0_011110111111));
wire t0_0111101111110, t0_0111101111111;
mixer mix_t0_011111 (.a(t0_0111110), .b(t0_0111111), .y(t0_011111));
wire t0_0111110, t0_0111111;
mixer mix_t0_0111110 (.a(t0_01111100), .b(t0_01111101), .y(t0_0111110));
wire t0_01111100, t0_01111101;
mixer mix_t0_01111100 (.a(t0_011111000), .b(t0_011111001), .y(t0_01111100));
wire t0_011111000, t0_011111001;
mixer mix_t0_011111000 (.a(t0_0111110000), .b(t0_0111110001), .y(t0_011111000));
wire t0_0111110000, t0_0111110001;
mixer mix_t0_0111110000 (.a(t0_01111100000), .b(t0_01111100001), .y(t0_0111110000));
wire t0_01111100000, t0_01111100001;
mixer mix_t0_01111100000 (.a(t0_011111000000), .b(t0_011111000001), .y(t0_01111100000));
wire t0_011111000000, t0_011111000001;
mixer mix_t0_011111000000 (.a(t0_0111110000000), .b(t0_0111110000001), .y(t0_011111000000));
wire t0_0111110000000, t0_0111110000001;
mixer mix_t0_011111000001 (.a(t0_0111110000010), .b(t0_0111110000011), .y(t0_011111000001));
wire t0_0111110000010, t0_0111110000011;
mixer mix_t0_01111100001 (.a(t0_011111000010), .b(t0_011111000011), .y(t0_01111100001));
wire t0_011111000010, t0_011111000011;
mixer mix_t0_011111000010 (.a(t0_0111110000100), .b(t0_0111110000101), .y(t0_011111000010));
wire t0_0111110000100, t0_0111110000101;
mixer mix_t0_011111000011 (.a(t0_0111110000110), .b(t0_0111110000111), .y(t0_011111000011));
wire t0_0111110000110, t0_0111110000111;
mixer mix_t0_0111110001 (.a(t0_01111100010), .b(t0_01111100011), .y(t0_0111110001));
wire t0_01111100010, t0_01111100011;
mixer mix_t0_01111100010 (.a(t0_011111000100), .b(t0_011111000101), .y(t0_01111100010));
wire t0_011111000100, t0_011111000101;
mixer mix_t0_011111000100 (.a(t0_0111110001000), .b(t0_0111110001001), .y(t0_011111000100));
wire t0_0111110001000, t0_0111110001001;
mixer mix_t0_011111000101 (.a(t0_0111110001010), .b(t0_0111110001011), .y(t0_011111000101));
wire t0_0111110001010, t0_0111110001011;
mixer mix_t0_01111100011 (.a(t0_011111000110), .b(t0_011111000111), .y(t0_01111100011));
wire t0_011111000110, t0_011111000111;
mixer mix_t0_011111000110 (.a(t0_0111110001100), .b(t0_0111110001101), .y(t0_011111000110));
wire t0_0111110001100, t0_0111110001101;
mixer mix_t0_011111000111 (.a(t0_0111110001110), .b(t0_0111110001111), .y(t0_011111000111));
wire t0_0111110001110, t0_0111110001111;
mixer mix_t0_011111001 (.a(t0_0111110010), .b(t0_0111110011), .y(t0_011111001));
wire t0_0111110010, t0_0111110011;
mixer mix_t0_0111110010 (.a(t0_01111100100), .b(t0_01111100101), .y(t0_0111110010));
wire t0_01111100100, t0_01111100101;
mixer mix_t0_01111100100 (.a(t0_011111001000), .b(t0_011111001001), .y(t0_01111100100));
wire t0_011111001000, t0_011111001001;
mixer mix_t0_011111001000 (.a(t0_0111110010000), .b(t0_0111110010001), .y(t0_011111001000));
wire t0_0111110010000, t0_0111110010001;
mixer mix_t0_011111001001 (.a(t0_0111110010010), .b(t0_0111110010011), .y(t0_011111001001));
wire t0_0111110010010, t0_0111110010011;
mixer mix_t0_01111100101 (.a(t0_011111001010), .b(t0_011111001011), .y(t0_01111100101));
wire t0_011111001010, t0_011111001011;
mixer mix_t0_011111001010 (.a(t0_0111110010100), .b(t0_0111110010101), .y(t0_011111001010));
wire t0_0111110010100, t0_0111110010101;
mixer mix_t0_011111001011 (.a(t0_0111110010110), .b(t0_0111110010111), .y(t0_011111001011));
wire t0_0111110010110, t0_0111110010111;
mixer mix_t0_0111110011 (.a(t0_01111100110), .b(t0_01111100111), .y(t0_0111110011));
wire t0_01111100110, t0_01111100111;
mixer mix_t0_01111100110 (.a(t0_011111001100), .b(t0_011111001101), .y(t0_01111100110));
wire t0_011111001100, t0_011111001101;
mixer mix_t0_011111001100 (.a(t0_0111110011000), .b(t0_0111110011001), .y(t0_011111001100));
wire t0_0111110011000, t0_0111110011001;
mixer mix_t0_011111001101 (.a(t0_0111110011010), .b(t0_0111110011011), .y(t0_011111001101));
wire t0_0111110011010, t0_0111110011011;
mixer mix_t0_01111100111 (.a(t0_011111001110), .b(t0_011111001111), .y(t0_01111100111));
wire t0_011111001110, t0_011111001111;
mixer mix_t0_011111001110 (.a(t0_0111110011100), .b(t0_0111110011101), .y(t0_011111001110));
wire t0_0111110011100, t0_0111110011101;
mixer mix_t0_011111001111 (.a(t0_0111110011110), .b(t0_0111110011111), .y(t0_011111001111));
wire t0_0111110011110, t0_0111110011111;
mixer mix_t0_01111101 (.a(t0_011111010), .b(t0_011111011), .y(t0_01111101));
wire t0_011111010, t0_011111011;
mixer mix_t0_011111010 (.a(t0_0111110100), .b(t0_0111110101), .y(t0_011111010));
wire t0_0111110100, t0_0111110101;
mixer mix_t0_0111110100 (.a(t0_01111101000), .b(t0_01111101001), .y(t0_0111110100));
wire t0_01111101000, t0_01111101001;
mixer mix_t0_01111101000 (.a(t0_011111010000), .b(t0_011111010001), .y(t0_01111101000));
wire t0_011111010000, t0_011111010001;
mixer mix_t0_011111010000 (.a(t0_0111110100000), .b(t0_0111110100001), .y(t0_011111010000));
wire t0_0111110100000, t0_0111110100001;
mixer mix_t0_011111010001 (.a(t0_0111110100010), .b(t0_0111110100011), .y(t0_011111010001));
wire t0_0111110100010, t0_0111110100011;
mixer mix_t0_01111101001 (.a(t0_011111010010), .b(t0_011111010011), .y(t0_01111101001));
wire t0_011111010010, t0_011111010011;
mixer mix_t0_011111010010 (.a(t0_0111110100100), .b(t0_0111110100101), .y(t0_011111010010));
wire t0_0111110100100, t0_0111110100101;
mixer mix_t0_011111010011 (.a(t0_0111110100110), .b(t0_0111110100111), .y(t0_011111010011));
wire t0_0111110100110, t0_0111110100111;
mixer mix_t0_0111110101 (.a(t0_01111101010), .b(t0_01111101011), .y(t0_0111110101));
wire t0_01111101010, t0_01111101011;
mixer mix_t0_01111101010 (.a(t0_011111010100), .b(t0_011111010101), .y(t0_01111101010));
wire t0_011111010100, t0_011111010101;
mixer mix_t0_011111010100 (.a(t0_0111110101000), .b(t0_0111110101001), .y(t0_011111010100));
wire t0_0111110101000, t0_0111110101001;
mixer mix_t0_011111010101 (.a(t0_0111110101010), .b(t0_0111110101011), .y(t0_011111010101));
wire t0_0111110101010, t0_0111110101011;
mixer mix_t0_01111101011 (.a(t0_011111010110), .b(t0_011111010111), .y(t0_01111101011));
wire t0_011111010110, t0_011111010111;
mixer mix_t0_011111010110 (.a(t0_0111110101100), .b(t0_0111110101101), .y(t0_011111010110));
wire t0_0111110101100, t0_0111110101101;
mixer mix_t0_011111010111 (.a(t0_0111110101110), .b(t0_0111110101111), .y(t0_011111010111));
wire t0_0111110101110, t0_0111110101111;
mixer mix_t0_011111011 (.a(t0_0111110110), .b(t0_0111110111), .y(t0_011111011));
wire t0_0111110110, t0_0111110111;
mixer mix_t0_0111110110 (.a(t0_01111101100), .b(t0_01111101101), .y(t0_0111110110));
wire t0_01111101100, t0_01111101101;
mixer mix_t0_01111101100 (.a(t0_011111011000), .b(t0_011111011001), .y(t0_01111101100));
wire t0_011111011000, t0_011111011001;
mixer mix_t0_011111011000 (.a(t0_0111110110000), .b(t0_0111110110001), .y(t0_011111011000));
wire t0_0111110110000, t0_0111110110001;
mixer mix_t0_011111011001 (.a(t0_0111110110010), .b(t0_0111110110011), .y(t0_011111011001));
wire t0_0111110110010, t0_0111110110011;
mixer mix_t0_01111101101 (.a(t0_011111011010), .b(t0_011111011011), .y(t0_01111101101));
wire t0_011111011010, t0_011111011011;
mixer mix_t0_011111011010 (.a(t0_0111110110100), .b(t0_0111110110101), .y(t0_011111011010));
wire t0_0111110110100, t0_0111110110101;
mixer mix_t0_011111011011 (.a(t0_0111110110110), .b(t0_0111110110111), .y(t0_011111011011));
wire t0_0111110110110, t0_0111110110111;
mixer mix_t0_0111110111 (.a(t0_01111101110), .b(t0_01111101111), .y(t0_0111110111));
wire t0_01111101110, t0_01111101111;
mixer mix_t0_01111101110 (.a(t0_011111011100), .b(t0_011111011101), .y(t0_01111101110));
wire t0_011111011100, t0_011111011101;
mixer mix_t0_011111011100 (.a(t0_0111110111000), .b(t0_0111110111001), .y(t0_011111011100));
wire t0_0111110111000, t0_0111110111001;
mixer mix_t0_011111011101 (.a(t0_0111110111010), .b(t0_0111110111011), .y(t0_011111011101));
wire t0_0111110111010, t0_0111110111011;
mixer mix_t0_01111101111 (.a(t0_011111011110), .b(t0_011111011111), .y(t0_01111101111));
wire t0_011111011110, t0_011111011111;
mixer mix_t0_011111011110 (.a(t0_0111110111100), .b(t0_0111110111101), .y(t0_011111011110));
wire t0_0111110111100, t0_0111110111101;
mixer mix_t0_011111011111 (.a(t0_0111110111110), .b(t0_0111110111111), .y(t0_011111011111));
wire t0_0111110111110, t0_0111110111111;
mixer mix_t0_0111111 (.a(t0_01111110), .b(t0_01111111), .y(t0_0111111));
wire t0_01111110, t0_01111111;
mixer mix_t0_01111110 (.a(t0_011111100), .b(t0_011111101), .y(t0_01111110));
wire t0_011111100, t0_011111101;
mixer mix_t0_011111100 (.a(t0_0111111000), .b(t0_0111111001), .y(t0_011111100));
wire t0_0111111000, t0_0111111001;
mixer mix_t0_0111111000 (.a(t0_01111110000), .b(t0_01111110001), .y(t0_0111111000));
wire t0_01111110000, t0_01111110001;
mixer mix_t0_01111110000 (.a(t0_011111100000), .b(t0_011111100001), .y(t0_01111110000));
wire t0_011111100000, t0_011111100001;
mixer mix_t0_011111100000 (.a(t0_0111111000000), .b(t0_0111111000001), .y(t0_011111100000));
wire t0_0111111000000, t0_0111111000001;
mixer mix_t0_011111100001 (.a(t0_0111111000010), .b(t0_0111111000011), .y(t0_011111100001));
wire t0_0111111000010, t0_0111111000011;
mixer mix_t0_01111110001 (.a(t0_011111100010), .b(t0_011111100011), .y(t0_01111110001));
wire t0_011111100010, t0_011111100011;
mixer mix_t0_011111100010 (.a(t0_0111111000100), .b(t0_0111111000101), .y(t0_011111100010));
wire t0_0111111000100, t0_0111111000101;
mixer mix_t0_011111100011 (.a(t0_0111111000110), .b(t0_0111111000111), .y(t0_011111100011));
wire t0_0111111000110, t0_0111111000111;
mixer mix_t0_0111111001 (.a(t0_01111110010), .b(t0_01111110011), .y(t0_0111111001));
wire t0_01111110010, t0_01111110011;
mixer mix_t0_01111110010 (.a(t0_011111100100), .b(t0_011111100101), .y(t0_01111110010));
wire t0_011111100100, t0_011111100101;
mixer mix_t0_011111100100 (.a(t0_0111111001000), .b(t0_0111111001001), .y(t0_011111100100));
wire t0_0111111001000, t0_0111111001001;
mixer mix_t0_011111100101 (.a(t0_0111111001010), .b(t0_0111111001011), .y(t0_011111100101));
wire t0_0111111001010, t0_0111111001011;
mixer mix_t0_01111110011 (.a(t0_011111100110), .b(t0_011111100111), .y(t0_01111110011));
wire t0_011111100110, t0_011111100111;
mixer mix_t0_011111100110 (.a(t0_0111111001100), .b(t0_0111111001101), .y(t0_011111100110));
wire t0_0111111001100, t0_0111111001101;
mixer mix_t0_011111100111 (.a(t0_0111111001110), .b(t0_0111111001111), .y(t0_011111100111));
wire t0_0111111001110, t0_0111111001111;
mixer mix_t0_011111101 (.a(t0_0111111010), .b(t0_0111111011), .y(t0_011111101));
wire t0_0111111010, t0_0111111011;
mixer mix_t0_0111111010 (.a(t0_01111110100), .b(t0_01111110101), .y(t0_0111111010));
wire t0_01111110100, t0_01111110101;
mixer mix_t0_01111110100 (.a(t0_011111101000), .b(t0_011111101001), .y(t0_01111110100));
wire t0_011111101000, t0_011111101001;
mixer mix_t0_011111101000 (.a(t0_0111111010000), .b(t0_0111111010001), .y(t0_011111101000));
wire t0_0111111010000, t0_0111111010001;
mixer mix_t0_011111101001 (.a(t0_0111111010010), .b(t0_0111111010011), .y(t0_011111101001));
wire t0_0111111010010, t0_0111111010011;
mixer mix_t0_01111110101 (.a(t0_011111101010), .b(t0_011111101011), .y(t0_01111110101));
wire t0_011111101010, t0_011111101011;
mixer mix_t0_011111101010 (.a(t0_0111111010100), .b(t0_0111111010101), .y(t0_011111101010));
wire t0_0111111010100, t0_0111111010101;
mixer mix_t0_011111101011 (.a(t0_0111111010110), .b(t0_0111111010111), .y(t0_011111101011));
wire t0_0111111010110, t0_0111111010111;
mixer mix_t0_0111111011 (.a(t0_01111110110), .b(t0_01111110111), .y(t0_0111111011));
wire t0_01111110110, t0_01111110111;
mixer mix_t0_01111110110 (.a(t0_011111101100), .b(t0_011111101101), .y(t0_01111110110));
wire t0_011111101100, t0_011111101101;
mixer mix_t0_011111101100 (.a(t0_0111111011000), .b(t0_0111111011001), .y(t0_011111101100));
wire t0_0111111011000, t0_0111111011001;
mixer mix_t0_011111101101 (.a(t0_0111111011010), .b(t0_0111111011011), .y(t0_011111101101));
wire t0_0111111011010, t0_0111111011011;
mixer mix_t0_01111110111 (.a(t0_011111101110), .b(t0_011111101111), .y(t0_01111110111));
wire t0_011111101110, t0_011111101111;
mixer mix_t0_011111101110 (.a(t0_0111111011100), .b(t0_0111111011101), .y(t0_011111101110));
wire t0_0111111011100, t0_0111111011101;
mixer mix_t0_011111101111 (.a(t0_0111111011110), .b(t0_0111111011111), .y(t0_011111101111));
wire t0_0111111011110, t0_0111111011111;
mixer mix_t0_01111111 (.a(t0_011111110), .b(t0_011111111), .y(t0_01111111));
wire t0_011111110, t0_011111111;
mixer mix_t0_011111110 (.a(t0_0111111100), .b(t0_0111111101), .y(t0_011111110));
wire t0_0111111100, t0_0111111101;
mixer mix_t0_0111111100 (.a(t0_01111111000), .b(t0_01111111001), .y(t0_0111111100));
wire t0_01111111000, t0_01111111001;
mixer mix_t0_01111111000 (.a(t0_011111110000), .b(t0_011111110001), .y(t0_01111111000));
wire t0_011111110000, t0_011111110001;
mixer mix_t0_011111110000 (.a(t0_0111111100000), .b(t0_0111111100001), .y(t0_011111110000));
wire t0_0111111100000, t0_0111111100001;
mixer mix_t0_011111110001 (.a(t0_0111111100010), .b(t0_0111111100011), .y(t0_011111110001));
wire t0_0111111100010, t0_0111111100011;
mixer mix_t0_01111111001 (.a(t0_011111110010), .b(t0_011111110011), .y(t0_01111111001));
wire t0_011111110010, t0_011111110011;
mixer mix_t0_011111110010 (.a(t0_0111111100100), .b(t0_0111111100101), .y(t0_011111110010));
wire t0_0111111100100, t0_0111111100101;
mixer mix_t0_011111110011 (.a(t0_0111111100110), .b(t0_0111111100111), .y(t0_011111110011));
wire t0_0111111100110, t0_0111111100111;
mixer mix_t0_0111111101 (.a(t0_01111111010), .b(t0_01111111011), .y(t0_0111111101));
wire t0_01111111010, t0_01111111011;
mixer mix_t0_01111111010 (.a(t0_011111110100), .b(t0_011111110101), .y(t0_01111111010));
wire t0_011111110100, t0_011111110101;
mixer mix_t0_011111110100 (.a(t0_0111111101000), .b(t0_0111111101001), .y(t0_011111110100));
wire t0_0111111101000, t0_0111111101001;
mixer mix_t0_011111110101 (.a(t0_0111111101010), .b(t0_0111111101011), .y(t0_011111110101));
wire t0_0111111101010, t0_0111111101011;
mixer mix_t0_01111111011 (.a(t0_011111110110), .b(t0_011111110111), .y(t0_01111111011));
wire t0_011111110110, t0_011111110111;
mixer mix_t0_011111110110 (.a(t0_0111111101100), .b(t0_0111111101101), .y(t0_011111110110));
wire t0_0111111101100, t0_0111111101101;
mixer mix_t0_011111110111 (.a(t0_0111111101110), .b(t0_0111111101111), .y(t0_011111110111));
wire t0_0111111101110, t0_0111111101111;
mixer mix_t0_011111111 (.a(t0_0111111110), .b(t0_0111111111), .y(t0_011111111));
wire t0_0111111110, t0_0111111111;
mixer mix_t0_0111111110 (.a(t0_01111111100), .b(t0_01111111101), .y(t0_0111111110));
wire t0_01111111100, t0_01111111101;
mixer mix_t0_01111111100 (.a(t0_011111111000), .b(t0_011111111001), .y(t0_01111111100));
wire t0_011111111000, t0_011111111001;
mixer mix_t0_011111111000 (.a(t0_0111111110000), .b(t0_0111111110001), .y(t0_011111111000));
wire t0_0111111110000, t0_0111111110001;
mixer mix_t0_011111111001 (.a(t0_0111111110010), .b(t0_0111111110011), .y(t0_011111111001));
wire t0_0111111110010, t0_0111111110011;
mixer mix_t0_01111111101 (.a(t0_011111111010), .b(t0_011111111011), .y(t0_01111111101));
wire t0_011111111010, t0_011111111011;
mixer mix_t0_011111111010 (.a(t0_0111111110100), .b(t0_0111111110101), .y(t0_011111111010));
wire t0_0111111110100, t0_0111111110101;
mixer mix_t0_011111111011 (.a(t0_0111111110110), .b(t0_0111111110111), .y(t0_011111111011));
wire t0_0111111110110, t0_0111111110111;
mixer mix_t0_0111111111 (.a(t0_01111111110), .b(t0_01111111111), .y(t0_0111111111));
wire t0_01111111110, t0_01111111111;
mixer mix_t0_01111111110 (.a(t0_011111111100), .b(t0_011111111101), .y(t0_01111111110));
wire t0_011111111100, t0_011111111101;
mixer mix_t0_011111111100 (.a(t0_0111111111000), .b(t0_0111111111001), .y(t0_011111111100));
wire t0_0111111111000, t0_0111111111001;
mixer mix_t0_011111111101 (.a(t0_0111111111010), .b(t0_0111111111011), .y(t0_011111111101));
wire t0_0111111111010, t0_0111111111011;
mixer mix_t0_01111111111 (.a(t0_011111111110), .b(t0_011111111111), .y(t0_01111111111));
wire t0_011111111110, t0_011111111111;
mixer mix_t0_011111111110 (.a(t0_0111111111100), .b(t0_0111111111101), .y(t0_011111111110));
wire t0_0111111111100, t0_0111111111101;
mixer mix_t0_011111111111 (.a(t0_0111111111110), .b(t0_0111111111111), .y(t0_011111111111));
wire t0_0111111111110, t0_0111111111111;
wire t0_0;
assign out_0 = t0_0;
assign input_0 = t0_0000000000000;
assign input_1 = t0_0000000000001;
assign input_2 = t0_0000000000010;
assign input_3 = t0_0000000000011;
assign input_4 = t0_0000000000100;
assign input_5 = t0_0000000000101;
assign input_6 = t0_0000000000110;
assign input_7 = t0_0000000000111;
assign input_8 = t0_0000000001000;
assign input_9 = t0_0000000001001;
assign input_10 = t0_0000000001010;
assign input_11 = t0_0000000001011;
assign input_12 = t0_0000000001100;
assign input_13 = t0_0000000001101;
assign input_14 = t0_0000000001110;
assign input_15 = t0_0000000001111;
assign input_16 = t0_0000000010000;
assign input_17 = t0_0000000010001;
assign input_18 = t0_0000000010010;
assign input_19 = t0_0000000010011;
assign input_20 = t0_0000000010100;
assign input_21 = t0_0000000010101;
assign input_22 = t0_0000000010110;
assign input_23 = t0_0000000010111;
assign input_24 = t0_0000000011000;
assign input_25 = t0_0000000011001;
assign input_26 = t0_0000000011010;
assign input_27 = t0_0000000011011;
assign input_28 = t0_0000000011100;
assign input_29 = t0_0000000011101;
assign input_30 = t0_0000000011110;
assign input_31 = t0_0000000011111;
assign input_32 = t0_0000000100000;
assign input_33 = t0_0000000100001;
assign input_34 = t0_0000000100010;
assign input_35 = t0_0000000100011;
assign input_36 = t0_0000000100100;
assign input_37 = t0_0000000100101;
assign input_38 = t0_0000000100110;
assign input_39 = t0_0000000100111;
assign input_40 = t0_0000000101000;
assign input_41 = t0_0000000101001;
assign input_42 = t0_0000000101010;
assign input_43 = t0_0000000101011;
assign input_44 = t0_0000000101100;
assign input_45 = t0_0000000101101;
assign input_46 = t0_0000000101110;
assign input_47 = t0_0000000101111;
assign input_48 = t0_0000000110000;
assign input_49 = t0_0000000110001;
assign input_50 = t0_0000000110010;
assign input_51 = t0_0000000110011;
assign input_52 = t0_0000000110100;
assign input_53 = t0_0000000110101;
assign input_54 = t0_0000000110110;
assign input_55 = t0_0000000110111;
assign input_56 = t0_0000000111000;
assign input_57 = t0_0000000111001;
assign input_58 = t0_0000000111010;
assign input_59 = t0_0000000111011;
assign input_60 = t0_0000000111100;
assign input_61 = t0_0000000111101;
assign input_62 = t0_0000000111110;
assign input_63 = t0_0000000111111;
assign input_64 = t0_0000001000000;
assign input_65 = t0_0000001000001;
assign input_66 = t0_0000001000010;
assign input_67 = t0_0000001000011;
assign input_68 = t0_0000001000100;
assign input_69 = t0_0000001000101;
assign input_70 = t0_0000001000110;
assign input_71 = t0_0000001000111;
assign input_72 = t0_0000001001000;
assign input_73 = t0_0000001001001;
assign input_74 = t0_0000001001010;
assign input_75 = t0_0000001001011;
assign input_76 = t0_0000001001100;
assign input_77 = t0_0000001001101;
assign input_78 = t0_0000001001110;
assign input_79 = t0_0000001001111;
assign input_80 = t0_0000001010000;
assign input_81 = t0_0000001010001;
assign input_82 = t0_0000001010010;
assign input_83 = t0_0000001010011;
assign input_84 = t0_0000001010100;
assign input_85 = t0_0000001010101;
assign input_86 = t0_0000001010110;
assign input_87 = t0_0000001010111;
assign input_88 = t0_0000001011000;
assign input_89 = t0_0000001011001;
assign input_90 = t0_0000001011010;
assign input_91 = t0_0000001011011;
assign input_92 = t0_0000001011100;
assign input_93 = t0_0000001011101;
assign input_94 = t0_0000001011110;
assign input_95 = t0_0000001011111;
assign input_96 = t0_0000001100000;
assign input_97 = t0_0000001100001;
assign input_98 = t0_0000001100010;
assign input_99 = t0_0000001100011;
assign input_100 = t0_0000001100100;
assign input_101 = t0_0000001100101;
assign input_102 = t0_0000001100110;
assign input_103 = t0_0000001100111;
assign input_104 = t0_0000001101000;
assign input_105 = t0_0000001101001;
assign input_106 = t0_0000001101010;
assign input_107 = t0_0000001101011;
assign input_108 = t0_0000001101100;
assign input_109 = t0_0000001101101;
assign input_110 = t0_0000001101110;
assign input_111 = t0_0000001101111;
assign input_112 = t0_0000001110000;
assign input_113 = t0_0000001110001;
assign input_114 = t0_0000001110010;
assign input_115 = t0_0000001110011;
assign input_116 = t0_0000001110100;
assign input_117 = t0_0000001110101;
assign input_118 = t0_0000001110110;
assign input_119 = t0_0000001110111;
assign input_120 = t0_0000001111000;
assign input_121 = t0_0000001111001;
assign input_122 = t0_0000001111010;
assign input_123 = t0_0000001111011;
assign input_124 = t0_0000001111100;
assign input_125 = t0_0000001111101;
assign input_126 = t0_0000001111110;
assign input_127 = t0_0000001111111;
assign input_128 = t0_0000010000000;
assign input_129 = t0_0000010000001;
assign input_130 = t0_0000010000010;
assign input_131 = t0_0000010000011;
assign input_132 = t0_0000010000100;
assign input_133 = t0_0000010000101;
assign input_134 = t0_0000010000110;
assign input_135 = t0_0000010000111;
assign input_136 = t0_0000010001000;
assign input_137 = t0_0000010001001;
assign input_138 = t0_0000010001010;
assign input_139 = t0_0000010001011;
assign input_140 = t0_0000010001100;
assign input_141 = t0_0000010001101;
assign input_142 = t0_0000010001110;
assign input_143 = t0_0000010001111;
assign input_144 = t0_0000010010000;
assign input_145 = t0_0000010010001;
assign input_146 = t0_0000010010010;
assign input_147 = t0_0000010010011;
assign input_148 = t0_0000010010100;
assign input_149 = t0_0000010010101;
assign input_150 = t0_0000010010110;
assign input_151 = t0_0000010010111;
assign input_152 = t0_0000010011000;
assign input_153 = t0_0000010011001;
assign input_154 = t0_0000010011010;
assign input_155 = t0_0000010011011;
assign input_156 = t0_0000010011100;
assign input_157 = t0_0000010011101;
assign input_158 = t0_0000010011110;
assign input_159 = t0_0000010011111;
assign input_160 = t0_0000010100000;
assign input_161 = t0_0000010100001;
assign input_162 = t0_0000010100010;
assign input_163 = t0_0000010100011;
assign input_164 = t0_0000010100100;
assign input_165 = t0_0000010100101;
assign input_166 = t0_0000010100110;
assign input_167 = t0_0000010100111;
assign input_168 = t0_0000010101000;
assign input_169 = t0_0000010101001;
assign input_170 = t0_0000010101010;
assign input_171 = t0_0000010101011;
assign input_172 = t0_0000010101100;
assign input_173 = t0_0000010101101;
assign input_174 = t0_0000010101110;
assign input_175 = t0_0000010101111;
assign input_176 = t0_0000010110000;
assign input_177 = t0_0000010110001;
assign input_178 = t0_0000010110010;
assign input_179 = t0_0000010110011;
assign input_180 = t0_0000010110100;
assign input_181 = t0_0000010110101;
assign input_182 = t0_0000010110110;
assign input_183 = t0_0000010110111;
assign input_184 = t0_0000010111000;
assign input_185 = t0_0000010111001;
assign input_186 = t0_0000010111010;
assign input_187 = t0_0000010111011;
assign input_188 = t0_0000010111100;
assign input_189 = t0_0000010111101;
assign input_190 = t0_0000010111110;
assign input_191 = t0_0000010111111;
assign input_192 = t0_0000011000000;
assign input_193 = t0_0000011000001;
assign input_194 = t0_0000011000010;
assign input_195 = t0_0000011000011;
assign input_196 = t0_0000011000100;
assign input_197 = t0_0000011000101;
assign input_198 = t0_0000011000110;
assign input_199 = t0_0000011000111;
assign input_200 = t0_0000011001000;
assign input_201 = t0_0000011001001;
assign input_202 = t0_0000011001010;
assign input_203 = t0_0000011001011;
assign input_204 = t0_0000011001100;
assign input_205 = t0_0000011001101;
assign input_206 = t0_0000011001110;
assign input_207 = t0_0000011001111;
assign input_208 = t0_0000011010000;
assign input_209 = t0_0000011010001;
assign input_210 = t0_0000011010010;
assign input_211 = t0_0000011010011;
assign input_212 = t0_0000011010100;
assign input_213 = t0_0000011010101;
assign input_214 = t0_0000011010110;
assign input_215 = t0_0000011010111;
assign input_216 = t0_0000011011000;
assign input_217 = t0_0000011011001;
assign input_218 = t0_0000011011010;
assign input_219 = t0_0000011011011;
assign input_220 = t0_0000011011100;
assign input_221 = t0_0000011011101;
assign input_222 = t0_0000011011110;
assign input_223 = t0_0000011011111;
assign input_224 = t0_0000011100000;
assign input_225 = t0_0000011100001;
assign input_226 = t0_0000011100010;
assign input_227 = t0_0000011100011;
assign input_228 = t0_0000011100100;
assign input_229 = t0_0000011100101;
assign input_230 = t0_0000011100110;
assign input_231 = t0_0000011100111;
assign input_232 = t0_0000011101000;
assign input_233 = t0_0000011101001;
assign input_234 = t0_0000011101010;
assign input_235 = t0_0000011101011;
assign input_236 = t0_0000011101100;
assign input_237 = t0_0000011101101;
assign input_238 = t0_0000011101110;
assign input_239 = t0_0000011101111;
assign input_240 = t0_0000011110000;
assign input_241 = t0_0000011110001;
assign input_242 = t0_0000011110010;
assign input_243 = t0_0000011110011;
assign input_244 = t0_0000011110100;
assign input_245 = t0_0000011110101;
assign input_246 = t0_0000011110110;
assign input_247 = t0_0000011110111;
assign input_248 = t0_0000011111000;
assign input_249 = t0_0000011111001;
assign input_250 = t0_0000011111010;
assign input_251 = t0_0000011111011;
assign input_252 = t0_0000011111100;
assign input_253 = t0_0000011111101;
assign input_254 = t0_0000011111110;
assign input_255 = t0_0000011111111;
assign input_256 = t0_0000100000000;
assign input_257 = t0_0000100000001;
assign input_258 = t0_0000100000010;
assign input_259 = t0_0000100000011;
assign input_260 = t0_0000100000100;
assign input_261 = t0_0000100000101;
assign input_262 = t0_0000100000110;
assign input_263 = t0_0000100000111;
assign input_264 = t0_0000100001000;
assign input_265 = t0_0000100001001;
assign input_266 = t0_0000100001010;
assign input_267 = t0_0000100001011;
assign input_268 = t0_0000100001100;
assign input_269 = t0_0000100001101;
assign input_270 = t0_0000100001110;
assign input_271 = t0_0000100001111;
assign input_272 = t0_0000100010000;
assign input_273 = t0_0000100010001;
assign input_274 = t0_0000100010010;
assign input_275 = t0_0000100010011;
assign input_276 = t0_0000100010100;
assign input_277 = t0_0000100010101;
assign input_278 = t0_0000100010110;
assign input_279 = t0_0000100010111;
assign input_280 = t0_0000100011000;
assign input_281 = t0_0000100011001;
assign input_282 = t0_0000100011010;
assign input_283 = t0_0000100011011;
assign input_284 = t0_0000100011100;
assign input_285 = t0_0000100011101;
assign input_286 = t0_0000100011110;
assign input_287 = t0_0000100011111;
assign input_288 = t0_0000100100000;
assign input_289 = t0_0000100100001;
assign input_290 = t0_0000100100010;
assign input_291 = t0_0000100100011;
assign input_292 = t0_0000100100100;
assign input_293 = t0_0000100100101;
assign input_294 = t0_0000100100110;
assign input_295 = t0_0000100100111;
assign input_296 = t0_0000100101000;
assign input_297 = t0_0000100101001;
assign input_298 = t0_0000100101010;
assign input_299 = t0_0000100101011;
assign input_300 = t0_0000100101100;
assign input_301 = t0_0000100101101;
assign input_302 = t0_0000100101110;
assign input_303 = t0_0000100101111;
assign input_304 = t0_0000100110000;
assign input_305 = t0_0000100110001;
assign input_306 = t0_0000100110010;
assign input_307 = t0_0000100110011;
assign input_308 = t0_0000100110100;
assign input_309 = t0_0000100110101;
assign input_310 = t0_0000100110110;
assign input_311 = t0_0000100110111;
assign input_312 = t0_0000100111000;
assign input_313 = t0_0000100111001;
assign input_314 = t0_0000100111010;
assign input_315 = t0_0000100111011;
assign input_316 = t0_0000100111100;
assign input_317 = t0_0000100111101;
assign input_318 = t0_0000100111110;
assign input_319 = t0_0000100111111;
assign input_320 = t0_0000101000000;
assign input_321 = t0_0000101000001;
assign input_322 = t0_0000101000010;
assign input_323 = t0_0000101000011;
assign input_324 = t0_0000101000100;
assign input_325 = t0_0000101000101;
assign input_326 = t0_0000101000110;
assign input_327 = t0_0000101000111;
assign input_328 = t0_0000101001000;
assign input_329 = t0_0000101001001;
assign input_330 = t0_0000101001010;
assign input_331 = t0_0000101001011;
assign input_332 = t0_0000101001100;
assign input_333 = t0_0000101001101;
assign input_334 = t0_0000101001110;
assign input_335 = t0_0000101001111;
assign input_336 = t0_0000101010000;
assign input_337 = t0_0000101010001;
assign input_338 = t0_0000101010010;
assign input_339 = t0_0000101010011;
assign input_340 = t0_0000101010100;
assign input_341 = t0_0000101010101;
assign input_342 = t0_0000101010110;
assign input_343 = t0_0000101010111;
assign input_344 = t0_0000101011000;
assign input_345 = t0_0000101011001;
assign input_346 = t0_0000101011010;
assign input_347 = t0_0000101011011;
assign input_348 = t0_0000101011100;
assign input_349 = t0_0000101011101;
assign input_350 = t0_0000101011110;
assign input_351 = t0_0000101011111;
assign input_352 = t0_0000101100000;
assign input_353 = t0_0000101100001;
assign input_354 = t0_0000101100010;
assign input_355 = t0_0000101100011;
assign input_356 = t0_0000101100100;
assign input_357 = t0_0000101100101;
assign input_358 = t0_0000101100110;
assign input_359 = t0_0000101100111;
assign input_360 = t0_0000101101000;
assign input_361 = t0_0000101101001;
assign input_362 = t0_0000101101010;
assign input_363 = t0_0000101101011;
assign input_364 = t0_0000101101100;
assign input_365 = t0_0000101101101;
assign input_366 = t0_0000101101110;
assign input_367 = t0_0000101101111;
assign input_368 = t0_0000101110000;
assign input_369 = t0_0000101110001;
assign input_370 = t0_0000101110010;
assign input_371 = t0_0000101110011;
assign input_372 = t0_0000101110100;
assign input_373 = t0_0000101110101;
assign input_374 = t0_0000101110110;
assign input_375 = t0_0000101110111;
assign input_376 = t0_0000101111000;
assign input_377 = t0_0000101111001;
assign input_378 = t0_0000101111010;
assign input_379 = t0_0000101111011;
assign input_380 = t0_0000101111100;
assign input_381 = t0_0000101111101;
assign input_382 = t0_0000101111110;
assign input_383 = t0_0000101111111;
assign input_384 = t0_0000110000000;
assign input_385 = t0_0000110000001;
assign input_386 = t0_0000110000010;
assign input_387 = t0_0000110000011;
assign input_388 = t0_0000110000100;
assign input_389 = t0_0000110000101;
assign input_390 = t0_0000110000110;
assign input_391 = t0_0000110000111;
assign input_392 = t0_0000110001000;
assign input_393 = t0_0000110001001;
assign input_394 = t0_0000110001010;
assign input_395 = t0_0000110001011;
assign input_396 = t0_0000110001100;
assign input_397 = t0_0000110001101;
assign input_398 = t0_0000110001110;
assign input_399 = t0_0000110001111;
assign input_400 = t0_0000110010000;
assign input_401 = t0_0000110010001;
assign input_402 = t0_0000110010010;
assign input_403 = t0_0000110010011;
assign input_404 = t0_0000110010100;
assign input_405 = t0_0000110010101;
assign input_406 = t0_0000110010110;
assign input_407 = t0_0000110010111;
assign input_408 = t0_0000110011000;
assign input_409 = t0_0000110011001;
assign input_410 = t0_0000110011010;
assign input_411 = t0_0000110011011;
assign input_412 = t0_0000110011100;
assign input_413 = t0_0000110011101;
assign input_414 = t0_0000110011110;
assign input_415 = t0_0000110011111;
assign input_416 = t0_0000110100000;
assign input_417 = t0_0000110100001;
assign input_418 = t0_0000110100010;
assign input_419 = t0_0000110100011;
assign input_420 = t0_0000110100100;
assign input_421 = t0_0000110100101;
assign input_422 = t0_0000110100110;
assign input_423 = t0_0000110100111;
assign input_424 = t0_0000110101000;
assign input_425 = t0_0000110101001;
assign input_426 = t0_0000110101010;
assign input_427 = t0_0000110101011;
assign input_428 = t0_0000110101100;
assign input_429 = t0_0000110101101;
assign input_430 = t0_0000110101110;
assign input_431 = t0_0000110101111;
assign input_432 = t0_0000110110000;
assign input_433 = t0_0000110110001;
assign input_434 = t0_0000110110010;
assign input_435 = t0_0000110110011;
assign input_436 = t0_0000110110100;
assign input_437 = t0_0000110110101;
assign input_438 = t0_0000110110110;
assign input_439 = t0_0000110110111;
assign input_440 = t0_0000110111000;
assign input_441 = t0_0000110111001;
assign input_442 = t0_0000110111010;
assign input_443 = t0_0000110111011;
assign input_444 = t0_0000110111100;
assign input_445 = t0_0000110111101;
assign input_446 = t0_0000110111110;
assign input_447 = t0_0000110111111;
assign input_448 = t0_0000111000000;
assign input_449 = t0_0000111000001;
assign input_450 = t0_0000111000010;
assign input_451 = t0_0000111000011;
assign input_452 = t0_0000111000100;
assign input_453 = t0_0000111000101;
assign input_454 = t0_0000111000110;
assign input_455 = t0_0000111000111;
assign input_456 = t0_0000111001000;
assign input_457 = t0_0000111001001;
assign input_458 = t0_0000111001010;
assign input_459 = t0_0000111001011;
assign input_460 = t0_0000111001100;
assign input_461 = t0_0000111001101;
assign input_462 = t0_0000111001110;
assign input_463 = t0_0000111001111;
assign input_464 = t0_0000111010000;
assign input_465 = t0_0000111010001;
assign input_466 = t0_0000111010010;
assign input_467 = t0_0000111010011;
assign input_468 = t0_0000111010100;
assign input_469 = t0_0000111010101;
assign input_470 = t0_0000111010110;
assign input_471 = t0_0000111010111;
assign input_472 = t0_0000111011000;
assign input_473 = t0_0000111011001;
assign input_474 = t0_0000111011010;
assign input_475 = t0_0000111011011;
assign input_476 = t0_0000111011100;
assign input_477 = t0_0000111011101;
assign input_478 = t0_0000111011110;
assign input_479 = t0_0000111011111;
assign input_480 = t0_0000111100000;
assign input_481 = t0_0000111100001;
assign input_482 = t0_0000111100010;
assign input_483 = t0_0000111100011;
assign input_484 = t0_0000111100100;
assign input_485 = t0_0000111100101;
assign input_486 = t0_0000111100110;
assign input_487 = t0_0000111100111;
assign input_488 = t0_0000111101000;
assign input_489 = t0_0000111101001;
assign input_490 = t0_0000111101010;
assign input_491 = t0_0000111101011;
assign input_492 = t0_0000111101100;
assign input_493 = t0_0000111101101;
assign input_494 = t0_0000111101110;
assign input_495 = t0_0000111101111;
assign input_496 = t0_0000111110000;
assign input_497 = t0_0000111110001;
assign input_498 = t0_0000111110010;
assign input_499 = t0_0000111110011;
assign input_500 = t0_0000111110100;
assign input_501 = t0_0000111110101;
assign input_502 = t0_0000111110110;
assign input_503 = t0_0000111110111;
assign input_504 = t0_0000111111000;
assign input_505 = t0_0000111111001;
assign input_506 = t0_0000111111010;
assign input_507 = t0_0000111111011;
assign input_508 = t0_0000111111100;
assign input_509 = t0_0000111111101;
assign input_510 = t0_0000111111110;
assign input_511 = t0_0000111111111;
assign input_512 = t0_0001000000000;
assign input_513 = t0_0001000000001;
assign input_514 = t0_0001000000010;
assign input_515 = t0_0001000000011;
assign input_516 = t0_0001000000100;
assign input_517 = t0_0001000000101;
assign input_518 = t0_0001000000110;
assign input_519 = t0_0001000000111;
assign input_520 = t0_0001000001000;
assign input_521 = t0_0001000001001;
assign input_522 = t0_0001000001010;
assign input_523 = t0_0001000001011;
assign input_524 = t0_0001000001100;
assign input_525 = t0_0001000001101;
assign input_526 = t0_0001000001110;
assign input_527 = t0_0001000001111;
assign input_528 = t0_0001000010000;
assign input_529 = t0_0001000010001;
assign input_530 = t0_0001000010010;
assign input_531 = t0_0001000010011;
assign input_532 = t0_0001000010100;
assign input_533 = t0_0001000010101;
assign input_534 = t0_0001000010110;
assign input_535 = t0_0001000010111;
assign input_536 = t0_0001000011000;
assign input_537 = t0_0001000011001;
assign input_538 = t0_0001000011010;
assign input_539 = t0_0001000011011;
assign input_540 = t0_0001000011100;
assign input_541 = t0_0001000011101;
assign input_542 = t0_0001000011110;
assign input_543 = t0_0001000011111;
assign input_544 = t0_0001000100000;
assign input_545 = t0_0001000100001;
assign input_546 = t0_0001000100010;
assign input_547 = t0_0001000100011;
assign input_548 = t0_0001000100100;
assign input_549 = t0_0001000100101;
assign input_550 = t0_0001000100110;
assign input_551 = t0_0001000100111;
assign input_552 = t0_0001000101000;
assign input_553 = t0_0001000101001;
assign input_554 = t0_0001000101010;
assign input_555 = t0_0001000101011;
assign input_556 = t0_0001000101100;
assign input_557 = t0_0001000101101;
assign input_558 = t0_0001000101110;
assign input_559 = t0_0001000101111;
assign input_560 = t0_0001000110000;
assign input_561 = t0_0001000110001;
assign input_562 = t0_0001000110010;
assign input_563 = t0_0001000110011;
assign input_564 = t0_0001000110100;
assign input_565 = t0_0001000110101;
assign input_566 = t0_0001000110110;
assign input_567 = t0_0001000110111;
assign input_568 = t0_0001000111000;
assign input_569 = t0_0001000111001;
assign input_570 = t0_0001000111010;
assign input_571 = t0_0001000111011;
assign input_572 = t0_0001000111100;
assign input_573 = t0_0001000111101;
assign input_574 = t0_0001000111110;
assign input_575 = t0_0001000111111;
assign input_576 = t0_0001001000000;
assign input_577 = t0_0001001000001;
assign input_578 = t0_0001001000010;
assign input_579 = t0_0001001000011;
assign input_580 = t0_0001001000100;
assign input_581 = t0_0001001000101;
assign input_582 = t0_0001001000110;
assign input_583 = t0_0001001000111;
assign input_584 = t0_0001001001000;
assign input_585 = t0_0001001001001;
assign input_586 = t0_0001001001010;
assign input_587 = t0_0001001001011;
assign input_588 = t0_0001001001100;
assign input_589 = t0_0001001001101;
assign input_590 = t0_0001001001110;
assign input_591 = t0_0001001001111;
assign input_592 = t0_0001001010000;
assign input_593 = t0_0001001010001;
assign input_594 = t0_0001001010010;
assign input_595 = t0_0001001010011;
assign input_596 = t0_0001001010100;
assign input_597 = t0_0001001010101;
assign input_598 = t0_0001001010110;
assign input_599 = t0_0001001010111;
assign input_600 = t0_0001001011000;
assign input_601 = t0_0001001011001;
assign input_602 = t0_0001001011010;
assign input_603 = t0_0001001011011;
assign input_604 = t0_0001001011100;
assign input_605 = t0_0001001011101;
assign input_606 = t0_0001001011110;
assign input_607 = t0_0001001011111;
assign input_608 = t0_0001001100000;
assign input_609 = t0_0001001100001;
assign input_610 = t0_0001001100010;
assign input_611 = t0_0001001100011;
assign input_612 = t0_0001001100100;
assign input_613 = t0_0001001100101;
assign input_614 = t0_0001001100110;
assign input_615 = t0_0001001100111;
assign input_616 = t0_0001001101000;
assign input_617 = t0_0001001101001;
assign input_618 = t0_0001001101010;
assign input_619 = t0_0001001101011;
assign input_620 = t0_0001001101100;
assign input_621 = t0_0001001101101;
assign input_622 = t0_0001001101110;
assign input_623 = t0_0001001101111;
assign input_624 = t0_0001001110000;
assign input_625 = t0_0001001110001;
assign input_626 = t0_0001001110010;
assign input_627 = t0_0001001110011;
assign input_628 = t0_0001001110100;
assign input_629 = t0_0001001110101;
assign input_630 = t0_0001001110110;
assign input_631 = t0_0001001110111;
assign input_632 = t0_0001001111000;
assign input_633 = t0_0001001111001;
assign input_634 = t0_0001001111010;
assign input_635 = t0_0001001111011;
assign input_636 = t0_0001001111100;
assign input_637 = t0_0001001111101;
assign input_638 = t0_0001001111110;
assign input_639 = t0_0001001111111;
assign input_640 = t0_0001010000000;
assign input_641 = t0_0001010000001;
assign input_642 = t0_0001010000010;
assign input_643 = t0_0001010000011;
assign input_644 = t0_0001010000100;
assign input_645 = t0_0001010000101;
assign input_646 = t0_0001010000110;
assign input_647 = t0_0001010000111;
assign input_648 = t0_0001010001000;
assign input_649 = t0_0001010001001;
assign input_650 = t0_0001010001010;
assign input_651 = t0_0001010001011;
assign input_652 = t0_0001010001100;
assign input_653 = t0_0001010001101;
assign input_654 = t0_0001010001110;
assign input_655 = t0_0001010001111;
assign input_656 = t0_0001010010000;
assign input_657 = t0_0001010010001;
assign input_658 = t0_0001010010010;
assign input_659 = t0_0001010010011;
assign input_660 = t0_0001010010100;
assign input_661 = t0_0001010010101;
assign input_662 = t0_0001010010110;
assign input_663 = t0_0001010010111;
assign input_664 = t0_0001010011000;
assign input_665 = t0_0001010011001;
assign input_666 = t0_0001010011010;
assign input_667 = t0_0001010011011;
assign input_668 = t0_0001010011100;
assign input_669 = t0_0001010011101;
assign input_670 = t0_0001010011110;
assign input_671 = t0_0001010011111;
assign input_672 = t0_0001010100000;
assign input_673 = t0_0001010100001;
assign input_674 = t0_0001010100010;
assign input_675 = t0_0001010100011;
assign input_676 = t0_0001010100100;
assign input_677 = t0_0001010100101;
assign input_678 = t0_0001010100110;
assign input_679 = t0_0001010100111;
assign input_680 = t0_0001010101000;
assign input_681 = t0_0001010101001;
assign input_682 = t0_0001010101010;
assign input_683 = t0_0001010101011;
assign input_684 = t0_0001010101100;
assign input_685 = t0_0001010101101;
assign input_686 = t0_0001010101110;
assign input_687 = t0_0001010101111;
assign input_688 = t0_0001010110000;
assign input_689 = t0_0001010110001;
assign input_690 = t0_0001010110010;
assign input_691 = t0_0001010110011;
assign input_692 = t0_0001010110100;
assign input_693 = t0_0001010110101;
assign input_694 = t0_0001010110110;
assign input_695 = t0_0001010110111;
assign input_696 = t0_0001010111000;
assign input_697 = t0_0001010111001;
assign input_698 = t0_0001010111010;
assign input_699 = t0_0001010111011;
assign input_700 = t0_0001010111100;
assign input_701 = t0_0001010111101;
assign input_702 = t0_0001010111110;
assign input_703 = t0_0001010111111;
assign input_704 = t0_0001011000000;
assign input_705 = t0_0001011000001;
assign input_706 = t0_0001011000010;
assign input_707 = t0_0001011000011;
assign input_708 = t0_0001011000100;
assign input_709 = t0_0001011000101;
assign input_710 = t0_0001011000110;
assign input_711 = t0_0001011000111;
assign input_712 = t0_0001011001000;
assign input_713 = t0_0001011001001;
assign input_714 = t0_0001011001010;
assign input_715 = t0_0001011001011;
assign input_716 = t0_0001011001100;
assign input_717 = t0_0001011001101;
assign input_718 = t0_0001011001110;
assign input_719 = t0_0001011001111;
assign input_720 = t0_0001011010000;
assign input_721 = t0_0001011010001;
assign input_722 = t0_0001011010010;
assign input_723 = t0_0001011010011;
assign input_724 = t0_0001011010100;
assign input_725 = t0_0001011010101;
assign input_726 = t0_0001011010110;
assign input_727 = t0_0001011010111;
assign input_728 = t0_0001011011000;
assign input_729 = t0_0001011011001;
assign input_730 = t0_0001011011010;
assign input_731 = t0_0001011011011;
assign input_732 = t0_0001011011100;
assign input_733 = t0_0001011011101;
assign input_734 = t0_0001011011110;
assign input_735 = t0_0001011011111;
assign input_736 = t0_0001011100000;
assign input_737 = t0_0001011100001;
assign input_738 = t0_0001011100010;
assign input_739 = t0_0001011100011;
assign input_740 = t0_0001011100100;
assign input_741 = t0_0001011100101;
assign input_742 = t0_0001011100110;
assign input_743 = t0_0001011100111;
assign input_744 = t0_0001011101000;
assign input_745 = t0_0001011101001;
assign input_746 = t0_0001011101010;
assign input_747 = t0_0001011101011;
assign input_748 = t0_0001011101100;
assign input_749 = t0_0001011101101;
assign input_750 = t0_0001011101110;
assign input_751 = t0_0001011101111;
assign input_752 = t0_0001011110000;
assign input_753 = t0_0001011110001;
assign input_754 = t0_0001011110010;
assign input_755 = t0_0001011110011;
assign input_756 = t0_0001011110100;
assign input_757 = t0_0001011110101;
assign input_758 = t0_0001011110110;
assign input_759 = t0_0001011110111;
assign input_760 = t0_0001011111000;
assign input_761 = t0_0001011111001;
assign input_762 = t0_0001011111010;
assign input_763 = t0_0001011111011;
assign input_764 = t0_0001011111100;
assign input_765 = t0_0001011111101;
assign input_766 = t0_0001011111110;
assign input_767 = t0_0001011111111;
assign input_768 = t0_0001100000000;
assign input_769 = t0_0001100000001;
assign input_770 = t0_0001100000010;
assign input_771 = t0_0001100000011;
assign input_772 = t0_0001100000100;
assign input_773 = t0_0001100000101;
assign input_774 = t0_0001100000110;
assign input_775 = t0_0001100000111;
assign input_776 = t0_0001100001000;
assign input_777 = t0_0001100001001;
assign input_778 = t0_0001100001010;
assign input_779 = t0_0001100001011;
assign input_780 = t0_0001100001100;
assign input_781 = t0_0001100001101;
assign input_782 = t0_0001100001110;
assign input_783 = t0_0001100001111;
assign input_784 = t0_0001100010000;
assign input_785 = t0_0001100010001;
assign input_786 = t0_0001100010010;
assign input_787 = t0_0001100010011;
assign input_788 = t0_0001100010100;
assign input_789 = t0_0001100010101;
assign input_790 = t0_0001100010110;
assign input_791 = t0_0001100010111;
assign input_792 = t0_0001100011000;
assign input_793 = t0_0001100011001;
assign input_794 = t0_0001100011010;
assign input_795 = t0_0001100011011;
assign input_796 = t0_0001100011100;
assign input_797 = t0_0001100011101;
assign input_798 = t0_0001100011110;
assign input_799 = t0_0001100011111;
assign input_800 = t0_0001100100000;
assign input_801 = t0_0001100100001;
assign input_802 = t0_0001100100010;
assign input_803 = t0_0001100100011;
assign input_804 = t0_0001100100100;
assign input_805 = t0_0001100100101;
assign input_806 = t0_0001100100110;
assign input_807 = t0_0001100100111;
assign input_808 = t0_0001100101000;
assign input_809 = t0_0001100101001;
assign input_810 = t0_0001100101010;
assign input_811 = t0_0001100101011;
assign input_812 = t0_0001100101100;
assign input_813 = t0_0001100101101;
assign input_814 = t0_0001100101110;
assign input_815 = t0_0001100101111;
assign input_816 = t0_0001100110000;
assign input_817 = t0_0001100110001;
assign input_818 = t0_0001100110010;
assign input_819 = t0_0001100110011;
assign input_820 = t0_0001100110100;
assign input_821 = t0_0001100110101;
assign input_822 = t0_0001100110110;
assign input_823 = t0_0001100110111;
assign input_824 = t0_0001100111000;
assign input_825 = t0_0001100111001;
assign input_826 = t0_0001100111010;
assign input_827 = t0_0001100111011;
assign input_828 = t0_0001100111100;
assign input_829 = t0_0001100111101;
assign input_830 = t0_0001100111110;
assign input_831 = t0_0001100111111;
assign input_832 = t0_0001101000000;
assign input_833 = t0_0001101000001;
assign input_834 = t0_0001101000010;
assign input_835 = t0_0001101000011;
assign input_836 = t0_0001101000100;
assign input_837 = t0_0001101000101;
assign input_838 = t0_0001101000110;
assign input_839 = t0_0001101000111;
assign input_840 = t0_0001101001000;
assign input_841 = t0_0001101001001;
assign input_842 = t0_0001101001010;
assign input_843 = t0_0001101001011;
assign input_844 = t0_0001101001100;
assign input_845 = t0_0001101001101;
assign input_846 = t0_0001101001110;
assign input_847 = t0_0001101001111;
assign input_848 = t0_0001101010000;
assign input_849 = t0_0001101010001;
assign input_850 = t0_0001101010010;
assign input_851 = t0_0001101010011;
assign input_852 = t0_0001101010100;
assign input_853 = t0_0001101010101;
assign input_854 = t0_0001101010110;
assign input_855 = t0_0001101010111;
assign input_856 = t0_0001101011000;
assign input_857 = t0_0001101011001;
assign input_858 = t0_0001101011010;
assign input_859 = t0_0001101011011;
assign input_860 = t0_0001101011100;
assign input_861 = t0_0001101011101;
assign input_862 = t0_0001101011110;
assign input_863 = t0_0001101011111;
assign input_864 = t0_0001101100000;
assign input_865 = t0_0001101100001;
assign input_866 = t0_0001101100010;
assign input_867 = t0_0001101100011;
assign input_868 = t0_0001101100100;
assign input_869 = t0_0001101100101;
assign input_870 = t0_0001101100110;
assign input_871 = t0_0001101100111;
assign input_872 = t0_0001101101000;
assign input_873 = t0_0001101101001;
assign input_874 = t0_0001101101010;
assign input_875 = t0_0001101101011;
assign input_876 = t0_0001101101100;
assign input_877 = t0_0001101101101;
assign input_878 = t0_0001101101110;
assign input_879 = t0_0001101101111;
assign input_880 = t0_0001101110000;
assign input_881 = t0_0001101110001;
assign input_882 = t0_0001101110010;
assign input_883 = t0_0001101110011;
assign input_884 = t0_0001101110100;
assign input_885 = t0_0001101110101;
assign input_886 = t0_0001101110110;
assign input_887 = t0_0001101110111;
assign input_888 = t0_0001101111000;
assign input_889 = t0_0001101111001;
assign input_890 = t0_0001101111010;
assign input_891 = t0_0001101111011;
assign input_892 = t0_0001101111100;
assign input_893 = t0_0001101111101;
assign input_894 = t0_0001101111110;
assign input_895 = t0_0001101111111;
assign input_896 = t0_0001110000000;
assign input_897 = t0_0001110000001;
assign input_898 = t0_0001110000010;
assign input_899 = t0_0001110000011;
assign input_900 = t0_0001110000100;
assign input_901 = t0_0001110000101;
assign input_902 = t0_0001110000110;
assign input_903 = t0_0001110000111;
assign input_904 = t0_0001110001000;
assign input_905 = t0_0001110001001;
assign input_906 = t0_0001110001010;
assign input_907 = t0_0001110001011;
assign input_908 = t0_0001110001100;
assign input_909 = t0_0001110001101;
assign input_910 = t0_0001110001110;
assign input_911 = t0_0001110001111;
assign input_912 = t0_0001110010000;
assign input_913 = t0_0001110010001;
assign input_914 = t0_0001110010010;
assign input_915 = t0_0001110010011;
assign input_916 = t0_0001110010100;
assign input_917 = t0_0001110010101;
assign input_918 = t0_0001110010110;
assign input_919 = t0_0001110010111;
assign input_920 = t0_0001110011000;
assign input_921 = t0_0001110011001;
assign input_922 = t0_0001110011010;
assign input_923 = t0_0001110011011;
assign input_924 = t0_0001110011100;
assign input_925 = t0_0001110011101;
assign input_926 = t0_0001110011110;
assign input_927 = t0_0001110011111;
assign input_928 = t0_0001110100000;
assign input_929 = t0_0001110100001;
assign input_930 = t0_0001110100010;
assign input_931 = t0_0001110100011;
assign input_932 = t0_0001110100100;
assign input_933 = t0_0001110100101;
assign input_934 = t0_0001110100110;
assign input_935 = t0_0001110100111;
assign input_936 = t0_0001110101000;
assign input_937 = t0_0001110101001;
assign input_938 = t0_0001110101010;
assign input_939 = t0_0001110101011;
assign input_940 = t0_0001110101100;
assign input_941 = t0_0001110101101;
assign input_942 = t0_0001110101110;
assign input_943 = t0_0001110101111;
assign input_944 = t0_0001110110000;
assign input_945 = t0_0001110110001;
assign input_946 = t0_0001110110010;
assign input_947 = t0_0001110110011;
assign input_948 = t0_0001110110100;
assign input_949 = t0_0001110110101;
assign input_950 = t0_0001110110110;
assign input_951 = t0_0001110110111;
assign input_952 = t0_0001110111000;
assign input_953 = t0_0001110111001;
assign input_954 = t0_0001110111010;
assign input_955 = t0_0001110111011;
assign input_956 = t0_0001110111100;
assign input_957 = t0_0001110111101;
assign input_958 = t0_0001110111110;
assign input_959 = t0_0001110111111;
assign input_960 = t0_0001111000000;
assign input_961 = t0_0001111000001;
assign input_962 = t0_0001111000010;
assign input_963 = t0_0001111000011;
assign input_964 = t0_0001111000100;
assign input_965 = t0_0001111000101;
assign input_966 = t0_0001111000110;
assign input_967 = t0_0001111000111;
assign input_968 = t0_0001111001000;
assign input_969 = t0_0001111001001;
assign input_970 = t0_0001111001010;
assign input_971 = t0_0001111001011;
assign input_972 = t0_0001111001100;
assign input_973 = t0_0001111001101;
assign input_974 = t0_0001111001110;
assign input_975 = t0_0001111001111;
assign input_976 = t0_0001111010000;
assign input_977 = t0_0001111010001;
assign input_978 = t0_0001111010010;
assign input_979 = t0_0001111010011;
assign input_980 = t0_0001111010100;
assign input_981 = t0_0001111010101;
assign input_982 = t0_0001111010110;
assign input_983 = t0_0001111010111;
assign input_984 = t0_0001111011000;
assign input_985 = t0_0001111011001;
assign input_986 = t0_0001111011010;
assign input_987 = t0_0001111011011;
assign input_988 = t0_0001111011100;
assign input_989 = t0_0001111011101;
assign input_990 = t0_0001111011110;
assign input_991 = t0_0001111011111;
assign input_992 = t0_0001111100000;
assign input_993 = t0_0001111100001;
assign input_994 = t0_0001111100010;
assign input_995 = t0_0001111100011;
assign input_996 = t0_0001111100100;
assign input_997 = t0_0001111100101;
assign input_998 = t0_0001111100110;
assign input_999 = t0_0001111100111;
assign input_1000 = t0_0001111101000;
assign input_1001 = t0_0001111101001;
assign input_1002 = t0_0001111101010;
assign input_1003 = t0_0001111101011;
assign input_1004 = t0_0001111101100;
assign input_1005 = t0_0001111101101;
assign input_1006 = t0_0001111101110;
assign input_1007 = t0_0001111101111;
assign input_1008 = t0_0001111110000;
assign input_1009 = t0_0001111110001;
assign input_1010 = t0_0001111110010;
assign input_1011 = t0_0001111110011;
assign input_1012 = t0_0001111110100;
assign input_1013 = t0_0001111110101;
assign input_1014 = t0_0001111110110;
assign input_1015 = t0_0001111110111;
assign input_1016 = t0_0001111111000;
assign input_1017 = t0_0001111111001;
assign input_1018 = t0_0001111111010;
assign input_1019 = t0_0001111111011;
assign input_1020 = t0_0001111111100;
assign input_1021 = t0_0001111111101;
assign input_1022 = t0_0001111111110;
assign input_1023 = t0_0001111111111;
assign input_1024 = t0_0010000000000;
assign input_1025 = t0_0010000000001;
assign input_1026 = t0_0010000000010;
assign input_1027 = t0_0010000000011;
assign input_1028 = t0_0010000000100;
assign input_1029 = t0_0010000000101;
assign input_1030 = t0_0010000000110;
assign input_1031 = t0_0010000000111;
assign input_1032 = t0_0010000001000;
assign input_1033 = t0_0010000001001;
assign input_1034 = t0_0010000001010;
assign input_1035 = t0_0010000001011;
assign input_1036 = t0_0010000001100;
assign input_1037 = t0_0010000001101;
assign input_1038 = t0_0010000001110;
assign input_1039 = t0_0010000001111;
assign input_1040 = t0_0010000010000;
assign input_1041 = t0_0010000010001;
assign input_1042 = t0_0010000010010;
assign input_1043 = t0_0010000010011;
assign input_1044 = t0_0010000010100;
assign input_1045 = t0_0010000010101;
assign input_1046 = t0_0010000010110;
assign input_1047 = t0_0010000010111;
assign input_1048 = t0_0010000011000;
assign input_1049 = t0_0010000011001;
assign input_1050 = t0_0010000011010;
assign input_1051 = t0_0010000011011;
assign input_1052 = t0_0010000011100;
assign input_1053 = t0_0010000011101;
assign input_1054 = t0_0010000011110;
assign input_1055 = t0_0010000011111;
assign input_1056 = t0_0010000100000;
assign input_1057 = t0_0010000100001;
assign input_1058 = t0_0010000100010;
assign input_1059 = t0_0010000100011;
assign input_1060 = t0_0010000100100;
assign input_1061 = t0_0010000100101;
assign input_1062 = t0_0010000100110;
assign input_1063 = t0_0010000100111;
assign input_1064 = t0_0010000101000;
assign input_1065 = t0_0010000101001;
assign input_1066 = t0_0010000101010;
assign input_1067 = t0_0010000101011;
assign input_1068 = t0_0010000101100;
assign input_1069 = t0_0010000101101;
assign input_1070 = t0_0010000101110;
assign input_1071 = t0_0010000101111;
assign input_1072 = t0_0010000110000;
assign input_1073 = t0_0010000110001;
assign input_1074 = t0_0010000110010;
assign input_1075 = t0_0010000110011;
assign input_1076 = t0_0010000110100;
assign input_1077 = t0_0010000110101;
assign input_1078 = t0_0010000110110;
assign input_1079 = t0_0010000110111;
assign input_1080 = t0_0010000111000;
assign input_1081 = t0_0010000111001;
assign input_1082 = t0_0010000111010;
assign input_1083 = t0_0010000111011;
assign input_1084 = t0_0010000111100;
assign input_1085 = t0_0010000111101;
assign input_1086 = t0_0010000111110;
assign input_1087 = t0_0010000111111;
assign input_1088 = t0_0010001000000;
assign input_1089 = t0_0010001000001;
assign input_1090 = t0_0010001000010;
assign input_1091 = t0_0010001000011;
assign input_1092 = t0_0010001000100;
assign input_1093 = t0_0010001000101;
assign input_1094 = t0_0010001000110;
assign input_1095 = t0_0010001000111;
assign input_1096 = t0_0010001001000;
assign input_1097 = t0_0010001001001;
assign input_1098 = t0_0010001001010;
assign input_1099 = t0_0010001001011;
assign input_1100 = t0_0010001001100;
assign input_1101 = t0_0010001001101;
assign input_1102 = t0_0010001001110;
assign input_1103 = t0_0010001001111;
assign input_1104 = t0_0010001010000;
assign input_1105 = t0_0010001010001;
assign input_1106 = t0_0010001010010;
assign input_1107 = t0_0010001010011;
assign input_1108 = t0_0010001010100;
assign input_1109 = t0_0010001010101;
assign input_1110 = t0_0010001010110;
assign input_1111 = t0_0010001010111;
assign input_1112 = t0_0010001011000;
assign input_1113 = t0_0010001011001;
assign input_1114 = t0_0010001011010;
assign input_1115 = t0_0010001011011;
assign input_1116 = t0_0010001011100;
assign input_1117 = t0_0010001011101;
assign input_1118 = t0_0010001011110;
assign input_1119 = t0_0010001011111;
assign input_1120 = t0_0010001100000;
assign input_1121 = t0_0010001100001;
assign input_1122 = t0_0010001100010;
assign input_1123 = t0_0010001100011;
assign input_1124 = t0_0010001100100;
assign input_1125 = t0_0010001100101;
assign input_1126 = t0_0010001100110;
assign input_1127 = t0_0010001100111;
assign input_1128 = t0_0010001101000;
assign input_1129 = t0_0010001101001;
assign input_1130 = t0_0010001101010;
assign input_1131 = t0_0010001101011;
assign input_1132 = t0_0010001101100;
assign input_1133 = t0_0010001101101;
assign input_1134 = t0_0010001101110;
assign input_1135 = t0_0010001101111;
assign input_1136 = t0_0010001110000;
assign input_1137 = t0_0010001110001;
assign input_1138 = t0_0010001110010;
assign input_1139 = t0_0010001110011;
assign input_1140 = t0_0010001110100;
assign input_1141 = t0_0010001110101;
assign input_1142 = t0_0010001110110;
assign input_1143 = t0_0010001110111;
assign input_1144 = t0_0010001111000;
assign input_1145 = t0_0010001111001;
assign input_1146 = t0_0010001111010;
assign input_1147 = t0_0010001111011;
assign input_1148 = t0_0010001111100;
assign input_1149 = t0_0010001111101;
assign input_1150 = t0_0010001111110;
assign input_1151 = t0_0010001111111;
assign input_1152 = t0_0010010000000;
assign input_1153 = t0_0010010000001;
assign input_1154 = t0_0010010000010;
assign input_1155 = t0_0010010000011;
assign input_1156 = t0_0010010000100;
assign input_1157 = t0_0010010000101;
assign input_1158 = t0_0010010000110;
assign input_1159 = t0_0010010000111;
assign input_1160 = t0_0010010001000;
assign input_1161 = t0_0010010001001;
assign input_1162 = t0_0010010001010;
assign input_1163 = t0_0010010001011;
assign input_1164 = t0_0010010001100;
assign input_1165 = t0_0010010001101;
assign input_1166 = t0_0010010001110;
assign input_1167 = t0_0010010001111;
assign input_1168 = t0_0010010010000;
assign input_1169 = t0_0010010010001;
assign input_1170 = t0_0010010010010;
assign input_1171 = t0_0010010010011;
assign input_1172 = t0_0010010010100;
assign input_1173 = t0_0010010010101;
assign input_1174 = t0_0010010010110;
assign input_1175 = t0_0010010010111;
assign input_1176 = t0_0010010011000;
assign input_1177 = t0_0010010011001;
assign input_1178 = t0_0010010011010;
assign input_1179 = t0_0010010011011;
assign input_1180 = t0_0010010011100;
assign input_1181 = t0_0010010011101;
assign input_1182 = t0_0010010011110;
assign input_1183 = t0_0010010011111;
assign input_1184 = t0_0010010100000;
assign input_1185 = t0_0010010100001;
assign input_1186 = t0_0010010100010;
assign input_1187 = t0_0010010100011;
assign input_1188 = t0_0010010100100;
assign input_1189 = t0_0010010100101;
assign input_1190 = t0_0010010100110;
assign input_1191 = t0_0010010100111;
assign input_1192 = t0_0010010101000;
assign input_1193 = t0_0010010101001;
assign input_1194 = t0_0010010101010;
assign input_1195 = t0_0010010101011;
assign input_1196 = t0_0010010101100;
assign input_1197 = t0_0010010101101;
assign input_1198 = t0_0010010101110;
assign input_1199 = t0_0010010101111;
assign input_1200 = t0_0010010110000;
assign input_1201 = t0_0010010110001;
assign input_1202 = t0_0010010110010;
assign input_1203 = t0_0010010110011;
assign input_1204 = t0_0010010110100;
assign input_1205 = t0_0010010110101;
assign input_1206 = t0_0010010110110;
assign input_1207 = t0_0010010110111;
assign input_1208 = t0_0010010111000;
assign input_1209 = t0_0010010111001;
assign input_1210 = t0_0010010111010;
assign input_1211 = t0_0010010111011;
assign input_1212 = t0_0010010111100;
assign input_1213 = t0_0010010111101;
assign input_1214 = t0_0010010111110;
assign input_1215 = t0_0010010111111;
assign input_1216 = t0_0010011000000;
assign input_1217 = t0_0010011000001;
assign input_1218 = t0_0010011000010;
assign input_1219 = t0_0010011000011;
assign input_1220 = t0_0010011000100;
assign input_1221 = t0_0010011000101;
assign input_1222 = t0_0010011000110;
assign input_1223 = t0_0010011000111;
assign input_1224 = t0_0010011001000;
assign input_1225 = t0_0010011001001;
assign input_1226 = t0_0010011001010;
assign input_1227 = t0_0010011001011;
assign input_1228 = t0_0010011001100;
assign input_1229 = t0_0010011001101;
assign input_1230 = t0_0010011001110;
assign input_1231 = t0_0010011001111;
assign input_1232 = t0_0010011010000;
assign input_1233 = t0_0010011010001;
assign input_1234 = t0_0010011010010;
assign input_1235 = t0_0010011010011;
assign input_1236 = t0_0010011010100;
assign input_1237 = t0_0010011010101;
assign input_1238 = t0_0010011010110;
assign input_1239 = t0_0010011010111;
assign input_1240 = t0_0010011011000;
assign input_1241 = t0_0010011011001;
assign input_1242 = t0_0010011011010;
assign input_1243 = t0_0010011011011;
assign input_1244 = t0_0010011011100;
assign input_1245 = t0_0010011011101;
assign input_1246 = t0_0010011011110;
assign input_1247 = t0_0010011011111;
assign input_1248 = t0_0010011100000;
assign input_1249 = t0_0010011100001;
assign input_1250 = t0_0010011100010;
assign input_1251 = t0_0010011100011;
assign input_1252 = t0_0010011100100;
assign input_1253 = t0_0010011100101;
assign input_1254 = t0_0010011100110;
assign input_1255 = t0_0010011100111;
assign input_1256 = t0_0010011101000;
assign input_1257 = t0_0010011101001;
assign input_1258 = t0_0010011101010;
assign input_1259 = t0_0010011101011;
assign input_1260 = t0_0010011101100;
assign input_1261 = t0_0010011101101;
assign input_1262 = t0_0010011101110;
assign input_1263 = t0_0010011101111;
assign input_1264 = t0_0010011110000;
assign input_1265 = t0_0010011110001;
assign input_1266 = t0_0010011110010;
assign input_1267 = t0_0010011110011;
assign input_1268 = t0_0010011110100;
assign input_1269 = t0_0010011110101;
assign input_1270 = t0_0010011110110;
assign input_1271 = t0_0010011110111;
assign input_1272 = t0_0010011111000;
assign input_1273 = t0_0010011111001;
assign input_1274 = t0_0010011111010;
assign input_1275 = t0_0010011111011;
assign input_1276 = t0_0010011111100;
assign input_1277 = t0_0010011111101;
assign input_1278 = t0_0010011111110;
assign input_1279 = t0_0010011111111;
assign input_1280 = t0_0010100000000;
assign input_1281 = t0_0010100000001;
assign input_1282 = t0_0010100000010;
assign input_1283 = t0_0010100000011;
assign input_1284 = t0_0010100000100;
assign input_1285 = t0_0010100000101;
assign input_1286 = t0_0010100000110;
assign input_1287 = t0_0010100000111;
assign input_1288 = t0_0010100001000;
assign input_1289 = t0_0010100001001;
assign input_1290 = t0_0010100001010;
assign input_1291 = t0_0010100001011;
assign input_1292 = t0_0010100001100;
assign input_1293 = t0_0010100001101;
assign input_1294 = t0_0010100001110;
assign input_1295 = t0_0010100001111;
assign input_1296 = t0_0010100010000;
assign input_1297 = t0_0010100010001;
assign input_1298 = t0_0010100010010;
assign input_1299 = t0_0010100010011;
assign input_1300 = t0_0010100010100;
assign input_1301 = t0_0010100010101;
assign input_1302 = t0_0010100010110;
assign input_1303 = t0_0010100010111;
assign input_1304 = t0_0010100011000;
assign input_1305 = t0_0010100011001;
assign input_1306 = t0_0010100011010;
assign input_1307 = t0_0010100011011;
assign input_1308 = t0_0010100011100;
assign input_1309 = t0_0010100011101;
assign input_1310 = t0_0010100011110;
assign input_1311 = t0_0010100011111;
assign input_1312 = t0_0010100100000;
assign input_1313 = t0_0010100100001;
assign input_1314 = t0_0010100100010;
assign input_1315 = t0_0010100100011;
assign input_1316 = t0_0010100100100;
assign input_1317 = t0_0010100100101;
assign input_1318 = t0_0010100100110;
assign input_1319 = t0_0010100100111;
assign input_1320 = t0_0010100101000;
assign input_1321 = t0_0010100101001;
assign input_1322 = t0_0010100101010;
assign input_1323 = t0_0010100101011;
assign input_1324 = t0_0010100101100;
assign input_1325 = t0_0010100101101;
assign input_1326 = t0_0010100101110;
assign input_1327 = t0_0010100101111;
assign input_1328 = t0_0010100110000;
assign input_1329 = t0_0010100110001;
assign input_1330 = t0_0010100110010;
assign input_1331 = t0_0010100110011;
assign input_1332 = t0_0010100110100;
assign input_1333 = t0_0010100110101;
assign input_1334 = t0_0010100110110;
assign input_1335 = t0_0010100110111;
assign input_1336 = t0_0010100111000;
assign input_1337 = t0_0010100111001;
assign input_1338 = t0_0010100111010;
assign input_1339 = t0_0010100111011;
assign input_1340 = t0_0010100111100;
assign input_1341 = t0_0010100111101;
assign input_1342 = t0_0010100111110;
assign input_1343 = t0_0010100111111;
assign input_1344 = t0_0010101000000;
assign input_1345 = t0_0010101000001;
assign input_1346 = t0_0010101000010;
assign input_1347 = t0_0010101000011;
assign input_1348 = t0_0010101000100;
assign input_1349 = t0_0010101000101;
assign input_1350 = t0_0010101000110;
assign input_1351 = t0_0010101000111;
assign input_1352 = t0_0010101001000;
assign input_1353 = t0_0010101001001;
assign input_1354 = t0_0010101001010;
assign input_1355 = t0_0010101001011;
assign input_1356 = t0_0010101001100;
assign input_1357 = t0_0010101001101;
assign input_1358 = t0_0010101001110;
assign input_1359 = t0_0010101001111;
assign input_1360 = t0_0010101010000;
assign input_1361 = t0_0010101010001;
assign input_1362 = t0_0010101010010;
assign input_1363 = t0_0010101010011;
assign input_1364 = t0_0010101010100;
assign input_1365 = t0_0010101010101;
assign input_1366 = t0_0010101010110;
assign input_1367 = t0_0010101010111;
assign input_1368 = t0_0010101011000;
assign input_1369 = t0_0010101011001;
assign input_1370 = t0_0010101011010;
assign input_1371 = t0_0010101011011;
assign input_1372 = t0_0010101011100;
assign input_1373 = t0_0010101011101;
assign input_1374 = t0_0010101011110;
assign input_1375 = t0_0010101011111;
assign input_1376 = t0_0010101100000;
assign input_1377 = t0_0010101100001;
assign input_1378 = t0_0010101100010;
assign input_1379 = t0_0010101100011;
assign input_1380 = t0_0010101100100;
assign input_1381 = t0_0010101100101;
assign input_1382 = t0_0010101100110;
assign input_1383 = t0_0010101100111;
assign input_1384 = t0_0010101101000;
assign input_1385 = t0_0010101101001;
assign input_1386 = t0_0010101101010;
assign input_1387 = t0_0010101101011;
assign input_1388 = t0_0010101101100;
assign input_1389 = t0_0010101101101;
assign input_1390 = t0_0010101101110;
assign input_1391 = t0_0010101101111;
assign input_1392 = t0_0010101110000;
assign input_1393 = t0_0010101110001;
assign input_1394 = t0_0010101110010;
assign input_1395 = t0_0010101110011;
assign input_1396 = t0_0010101110100;
assign input_1397 = t0_0010101110101;
assign input_1398 = t0_0010101110110;
assign input_1399 = t0_0010101110111;
assign input_1400 = t0_0010101111000;
assign input_1401 = t0_0010101111001;
assign input_1402 = t0_0010101111010;
assign input_1403 = t0_0010101111011;
assign input_1404 = t0_0010101111100;
assign input_1405 = t0_0010101111101;
assign input_1406 = t0_0010101111110;
assign input_1407 = t0_0010101111111;
assign input_1408 = t0_0010110000000;
assign input_1409 = t0_0010110000001;
assign input_1410 = t0_0010110000010;
assign input_1411 = t0_0010110000011;
assign input_1412 = t0_0010110000100;
assign input_1413 = t0_0010110000101;
assign input_1414 = t0_0010110000110;
assign input_1415 = t0_0010110000111;
assign input_1416 = t0_0010110001000;
assign input_1417 = t0_0010110001001;
assign input_1418 = t0_0010110001010;
assign input_1419 = t0_0010110001011;
assign input_1420 = t0_0010110001100;
assign input_1421 = t0_0010110001101;
assign input_1422 = t0_0010110001110;
assign input_1423 = t0_0010110001111;
assign input_1424 = t0_0010110010000;
assign input_1425 = t0_0010110010001;
assign input_1426 = t0_0010110010010;
assign input_1427 = t0_0010110010011;
assign input_1428 = t0_0010110010100;
assign input_1429 = t0_0010110010101;
assign input_1430 = t0_0010110010110;
assign input_1431 = t0_0010110010111;
assign input_1432 = t0_0010110011000;
assign input_1433 = t0_0010110011001;
assign input_1434 = t0_0010110011010;
assign input_1435 = t0_0010110011011;
assign input_1436 = t0_0010110011100;
assign input_1437 = t0_0010110011101;
assign input_1438 = t0_0010110011110;
assign input_1439 = t0_0010110011111;
assign input_1440 = t0_0010110100000;
assign input_1441 = t0_0010110100001;
assign input_1442 = t0_0010110100010;
assign input_1443 = t0_0010110100011;
assign input_1444 = t0_0010110100100;
assign input_1445 = t0_0010110100101;
assign input_1446 = t0_0010110100110;
assign input_1447 = t0_0010110100111;
assign input_1448 = t0_0010110101000;
assign input_1449 = t0_0010110101001;
assign input_1450 = t0_0010110101010;
assign input_1451 = t0_0010110101011;
assign input_1452 = t0_0010110101100;
assign input_1453 = t0_0010110101101;
assign input_1454 = t0_0010110101110;
assign input_1455 = t0_0010110101111;
assign input_1456 = t0_0010110110000;
assign input_1457 = t0_0010110110001;
assign input_1458 = t0_0010110110010;
assign input_1459 = t0_0010110110011;
assign input_1460 = t0_0010110110100;
assign input_1461 = t0_0010110110101;
assign input_1462 = t0_0010110110110;
assign input_1463 = t0_0010110110111;
assign input_1464 = t0_0010110111000;
assign input_1465 = t0_0010110111001;
assign input_1466 = t0_0010110111010;
assign input_1467 = t0_0010110111011;
assign input_1468 = t0_0010110111100;
assign input_1469 = t0_0010110111101;
assign input_1470 = t0_0010110111110;
assign input_1471 = t0_0010110111111;
assign input_1472 = t0_0010111000000;
assign input_1473 = t0_0010111000001;
assign input_1474 = t0_0010111000010;
assign input_1475 = t0_0010111000011;
assign input_1476 = t0_0010111000100;
assign input_1477 = t0_0010111000101;
assign input_1478 = t0_0010111000110;
assign input_1479 = t0_0010111000111;
assign input_1480 = t0_0010111001000;
assign input_1481 = t0_0010111001001;
assign input_1482 = t0_0010111001010;
assign input_1483 = t0_0010111001011;
assign input_1484 = t0_0010111001100;
assign input_1485 = t0_0010111001101;
assign input_1486 = t0_0010111001110;
assign input_1487 = t0_0010111001111;
assign input_1488 = t0_0010111010000;
assign input_1489 = t0_0010111010001;
assign input_1490 = t0_0010111010010;
assign input_1491 = t0_0010111010011;
assign input_1492 = t0_0010111010100;
assign input_1493 = t0_0010111010101;
assign input_1494 = t0_0010111010110;
assign input_1495 = t0_0010111010111;
assign input_1496 = t0_0010111011000;
assign input_1497 = t0_0010111011001;
assign input_1498 = t0_0010111011010;
assign input_1499 = t0_0010111011011;
assign input_1500 = t0_0010111011100;
assign input_1501 = t0_0010111011101;
assign input_1502 = t0_0010111011110;
assign input_1503 = t0_0010111011111;
assign input_1504 = t0_0010111100000;
assign input_1505 = t0_0010111100001;
assign input_1506 = t0_0010111100010;
assign input_1507 = t0_0010111100011;
assign input_1508 = t0_0010111100100;
assign input_1509 = t0_0010111100101;
assign input_1510 = t0_0010111100110;
assign input_1511 = t0_0010111100111;
assign input_1512 = t0_0010111101000;
assign input_1513 = t0_0010111101001;
assign input_1514 = t0_0010111101010;
assign input_1515 = t0_0010111101011;
assign input_1516 = t0_0010111101100;
assign input_1517 = t0_0010111101101;
assign input_1518 = t0_0010111101110;
assign input_1519 = t0_0010111101111;
assign input_1520 = t0_0010111110000;
assign input_1521 = t0_0010111110001;
assign input_1522 = t0_0010111110010;
assign input_1523 = t0_0010111110011;
assign input_1524 = t0_0010111110100;
assign input_1525 = t0_0010111110101;
assign input_1526 = t0_0010111110110;
assign input_1527 = t0_0010111110111;
assign input_1528 = t0_0010111111000;
assign input_1529 = t0_0010111111001;
assign input_1530 = t0_0010111111010;
assign input_1531 = t0_0010111111011;
assign input_1532 = t0_0010111111100;
assign input_1533 = t0_0010111111101;
assign input_1534 = t0_0010111111110;
assign input_1535 = t0_0010111111111;
assign input_1536 = t0_0011000000000;
assign input_1537 = t0_0011000000001;
assign input_1538 = t0_0011000000010;
assign input_1539 = t0_0011000000011;
assign input_1540 = t0_0011000000100;
assign input_1541 = t0_0011000000101;
assign input_1542 = t0_0011000000110;
assign input_1543 = t0_0011000000111;
assign input_1544 = t0_0011000001000;
assign input_1545 = t0_0011000001001;
assign input_1546 = t0_0011000001010;
assign input_1547 = t0_0011000001011;
assign input_1548 = t0_0011000001100;
assign input_1549 = t0_0011000001101;
assign input_1550 = t0_0011000001110;
assign input_1551 = t0_0011000001111;
assign input_1552 = t0_0011000010000;
assign input_1553 = t0_0011000010001;
assign input_1554 = t0_0011000010010;
assign input_1555 = t0_0011000010011;
assign input_1556 = t0_0011000010100;
assign input_1557 = t0_0011000010101;
assign input_1558 = t0_0011000010110;
assign input_1559 = t0_0011000010111;
assign input_1560 = t0_0011000011000;
assign input_1561 = t0_0011000011001;
assign input_1562 = t0_0011000011010;
assign input_1563 = t0_0011000011011;
assign input_1564 = t0_0011000011100;
assign input_1565 = t0_0011000011101;
assign input_1566 = t0_0011000011110;
assign input_1567 = t0_0011000011111;
assign input_1568 = t0_0011000100000;
assign input_1569 = t0_0011000100001;
assign input_1570 = t0_0011000100010;
assign input_1571 = t0_0011000100011;
assign input_1572 = t0_0011000100100;
assign input_1573 = t0_0011000100101;
assign input_1574 = t0_0011000100110;
assign input_1575 = t0_0011000100111;
assign input_1576 = t0_0011000101000;
assign input_1577 = t0_0011000101001;
assign input_1578 = t0_0011000101010;
assign input_1579 = t0_0011000101011;
assign input_1580 = t0_0011000101100;
assign input_1581 = t0_0011000101101;
assign input_1582 = t0_0011000101110;
assign input_1583 = t0_0011000101111;
assign input_1584 = t0_0011000110000;
assign input_1585 = t0_0011000110001;
assign input_1586 = t0_0011000110010;
assign input_1587 = t0_0011000110011;
assign input_1588 = t0_0011000110100;
assign input_1589 = t0_0011000110101;
assign input_1590 = t0_0011000110110;
assign input_1591 = t0_0011000110111;
assign input_1592 = t0_0011000111000;
assign input_1593 = t0_0011000111001;
assign input_1594 = t0_0011000111010;
assign input_1595 = t0_0011000111011;
assign input_1596 = t0_0011000111100;
assign input_1597 = t0_0011000111101;
assign input_1598 = t0_0011000111110;
assign input_1599 = t0_0011000111111;
assign input_1600 = t0_0011001000000;
assign input_1601 = t0_0011001000001;
assign input_1602 = t0_0011001000010;
assign input_1603 = t0_0011001000011;
assign input_1604 = t0_0011001000100;
assign input_1605 = t0_0011001000101;
assign input_1606 = t0_0011001000110;
assign input_1607 = t0_0011001000111;
assign input_1608 = t0_0011001001000;
assign input_1609 = t0_0011001001001;
assign input_1610 = t0_0011001001010;
assign input_1611 = t0_0011001001011;
assign input_1612 = t0_0011001001100;
assign input_1613 = t0_0011001001101;
assign input_1614 = t0_0011001001110;
assign input_1615 = t0_0011001001111;
assign input_1616 = t0_0011001010000;
assign input_1617 = t0_0011001010001;
assign input_1618 = t0_0011001010010;
assign input_1619 = t0_0011001010011;
assign input_1620 = t0_0011001010100;
assign input_1621 = t0_0011001010101;
assign input_1622 = t0_0011001010110;
assign input_1623 = t0_0011001010111;
assign input_1624 = t0_0011001011000;
assign input_1625 = t0_0011001011001;
assign input_1626 = t0_0011001011010;
assign input_1627 = t0_0011001011011;
assign input_1628 = t0_0011001011100;
assign input_1629 = t0_0011001011101;
assign input_1630 = t0_0011001011110;
assign input_1631 = t0_0011001011111;
assign input_1632 = t0_0011001100000;
assign input_1633 = t0_0011001100001;
assign input_1634 = t0_0011001100010;
assign input_1635 = t0_0011001100011;
assign input_1636 = t0_0011001100100;
assign input_1637 = t0_0011001100101;
assign input_1638 = t0_0011001100110;
assign input_1639 = t0_0011001100111;
assign input_1640 = t0_0011001101000;
assign input_1641 = t0_0011001101001;
assign input_1642 = t0_0011001101010;
assign input_1643 = t0_0011001101011;
assign input_1644 = t0_0011001101100;
assign input_1645 = t0_0011001101101;
assign input_1646 = t0_0011001101110;
assign input_1647 = t0_0011001101111;
assign input_1648 = t0_0011001110000;
assign input_1649 = t0_0011001110001;
assign input_1650 = t0_0011001110010;
assign input_1651 = t0_0011001110011;
assign input_1652 = t0_0011001110100;
assign input_1653 = t0_0011001110101;
assign input_1654 = t0_0011001110110;
assign input_1655 = t0_0011001110111;
assign input_1656 = t0_0011001111000;
assign input_1657 = t0_0011001111001;
assign input_1658 = t0_0011001111010;
assign input_1659 = t0_0011001111011;
assign input_1660 = t0_0011001111100;
assign input_1661 = t0_0011001111101;
assign input_1662 = t0_0011001111110;
assign input_1663 = t0_0011001111111;
assign input_1664 = t0_0011010000000;
assign input_1665 = t0_0011010000001;
assign input_1666 = t0_0011010000010;
assign input_1667 = t0_0011010000011;
assign input_1668 = t0_0011010000100;
assign input_1669 = t0_0011010000101;
assign input_1670 = t0_0011010000110;
assign input_1671 = t0_0011010000111;
assign input_1672 = t0_0011010001000;
assign input_1673 = t0_0011010001001;
assign input_1674 = t0_0011010001010;
assign input_1675 = t0_0011010001011;
assign input_1676 = t0_0011010001100;
assign input_1677 = t0_0011010001101;
assign input_1678 = t0_0011010001110;
assign input_1679 = t0_0011010001111;
assign input_1680 = t0_0011010010000;
assign input_1681 = t0_0011010010001;
assign input_1682 = t0_0011010010010;
assign input_1683 = t0_0011010010011;
assign input_1684 = t0_0011010010100;
assign input_1685 = t0_0011010010101;
assign input_1686 = t0_0011010010110;
assign input_1687 = t0_0011010010111;
assign input_1688 = t0_0011010011000;
assign input_1689 = t0_0011010011001;
assign input_1690 = t0_0011010011010;
assign input_1691 = t0_0011010011011;
assign input_1692 = t0_0011010011100;
assign input_1693 = t0_0011010011101;
assign input_1694 = t0_0011010011110;
assign input_1695 = t0_0011010011111;
assign input_1696 = t0_0011010100000;
assign input_1697 = t0_0011010100001;
assign input_1698 = t0_0011010100010;
assign input_1699 = t0_0011010100011;
assign input_1700 = t0_0011010100100;
assign input_1701 = t0_0011010100101;
assign input_1702 = t0_0011010100110;
assign input_1703 = t0_0011010100111;
assign input_1704 = t0_0011010101000;
assign input_1705 = t0_0011010101001;
assign input_1706 = t0_0011010101010;
assign input_1707 = t0_0011010101011;
assign input_1708 = t0_0011010101100;
assign input_1709 = t0_0011010101101;
assign input_1710 = t0_0011010101110;
assign input_1711 = t0_0011010101111;
assign input_1712 = t0_0011010110000;
assign input_1713 = t0_0011010110001;
assign input_1714 = t0_0011010110010;
assign input_1715 = t0_0011010110011;
assign input_1716 = t0_0011010110100;
assign input_1717 = t0_0011010110101;
assign input_1718 = t0_0011010110110;
assign input_1719 = t0_0011010110111;
assign input_1720 = t0_0011010111000;
assign input_1721 = t0_0011010111001;
assign input_1722 = t0_0011010111010;
assign input_1723 = t0_0011010111011;
assign input_1724 = t0_0011010111100;
assign input_1725 = t0_0011010111101;
assign input_1726 = t0_0011010111110;
assign input_1727 = t0_0011010111111;
assign input_1728 = t0_0011011000000;
assign input_1729 = t0_0011011000001;
assign input_1730 = t0_0011011000010;
assign input_1731 = t0_0011011000011;
assign input_1732 = t0_0011011000100;
assign input_1733 = t0_0011011000101;
assign input_1734 = t0_0011011000110;
assign input_1735 = t0_0011011000111;
assign input_1736 = t0_0011011001000;
assign input_1737 = t0_0011011001001;
assign input_1738 = t0_0011011001010;
assign input_1739 = t0_0011011001011;
assign input_1740 = t0_0011011001100;
assign input_1741 = t0_0011011001101;
assign input_1742 = t0_0011011001110;
assign input_1743 = t0_0011011001111;
assign input_1744 = t0_0011011010000;
assign input_1745 = t0_0011011010001;
assign input_1746 = t0_0011011010010;
assign input_1747 = t0_0011011010011;
assign input_1748 = t0_0011011010100;
assign input_1749 = t0_0011011010101;
assign input_1750 = t0_0011011010110;
assign input_1751 = t0_0011011010111;
assign input_1752 = t0_0011011011000;
assign input_1753 = t0_0011011011001;
assign input_1754 = t0_0011011011010;
assign input_1755 = t0_0011011011011;
assign input_1756 = t0_0011011011100;
assign input_1757 = t0_0011011011101;
assign input_1758 = t0_0011011011110;
assign input_1759 = t0_0011011011111;
assign input_1760 = t0_0011011100000;
assign input_1761 = t0_0011011100001;
assign input_1762 = t0_0011011100010;
assign input_1763 = t0_0011011100011;
assign input_1764 = t0_0011011100100;
assign input_1765 = t0_0011011100101;
assign input_1766 = t0_0011011100110;
assign input_1767 = t0_0011011100111;
assign input_1768 = t0_0011011101000;
assign input_1769 = t0_0011011101001;
assign input_1770 = t0_0011011101010;
assign input_1771 = t0_0011011101011;
assign input_1772 = t0_0011011101100;
assign input_1773 = t0_0011011101101;
assign input_1774 = t0_0011011101110;
assign input_1775 = t0_0011011101111;
assign input_1776 = t0_0011011110000;
assign input_1777 = t0_0011011110001;
assign input_1778 = t0_0011011110010;
assign input_1779 = t0_0011011110011;
assign input_1780 = t0_0011011110100;
assign input_1781 = t0_0011011110101;
assign input_1782 = t0_0011011110110;
assign input_1783 = t0_0011011110111;
assign input_1784 = t0_0011011111000;
assign input_1785 = t0_0011011111001;
assign input_1786 = t0_0011011111010;
assign input_1787 = t0_0011011111011;
assign input_1788 = t0_0011011111100;
assign input_1789 = t0_0011011111101;
assign input_1790 = t0_0011011111110;
assign input_1791 = t0_0011011111111;
assign input_1792 = t0_0011100000000;
assign input_1793 = t0_0011100000001;
assign input_1794 = t0_0011100000010;
assign input_1795 = t0_0011100000011;
assign input_1796 = t0_0011100000100;
assign input_1797 = t0_0011100000101;
assign input_1798 = t0_0011100000110;
assign input_1799 = t0_0011100000111;
assign input_1800 = t0_0011100001000;
assign input_1801 = t0_0011100001001;
assign input_1802 = t0_0011100001010;
assign input_1803 = t0_0011100001011;
assign input_1804 = t0_0011100001100;
assign input_1805 = t0_0011100001101;
assign input_1806 = t0_0011100001110;
assign input_1807 = t0_0011100001111;
assign input_1808 = t0_0011100010000;
assign input_1809 = t0_0011100010001;
assign input_1810 = t0_0011100010010;
assign input_1811 = t0_0011100010011;
assign input_1812 = t0_0011100010100;
assign input_1813 = t0_0011100010101;
assign input_1814 = t0_0011100010110;
assign input_1815 = t0_0011100010111;
assign input_1816 = t0_0011100011000;
assign input_1817 = t0_0011100011001;
assign input_1818 = t0_0011100011010;
assign input_1819 = t0_0011100011011;
assign input_1820 = t0_0011100011100;
assign input_1821 = t0_0011100011101;
assign input_1822 = t0_0011100011110;
assign input_1823 = t0_0011100011111;
assign input_1824 = t0_0011100100000;
assign input_1825 = t0_0011100100001;
assign input_1826 = t0_0011100100010;
assign input_1827 = t0_0011100100011;
assign input_1828 = t0_0011100100100;
assign input_1829 = t0_0011100100101;
assign input_1830 = t0_0011100100110;
assign input_1831 = t0_0011100100111;
assign input_1832 = t0_0011100101000;
assign input_1833 = t0_0011100101001;
assign input_1834 = t0_0011100101010;
assign input_1835 = t0_0011100101011;
assign input_1836 = t0_0011100101100;
assign input_1837 = t0_0011100101101;
assign input_1838 = t0_0011100101110;
assign input_1839 = t0_0011100101111;
assign input_1840 = t0_0011100110000;
assign input_1841 = t0_0011100110001;
assign input_1842 = t0_0011100110010;
assign input_1843 = t0_0011100110011;
assign input_1844 = t0_0011100110100;
assign input_1845 = t0_0011100110101;
assign input_1846 = t0_0011100110110;
assign input_1847 = t0_0011100110111;
assign input_1848 = t0_0011100111000;
assign input_1849 = t0_0011100111001;
assign input_1850 = t0_0011100111010;
assign input_1851 = t0_0011100111011;
assign input_1852 = t0_0011100111100;
assign input_1853 = t0_0011100111101;
assign input_1854 = t0_0011100111110;
assign input_1855 = t0_0011100111111;
assign input_1856 = t0_0011101000000;
assign input_1857 = t0_0011101000001;
assign input_1858 = t0_0011101000010;
assign input_1859 = t0_0011101000011;
assign input_1860 = t0_0011101000100;
assign input_1861 = t0_0011101000101;
assign input_1862 = t0_0011101000110;
assign input_1863 = t0_0011101000111;
assign input_1864 = t0_0011101001000;
assign input_1865 = t0_0011101001001;
assign input_1866 = t0_0011101001010;
assign input_1867 = t0_0011101001011;
assign input_1868 = t0_0011101001100;
assign input_1869 = t0_0011101001101;
assign input_1870 = t0_0011101001110;
assign input_1871 = t0_0011101001111;
assign input_1872 = t0_0011101010000;
assign input_1873 = t0_0011101010001;
assign input_1874 = t0_0011101010010;
assign input_1875 = t0_0011101010011;
assign input_1876 = t0_0011101010100;
assign input_1877 = t0_0011101010101;
assign input_1878 = t0_0011101010110;
assign input_1879 = t0_0011101010111;
assign input_1880 = t0_0011101011000;
assign input_1881 = t0_0011101011001;
assign input_1882 = t0_0011101011010;
assign input_1883 = t0_0011101011011;
assign input_1884 = t0_0011101011100;
assign input_1885 = t0_0011101011101;
assign input_1886 = t0_0011101011110;
assign input_1887 = t0_0011101011111;
assign input_1888 = t0_0011101100000;
assign input_1889 = t0_0011101100001;
assign input_1890 = t0_0011101100010;
assign input_1891 = t0_0011101100011;
assign input_1892 = t0_0011101100100;
assign input_1893 = t0_0011101100101;
assign input_1894 = t0_0011101100110;
assign input_1895 = t0_0011101100111;
assign input_1896 = t0_0011101101000;
assign input_1897 = t0_0011101101001;
assign input_1898 = t0_0011101101010;
assign input_1899 = t0_0011101101011;
assign input_1900 = t0_0011101101100;
assign input_1901 = t0_0011101101101;
assign input_1902 = t0_0011101101110;
assign input_1903 = t0_0011101101111;
assign input_1904 = t0_0011101110000;
assign input_1905 = t0_0011101110001;
assign input_1906 = t0_0011101110010;
assign input_1907 = t0_0011101110011;
assign input_1908 = t0_0011101110100;
assign input_1909 = t0_0011101110101;
assign input_1910 = t0_0011101110110;
assign input_1911 = t0_0011101110111;
assign input_1912 = t0_0011101111000;
assign input_1913 = t0_0011101111001;
assign input_1914 = t0_0011101111010;
assign input_1915 = t0_0011101111011;
assign input_1916 = t0_0011101111100;
assign input_1917 = t0_0011101111101;
assign input_1918 = t0_0011101111110;
assign input_1919 = t0_0011101111111;
assign input_1920 = t0_0011110000000;
assign input_1921 = t0_0011110000001;
assign input_1922 = t0_0011110000010;
assign input_1923 = t0_0011110000011;
assign input_1924 = t0_0011110000100;
assign input_1925 = t0_0011110000101;
assign input_1926 = t0_0011110000110;
assign input_1927 = t0_0011110000111;
assign input_1928 = t0_0011110001000;
assign input_1929 = t0_0011110001001;
assign input_1930 = t0_0011110001010;
assign input_1931 = t0_0011110001011;
assign input_1932 = t0_0011110001100;
assign input_1933 = t0_0011110001101;
assign input_1934 = t0_0011110001110;
assign input_1935 = t0_0011110001111;
assign input_1936 = t0_0011110010000;
assign input_1937 = t0_0011110010001;
assign input_1938 = t0_0011110010010;
assign input_1939 = t0_0011110010011;
assign input_1940 = t0_0011110010100;
assign input_1941 = t0_0011110010101;
assign input_1942 = t0_0011110010110;
assign input_1943 = t0_0011110010111;
assign input_1944 = t0_0011110011000;
assign input_1945 = t0_0011110011001;
assign input_1946 = t0_0011110011010;
assign input_1947 = t0_0011110011011;
assign input_1948 = t0_0011110011100;
assign input_1949 = t0_0011110011101;
assign input_1950 = t0_0011110011110;
assign input_1951 = t0_0011110011111;
assign input_1952 = t0_0011110100000;
assign input_1953 = t0_0011110100001;
assign input_1954 = t0_0011110100010;
assign input_1955 = t0_0011110100011;
assign input_1956 = t0_0011110100100;
assign input_1957 = t0_0011110100101;
assign input_1958 = t0_0011110100110;
assign input_1959 = t0_0011110100111;
assign input_1960 = t0_0011110101000;
assign input_1961 = t0_0011110101001;
assign input_1962 = t0_0011110101010;
assign input_1963 = t0_0011110101011;
assign input_1964 = t0_0011110101100;
assign input_1965 = t0_0011110101101;
assign input_1966 = t0_0011110101110;
assign input_1967 = t0_0011110101111;
assign input_1968 = t0_0011110110000;
assign input_1969 = t0_0011110110001;
assign input_1970 = t0_0011110110010;
assign input_1971 = t0_0011110110011;
assign input_1972 = t0_0011110110100;
assign input_1973 = t0_0011110110101;
assign input_1974 = t0_0011110110110;
assign input_1975 = t0_0011110110111;
assign input_1976 = t0_0011110111000;
assign input_1977 = t0_0011110111001;
assign input_1978 = t0_0011110111010;
assign input_1979 = t0_0011110111011;
assign input_1980 = t0_0011110111100;
assign input_1981 = t0_0011110111101;
assign input_1982 = t0_0011110111110;
assign input_1983 = t0_0011110111111;
assign input_1984 = t0_0011111000000;
assign input_1985 = t0_0011111000001;
assign input_1986 = t0_0011111000010;
assign input_1987 = t0_0011111000011;
assign input_1988 = t0_0011111000100;
assign input_1989 = t0_0011111000101;
assign input_1990 = t0_0011111000110;
assign input_1991 = t0_0011111000111;
assign input_1992 = t0_0011111001000;
assign input_1993 = t0_0011111001001;
assign input_1994 = t0_0011111001010;
assign input_1995 = t0_0011111001011;
assign input_1996 = t0_0011111001100;
assign input_1997 = t0_0011111001101;
assign input_1998 = t0_0011111001110;
assign input_1999 = t0_0011111001111;
assign input_2000 = t0_0011111010000;
assign input_2001 = t0_0011111010001;
assign input_2002 = t0_0011111010010;
assign input_2003 = t0_0011111010011;
assign input_2004 = t0_0011111010100;
assign input_2005 = t0_0011111010101;
assign input_2006 = t0_0011111010110;
assign input_2007 = t0_0011111010111;
assign input_2008 = t0_0011111011000;
assign input_2009 = t0_0011111011001;
assign input_2010 = t0_0011111011010;
assign input_2011 = t0_0011111011011;
assign input_2012 = t0_0011111011100;
assign input_2013 = t0_0011111011101;
assign input_2014 = t0_0011111011110;
assign input_2015 = t0_0011111011111;
assign input_2016 = t0_0011111100000;
assign input_2017 = t0_0011111100001;
assign input_2018 = t0_0011111100010;
assign input_2019 = t0_0011111100011;
assign input_2020 = t0_0011111100100;
assign input_2021 = t0_0011111100101;
assign input_2022 = t0_0011111100110;
assign input_2023 = t0_0011111100111;
assign input_2024 = t0_0011111101000;
assign input_2025 = t0_0011111101001;
assign input_2026 = t0_0011111101010;
assign input_2027 = t0_0011111101011;
assign input_2028 = t0_0011111101100;
assign input_2029 = t0_0011111101101;
assign input_2030 = t0_0011111101110;
assign input_2031 = t0_0011111101111;
assign input_2032 = t0_0011111110000;
assign input_2033 = t0_0011111110001;
assign input_2034 = t0_0011111110010;
assign input_2035 = t0_0011111110011;
assign input_2036 = t0_0011111110100;
assign input_2037 = t0_0011111110101;
assign input_2038 = t0_0011111110110;
assign input_2039 = t0_0011111110111;
assign input_2040 = t0_0011111111000;
assign input_2041 = t0_0011111111001;
assign input_2042 = t0_0011111111010;
assign input_2043 = t0_0011111111011;
assign input_2044 = t0_0011111111100;
assign input_2045 = t0_0011111111101;
assign input_2046 = t0_0011111111110;
assign input_2047 = t0_0011111111111;
assign input_2048 = t0_0100000000000;
assign input_2049 = t0_0100000000001;
assign input_2050 = t0_0100000000010;
assign input_2051 = t0_0100000000011;
assign input_2052 = t0_0100000000100;
assign input_2053 = t0_0100000000101;
assign input_2054 = t0_0100000000110;
assign input_2055 = t0_0100000000111;
assign input_2056 = t0_0100000001000;
assign input_2057 = t0_0100000001001;
assign input_2058 = t0_0100000001010;
assign input_2059 = t0_0100000001011;
assign input_2060 = t0_0100000001100;
assign input_2061 = t0_0100000001101;
assign input_2062 = t0_0100000001110;
assign input_2063 = t0_0100000001111;
assign input_2064 = t0_0100000010000;
assign input_2065 = t0_0100000010001;
assign input_2066 = t0_0100000010010;
assign input_2067 = t0_0100000010011;
assign input_2068 = t0_0100000010100;
assign input_2069 = t0_0100000010101;
assign input_2070 = t0_0100000010110;
assign input_2071 = t0_0100000010111;
assign input_2072 = t0_0100000011000;
assign input_2073 = t0_0100000011001;
assign input_2074 = t0_0100000011010;
assign input_2075 = t0_0100000011011;
assign input_2076 = t0_0100000011100;
assign input_2077 = t0_0100000011101;
assign input_2078 = t0_0100000011110;
assign input_2079 = t0_0100000011111;
assign input_2080 = t0_0100000100000;
assign input_2081 = t0_0100000100001;
assign input_2082 = t0_0100000100010;
assign input_2083 = t0_0100000100011;
assign input_2084 = t0_0100000100100;
assign input_2085 = t0_0100000100101;
assign input_2086 = t0_0100000100110;
assign input_2087 = t0_0100000100111;
assign input_2088 = t0_0100000101000;
assign input_2089 = t0_0100000101001;
assign input_2090 = t0_0100000101010;
assign input_2091 = t0_0100000101011;
assign input_2092 = t0_0100000101100;
assign input_2093 = t0_0100000101101;
assign input_2094 = t0_0100000101110;
assign input_2095 = t0_0100000101111;
assign input_2096 = t0_0100000110000;
assign input_2097 = t0_0100000110001;
assign input_2098 = t0_0100000110010;
assign input_2099 = t0_0100000110011;
assign input_2100 = t0_0100000110100;
assign input_2101 = t0_0100000110101;
assign input_2102 = t0_0100000110110;
assign input_2103 = t0_0100000110111;
assign input_2104 = t0_0100000111000;
assign input_2105 = t0_0100000111001;
assign input_2106 = t0_0100000111010;
assign input_2107 = t0_0100000111011;
assign input_2108 = t0_0100000111100;
assign input_2109 = t0_0100000111101;
assign input_2110 = t0_0100000111110;
assign input_2111 = t0_0100000111111;
assign input_2112 = t0_0100001000000;
assign input_2113 = t0_0100001000001;
assign input_2114 = t0_0100001000010;
assign input_2115 = t0_0100001000011;
assign input_2116 = t0_0100001000100;
assign input_2117 = t0_0100001000101;
assign input_2118 = t0_0100001000110;
assign input_2119 = t0_0100001000111;
assign input_2120 = t0_0100001001000;
assign input_2121 = t0_0100001001001;
assign input_2122 = t0_0100001001010;
assign input_2123 = t0_0100001001011;
assign input_2124 = t0_0100001001100;
assign input_2125 = t0_0100001001101;
assign input_2126 = t0_0100001001110;
assign input_2127 = t0_0100001001111;
assign input_2128 = t0_0100001010000;
assign input_2129 = t0_0100001010001;
assign input_2130 = t0_0100001010010;
assign input_2131 = t0_0100001010011;
assign input_2132 = t0_0100001010100;
assign input_2133 = t0_0100001010101;
assign input_2134 = t0_0100001010110;
assign input_2135 = t0_0100001010111;
assign input_2136 = t0_0100001011000;
assign input_2137 = t0_0100001011001;
assign input_2138 = t0_0100001011010;
assign input_2139 = t0_0100001011011;
assign input_2140 = t0_0100001011100;
assign input_2141 = t0_0100001011101;
assign input_2142 = t0_0100001011110;
assign input_2143 = t0_0100001011111;
assign input_2144 = t0_0100001100000;
assign input_2145 = t0_0100001100001;
assign input_2146 = t0_0100001100010;
assign input_2147 = t0_0100001100011;
assign input_2148 = t0_0100001100100;
assign input_2149 = t0_0100001100101;
assign input_2150 = t0_0100001100110;
assign input_2151 = t0_0100001100111;
assign input_2152 = t0_0100001101000;
assign input_2153 = t0_0100001101001;
assign input_2154 = t0_0100001101010;
assign input_2155 = t0_0100001101011;
assign input_2156 = t0_0100001101100;
assign input_2157 = t0_0100001101101;
assign input_2158 = t0_0100001101110;
assign input_2159 = t0_0100001101111;
assign input_2160 = t0_0100001110000;
assign input_2161 = t0_0100001110001;
assign input_2162 = t0_0100001110010;
assign input_2163 = t0_0100001110011;
assign input_2164 = t0_0100001110100;
assign input_2165 = t0_0100001110101;
assign input_2166 = t0_0100001110110;
assign input_2167 = t0_0100001110111;
assign input_2168 = t0_0100001111000;
assign input_2169 = t0_0100001111001;
assign input_2170 = t0_0100001111010;
assign input_2171 = t0_0100001111011;
assign input_2172 = t0_0100001111100;
assign input_2173 = t0_0100001111101;
assign input_2174 = t0_0100001111110;
assign input_2175 = t0_0100001111111;
assign input_2176 = t0_0100010000000;
assign input_2177 = t0_0100010000001;
assign input_2178 = t0_0100010000010;
assign input_2179 = t0_0100010000011;
assign input_2180 = t0_0100010000100;
assign input_2181 = t0_0100010000101;
assign input_2182 = t0_0100010000110;
assign input_2183 = t0_0100010000111;
assign input_2184 = t0_0100010001000;
assign input_2185 = t0_0100010001001;
assign input_2186 = t0_0100010001010;
assign input_2187 = t0_0100010001011;
assign input_2188 = t0_0100010001100;
assign input_2189 = t0_0100010001101;
assign input_2190 = t0_0100010001110;
assign input_2191 = t0_0100010001111;
assign input_2192 = t0_0100010010000;
assign input_2193 = t0_0100010010001;
assign input_2194 = t0_0100010010010;
assign input_2195 = t0_0100010010011;
assign input_2196 = t0_0100010010100;
assign input_2197 = t0_0100010010101;
assign input_2198 = t0_0100010010110;
assign input_2199 = t0_0100010010111;
assign input_2200 = t0_0100010011000;
assign input_2201 = t0_0100010011001;
assign input_2202 = t0_0100010011010;
assign input_2203 = t0_0100010011011;
assign input_2204 = t0_0100010011100;
assign input_2205 = t0_0100010011101;
assign input_2206 = t0_0100010011110;
assign input_2207 = t0_0100010011111;
assign input_2208 = t0_0100010100000;
assign input_2209 = t0_0100010100001;
assign input_2210 = t0_0100010100010;
assign input_2211 = t0_0100010100011;
assign input_2212 = t0_0100010100100;
assign input_2213 = t0_0100010100101;
assign input_2214 = t0_0100010100110;
assign input_2215 = t0_0100010100111;
assign input_2216 = t0_0100010101000;
assign input_2217 = t0_0100010101001;
assign input_2218 = t0_0100010101010;
assign input_2219 = t0_0100010101011;
assign input_2220 = t0_0100010101100;
assign input_2221 = t0_0100010101101;
assign input_2222 = t0_0100010101110;
assign input_2223 = t0_0100010101111;
assign input_2224 = t0_0100010110000;
assign input_2225 = t0_0100010110001;
assign input_2226 = t0_0100010110010;
assign input_2227 = t0_0100010110011;
assign input_2228 = t0_0100010110100;
assign input_2229 = t0_0100010110101;
assign input_2230 = t0_0100010110110;
assign input_2231 = t0_0100010110111;
assign input_2232 = t0_0100010111000;
assign input_2233 = t0_0100010111001;
assign input_2234 = t0_0100010111010;
assign input_2235 = t0_0100010111011;
assign input_2236 = t0_0100010111100;
assign input_2237 = t0_0100010111101;
assign input_2238 = t0_0100010111110;
assign input_2239 = t0_0100010111111;
assign input_2240 = t0_0100011000000;
assign input_2241 = t0_0100011000001;
assign input_2242 = t0_0100011000010;
assign input_2243 = t0_0100011000011;
assign input_2244 = t0_0100011000100;
assign input_2245 = t0_0100011000101;
assign input_2246 = t0_0100011000110;
assign input_2247 = t0_0100011000111;
assign input_2248 = t0_0100011001000;
assign input_2249 = t0_0100011001001;
assign input_2250 = t0_0100011001010;
assign input_2251 = t0_0100011001011;
assign input_2252 = t0_0100011001100;
assign input_2253 = t0_0100011001101;
assign input_2254 = t0_0100011001110;
assign input_2255 = t0_0100011001111;
assign input_2256 = t0_0100011010000;
assign input_2257 = t0_0100011010001;
assign input_2258 = t0_0100011010010;
assign input_2259 = t0_0100011010011;
assign input_2260 = t0_0100011010100;
assign input_2261 = t0_0100011010101;
assign input_2262 = t0_0100011010110;
assign input_2263 = t0_0100011010111;
assign input_2264 = t0_0100011011000;
assign input_2265 = t0_0100011011001;
assign input_2266 = t0_0100011011010;
assign input_2267 = t0_0100011011011;
assign input_2268 = t0_0100011011100;
assign input_2269 = t0_0100011011101;
assign input_2270 = t0_0100011011110;
assign input_2271 = t0_0100011011111;
assign input_2272 = t0_0100011100000;
assign input_2273 = t0_0100011100001;
assign input_2274 = t0_0100011100010;
assign input_2275 = t0_0100011100011;
assign input_2276 = t0_0100011100100;
assign input_2277 = t0_0100011100101;
assign input_2278 = t0_0100011100110;
assign input_2279 = t0_0100011100111;
assign input_2280 = t0_0100011101000;
assign input_2281 = t0_0100011101001;
assign input_2282 = t0_0100011101010;
assign input_2283 = t0_0100011101011;
assign input_2284 = t0_0100011101100;
assign input_2285 = t0_0100011101101;
assign input_2286 = t0_0100011101110;
assign input_2287 = t0_0100011101111;
assign input_2288 = t0_0100011110000;
assign input_2289 = t0_0100011110001;
assign input_2290 = t0_0100011110010;
assign input_2291 = t0_0100011110011;
assign input_2292 = t0_0100011110100;
assign input_2293 = t0_0100011110101;
assign input_2294 = t0_0100011110110;
assign input_2295 = t0_0100011110111;
assign input_2296 = t0_0100011111000;
assign input_2297 = t0_0100011111001;
assign input_2298 = t0_0100011111010;
assign input_2299 = t0_0100011111011;
assign input_2300 = t0_0100011111100;
assign input_2301 = t0_0100011111101;
assign input_2302 = t0_0100011111110;
assign input_2303 = t0_0100011111111;
assign input_2304 = t0_0100100000000;
assign input_2305 = t0_0100100000001;
assign input_2306 = t0_0100100000010;
assign input_2307 = t0_0100100000011;
assign input_2308 = t0_0100100000100;
assign input_2309 = t0_0100100000101;
assign input_2310 = t0_0100100000110;
assign input_2311 = t0_0100100000111;
assign input_2312 = t0_0100100001000;
assign input_2313 = t0_0100100001001;
assign input_2314 = t0_0100100001010;
assign input_2315 = t0_0100100001011;
assign input_2316 = t0_0100100001100;
assign input_2317 = t0_0100100001101;
assign input_2318 = t0_0100100001110;
assign input_2319 = t0_0100100001111;
assign input_2320 = t0_0100100010000;
assign input_2321 = t0_0100100010001;
assign input_2322 = t0_0100100010010;
assign input_2323 = t0_0100100010011;
assign input_2324 = t0_0100100010100;
assign input_2325 = t0_0100100010101;
assign input_2326 = t0_0100100010110;
assign input_2327 = t0_0100100010111;
assign input_2328 = t0_0100100011000;
assign input_2329 = t0_0100100011001;
assign input_2330 = t0_0100100011010;
assign input_2331 = t0_0100100011011;
assign input_2332 = t0_0100100011100;
assign input_2333 = t0_0100100011101;
assign input_2334 = t0_0100100011110;
assign input_2335 = t0_0100100011111;
assign input_2336 = t0_0100100100000;
assign input_2337 = t0_0100100100001;
assign input_2338 = t0_0100100100010;
assign input_2339 = t0_0100100100011;
assign input_2340 = t0_0100100100100;
assign input_2341 = t0_0100100100101;
assign input_2342 = t0_0100100100110;
assign input_2343 = t0_0100100100111;
assign input_2344 = t0_0100100101000;
assign input_2345 = t0_0100100101001;
assign input_2346 = t0_0100100101010;
assign input_2347 = t0_0100100101011;
assign input_2348 = t0_0100100101100;
assign input_2349 = t0_0100100101101;
assign input_2350 = t0_0100100101110;
assign input_2351 = t0_0100100101111;
assign input_2352 = t0_0100100110000;
assign input_2353 = t0_0100100110001;
assign input_2354 = t0_0100100110010;
assign input_2355 = t0_0100100110011;
assign input_2356 = t0_0100100110100;
assign input_2357 = t0_0100100110101;
assign input_2358 = t0_0100100110110;
assign input_2359 = t0_0100100110111;
assign input_2360 = t0_0100100111000;
assign input_2361 = t0_0100100111001;
assign input_2362 = t0_0100100111010;
assign input_2363 = t0_0100100111011;
assign input_2364 = t0_0100100111100;
assign input_2365 = t0_0100100111101;
assign input_2366 = t0_0100100111110;
assign input_2367 = t0_0100100111111;
assign input_2368 = t0_0100101000000;
assign input_2369 = t0_0100101000001;
assign input_2370 = t0_0100101000010;
assign input_2371 = t0_0100101000011;
assign input_2372 = t0_0100101000100;
assign input_2373 = t0_0100101000101;
assign input_2374 = t0_0100101000110;
assign input_2375 = t0_0100101000111;
assign input_2376 = t0_0100101001000;
assign input_2377 = t0_0100101001001;
assign input_2378 = t0_0100101001010;
assign input_2379 = t0_0100101001011;
assign input_2380 = t0_0100101001100;
assign input_2381 = t0_0100101001101;
assign input_2382 = t0_0100101001110;
assign input_2383 = t0_0100101001111;
assign input_2384 = t0_0100101010000;
assign input_2385 = t0_0100101010001;
assign input_2386 = t0_0100101010010;
assign input_2387 = t0_0100101010011;
assign input_2388 = t0_0100101010100;
assign input_2389 = t0_0100101010101;
assign input_2390 = t0_0100101010110;
assign input_2391 = t0_0100101010111;
assign input_2392 = t0_0100101011000;
assign input_2393 = t0_0100101011001;
assign input_2394 = t0_0100101011010;
assign input_2395 = t0_0100101011011;
assign input_2396 = t0_0100101011100;
assign input_2397 = t0_0100101011101;
assign input_2398 = t0_0100101011110;
assign input_2399 = t0_0100101011111;
assign input_2400 = t0_0100101100000;
assign input_2401 = t0_0100101100001;
assign input_2402 = t0_0100101100010;
assign input_2403 = t0_0100101100011;
assign input_2404 = t0_0100101100100;
assign input_2405 = t0_0100101100101;
assign input_2406 = t0_0100101100110;
assign input_2407 = t0_0100101100111;
assign input_2408 = t0_0100101101000;
assign input_2409 = t0_0100101101001;
assign input_2410 = t0_0100101101010;
assign input_2411 = t0_0100101101011;
assign input_2412 = t0_0100101101100;
assign input_2413 = t0_0100101101101;
assign input_2414 = t0_0100101101110;
assign input_2415 = t0_0100101101111;
assign input_2416 = t0_0100101110000;
assign input_2417 = t0_0100101110001;
assign input_2418 = t0_0100101110010;
assign input_2419 = t0_0100101110011;
assign input_2420 = t0_0100101110100;
assign input_2421 = t0_0100101110101;
assign input_2422 = t0_0100101110110;
assign input_2423 = t0_0100101110111;
assign input_2424 = t0_0100101111000;
assign input_2425 = t0_0100101111001;
assign input_2426 = t0_0100101111010;
assign input_2427 = t0_0100101111011;
assign input_2428 = t0_0100101111100;
assign input_2429 = t0_0100101111101;
assign input_2430 = t0_0100101111110;
assign input_2431 = t0_0100101111111;
assign input_2432 = t0_0100110000000;
assign input_2433 = t0_0100110000001;
assign input_2434 = t0_0100110000010;
assign input_2435 = t0_0100110000011;
assign input_2436 = t0_0100110000100;
assign input_2437 = t0_0100110000101;
assign input_2438 = t0_0100110000110;
assign input_2439 = t0_0100110000111;
assign input_2440 = t0_0100110001000;
assign input_2441 = t0_0100110001001;
assign input_2442 = t0_0100110001010;
assign input_2443 = t0_0100110001011;
assign input_2444 = t0_0100110001100;
assign input_2445 = t0_0100110001101;
assign input_2446 = t0_0100110001110;
assign input_2447 = t0_0100110001111;
assign input_2448 = t0_0100110010000;
assign input_2449 = t0_0100110010001;
assign input_2450 = t0_0100110010010;
assign input_2451 = t0_0100110010011;
assign input_2452 = t0_0100110010100;
assign input_2453 = t0_0100110010101;
assign input_2454 = t0_0100110010110;
assign input_2455 = t0_0100110010111;
assign input_2456 = t0_0100110011000;
assign input_2457 = t0_0100110011001;
assign input_2458 = t0_0100110011010;
assign input_2459 = t0_0100110011011;
assign input_2460 = t0_0100110011100;
assign input_2461 = t0_0100110011101;
assign input_2462 = t0_0100110011110;
assign input_2463 = t0_0100110011111;
assign input_2464 = t0_0100110100000;
assign input_2465 = t0_0100110100001;
assign input_2466 = t0_0100110100010;
assign input_2467 = t0_0100110100011;
assign input_2468 = t0_0100110100100;
assign input_2469 = t0_0100110100101;
assign input_2470 = t0_0100110100110;
assign input_2471 = t0_0100110100111;
assign input_2472 = t0_0100110101000;
assign input_2473 = t0_0100110101001;
assign input_2474 = t0_0100110101010;
assign input_2475 = t0_0100110101011;
assign input_2476 = t0_0100110101100;
assign input_2477 = t0_0100110101101;
assign input_2478 = t0_0100110101110;
assign input_2479 = t0_0100110101111;
assign input_2480 = t0_0100110110000;
assign input_2481 = t0_0100110110001;
assign input_2482 = t0_0100110110010;
assign input_2483 = t0_0100110110011;
assign input_2484 = t0_0100110110100;
assign input_2485 = t0_0100110110101;
assign input_2486 = t0_0100110110110;
assign input_2487 = t0_0100110110111;
assign input_2488 = t0_0100110111000;
assign input_2489 = t0_0100110111001;
assign input_2490 = t0_0100110111010;
assign input_2491 = t0_0100110111011;
assign input_2492 = t0_0100110111100;
assign input_2493 = t0_0100110111101;
assign input_2494 = t0_0100110111110;
assign input_2495 = t0_0100110111111;
assign input_2496 = t0_0100111000000;
assign input_2497 = t0_0100111000001;
assign input_2498 = t0_0100111000010;
assign input_2499 = t0_0100111000011;
assign input_2500 = t0_0100111000100;
assign input_2501 = t0_0100111000101;
assign input_2502 = t0_0100111000110;
assign input_2503 = t0_0100111000111;
assign input_2504 = t0_0100111001000;
assign input_2505 = t0_0100111001001;
assign input_2506 = t0_0100111001010;
assign input_2507 = t0_0100111001011;
assign input_2508 = t0_0100111001100;
assign input_2509 = t0_0100111001101;
assign input_2510 = t0_0100111001110;
assign input_2511 = t0_0100111001111;
assign input_2512 = t0_0100111010000;
assign input_2513 = t0_0100111010001;
assign input_2514 = t0_0100111010010;
assign input_2515 = t0_0100111010011;
assign input_2516 = t0_0100111010100;
assign input_2517 = t0_0100111010101;
assign input_2518 = t0_0100111010110;
assign input_2519 = t0_0100111010111;
assign input_2520 = t0_0100111011000;
assign input_2521 = t0_0100111011001;
assign input_2522 = t0_0100111011010;
assign input_2523 = t0_0100111011011;
assign input_2524 = t0_0100111011100;
assign input_2525 = t0_0100111011101;
assign input_2526 = t0_0100111011110;
assign input_2527 = t0_0100111011111;
assign input_2528 = t0_0100111100000;
assign input_2529 = t0_0100111100001;
assign input_2530 = t0_0100111100010;
assign input_2531 = t0_0100111100011;
assign input_2532 = t0_0100111100100;
assign input_2533 = t0_0100111100101;
assign input_2534 = t0_0100111100110;
assign input_2535 = t0_0100111100111;
assign input_2536 = t0_0100111101000;
assign input_2537 = t0_0100111101001;
assign input_2538 = t0_0100111101010;
assign input_2539 = t0_0100111101011;
assign input_2540 = t0_0100111101100;
assign input_2541 = t0_0100111101101;
assign input_2542 = t0_0100111101110;
assign input_2543 = t0_0100111101111;
assign input_2544 = t0_0100111110000;
assign input_2545 = t0_0100111110001;
assign input_2546 = t0_0100111110010;
assign input_2547 = t0_0100111110011;
assign input_2548 = t0_0100111110100;
assign input_2549 = t0_0100111110101;
assign input_2550 = t0_0100111110110;
assign input_2551 = t0_0100111110111;
assign input_2552 = t0_0100111111000;
assign input_2553 = t0_0100111111001;
assign input_2554 = t0_0100111111010;
assign input_2555 = t0_0100111111011;
assign input_2556 = t0_0100111111100;
assign input_2557 = t0_0100111111101;
assign input_2558 = t0_0100111111110;
assign input_2559 = t0_0100111111111;
assign input_2560 = t0_0101000000000;
assign input_2561 = t0_0101000000001;
assign input_2562 = t0_0101000000010;
assign input_2563 = t0_0101000000011;
assign input_2564 = t0_0101000000100;
assign input_2565 = t0_0101000000101;
assign input_2566 = t0_0101000000110;
assign input_2567 = t0_0101000000111;
assign input_2568 = t0_0101000001000;
assign input_2569 = t0_0101000001001;
assign input_2570 = t0_0101000001010;
assign input_2571 = t0_0101000001011;
assign input_2572 = t0_0101000001100;
assign input_2573 = t0_0101000001101;
assign input_2574 = t0_0101000001110;
assign input_2575 = t0_0101000001111;
assign input_2576 = t0_0101000010000;
assign input_2577 = t0_0101000010001;
assign input_2578 = t0_0101000010010;
assign input_2579 = t0_0101000010011;
assign input_2580 = t0_0101000010100;
assign input_2581 = t0_0101000010101;
assign input_2582 = t0_0101000010110;
assign input_2583 = t0_0101000010111;
assign input_2584 = t0_0101000011000;
assign input_2585 = t0_0101000011001;
assign input_2586 = t0_0101000011010;
assign input_2587 = t0_0101000011011;
assign input_2588 = t0_0101000011100;
assign input_2589 = t0_0101000011101;
assign input_2590 = t0_0101000011110;
assign input_2591 = t0_0101000011111;
assign input_2592 = t0_0101000100000;
assign input_2593 = t0_0101000100001;
assign input_2594 = t0_0101000100010;
assign input_2595 = t0_0101000100011;
assign input_2596 = t0_0101000100100;
assign input_2597 = t0_0101000100101;
assign input_2598 = t0_0101000100110;
assign input_2599 = t0_0101000100111;
assign input_2600 = t0_0101000101000;
assign input_2601 = t0_0101000101001;
assign input_2602 = t0_0101000101010;
assign input_2603 = t0_0101000101011;
assign input_2604 = t0_0101000101100;
assign input_2605 = t0_0101000101101;
assign input_2606 = t0_0101000101110;
assign input_2607 = t0_0101000101111;
assign input_2608 = t0_0101000110000;
assign input_2609 = t0_0101000110001;
assign input_2610 = t0_0101000110010;
assign input_2611 = t0_0101000110011;
assign input_2612 = t0_0101000110100;
assign input_2613 = t0_0101000110101;
assign input_2614 = t0_0101000110110;
assign input_2615 = t0_0101000110111;
assign input_2616 = t0_0101000111000;
assign input_2617 = t0_0101000111001;
assign input_2618 = t0_0101000111010;
assign input_2619 = t0_0101000111011;
assign input_2620 = t0_0101000111100;
assign input_2621 = t0_0101000111101;
assign input_2622 = t0_0101000111110;
assign input_2623 = t0_0101000111111;
assign input_2624 = t0_0101001000000;
assign input_2625 = t0_0101001000001;
assign input_2626 = t0_0101001000010;
assign input_2627 = t0_0101001000011;
assign input_2628 = t0_0101001000100;
assign input_2629 = t0_0101001000101;
assign input_2630 = t0_0101001000110;
assign input_2631 = t0_0101001000111;
assign input_2632 = t0_0101001001000;
assign input_2633 = t0_0101001001001;
assign input_2634 = t0_0101001001010;
assign input_2635 = t0_0101001001011;
assign input_2636 = t0_0101001001100;
assign input_2637 = t0_0101001001101;
assign input_2638 = t0_0101001001110;
assign input_2639 = t0_0101001001111;
assign input_2640 = t0_0101001010000;
assign input_2641 = t0_0101001010001;
assign input_2642 = t0_0101001010010;
assign input_2643 = t0_0101001010011;
assign input_2644 = t0_0101001010100;
assign input_2645 = t0_0101001010101;
assign input_2646 = t0_0101001010110;
assign input_2647 = t0_0101001010111;
assign input_2648 = t0_0101001011000;
assign input_2649 = t0_0101001011001;
assign input_2650 = t0_0101001011010;
assign input_2651 = t0_0101001011011;
assign input_2652 = t0_0101001011100;
assign input_2653 = t0_0101001011101;
assign input_2654 = t0_0101001011110;
assign input_2655 = t0_0101001011111;
assign input_2656 = t0_0101001100000;
assign input_2657 = t0_0101001100001;
assign input_2658 = t0_0101001100010;
assign input_2659 = t0_0101001100011;
assign input_2660 = t0_0101001100100;
assign input_2661 = t0_0101001100101;
assign input_2662 = t0_0101001100110;
assign input_2663 = t0_0101001100111;
assign input_2664 = t0_0101001101000;
assign input_2665 = t0_0101001101001;
assign input_2666 = t0_0101001101010;
assign input_2667 = t0_0101001101011;
assign input_2668 = t0_0101001101100;
assign input_2669 = t0_0101001101101;
assign input_2670 = t0_0101001101110;
assign input_2671 = t0_0101001101111;
assign input_2672 = t0_0101001110000;
assign input_2673 = t0_0101001110001;
assign input_2674 = t0_0101001110010;
assign input_2675 = t0_0101001110011;
assign input_2676 = t0_0101001110100;
assign input_2677 = t0_0101001110101;
assign input_2678 = t0_0101001110110;
assign input_2679 = t0_0101001110111;
assign input_2680 = t0_0101001111000;
assign input_2681 = t0_0101001111001;
assign input_2682 = t0_0101001111010;
assign input_2683 = t0_0101001111011;
assign input_2684 = t0_0101001111100;
assign input_2685 = t0_0101001111101;
assign input_2686 = t0_0101001111110;
assign input_2687 = t0_0101001111111;
assign input_2688 = t0_0101010000000;
assign input_2689 = t0_0101010000001;
assign input_2690 = t0_0101010000010;
assign input_2691 = t0_0101010000011;
assign input_2692 = t0_0101010000100;
assign input_2693 = t0_0101010000101;
assign input_2694 = t0_0101010000110;
assign input_2695 = t0_0101010000111;
assign input_2696 = t0_0101010001000;
assign input_2697 = t0_0101010001001;
assign input_2698 = t0_0101010001010;
assign input_2699 = t0_0101010001011;
assign input_2700 = t0_0101010001100;
assign input_2701 = t0_0101010001101;
assign input_2702 = t0_0101010001110;
assign input_2703 = t0_0101010001111;
assign input_2704 = t0_0101010010000;
assign input_2705 = t0_0101010010001;
assign input_2706 = t0_0101010010010;
assign input_2707 = t0_0101010010011;
assign input_2708 = t0_0101010010100;
assign input_2709 = t0_0101010010101;
assign input_2710 = t0_0101010010110;
assign input_2711 = t0_0101010010111;
assign input_2712 = t0_0101010011000;
assign input_2713 = t0_0101010011001;
assign input_2714 = t0_0101010011010;
assign input_2715 = t0_0101010011011;
assign input_2716 = t0_0101010011100;
assign input_2717 = t0_0101010011101;
assign input_2718 = t0_0101010011110;
assign input_2719 = t0_0101010011111;
assign input_2720 = t0_0101010100000;
assign input_2721 = t0_0101010100001;
assign input_2722 = t0_0101010100010;
assign input_2723 = t0_0101010100011;
assign input_2724 = t0_0101010100100;
assign input_2725 = t0_0101010100101;
assign input_2726 = t0_0101010100110;
assign input_2727 = t0_0101010100111;
assign input_2728 = t0_0101010101000;
assign input_2729 = t0_0101010101001;
assign input_2730 = t0_0101010101010;
assign input_2731 = t0_0101010101011;
assign input_2732 = t0_0101010101100;
assign input_2733 = t0_0101010101101;
assign input_2734 = t0_0101010101110;
assign input_2735 = t0_0101010101111;
assign input_2736 = t0_0101010110000;
assign input_2737 = t0_0101010110001;
assign input_2738 = t0_0101010110010;
assign input_2739 = t0_0101010110011;
assign input_2740 = t0_0101010110100;
assign input_2741 = t0_0101010110101;
assign input_2742 = t0_0101010110110;
assign input_2743 = t0_0101010110111;
assign input_2744 = t0_0101010111000;
assign input_2745 = t0_0101010111001;
assign input_2746 = t0_0101010111010;
assign input_2747 = t0_0101010111011;
assign input_2748 = t0_0101010111100;
assign input_2749 = t0_0101010111101;
assign input_2750 = t0_0101010111110;
assign input_2751 = t0_0101010111111;
assign input_2752 = t0_0101011000000;
assign input_2753 = t0_0101011000001;
assign input_2754 = t0_0101011000010;
assign input_2755 = t0_0101011000011;
assign input_2756 = t0_0101011000100;
assign input_2757 = t0_0101011000101;
assign input_2758 = t0_0101011000110;
assign input_2759 = t0_0101011000111;
assign input_2760 = t0_0101011001000;
assign input_2761 = t0_0101011001001;
assign input_2762 = t0_0101011001010;
assign input_2763 = t0_0101011001011;
assign input_2764 = t0_0101011001100;
assign input_2765 = t0_0101011001101;
assign input_2766 = t0_0101011001110;
assign input_2767 = t0_0101011001111;
assign input_2768 = t0_0101011010000;
assign input_2769 = t0_0101011010001;
assign input_2770 = t0_0101011010010;
assign input_2771 = t0_0101011010011;
assign input_2772 = t0_0101011010100;
assign input_2773 = t0_0101011010101;
assign input_2774 = t0_0101011010110;
assign input_2775 = t0_0101011010111;
assign input_2776 = t0_0101011011000;
assign input_2777 = t0_0101011011001;
assign input_2778 = t0_0101011011010;
assign input_2779 = t0_0101011011011;
assign input_2780 = t0_0101011011100;
assign input_2781 = t0_0101011011101;
assign input_2782 = t0_0101011011110;
assign input_2783 = t0_0101011011111;
assign input_2784 = t0_0101011100000;
assign input_2785 = t0_0101011100001;
assign input_2786 = t0_0101011100010;
assign input_2787 = t0_0101011100011;
assign input_2788 = t0_0101011100100;
assign input_2789 = t0_0101011100101;
assign input_2790 = t0_0101011100110;
assign input_2791 = t0_0101011100111;
assign input_2792 = t0_0101011101000;
assign input_2793 = t0_0101011101001;
assign input_2794 = t0_0101011101010;
assign input_2795 = t0_0101011101011;
assign input_2796 = t0_0101011101100;
assign input_2797 = t0_0101011101101;
assign input_2798 = t0_0101011101110;
assign input_2799 = t0_0101011101111;
assign input_2800 = t0_0101011110000;
assign input_2801 = t0_0101011110001;
assign input_2802 = t0_0101011110010;
assign input_2803 = t0_0101011110011;
assign input_2804 = t0_0101011110100;
assign input_2805 = t0_0101011110101;
assign input_2806 = t0_0101011110110;
assign input_2807 = t0_0101011110111;
assign input_2808 = t0_0101011111000;
assign input_2809 = t0_0101011111001;
assign input_2810 = t0_0101011111010;
assign input_2811 = t0_0101011111011;
assign input_2812 = t0_0101011111100;
assign input_2813 = t0_0101011111101;
assign input_2814 = t0_0101011111110;
assign input_2815 = t0_0101011111111;
assign input_2816 = t0_0101100000000;
assign input_2817 = t0_0101100000001;
assign input_2818 = t0_0101100000010;
assign input_2819 = t0_0101100000011;
assign input_2820 = t0_0101100000100;
assign input_2821 = t0_0101100000101;
assign input_2822 = t0_0101100000110;
assign input_2823 = t0_0101100000111;
assign input_2824 = t0_0101100001000;
assign input_2825 = t0_0101100001001;
assign input_2826 = t0_0101100001010;
assign input_2827 = t0_0101100001011;
assign input_2828 = t0_0101100001100;
assign input_2829 = t0_0101100001101;
assign input_2830 = t0_0101100001110;
assign input_2831 = t0_0101100001111;
assign input_2832 = t0_0101100010000;
assign input_2833 = t0_0101100010001;
assign input_2834 = t0_0101100010010;
assign input_2835 = t0_0101100010011;
assign input_2836 = t0_0101100010100;
assign input_2837 = t0_0101100010101;
assign input_2838 = t0_0101100010110;
assign input_2839 = t0_0101100010111;
assign input_2840 = t0_0101100011000;
assign input_2841 = t0_0101100011001;
assign input_2842 = t0_0101100011010;
assign input_2843 = t0_0101100011011;
assign input_2844 = t0_0101100011100;
assign input_2845 = t0_0101100011101;
assign input_2846 = t0_0101100011110;
assign input_2847 = t0_0101100011111;
assign input_2848 = t0_0101100100000;
assign input_2849 = t0_0101100100001;
assign input_2850 = t0_0101100100010;
assign input_2851 = t0_0101100100011;
assign input_2852 = t0_0101100100100;
assign input_2853 = t0_0101100100101;
assign input_2854 = t0_0101100100110;
assign input_2855 = t0_0101100100111;
assign input_2856 = t0_0101100101000;
assign input_2857 = t0_0101100101001;
assign input_2858 = t0_0101100101010;
assign input_2859 = t0_0101100101011;
assign input_2860 = t0_0101100101100;
assign input_2861 = t0_0101100101101;
assign input_2862 = t0_0101100101110;
assign input_2863 = t0_0101100101111;
assign input_2864 = t0_0101100110000;
assign input_2865 = t0_0101100110001;
assign input_2866 = t0_0101100110010;
assign input_2867 = t0_0101100110011;
assign input_2868 = t0_0101100110100;
assign input_2869 = t0_0101100110101;
assign input_2870 = t0_0101100110110;
assign input_2871 = t0_0101100110111;
assign input_2872 = t0_0101100111000;
assign input_2873 = t0_0101100111001;
assign input_2874 = t0_0101100111010;
assign input_2875 = t0_0101100111011;
assign input_2876 = t0_0101100111100;
assign input_2877 = t0_0101100111101;
assign input_2878 = t0_0101100111110;
assign input_2879 = t0_0101100111111;
assign input_2880 = t0_0101101000000;
assign input_2881 = t0_0101101000001;
assign input_2882 = t0_0101101000010;
assign input_2883 = t0_0101101000011;
assign input_2884 = t0_0101101000100;
assign input_2885 = t0_0101101000101;
assign input_2886 = t0_0101101000110;
assign input_2887 = t0_0101101000111;
assign input_2888 = t0_0101101001000;
assign input_2889 = t0_0101101001001;
assign input_2890 = t0_0101101001010;
assign input_2891 = t0_0101101001011;
assign input_2892 = t0_0101101001100;
assign input_2893 = t0_0101101001101;
assign input_2894 = t0_0101101001110;
assign input_2895 = t0_0101101001111;
assign input_2896 = t0_0101101010000;
assign input_2897 = t0_0101101010001;
assign input_2898 = t0_0101101010010;
assign input_2899 = t0_0101101010011;
assign input_2900 = t0_0101101010100;
assign input_2901 = t0_0101101010101;
assign input_2902 = t0_0101101010110;
assign input_2903 = t0_0101101010111;
assign input_2904 = t0_0101101011000;
assign input_2905 = t0_0101101011001;
assign input_2906 = t0_0101101011010;
assign input_2907 = t0_0101101011011;
assign input_2908 = t0_0101101011100;
assign input_2909 = t0_0101101011101;
assign input_2910 = t0_0101101011110;
assign input_2911 = t0_0101101011111;
assign input_2912 = t0_0101101100000;
assign input_2913 = t0_0101101100001;
assign input_2914 = t0_0101101100010;
assign input_2915 = t0_0101101100011;
assign input_2916 = t0_0101101100100;
assign input_2917 = t0_0101101100101;
assign input_2918 = t0_0101101100110;
assign input_2919 = t0_0101101100111;
assign input_2920 = t0_0101101101000;
assign input_2921 = t0_0101101101001;
assign input_2922 = t0_0101101101010;
assign input_2923 = t0_0101101101011;
assign input_2924 = t0_0101101101100;
assign input_2925 = t0_0101101101101;
assign input_2926 = t0_0101101101110;
assign input_2927 = t0_0101101101111;
assign input_2928 = t0_0101101110000;
assign input_2929 = t0_0101101110001;
assign input_2930 = t0_0101101110010;
assign input_2931 = t0_0101101110011;
assign input_2932 = t0_0101101110100;
assign input_2933 = t0_0101101110101;
assign input_2934 = t0_0101101110110;
assign input_2935 = t0_0101101110111;
assign input_2936 = t0_0101101111000;
assign input_2937 = t0_0101101111001;
assign input_2938 = t0_0101101111010;
assign input_2939 = t0_0101101111011;
assign input_2940 = t0_0101101111100;
assign input_2941 = t0_0101101111101;
assign input_2942 = t0_0101101111110;
assign input_2943 = t0_0101101111111;
assign input_2944 = t0_0101110000000;
assign input_2945 = t0_0101110000001;
assign input_2946 = t0_0101110000010;
assign input_2947 = t0_0101110000011;
assign input_2948 = t0_0101110000100;
assign input_2949 = t0_0101110000101;
assign input_2950 = t0_0101110000110;
assign input_2951 = t0_0101110000111;
assign input_2952 = t0_0101110001000;
assign input_2953 = t0_0101110001001;
assign input_2954 = t0_0101110001010;
assign input_2955 = t0_0101110001011;
assign input_2956 = t0_0101110001100;
assign input_2957 = t0_0101110001101;
assign input_2958 = t0_0101110001110;
assign input_2959 = t0_0101110001111;
assign input_2960 = t0_0101110010000;
assign input_2961 = t0_0101110010001;
assign input_2962 = t0_0101110010010;
assign input_2963 = t0_0101110010011;
assign input_2964 = t0_0101110010100;
assign input_2965 = t0_0101110010101;
assign input_2966 = t0_0101110010110;
assign input_2967 = t0_0101110010111;
assign input_2968 = t0_0101110011000;
assign input_2969 = t0_0101110011001;
assign input_2970 = t0_0101110011010;
assign input_2971 = t0_0101110011011;
assign input_2972 = t0_0101110011100;
assign input_2973 = t0_0101110011101;
assign input_2974 = t0_0101110011110;
assign input_2975 = t0_0101110011111;
assign input_2976 = t0_0101110100000;
assign input_2977 = t0_0101110100001;
assign input_2978 = t0_0101110100010;
assign input_2979 = t0_0101110100011;
assign input_2980 = t0_0101110100100;
assign input_2981 = t0_0101110100101;
assign input_2982 = t0_0101110100110;
assign input_2983 = t0_0101110100111;
assign input_2984 = t0_0101110101000;
assign input_2985 = t0_0101110101001;
assign input_2986 = t0_0101110101010;
assign input_2987 = t0_0101110101011;
assign input_2988 = t0_0101110101100;
assign input_2989 = t0_0101110101101;
assign input_2990 = t0_0101110101110;
assign input_2991 = t0_0101110101111;
assign input_2992 = t0_0101110110000;
assign input_2993 = t0_0101110110001;
assign input_2994 = t0_0101110110010;
assign input_2995 = t0_0101110110011;
assign input_2996 = t0_0101110110100;
assign input_2997 = t0_0101110110101;
assign input_2998 = t0_0101110110110;
assign input_2999 = t0_0101110110111;
assign input_3000 = t0_0101110111000;
assign input_3001 = t0_0101110111001;
assign input_3002 = t0_0101110111010;
assign input_3003 = t0_0101110111011;
assign input_3004 = t0_0101110111100;
assign input_3005 = t0_0101110111101;
assign input_3006 = t0_0101110111110;
assign input_3007 = t0_0101110111111;
assign input_3008 = t0_0101111000000;
assign input_3009 = t0_0101111000001;
assign input_3010 = t0_0101111000010;
assign input_3011 = t0_0101111000011;
assign input_3012 = t0_0101111000100;
assign input_3013 = t0_0101111000101;
assign input_3014 = t0_0101111000110;
assign input_3015 = t0_0101111000111;
assign input_3016 = t0_0101111001000;
assign input_3017 = t0_0101111001001;
assign input_3018 = t0_0101111001010;
assign input_3019 = t0_0101111001011;
assign input_3020 = t0_0101111001100;
assign input_3021 = t0_0101111001101;
assign input_3022 = t0_0101111001110;
assign input_3023 = t0_0101111001111;
assign input_3024 = t0_0101111010000;
assign input_3025 = t0_0101111010001;
assign input_3026 = t0_0101111010010;
assign input_3027 = t0_0101111010011;
assign input_3028 = t0_0101111010100;
assign input_3029 = t0_0101111010101;
assign input_3030 = t0_0101111010110;
assign input_3031 = t0_0101111010111;
assign input_3032 = t0_0101111011000;
assign input_3033 = t0_0101111011001;
assign input_3034 = t0_0101111011010;
assign input_3035 = t0_0101111011011;
assign input_3036 = t0_0101111011100;
assign input_3037 = t0_0101111011101;
assign input_3038 = t0_0101111011110;
assign input_3039 = t0_0101111011111;
assign input_3040 = t0_0101111100000;
assign input_3041 = t0_0101111100001;
assign input_3042 = t0_0101111100010;
assign input_3043 = t0_0101111100011;
assign input_3044 = t0_0101111100100;
assign input_3045 = t0_0101111100101;
assign input_3046 = t0_0101111100110;
assign input_3047 = t0_0101111100111;
assign input_3048 = t0_0101111101000;
assign input_3049 = t0_0101111101001;
assign input_3050 = t0_0101111101010;
assign input_3051 = t0_0101111101011;
assign input_3052 = t0_0101111101100;
assign input_3053 = t0_0101111101101;
assign input_3054 = t0_0101111101110;
assign input_3055 = t0_0101111101111;
assign input_3056 = t0_0101111110000;
assign input_3057 = t0_0101111110001;
assign input_3058 = t0_0101111110010;
assign input_3059 = t0_0101111110011;
assign input_3060 = t0_0101111110100;
assign input_3061 = t0_0101111110101;
assign input_3062 = t0_0101111110110;
assign input_3063 = t0_0101111110111;
assign input_3064 = t0_0101111111000;
assign input_3065 = t0_0101111111001;
assign input_3066 = t0_0101111111010;
assign input_3067 = t0_0101111111011;
assign input_3068 = t0_0101111111100;
assign input_3069 = t0_0101111111101;
assign input_3070 = t0_0101111111110;
assign input_3071 = t0_0101111111111;
assign input_3072 = t0_0110000000000;
assign input_3073 = t0_0110000000001;
assign input_3074 = t0_0110000000010;
assign input_3075 = t0_0110000000011;
assign input_3076 = t0_0110000000100;
assign input_3077 = t0_0110000000101;
assign input_3078 = t0_0110000000110;
assign input_3079 = t0_0110000000111;
assign input_3080 = t0_0110000001000;
assign input_3081 = t0_0110000001001;
assign input_3082 = t0_0110000001010;
assign input_3083 = t0_0110000001011;
assign input_3084 = t0_0110000001100;
assign input_3085 = t0_0110000001101;
assign input_3086 = t0_0110000001110;
assign input_3087 = t0_0110000001111;
assign input_3088 = t0_0110000010000;
assign input_3089 = t0_0110000010001;
assign input_3090 = t0_0110000010010;
assign input_3091 = t0_0110000010011;
assign input_3092 = t0_0110000010100;
assign input_3093 = t0_0110000010101;
assign input_3094 = t0_0110000010110;
assign input_3095 = t0_0110000010111;
assign input_3096 = t0_0110000011000;
assign input_3097 = t0_0110000011001;
assign input_3098 = t0_0110000011010;
assign input_3099 = t0_0110000011011;
assign input_3100 = t0_0110000011100;
assign input_3101 = t0_0110000011101;
assign input_3102 = t0_0110000011110;
assign input_3103 = t0_0110000011111;
assign input_3104 = t0_0110000100000;
assign input_3105 = t0_0110000100001;
assign input_3106 = t0_0110000100010;
assign input_3107 = t0_0110000100011;
assign input_3108 = t0_0110000100100;
assign input_3109 = t0_0110000100101;
assign input_3110 = t0_0110000100110;
assign input_3111 = t0_0110000100111;
assign input_3112 = t0_0110000101000;
assign input_3113 = t0_0110000101001;
assign input_3114 = t0_0110000101010;
assign input_3115 = t0_0110000101011;
assign input_3116 = t0_0110000101100;
assign input_3117 = t0_0110000101101;
assign input_3118 = t0_0110000101110;
assign input_3119 = t0_0110000101111;
assign input_3120 = t0_0110000110000;
assign input_3121 = t0_0110000110001;
assign input_3122 = t0_0110000110010;
assign input_3123 = t0_0110000110011;
assign input_3124 = t0_0110000110100;
assign input_3125 = t0_0110000110101;
assign input_3126 = t0_0110000110110;
assign input_3127 = t0_0110000110111;
assign input_3128 = t0_0110000111000;
assign input_3129 = t0_0110000111001;
assign input_3130 = t0_0110000111010;
assign input_3131 = t0_0110000111011;
assign input_3132 = t0_0110000111100;
assign input_3133 = t0_0110000111101;
assign input_3134 = t0_0110000111110;
assign input_3135 = t0_0110000111111;
assign input_3136 = t0_0110001000000;
assign input_3137 = t0_0110001000001;
assign input_3138 = t0_0110001000010;
assign input_3139 = t0_0110001000011;
assign input_3140 = t0_0110001000100;
assign input_3141 = t0_0110001000101;
assign input_3142 = t0_0110001000110;
assign input_3143 = t0_0110001000111;
assign input_3144 = t0_0110001001000;
assign input_3145 = t0_0110001001001;
assign input_3146 = t0_0110001001010;
assign input_3147 = t0_0110001001011;
assign input_3148 = t0_0110001001100;
assign input_3149 = t0_0110001001101;
assign input_3150 = t0_0110001001110;
assign input_3151 = t0_0110001001111;
assign input_3152 = t0_0110001010000;
assign input_3153 = t0_0110001010001;
assign input_3154 = t0_0110001010010;
assign input_3155 = t0_0110001010011;
assign input_3156 = t0_0110001010100;
assign input_3157 = t0_0110001010101;
assign input_3158 = t0_0110001010110;
assign input_3159 = t0_0110001010111;
assign input_3160 = t0_0110001011000;
assign input_3161 = t0_0110001011001;
assign input_3162 = t0_0110001011010;
assign input_3163 = t0_0110001011011;
assign input_3164 = t0_0110001011100;
assign input_3165 = t0_0110001011101;
assign input_3166 = t0_0110001011110;
assign input_3167 = t0_0110001011111;
assign input_3168 = t0_0110001100000;
assign input_3169 = t0_0110001100001;
assign input_3170 = t0_0110001100010;
assign input_3171 = t0_0110001100011;
assign input_3172 = t0_0110001100100;
assign input_3173 = t0_0110001100101;
assign input_3174 = t0_0110001100110;
assign input_3175 = t0_0110001100111;
assign input_3176 = t0_0110001101000;
assign input_3177 = t0_0110001101001;
assign input_3178 = t0_0110001101010;
assign input_3179 = t0_0110001101011;
assign input_3180 = t0_0110001101100;
assign input_3181 = t0_0110001101101;
assign input_3182 = t0_0110001101110;
assign input_3183 = t0_0110001101111;
assign input_3184 = t0_0110001110000;
assign input_3185 = t0_0110001110001;
assign input_3186 = t0_0110001110010;
assign input_3187 = t0_0110001110011;
assign input_3188 = t0_0110001110100;
assign input_3189 = t0_0110001110101;
assign input_3190 = t0_0110001110110;
assign input_3191 = t0_0110001110111;
assign input_3192 = t0_0110001111000;
assign input_3193 = t0_0110001111001;
assign input_3194 = t0_0110001111010;
assign input_3195 = t0_0110001111011;
assign input_3196 = t0_0110001111100;
assign input_3197 = t0_0110001111101;
assign input_3198 = t0_0110001111110;
assign input_3199 = t0_0110001111111;
assign input_3200 = t0_0110010000000;
assign input_3201 = t0_0110010000001;
assign input_3202 = t0_0110010000010;
assign input_3203 = t0_0110010000011;
assign input_3204 = t0_0110010000100;
assign input_3205 = t0_0110010000101;
assign input_3206 = t0_0110010000110;
assign input_3207 = t0_0110010000111;
assign input_3208 = t0_0110010001000;
assign input_3209 = t0_0110010001001;
assign input_3210 = t0_0110010001010;
assign input_3211 = t0_0110010001011;
assign input_3212 = t0_0110010001100;
assign input_3213 = t0_0110010001101;
assign input_3214 = t0_0110010001110;
assign input_3215 = t0_0110010001111;
assign input_3216 = t0_0110010010000;
assign input_3217 = t0_0110010010001;
assign input_3218 = t0_0110010010010;
assign input_3219 = t0_0110010010011;
assign input_3220 = t0_0110010010100;
assign input_3221 = t0_0110010010101;
assign input_3222 = t0_0110010010110;
assign input_3223 = t0_0110010010111;
assign input_3224 = t0_0110010011000;
assign input_3225 = t0_0110010011001;
assign input_3226 = t0_0110010011010;
assign input_3227 = t0_0110010011011;
assign input_3228 = t0_0110010011100;
assign input_3229 = t0_0110010011101;
assign input_3230 = t0_0110010011110;
assign input_3231 = t0_0110010011111;
assign input_3232 = t0_0110010100000;
assign input_3233 = t0_0110010100001;
assign input_3234 = t0_0110010100010;
assign input_3235 = t0_0110010100011;
assign input_3236 = t0_0110010100100;
assign input_3237 = t0_0110010100101;
assign input_3238 = t0_0110010100110;
assign input_3239 = t0_0110010100111;
assign input_3240 = t0_0110010101000;
assign input_3241 = t0_0110010101001;
assign input_3242 = t0_0110010101010;
assign input_3243 = t0_0110010101011;
assign input_3244 = t0_0110010101100;
assign input_3245 = t0_0110010101101;
assign input_3246 = t0_0110010101110;
assign input_3247 = t0_0110010101111;
assign input_3248 = t0_0110010110000;
assign input_3249 = t0_0110010110001;
assign input_3250 = t0_0110010110010;
assign input_3251 = t0_0110010110011;
assign input_3252 = t0_0110010110100;
assign input_3253 = t0_0110010110101;
assign input_3254 = t0_0110010110110;
assign input_3255 = t0_0110010110111;
assign input_3256 = t0_0110010111000;
assign input_3257 = t0_0110010111001;
assign input_3258 = t0_0110010111010;
assign input_3259 = t0_0110010111011;
assign input_3260 = t0_0110010111100;
assign input_3261 = t0_0110010111101;
assign input_3262 = t0_0110010111110;
assign input_3263 = t0_0110010111111;
assign input_3264 = t0_0110011000000;
assign input_3265 = t0_0110011000001;
assign input_3266 = t0_0110011000010;
assign input_3267 = t0_0110011000011;
assign input_3268 = t0_0110011000100;
assign input_3269 = t0_0110011000101;
assign input_3270 = t0_0110011000110;
assign input_3271 = t0_0110011000111;
assign input_3272 = t0_0110011001000;
assign input_3273 = t0_0110011001001;
assign input_3274 = t0_0110011001010;
assign input_3275 = t0_0110011001011;
assign input_3276 = t0_0110011001100;
assign input_3277 = t0_0110011001101;
assign input_3278 = t0_0110011001110;
assign input_3279 = t0_0110011001111;
assign input_3280 = t0_0110011010000;
assign input_3281 = t0_0110011010001;
assign input_3282 = t0_0110011010010;
assign input_3283 = t0_0110011010011;
assign input_3284 = t0_0110011010100;
assign input_3285 = t0_0110011010101;
assign input_3286 = t0_0110011010110;
assign input_3287 = t0_0110011010111;
assign input_3288 = t0_0110011011000;
assign input_3289 = t0_0110011011001;
assign input_3290 = t0_0110011011010;
assign input_3291 = t0_0110011011011;
assign input_3292 = t0_0110011011100;
assign input_3293 = t0_0110011011101;
assign input_3294 = t0_0110011011110;
assign input_3295 = t0_0110011011111;
assign input_3296 = t0_0110011100000;
assign input_3297 = t0_0110011100001;
assign input_3298 = t0_0110011100010;
assign input_3299 = t0_0110011100011;
assign input_3300 = t0_0110011100100;
assign input_3301 = t0_0110011100101;
assign input_3302 = t0_0110011100110;
assign input_3303 = t0_0110011100111;
assign input_3304 = t0_0110011101000;
assign input_3305 = t0_0110011101001;
assign input_3306 = t0_0110011101010;
assign input_3307 = t0_0110011101011;
assign input_3308 = t0_0110011101100;
assign input_3309 = t0_0110011101101;
assign input_3310 = t0_0110011101110;
assign input_3311 = t0_0110011101111;
assign input_3312 = t0_0110011110000;
assign input_3313 = t0_0110011110001;
assign input_3314 = t0_0110011110010;
assign input_3315 = t0_0110011110011;
assign input_3316 = t0_0110011110100;
assign input_3317 = t0_0110011110101;
assign input_3318 = t0_0110011110110;
assign input_3319 = t0_0110011110111;
assign input_3320 = t0_0110011111000;
assign input_3321 = t0_0110011111001;
assign input_3322 = t0_0110011111010;
assign input_3323 = t0_0110011111011;
assign input_3324 = t0_0110011111100;
assign input_3325 = t0_0110011111101;
assign input_3326 = t0_0110011111110;
assign input_3327 = t0_0110011111111;
assign input_3328 = t0_0110100000000;
assign input_3329 = t0_0110100000001;
assign input_3330 = t0_0110100000010;
assign input_3331 = t0_0110100000011;
assign input_3332 = t0_0110100000100;
assign input_3333 = t0_0110100000101;
assign input_3334 = t0_0110100000110;
assign input_3335 = t0_0110100000111;
assign input_3336 = t0_0110100001000;
assign input_3337 = t0_0110100001001;
assign input_3338 = t0_0110100001010;
assign input_3339 = t0_0110100001011;
assign input_3340 = t0_0110100001100;
assign input_3341 = t0_0110100001101;
assign input_3342 = t0_0110100001110;
assign input_3343 = t0_0110100001111;
assign input_3344 = t0_0110100010000;
assign input_3345 = t0_0110100010001;
assign input_3346 = t0_0110100010010;
assign input_3347 = t0_0110100010011;
assign input_3348 = t0_0110100010100;
assign input_3349 = t0_0110100010101;
assign input_3350 = t0_0110100010110;
assign input_3351 = t0_0110100010111;
assign input_3352 = t0_0110100011000;
assign input_3353 = t0_0110100011001;
assign input_3354 = t0_0110100011010;
assign input_3355 = t0_0110100011011;
assign input_3356 = t0_0110100011100;
assign input_3357 = t0_0110100011101;
assign input_3358 = t0_0110100011110;
assign input_3359 = t0_0110100011111;
assign input_3360 = t0_0110100100000;
assign input_3361 = t0_0110100100001;
assign input_3362 = t0_0110100100010;
assign input_3363 = t0_0110100100011;
assign input_3364 = t0_0110100100100;
assign input_3365 = t0_0110100100101;
assign input_3366 = t0_0110100100110;
assign input_3367 = t0_0110100100111;
assign input_3368 = t0_0110100101000;
assign input_3369 = t0_0110100101001;
assign input_3370 = t0_0110100101010;
assign input_3371 = t0_0110100101011;
assign input_3372 = t0_0110100101100;
assign input_3373 = t0_0110100101101;
assign input_3374 = t0_0110100101110;
assign input_3375 = t0_0110100101111;
assign input_3376 = t0_0110100110000;
assign input_3377 = t0_0110100110001;
assign input_3378 = t0_0110100110010;
assign input_3379 = t0_0110100110011;
assign input_3380 = t0_0110100110100;
assign input_3381 = t0_0110100110101;
assign input_3382 = t0_0110100110110;
assign input_3383 = t0_0110100110111;
assign input_3384 = t0_0110100111000;
assign input_3385 = t0_0110100111001;
assign input_3386 = t0_0110100111010;
assign input_3387 = t0_0110100111011;
assign input_3388 = t0_0110100111100;
assign input_3389 = t0_0110100111101;
assign input_3390 = t0_0110100111110;
assign input_3391 = t0_0110100111111;
assign input_3392 = t0_0110101000000;
assign input_3393 = t0_0110101000001;
assign input_3394 = t0_0110101000010;
assign input_3395 = t0_0110101000011;
assign input_3396 = t0_0110101000100;
assign input_3397 = t0_0110101000101;
assign input_3398 = t0_0110101000110;
assign input_3399 = t0_0110101000111;
assign input_3400 = t0_0110101001000;
assign input_3401 = t0_0110101001001;
assign input_3402 = t0_0110101001010;
assign input_3403 = t0_0110101001011;
assign input_3404 = t0_0110101001100;
assign input_3405 = t0_0110101001101;
assign input_3406 = t0_0110101001110;
assign input_3407 = t0_0110101001111;
assign input_3408 = t0_0110101010000;
assign input_3409 = t0_0110101010001;
assign input_3410 = t0_0110101010010;
assign input_3411 = t0_0110101010011;
assign input_3412 = t0_0110101010100;
assign input_3413 = t0_0110101010101;
assign input_3414 = t0_0110101010110;
assign input_3415 = t0_0110101010111;
assign input_3416 = t0_0110101011000;
assign input_3417 = t0_0110101011001;
assign input_3418 = t0_0110101011010;
assign input_3419 = t0_0110101011011;
assign input_3420 = t0_0110101011100;
assign input_3421 = t0_0110101011101;
assign input_3422 = t0_0110101011110;
assign input_3423 = t0_0110101011111;
assign input_3424 = t0_0110101100000;
assign input_3425 = t0_0110101100001;
assign input_3426 = t0_0110101100010;
assign input_3427 = t0_0110101100011;
assign input_3428 = t0_0110101100100;
assign input_3429 = t0_0110101100101;
assign input_3430 = t0_0110101100110;
assign input_3431 = t0_0110101100111;
assign input_3432 = t0_0110101101000;
assign input_3433 = t0_0110101101001;
assign input_3434 = t0_0110101101010;
assign input_3435 = t0_0110101101011;
assign input_3436 = t0_0110101101100;
assign input_3437 = t0_0110101101101;
assign input_3438 = t0_0110101101110;
assign input_3439 = t0_0110101101111;
assign input_3440 = t0_0110101110000;
assign input_3441 = t0_0110101110001;
assign input_3442 = t0_0110101110010;
assign input_3443 = t0_0110101110011;
assign input_3444 = t0_0110101110100;
assign input_3445 = t0_0110101110101;
assign input_3446 = t0_0110101110110;
assign input_3447 = t0_0110101110111;
assign input_3448 = t0_0110101111000;
assign input_3449 = t0_0110101111001;
assign input_3450 = t0_0110101111010;
assign input_3451 = t0_0110101111011;
assign input_3452 = t0_0110101111100;
assign input_3453 = t0_0110101111101;
assign input_3454 = t0_0110101111110;
assign input_3455 = t0_0110101111111;
assign input_3456 = t0_0110110000000;
assign input_3457 = t0_0110110000001;
assign input_3458 = t0_0110110000010;
assign input_3459 = t0_0110110000011;
assign input_3460 = t0_0110110000100;
assign input_3461 = t0_0110110000101;
assign input_3462 = t0_0110110000110;
assign input_3463 = t0_0110110000111;
assign input_3464 = t0_0110110001000;
assign input_3465 = t0_0110110001001;
assign input_3466 = t0_0110110001010;
assign input_3467 = t0_0110110001011;
assign input_3468 = t0_0110110001100;
assign input_3469 = t0_0110110001101;
assign input_3470 = t0_0110110001110;
assign input_3471 = t0_0110110001111;
assign input_3472 = t0_0110110010000;
assign input_3473 = t0_0110110010001;
assign input_3474 = t0_0110110010010;
assign input_3475 = t0_0110110010011;
assign input_3476 = t0_0110110010100;
assign input_3477 = t0_0110110010101;
assign input_3478 = t0_0110110010110;
assign input_3479 = t0_0110110010111;
assign input_3480 = t0_0110110011000;
assign input_3481 = t0_0110110011001;
assign input_3482 = t0_0110110011010;
assign input_3483 = t0_0110110011011;
assign input_3484 = t0_0110110011100;
assign input_3485 = t0_0110110011101;
assign input_3486 = t0_0110110011110;
assign input_3487 = t0_0110110011111;
assign input_3488 = t0_0110110100000;
assign input_3489 = t0_0110110100001;
assign input_3490 = t0_0110110100010;
assign input_3491 = t0_0110110100011;
assign input_3492 = t0_0110110100100;
assign input_3493 = t0_0110110100101;
assign input_3494 = t0_0110110100110;
assign input_3495 = t0_0110110100111;
assign input_3496 = t0_0110110101000;
assign input_3497 = t0_0110110101001;
assign input_3498 = t0_0110110101010;
assign input_3499 = t0_0110110101011;
assign input_3500 = t0_0110110101100;
assign input_3501 = t0_0110110101101;
assign input_3502 = t0_0110110101110;
assign input_3503 = t0_0110110101111;
assign input_3504 = t0_0110110110000;
assign input_3505 = t0_0110110110001;
assign input_3506 = t0_0110110110010;
assign input_3507 = t0_0110110110011;
assign input_3508 = t0_0110110110100;
assign input_3509 = t0_0110110110101;
assign input_3510 = t0_0110110110110;
assign input_3511 = t0_0110110110111;
assign input_3512 = t0_0110110111000;
assign input_3513 = t0_0110110111001;
assign input_3514 = t0_0110110111010;
assign input_3515 = t0_0110110111011;
assign input_3516 = t0_0110110111100;
assign input_3517 = t0_0110110111101;
assign input_3518 = t0_0110110111110;
assign input_3519 = t0_0110110111111;
assign input_3520 = t0_0110111000000;
assign input_3521 = t0_0110111000001;
assign input_3522 = t0_0110111000010;
assign input_3523 = t0_0110111000011;
assign input_3524 = t0_0110111000100;
assign input_3525 = t0_0110111000101;
assign input_3526 = t0_0110111000110;
assign input_3527 = t0_0110111000111;
assign input_3528 = t0_0110111001000;
assign input_3529 = t0_0110111001001;
assign input_3530 = t0_0110111001010;
assign input_3531 = t0_0110111001011;
assign input_3532 = t0_0110111001100;
assign input_3533 = t0_0110111001101;
assign input_3534 = t0_0110111001110;
assign input_3535 = t0_0110111001111;
assign input_3536 = t0_0110111010000;
assign input_3537 = t0_0110111010001;
assign input_3538 = t0_0110111010010;
assign input_3539 = t0_0110111010011;
assign input_3540 = t0_0110111010100;
assign input_3541 = t0_0110111010101;
assign input_3542 = t0_0110111010110;
assign input_3543 = t0_0110111010111;
assign input_3544 = t0_0110111011000;
assign input_3545 = t0_0110111011001;
assign input_3546 = t0_0110111011010;
assign input_3547 = t0_0110111011011;
assign input_3548 = t0_0110111011100;
assign input_3549 = t0_0110111011101;
assign input_3550 = t0_0110111011110;
assign input_3551 = t0_0110111011111;
assign input_3552 = t0_0110111100000;
assign input_3553 = t0_0110111100001;
assign input_3554 = t0_0110111100010;
assign input_3555 = t0_0110111100011;
assign input_3556 = t0_0110111100100;
assign input_3557 = t0_0110111100101;
assign input_3558 = t0_0110111100110;
assign input_3559 = t0_0110111100111;
assign input_3560 = t0_0110111101000;
assign input_3561 = t0_0110111101001;
assign input_3562 = t0_0110111101010;
assign input_3563 = t0_0110111101011;
assign input_3564 = t0_0110111101100;
assign input_3565 = t0_0110111101101;
assign input_3566 = t0_0110111101110;
assign input_3567 = t0_0110111101111;
assign input_3568 = t0_0110111110000;
assign input_3569 = t0_0110111110001;
assign input_3570 = t0_0110111110010;
assign input_3571 = t0_0110111110011;
assign input_3572 = t0_0110111110100;
assign input_3573 = t0_0110111110101;
assign input_3574 = t0_0110111110110;
assign input_3575 = t0_0110111110111;
assign input_3576 = t0_0110111111000;
assign input_3577 = t0_0110111111001;
assign input_3578 = t0_0110111111010;
assign input_3579 = t0_0110111111011;
assign input_3580 = t0_0110111111100;
assign input_3581 = t0_0110111111101;
assign input_3582 = t0_0110111111110;
assign input_3583 = t0_0110111111111;
assign input_3584 = t0_0111000000000;
assign input_3585 = t0_0111000000001;
assign input_3586 = t0_0111000000010;
assign input_3587 = t0_0111000000011;
assign input_3588 = t0_0111000000100;
assign input_3589 = t0_0111000000101;
assign input_3590 = t0_0111000000110;
assign input_3591 = t0_0111000000111;
assign input_3592 = t0_0111000001000;
assign input_3593 = t0_0111000001001;
assign input_3594 = t0_0111000001010;
assign input_3595 = t0_0111000001011;
assign input_3596 = t0_0111000001100;
assign input_3597 = t0_0111000001101;
assign input_3598 = t0_0111000001110;
assign input_3599 = t0_0111000001111;
assign input_3600 = t0_0111000010000;
assign input_3601 = t0_0111000010001;
assign input_3602 = t0_0111000010010;
assign input_3603 = t0_0111000010011;
assign input_3604 = t0_0111000010100;
assign input_3605 = t0_0111000010101;
assign input_3606 = t0_0111000010110;
assign input_3607 = t0_0111000010111;
assign input_3608 = t0_0111000011000;
assign input_3609 = t0_0111000011001;
assign input_3610 = t0_0111000011010;
assign input_3611 = t0_0111000011011;
assign input_3612 = t0_0111000011100;
assign input_3613 = t0_0111000011101;
assign input_3614 = t0_0111000011110;
assign input_3615 = t0_0111000011111;
assign input_3616 = t0_0111000100000;
assign input_3617 = t0_0111000100001;
assign input_3618 = t0_0111000100010;
assign input_3619 = t0_0111000100011;
assign input_3620 = t0_0111000100100;
assign input_3621 = t0_0111000100101;
assign input_3622 = t0_0111000100110;
assign input_3623 = t0_0111000100111;
assign input_3624 = t0_0111000101000;
assign input_3625 = t0_0111000101001;
assign input_3626 = t0_0111000101010;
assign input_3627 = t0_0111000101011;
assign input_3628 = t0_0111000101100;
assign input_3629 = t0_0111000101101;
assign input_3630 = t0_0111000101110;
assign input_3631 = t0_0111000101111;
assign input_3632 = t0_0111000110000;
assign input_3633 = t0_0111000110001;
assign input_3634 = t0_0111000110010;
assign input_3635 = t0_0111000110011;
assign input_3636 = t0_0111000110100;
assign input_3637 = t0_0111000110101;
assign input_3638 = t0_0111000110110;
assign input_3639 = t0_0111000110111;
assign input_3640 = t0_0111000111000;
assign input_3641 = t0_0111000111001;
assign input_3642 = t0_0111000111010;
assign input_3643 = t0_0111000111011;
assign input_3644 = t0_0111000111100;
assign input_3645 = t0_0111000111101;
assign input_3646 = t0_0111000111110;
assign input_3647 = t0_0111000111111;
assign input_3648 = t0_0111001000000;
assign input_3649 = t0_0111001000001;
assign input_3650 = t0_0111001000010;
assign input_3651 = t0_0111001000011;
assign input_3652 = t0_0111001000100;
assign input_3653 = t0_0111001000101;
assign input_3654 = t0_0111001000110;
assign input_3655 = t0_0111001000111;
assign input_3656 = t0_0111001001000;
assign input_3657 = t0_0111001001001;
assign input_3658 = t0_0111001001010;
assign input_3659 = t0_0111001001011;
assign input_3660 = t0_0111001001100;
assign input_3661 = t0_0111001001101;
assign input_3662 = t0_0111001001110;
assign input_3663 = t0_0111001001111;
assign input_3664 = t0_0111001010000;
assign input_3665 = t0_0111001010001;
assign input_3666 = t0_0111001010010;
assign input_3667 = t0_0111001010011;
assign input_3668 = t0_0111001010100;
assign input_3669 = t0_0111001010101;
assign input_3670 = t0_0111001010110;
assign input_3671 = t0_0111001010111;
assign input_3672 = t0_0111001011000;
assign input_3673 = t0_0111001011001;
assign input_3674 = t0_0111001011010;
assign input_3675 = t0_0111001011011;
assign input_3676 = t0_0111001011100;
assign input_3677 = t0_0111001011101;
assign input_3678 = t0_0111001011110;
assign input_3679 = t0_0111001011111;
assign input_3680 = t0_0111001100000;
assign input_3681 = t0_0111001100001;
assign input_3682 = t0_0111001100010;
assign input_3683 = t0_0111001100011;
assign input_3684 = t0_0111001100100;
assign input_3685 = t0_0111001100101;
assign input_3686 = t0_0111001100110;
assign input_3687 = t0_0111001100111;
assign input_3688 = t0_0111001101000;
assign input_3689 = t0_0111001101001;
assign input_3690 = t0_0111001101010;
assign input_3691 = t0_0111001101011;
assign input_3692 = t0_0111001101100;
assign input_3693 = t0_0111001101101;
assign input_3694 = t0_0111001101110;
assign input_3695 = t0_0111001101111;
assign input_3696 = t0_0111001110000;
assign input_3697 = t0_0111001110001;
assign input_3698 = t0_0111001110010;
assign input_3699 = t0_0111001110011;
assign input_3700 = t0_0111001110100;
assign input_3701 = t0_0111001110101;
assign input_3702 = t0_0111001110110;
assign input_3703 = t0_0111001110111;
assign input_3704 = t0_0111001111000;
assign input_3705 = t0_0111001111001;
assign input_3706 = t0_0111001111010;
assign input_3707 = t0_0111001111011;
assign input_3708 = t0_0111001111100;
assign input_3709 = t0_0111001111101;
assign input_3710 = t0_0111001111110;
assign input_3711 = t0_0111001111111;
assign input_3712 = t0_0111010000000;
assign input_3713 = t0_0111010000001;
assign input_3714 = t0_0111010000010;
assign input_3715 = t0_0111010000011;
assign input_3716 = t0_0111010000100;
assign input_3717 = t0_0111010000101;
assign input_3718 = t0_0111010000110;
assign input_3719 = t0_0111010000111;
assign input_3720 = t0_0111010001000;
assign input_3721 = t0_0111010001001;
assign input_3722 = t0_0111010001010;
assign input_3723 = t0_0111010001011;
assign input_3724 = t0_0111010001100;
assign input_3725 = t0_0111010001101;
assign input_3726 = t0_0111010001110;
assign input_3727 = t0_0111010001111;
assign input_3728 = t0_0111010010000;
assign input_3729 = t0_0111010010001;
assign input_3730 = t0_0111010010010;
assign input_3731 = t0_0111010010011;
assign input_3732 = t0_0111010010100;
assign input_3733 = t0_0111010010101;
assign input_3734 = t0_0111010010110;
assign input_3735 = t0_0111010010111;
assign input_3736 = t0_0111010011000;
assign input_3737 = t0_0111010011001;
assign input_3738 = t0_0111010011010;
assign input_3739 = t0_0111010011011;
assign input_3740 = t0_0111010011100;
assign input_3741 = t0_0111010011101;
assign input_3742 = t0_0111010011110;
assign input_3743 = t0_0111010011111;
assign input_3744 = t0_0111010100000;
assign input_3745 = t0_0111010100001;
assign input_3746 = t0_0111010100010;
assign input_3747 = t0_0111010100011;
assign input_3748 = t0_0111010100100;
assign input_3749 = t0_0111010100101;
assign input_3750 = t0_0111010100110;
assign input_3751 = t0_0111010100111;
assign input_3752 = t0_0111010101000;
assign input_3753 = t0_0111010101001;
assign input_3754 = t0_0111010101010;
assign input_3755 = t0_0111010101011;
assign input_3756 = t0_0111010101100;
assign input_3757 = t0_0111010101101;
assign input_3758 = t0_0111010101110;
assign input_3759 = t0_0111010101111;
assign input_3760 = t0_0111010110000;
assign input_3761 = t0_0111010110001;
assign input_3762 = t0_0111010110010;
assign input_3763 = t0_0111010110011;
assign input_3764 = t0_0111010110100;
assign input_3765 = t0_0111010110101;
assign input_3766 = t0_0111010110110;
assign input_3767 = t0_0111010110111;
assign input_3768 = t0_0111010111000;
assign input_3769 = t0_0111010111001;
assign input_3770 = t0_0111010111010;
assign input_3771 = t0_0111010111011;
assign input_3772 = t0_0111010111100;
assign input_3773 = t0_0111010111101;
assign input_3774 = t0_0111010111110;
assign input_3775 = t0_0111010111111;
assign input_3776 = t0_0111011000000;
assign input_3777 = t0_0111011000001;
assign input_3778 = t0_0111011000010;
assign input_3779 = t0_0111011000011;
assign input_3780 = t0_0111011000100;
assign input_3781 = t0_0111011000101;
assign input_3782 = t0_0111011000110;
assign input_3783 = t0_0111011000111;
assign input_3784 = t0_0111011001000;
assign input_3785 = t0_0111011001001;
assign input_3786 = t0_0111011001010;
assign input_3787 = t0_0111011001011;
assign input_3788 = t0_0111011001100;
assign input_3789 = t0_0111011001101;
assign input_3790 = t0_0111011001110;
assign input_3791 = t0_0111011001111;
assign input_3792 = t0_0111011010000;
assign input_3793 = t0_0111011010001;
assign input_3794 = t0_0111011010010;
assign input_3795 = t0_0111011010011;
assign input_3796 = t0_0111011010100;
assign input_3797 = t0_0111011010101;
assign input_3798 = t0_0111011010110;
assign input_3799 = t0_0111011010111;
assign input_3800 = t0_0111011011000;
assign input_3801 = t0_0111011011001;
assign input_3802 = t0_0111011011010;
assign input_3803 = t0_0111011011011;
assign input_3804 = t0_0111011011100;
assign input_3805 = t0_0111011011101;
assign input_3806 = t0_0111011011110;
assign input_3807 = t0_0111011011111;
assign input_3808 = t0_0111011100000;
assign input_3809 = t0_0111011100001;
assign input_3810 = t0_0111011100010;
assign input_3811 = t0_0111011100011;
assign input_3812 = t0_0111011100100;
assign input_3813 = t0_0111011100101;
assign input_3814 = t0_0111011100110;
assign input_3815 = t0_0111011100111;
assign input_3816 = t0_0111011101000;
assign input_3817 = t0_0111011101001;
assign input_3818 = t0_0111011101010;
assign input_3819 = t0_0111011101011;
assign input_3820 = t0_0111011101100;
assign input_3821 = t0_0111011101101;
assign input_3822 = t0_0111011101110;
assign input_3823 = t0_0111011101111;
assign input_3824 = t0_0111011110000;
assign input_3825 = t0_0111011110001;
assign input_3826 = t0_0111011110010;
assign input_3827 = t0_0111011110011;
assign input_3828 = t0_0111011110100;
assign input_3829 = t0_0111011110101;
assign input_3830 = t0_0111011110110;
assign input_3831 = t0_0111011110111;
assign input_3832 = t0_0111011111000;
assign input_3833 = t0_0111011111001;
assign input_3834 = t0_0111011111010;
assign input_3835 = t0_0111011111011;
assign input_3836 = t0_0111011111100;
assign input_3837 = t0_0111011111101;
assign input_3838 = t0_0111011111110;
assign input_3839 = t0_0111011111111;
assign input_3840 = t0_0111100000000;
assign input_3841 = t0_0111100000001;
assign input_3842 = t0_0111100000010;
assign input_3843 = t0_0111100000011;
assign input_3844 = t0_0111100000100;
assign input_3845 = t0_0111100000101;
assign input_3846 = t0_0111100000110;
assign input_3847 = t0_0111100000111;
assign input_3848 = t0_0111100001000;
assign input_3849 = t0_0111100001001;
assign input_3850 = t0_0111100001010;
assign input_3851 = t0_0111100001011;
assign input_3852 = t0_0111100001100;
assign input_3853 = t0_0111100001101;
assign input_3854 = t0_0111100001110;
assign input_3855 = t0_0111100001111;
assign input_3856 = t0_0111100010000;
assign input_3857 = t0_0111100010001;
assign input_3858 = t0_0111100010010;
assign input_3859 = t0_0111100010011;
assign input_3860 = t0_0111100010100;
assign input_3861 = t0_0111100010101;
assign input_3862 = t0_0111100010110;
assign input_3863 = t0_0111100010111;
assign input_3864 = t0_0111100011000;
assign input_3865 = t0_0111100011001;
assign input_3866 = t0_0111100011010;
assign input_3867 = t0_0111100011011;
assign input_3868 = t0_0111100011100;
assign input_3869 = t0_0111100011101;
assign input_3870 = t0_0111100011110;
assign input_3871 = t0_0111100011111;
assign input_3872 = t0_0111100100000;
assign input_3873 = t0_0111100100001;
assign input_3874 = t0_0111100100010;
assign input_3875 = t0_0111100100011;
assign input_3876 = t0_0111100100100;
assign input_3877 = t0_0111100100101;
assign input_3878 = t0_0111100100110;
assign input_3879 = t0_0111100100111;
assign input_3880 = t0_0111100101000;
assign input_3881 = t0_0111100101001;
assign input_3882 = t0_0111100101010;
assign input_3883 = t0_0111100101011;
assign input_3884 = t0_0111100101100;
assign input_3885 = t0_0111100101101;
assign input_3886 = t0_0111100101110;
assign input_3887 = t0_0111100101111;
assign input_3888 = t0_0111100110000;
assign input_3889 = t0_0111100110001;
assign input_3890 = t0_0111100110010;
assign input_3891 = t0_0111100110011;
assign input_3892 = t0_0111100110100;
assign input_3893 = t0_0111100110101;
assign input_3894 = t0_0111100110110;
assign input_3895 = t0_0111100110111;
assign input_3896 = t0_0111100111000;
assign input_3897 = t0_0111100111001;
assign input_3898 = t0_0111100111010;
assign input_3899 = t0_0111100111011;
assign input_3900 = t0_0111100111100;
assign input_3901 = t0_0111100111101;
assign input_3902 = t0_0111100111110;
assign input_3903 = t0_0111100111111;
assign input_3904 = t0_0111101000000;
assign input_3905 = t0_0111101000001;
assign input_3906 = t0_0111101000010;
assign input_3907 = t0_0111101000011;
assign input_3908 = t0_0111101000100;
assign input_3909 = t0_0111101000101;
assign input_3910 = t0_0111101000110;
assign input_3911 = t0_0111101000111;
assign input_3912 = t0_0111101001000;
assign input_3913 = t0_0111101001001;
assign input_3914 = t0_0111101001010;
assign input_3915 = t0_0111101001011;
assign input_3916 = t0_0111101001100;
assign input_3917 = t0_0111101001101;
assign input_3918 = t0_0111101001110;
assign input_3919 = t0_0111101001111;
assign input_3920 = t0_0111101010000;
assign input_3921 = t0_0111101010001;
assign input_3922 = t0_0111101010010;
assign input_3923 = t0_0111101010011;
assign input_3924 = t0_0111101010100;
assign input_3925 = t0_0111101010101;
assign input_3926 = t0_0111101010110;
assign input_3927 = t0_0111101010111;
assign input_3928 = t0_0111101011000;
assign input_3929 = t0_0111101011001;
assign input_3930 = t0_0111101011010;
assign input_3931 = t0_0111101011011;
assign input_3932 = t0_0111101011100;
assign input_3933 = t0_0111101011101;
assign input_3934 = t0_0111101011110;
assign input_3935 = t0_0111101011111;
assign input_3936 = t0_0111101100000;
assign input_3937 = t0_0111101100001;
assign input_3938 = t0_0111101100010;
assign input_3939 = t0_0111101100011;
assign input_3940 = t0_0111101100100;
assign input_3941 = t0_0111101100101;
assign input_3942 = t0_0111101100110;
assign input_3943 = t0_0111101100111;
assign input_3944 = t0_0111101101000;
assign input_3945 = t0_0111101101001;
assign input_3946 = t0_0111101101010;
assign input_3947 = t0_0111101101011;
assign input_3948 = t0_0111101101100;
assign input_3949 = t0_0111101101101;
assign input_3950 = t0_0111101101110;
assign input_3951 = t0_0111101101111;
assign input_3952 = t0_0111101110000;
assign input_3953 = t0_0111101110001;
assign input_3954 = t0_0111101110010;
assign input_3955 = t0_0111101110011;
assign input_3956 = t0_0111101110100;
assign input_3957 = t0_0111101110101;
assign input_3958 = t0_0111101110110;
assign input_3959 = t0_0111101110111;
assign input_3960 = t0_0111101111000;
assign input_3961 = t0_0111101111001;
assign input_3962 = t0_0111101111010;
assign input_3963 = t0_0111101111011;
assign input_3964 = t0_0111101111100;
assign input_3965 = t0_0111101111101;
assign input_3966 = t0_0111101111110;
assign input_3967 = t0_0111101111111;
assign input_3968 = t0_0111110000000;
assign input_3969 = t0_0111110000001;
assign input_3970 = t0_0111110000010;
assign input_3971 = t0_0111110000011;
assign input_3972 = t0_0111110000100;
assign input_3973 = t0_0111110000101;
assign input_3974 = t0_0111110000110;
assign input_3975 = t0_0111110000111;
assign input_3976 = t0_0111110001000;
assign input_3977 = t0_0111110001001;
assign input_3978 = t0_0111110001010;
assign input_3979 = t0_0111110001011;
assign input_3980 = t0_0111110001100;
assign input_3981 = t0_0111110001101;
assign input_3982 = t0_0111110001110;
assign input_3983 = t0_0111110001111;
assign input_3984 = t0_0111110010000;
assign input_3985 = t0_0111110010001;
assign input_3986 = t0_0111110010010;
assign input_3987 = t0_0111110010011;
assign input_3988 = t0_0111110010100;
assign input_3989 = t0_0111110010101;
assign input_3990 = t0_0111110010110;
assign input_3991 = t0_0111110010111;
assign input_3992 = t0_0111110011000;
assign input_3993 = t0_0111110011001;
assign input_3994 = t0_0111110011010;
assign input_3995 = t0_0111110011011;
assign input_3996 = t0_0111110011100;
assign input_3997 = t0_0111110011101;
assign input_3998 = t0_0111110011110;
assign input_3999 = t0_0111110011111;
assign input_4000 = t0_0111110100000;
assign input_4001 = t0_0111110100001;
assign input_4002 = t0_0111110100010;
assign input_4003 = t0_0111110100011;
assign input_4004 = t0_0111110100100;
assign input_4005 = t0_0111110100101;
assign input_4006 = t0_0111110100110;
assign input_4007 = t0_0111110100111;
assign input_4008 = t0_0111110101000;
assign input_4009 = t0_0111110101001;
assign input_4010 = t0_0111110101010;
assign input_4011 = t0_0111110101011;
assign input_4012 = t0_0111110101100;
assign input_4013 = t0_0111110101101;
assign input_4014 = t0_0111110101110;
assign input_4015 = t0_0111110101111;
assign input_4016 = t0_0111110110000;
assign input_4017 = t0_0111110110001;
assign input_4018 = t0_0111110110010;
assign input_4019 = t0_0111110110011;
assign input_4020 = t0_0111110110100;
assign input_4021 = t0_0111110110101;
assign input_4022 = t0_0111110110110;
assign input_4023 = t0_0111110110111;
assign input_4024 = t0_0111110111000;
assign input_4025 = t0_0111110111001;
assign input_4026 = t0_0111110111010;
assign input_4027 = t0_0111110111011;
assign input_4028 = t0_0111110111100;
assign input_4029 = t0_0111110111101;
assign input_4030 = t0_0111110111110;
assign input_4031 = t0_0111110111111;
assign input_4032 = t0_0111111000000;
assign input_4033 = t0_0111111000001;
assign input_4034 = t0_0111111000010;
assign input_4035 = t0_0111111000011;
assign input_4036 = t0_0111111000100;
assign input_4037 = t0_0111111000101;
assign input_4038 = t0_0111111000110;
assign input_4039 = t0_0111111000111;
assign input_4040 = t0_0111111001000;
assign input_4041 = t0_0111111001001;
assign input_4042 = t0_0111111001010;
assign input_4043 = t0_0111111001011;
assign input_4044 = t0_0111111001100;
assign input_4045 = t0_0111111001101;
assign input_4046 = t0_0111111001110;
assign input_4047 = t0_0111111001111;
assign input_4048 = t0_0111111010000;
assign input_4049 = t0_0111111010001;
assign input_4050 = t0_0111111010010;
assign input_4051 = t0_0111111010011;
assign input_4052 = t0_0111111010100;
assign input_4053 = t0_0111111010101;
assign input_4054 = t0_0111111010110;
assign input_4055 = t0_0111111010111;
assign input_4056 = t0_0111111011000;
assign input_4057 = t0_0111111011001;
assign input_4058 = t0_0111111011010;
assign input_4059 = t0_0111111011011;
assign input_4060 = t0_0111111011100;
assign input_4061 = t0_0111111011101;
assign input_4062 = t0_0111111011110;
assign input_4063 = t0_0111111011111;
assign input_4064 = t0_0111111100000;
assign input_4065 = t0_0111111100001;
assign input_4066 = t0_0111111100010;
assign input_4067 = t0_0111111100011;
assign input_4068 = t0_0111111100100;
assign input_4069 = t0_0111111100101;
assign input_4070 = t0_0111111100110;
assign input_4071 = t0_0111111100111;
assign input_4072 = t0_0111111101000;
assign input_4073 = t0_0111111101001;
assign input_4074 = t0_0111111101010;
assign input_4075 = t0_0111111101011;
assign input_4076 = t0_0111111101100;
assign input_4077 = t0_0111111101101;
assign input_4078 = t0_0111111101110;
assign input_4079 = t0_0111111101111;
assign input_4080 = t0_0111111110000;
assign input_4081 = t0_0111111110001;
assign input_4082 = t0_0111111110010;
assign input_4083 = t0_0111111110011;
assign input_4084 = t0_0111111110100;
assign input_4085 = t0_0111111110101;
assign input_4086 = t0_0111111110110;
assign input_4087 = t0_0111111110111;
assign input_4088 = t0_0111111111000;
assign input_4089 = t0_0111111111001;
assign input_4090 = t0_0111111111010;
assign input_4091 = t0_0111111111011;
assign input_4092 = t0_0111111111100;
assign input_4093 = t0_0111111111101;
assign input_4094 = t0_0111111111110;
assign input_4095 = t0_0111111111111;
endmodule
