module multiplexer_7 (
inout k_0_0,k_7_0,k_7_1,k_7_2,k_7_3,k_7_4,k_7_5,k_7_6,k_7_7,k_7_8,k_7_9,k_7_10,k_7_11,k_7_12,k_7_13,k_7_14,k_7_15,k_7_16,k_7_17,k_7_18,k_7_19,k_7_20,k_7_21,k_7_22,k_7_23,k_7_24,k_7_25,k_7_26,k_7_27,k_7_28,k_7_29,k_7_30,k_7_31,k_7_32,k_7_33,k_7_34,k_7_35,k_7_36,k_7_37,k_7_38,k_7_39,k_7_40,k_7_41,k_7_42,k_7_43,k_7_44,k_7_45,k_7_46,k_7_47,k_7_48,k_7_49,k_7_50,k_7_51,k_7_52,k_7_53,k_7_54,k_7_55,k_7_56,k_7_57,k_7_58,k_7_59,k_7_60,k_7_61,k_7_62,k_7_63,k_7_64,k_7_65,k_7_66,k_7_67,k_7_68,k_7_69,k_7_70,k_7_71,k_7_72,k_7_73,k_7_74,k_7_75,k_7_76,k_7_77,k_7_78,k_7_79,k_7_80,k_7_81,k_7_82,k_7_83,k_7_84,k_7_85,k_7_86,k_7_87,k_7_88,k_7_89,k_7_90,k_7_91,k_7_92,k_7_93,k_7_94,k_7_95,k_7_96,k_7_97,k_7_98,k_7_99,k_7_100,k_7_101,k_7_102,k_7_103,k_7_104,k_7_105,k_7_106,k_7_107,k_7_108,k_7_109,k_7_110,k_7_111,k_7_112,k_7_113,k_7_114,k_7_115,k_7_116,k_7_117,k_7_118,k_7_119,k_7_120,k_7_121,k_7_122,k_7_123,k_7_124,k_7_125,k_7_126,k_7_127,
input c_0_0, c_0_1,
input c_1_0, c_1_1,
input c_2_0, c_2_1,
input c_3_0, c_3_1,
input c_4_0, c_4_1,
input c_5_0, c_5_1,
input c_6_0, c_6_1,
input c_7_0, c_7_1
);
wire k_1_0,k_1_1;
wire k_2_0,k_2_1,k_2_2,k_2_3;
wire k_3_0,k_3_1,k_3_2,k_3_3,k_3_4,k_3_5,k_3_6,k_3_7;
wire k_4_0,k_4_1,k_4_2,k_4_3,k_4_4,k_4_5,k_4_6,k_4_7,k_4_8,k_4_9,k_4_10,k_4_11,k_4_12,k_4_13,k_4_14,k_4_15;
wire k_5_0,k_5_1,k_5_2,k_5_3,k_5_4,k_5_5,k_5_6,k_5_7,k_5_8,k_5_9,k_5_10,k_5_11,k_5_12,k_5_13,k_5_14,k_5_15,k_5_16,k_5_17,k_5_18,k_5_19,k_5_20,k_5_21,k_5_22,k_5_23,k_5_24,k_5_25,k_5_26,k_5_27,k_5_28,k_5_29,k_5_30,k_5_31;
wire k_6_0,k_6_1,k_6_2,k_6_3,k_6_4,k_6_5,k_6_6,k_6_7,k_6_8,k_6_9,k_6_10,k_6_11,k_6_12,k_6_13,k_6_14,k_6_15,k_6_16,k_6_17,k_6_18,k_6_19,k_6_20,k_6_21,k_6_22,k_6_23,k_6_24,k_6_25,k_6_26,k_6_27,k_6_28,k_6_29,k_6_30,k_6_31,k_6_32,k_6_33,k_6_34,k_6_35,k_6_36,k_6_37,k_6_38,k_6_39,k_6_40,k_6_41,k_6_42,k_6_43,k_6_44,k_6_45,k_6_46,k_6_47,k_6_48,k_6_49,k_6_50,k_6_51,k_6_52,k_6_53,k_6_54,k_6_55,k_6_56,k_6_57,k_6_58,k_6_59,k_6_60,k_6_61,k_6_62,k_6_63;
valve v_1_0 (.fluid_in(k_1_0), .fluid_out(k_0_0), .air_in(c_1_0));
valve v_1_1 (.fluid_in(k_1_1), .fluid_out(k_0_0), .air_in(c_1_1));
valve v_2_0 (.fluid_in(k_2_0), .fluid_out(k_1_0), .air_in(c_2_0));
valve v_2_1 (.fluid_in(k_2_1), .fluid_out(k_1_0), .air_in(c_2_1));
valve v_2_2 (.fluid_in(k_2_2), .fluid_out(k_1_1), .air_in(c_2_0));
valve v_2_3 (.fluid_in(k_2_3), .fluid_out(k_1_1), .air_in(c_2_1));
valve v_3_0 (.fluid_in(k_3_0), .fluid_out(k_2_0), .air_in(c_3_0));
valve v_3_1 (.fluid_in(k_3_1), .fluid_out(k_2_0), .air_in(c_3_1));
valve v_3_2 (.fluid_in(k_3_2), .fluid_out(k_2_1), .air_in(c_3_0));
valve v_3_3 (.fluid_in(k_3_3), .fluid_out(k_2_1), .air_in(c_3_1));
valve v_3_4 (.fluid_in(k_3_4), .fluid_out(k_2_2), .air_in(c_3_0));
valve v_3_5 (.fluid_in(k_3_5), .fluid_out(k_2_2), .air_in(c_3_1));
valve v_3_6 (.fluid_in(k_3_6), .fluid_out(k_2_3), .air_in(c_3_0));
valve v_3_7 (.fluid_in(k_3_7), .fluid_out(k_2_3), .air_in(c_3_1));
valve v_4_0 (.fluid_in(k_4_0), .fluid_out(k_3_0), .air_in(c_4_0));
valve v_4_1 (.fluid_in(k_4_1), .fluid_out(k_3_0), .air_in(c_4_1));
valve v_4_2 (.fluid_in(k_4_2), .fluid_out(k_3_1), .air_in(c_4_0));
valve v_4_3 (.fluid_in(k_4_3), .fluid_out(k_3_1), .air_in(c_4_1));
valve v_4_4 (.fluid_in(k_4_4), .fluid_out(k_3_2), .air_in(c_4_0));
valve v_4_5 (.fluid_in(k_4_5), .fluid_out(k_3_2), .air_in(c_4_1));
valve v_4_6 (.fluid_in(k_4_6), .fluid_out(k_3_3), .air_in(c_4_0));
valve v_4_7 (.fluid_in(k_4_7), .fluid_out(k_3_3), .air_in(c_4_1));
valve v_4_8 (.fluid_in(k_4_8), .fluid_out(k_3_4), .air_in(c_4_0));
valve v_4_9 (.fluid_in(k_4_9), .fluid_out(k_3_4), .air_in(c_4_1));
valve v_4_10 (.fluid_in(k_4_10), .fluid_out(k_3_5), .air_in(c_4_0));
valve v_4_11 (.fluid_in(k_4_11), .fluid_out(k_3_5), .air_in(c_4_1));
valve v_4_12 (.fluid_in(k_4_12), .fluid_out(k_3_6), .air_in(c_4_0));
valve v_4_13 (.fluid_in(k_4_13), .fluid_out(k_3_6), .air_in(c_4_1));
valve v_4_14 (.fluid_in(k_4_14), .fluid_out(k_3_7), .air_in(c_4_0));
valve v_4_15 (.fluid_in(k_4_15), .fluid_out(k_3_7), .air_in(c_4_1));
valve v_5_0 (.fluid_in(k_5_0), .fluid_out(k_4_0), .air_in(c_5_0));
valve v_5_1 (.fluid_in(k_5_1), .fluid_out(k_4_0), .air_in(c_5_1));
valve v_5_2 (.fluid_in(k_5_2), .fluid_out(k_4_1), .air_in(c_5_0));
valve v_5_3 (.fluid_in(k_5_3), .fluid_out(k_4_1), .air_in(c_5_1));
valve v_5_4 (.fluid_in(k_5_4), .fluid_out(k_4_2), .air_in(c_5_0));
valve v_5_5 (.fluid_in(k_5_5), .fluid_out(k_4_2), .air_in(c_5_1));
valve v_5_6 (.fluid_in(k_5_6), .fluid_out(k_4_3), .air_in(c_5_0));
valve v_5_7 (.fluid_in(k_5_7), .fluid_out(k_4_3), .air_in(c_5_1));
valve v_5_8 (.fluid_in(k_5_8), .fluid_out(k_4_4), .air_in(c_5_0));
valve v_5_9 (.fluid_in(k_5_9), .fluid_out(k_4_4), .air_in(c_5_1));
valve v_5_10 (.fluid_in(k_5_10), .fluid_out(k_4_5), .air_in(c_5_0));
valve v_5_11 (.fluid_in(k_5_11), .fluid_out(k_4_5), .air_in(c_5_1));
valve v_5_12 (.fluid_in(k_5_12), .fluid_out(k_4_6), .air_in(c_5_0));
valve v_5_13 (.fluid_in(k_5_13), .fluid_out(k_4_6), .air_in(c_5_1));
valve v_5_14 (.fluid_in(k_5_14), .fluid_out(k_4_7), .air_in(c_5_0));
valve v_5_15 (.fluid_in(k_5_15), .fluid_out(k_4_7), .air_in(c_5_1));
valve v_5_16 (.fluid_in(k_5_16), .fluid_out(k_4_8), .air_in(c_5_0));
valve v_5_17 (.fluid_in(k_5_17), .fluid_out(k_4_8), .air_in(c_5_1));
valve v_5_18 (.fluid_in(k_5_18), .fluid_out(k_4_9), .air_in(c_5_0));
valve v_5_19 (.fluid_in(k_5_19), .fluid_out(k_4_9), .air_in(c_5_1));
valve v_5_20 (.fluid_in(k_5_20), .fluid_out(k_4_10), .air_in(c_5_0));
valve v_5_21 (.fluid_in(k_5_21), .fluid_out(k_4_10), .air_in(c_5_1));
valve v_5_22 (.fluid_in(k_5_22), .fluid_out(k_4_11), .air_in(c_5_0));
valve v_5_23 (.fluid_in(k_5_23), .fluid_out(k_4_11), .air_in(c_5_1));
valve v_5_24 (.fluid_in(k_5_24), .fluid_out(k_4_12), .air_in(c_5_0));
valve v_5_25 (.fluid_in(k_5_25), .fluid_out(k_4_12), .air_in(c_5_1));
valve v_5_26 (.fluid_in(k_5_26), .fluid_out(k_4_13), .air_in(c_5_0));
valve v_5_27 (.fluid_in(k_5_27), .fluid_out(k_4_13), .air_in(c_5_1));
valve v_5_28 (.fluid_in(k_5_28), .fluid_out(k_4_14), .air_in(c_5_0));
valve v_5_29 (.fluid_in(k_5_29), .fluid_out(k_4_14), .air_in(c_5_1));
valve v_5_30 (.fluid_in(k_5_30), .fluid_out(k_4_15), .air_in(c_5_0));
valve v_5_31 (.fluid_in(k_5_31), .fluid_out(k_4_15), .air_in(c_5_1));
valve v_6_0 (.fluid_in(k_6_0), .fluid_out(k_5_0), .air_in(c_6_0));
valve v_6_1 (.fluid_in(k_6_1), .fluid_out(k_5_0), .air_in(c_6_1));
valve v_6_2 (.fluid_in(k_6_2), .fluid_out(k_5_1), .air_in(c_6_0));
valve v_6_3 (.fluid_in(k_6_3), .fluid_out(k_5_1), .air_in(c_6_1));
valve v_6_4 (.fluid_in(k_6_4), .fluid_out(k_5_2), .air_in(c_6_0));
valve v_6_5 (.fluid_in(k_6_5), .fluid_out(k_5_2), .air_in(c_6_1));
valve v_6_6 (.fluid_in(k_6_6), .fluid_out(k_5_3), .air_in(c_6_0));
valve v_6_7 (.fluid_in(k_6_7), .fluid_out(k_5_3), .air_in(c_6_1));
valve v_6_8 (.fluid_in(k_6_8), .fluid_out(k_5_4), .air_in(c_6_0));
valve v_6_9 (.fluid_in(k_6_9), .fluid_out(k_5_4), .air_in(c_6_1));
valve v_6_10 (.fluid_in(k_6_10), .fluid_out(k_5_5), .air_in(c_6_0));
valve v_6_11 (.fluid_in(k_6_11), .fluid_out(k_5_5), .air_in(c_6_1));
valve v_6_12 (.fluid_in(k_6_12), .fluid_out(k_5_6), .air_in(c_6_0));
valve v_6_13 (.fluid_in(k_6_13), .fluid_out(k_5_6), .air_in(c_6_1));
valve v_6_14 (.fluid_in(k_6_14), .fluid_out(k_5_7), .air_in(c_6_0));
valve v_6_15 (.fluid_in(k_6_15), .fluid_out(k_5_7), .air_in(c_6_1));
valve v_6_16 (.fluid_in(k_6_16), .fluid_out(k_5_8), .air_in(c_6_0));
valve v_6_17 (.fluid_in(k_6_17), .fluid_out(k_5_8), .air_in(c_6_1));
valve v_6_18 (.fluid_in(k_6_18), .fluid_out(k_5_9), .air_in(c_6_0));
valve v_6_19 (.fluid_in(k_6_19), .fluid_out(k_5_9), .air_in(c_6_1));
valve v_6_20 (.fluid_in(k_6_20), .fluid_out(k_5_10), .air_in(c_6_0));
valve v_6_21 (.fluid_in(k_6_21), .fluid_out(k_5_10), .air_in(c_6_1));
valve v_6_22 (.fluid_in(k_6_22), .fluid_out(k_5_11), .air_in(c_6_0));
valve v_6_23 (.fluid_in(k_6_23), .fluid_out(k_5_11), .air_in(c_6_1));
valve v_6_24 (.fluid_in(k_6_24), .fluid_out(k_5_12), .air_in(c_6_0));
valve v_6_25 (.fluid_in(k_6_25), .fluid_out(k_5_12), .air_in(c_6_1));
valve v_6_26 (.fluid_in(k_6_26), .fluid_out(k_5_13), .air_in(c_6_0));
valve v_6_27 (.fluid_in(k_6_27), .fluid_out(k_5_13), .air_in(c_6_1));
valve v_6_28 (.fluid_in(k_6_28), .fluid_out(k_5_14), .air_in(c_6_0));
valve v_6_29 (.fluid_in(k_6_29), .fluid_out(k_5_14), .air_in(c_6_1));
valve v_6_30 (.fluid_in(k_6_30), .fluid_out(k_5_15), .air_in(c_6_0));
valve v_6_31 (.fluid_in(k_6_31), .fluid_out(k_5_15), .air_in(c_6_1));
valve v_6_32 (.fluid_in(k_6_32), .fluid_out(k_5_16), .air_in(c_6_0));
valve v_6_33 (.fluid_in(k_6_33), .fluid_out(k_5_16), .air_in(c_6_1));
valve v_6_34 (.fluid_in(k_6_34), .fluid_out(k_5_17), .air_in(c_6_0));
valve v_6_35 (.fluid_in(k_6_35), .fluid_out(k_5_17), .air_in(c_6_1));
valve v_6_36 (.fluid_in(k_6_36), .fluid_out(k_5_18), .air_in(c_6_0));
valve v_6_37 (.fluid_in(k_6_37), .fluid_out(k_5_18), .air_in(c_6_1));
valve v_6_38 (.fluid_in(k_6_38), .fluid_out(k_5_19), .air_in(c_6_0));
valve v_6_39 (.fluid_in(k_6_39), .fluid_out(k_5_19), .air_in(c_6_1));
valve v_6_40 (.fluid_in(k_6_40), .fluid_out(k_5_20), .air_in(c_6_0));
valve v_6_41 (.fluid_in(k_6_41), .fluid_out(k_5_20), .air_in(c_6_1));
valve v_6_42 (.fluid_in(k_6_42), .fluid_out(k_5_21), .air_in(c_6_0));
valve v_6_43 (.fluid_in(k_6_43), .fluid_out(k_5_21), .air_in(c_6_1));
valve v_6_44 (.fluid_in(k_6_44), .fluid_out(k_5_22), .air_in(c_6_0));
valve v_6_45 (.fluid_in(k_6_45), .fluid_out(k_5_22), .air_in(c_6_1));
valve v_6_46 (.fluid_in(k_6_46), .fluid_out(k_5_23), .air_in(c_6_0));
valve v_6_47 (.fluid_in(k_6_47), .fluid_out(k_5_23), .air_in(c_6_1));
valve v_6_48 (.fluid_in(k_6_48), .fluid_out(k_5_24), .air_in(c_6_0));
valve v_6_49 (.fluid_in(k_6_49), .fluid_out(k_5_24), .air_in(c_6_1));
valve v_6_50 (.fluid_in(k_6_50), .fluid_out(k_5_25), .air_in(c_6_0));
valve v_6_51 (.fluid_in(k_6_51), .fluid_out(k_5_25), .air_in(c_6_1));
valve v_6_52 (.fluid_in(k_6_52), .fluid_out(k_5_26), .air_in(c_6_0));
valve v_6_53 (.fluid_in(k_6_53), .fluid_out(k_5_26), .air_in(c_6_1));
valve v_6_54 (.fluid_in(k_6_54), .fluid_out(k_5_27), .air_in(c_6_0));
valve v_6_55 (.fluid_in(k_6_55), .fluid_out(k_5_27), .air_in(c_6_1));
valve v_6_56 (.fluid_in(k_6_56), .fluid_out(k_5_28), .air_in(c_6_0));
valve v_6_57 (.fluid_in(k_6_57), .fluid_out(k_5_28), .air_in(c_6_1));
valve v_6_58 (.fluid_in(k_6_58), .fluid_out(k_5_29), .air_in(c_6_0));
valve v_6_59 (.fluid_in(k_6_59), .fluid_out(k_5_29), .air_in(c_6_1));
valve v_6_60 (.fluid_in(k_6_60), .fluid_out(k_5_30), .air_in(c_6_0));
valve v_6_61 (.fluid_in(k_6_61), .fluid_out(k_5_30), .air_in(c_6_1));
valve v_6_62 (.fluid_in(k_6_62), .fluid_out(k_5_31), .air_in(c_6_0));
valve v_6_63 (.fluid_in(k_6_63), .fluid_out(k_5_31), .air_in(c_6_1));
valve v_7_0 (.fluid_in(k_7_0), .fluid_out(k_6_0), .air_in(c_7_0));
valve v_7_1 (.fluid_in(k_7_1), .fluid_out(k_6_0), .air_in(c_7_1));
valve v_7_2 (.fluid_in(k_7_2), .fluid_out(k_6_1), .air_in(c_7_0));
valve v_7_3 (.fluid_in(k_7_3), .fluid_out(k_6_1), .air_in(c_7_1));
valve v_7_4 (.fluid_in(k_7_4), .fluid_out(k_6_2), .air_in(c_7_0));
valve v_7_5 (.fluid_in(k_7_5), .fluid_out(k_6_2), .air_in(c_7_1));
valve v_7_6 (.fluid_in(k_7_6), .fluid_out(k_6_3), .air_in(c_7_0));
valve v_7_7 (.fluid_in(k_7_7), .fluid_out(k_6_3), .air_in(c_7_1));
valve v_7_8 (.fluid_in(k_7_8), .fluid_out(k_6_4), .air_in(c_7_0));
valve v_7_9 (.fluid_in(k_7_9), .fluid_out(k_6_4), .air_in(c_7_1));
valve v_7_10 (.fluid_in(k_7_10), .fluid_out(k_6_5), .air_in(c_7_0));
valve v_7_11 (.fluid_in(k_7_11), .fluid_out(k_6_5), .air_in(c_7_1));
valve v_7_12 (.fluid_in(k_7_12), .fluid_out(k_6_6), .air_in(c_7_0));
valve v_7_13 (.fluid_in(k_7_13), .fluid_out(k_6_6), .air_in(c_7_1));
valve v_7_14 (.fluid_in(k_7_14), .fluid_out(k_6_7), .air_in(c_7_0));
valve v_7_15 (.fluid_in(k_7_15), .fluid_out(k_6_7), .air_in(c_7_1));
valve v_7_16 (.fluid_in(k_7_16), .fluid_out(k_6_8), .air_in(c_7_0));
valve v_7_17 (.fluid_in(k_7_17), .fluid_out(k_6_8), .air_in(c_7_1));
valve v_7_18 (.fluid_in(k_7_18), .fluid_out(k_6_9), .air_in(c_7_0));
valve v_7_19 (.fluid_in(k_7_19), .fluid_out(k_6_9), .air_in(c_7_1));
valve v_7_20 (.fluid_in(k_7_20), .fluid_out(k_6_10), .air_in(c_7_0));
valve v_7_21 (.fluid_in(k_7_21), .fluid_out(k_6_10), .air_in(c_7_1));
valve v_7_22 (.fluid_in(k_7_22), .fluid_out(k_6_11), .air_in(c_7_0));
valve v_7_23 (.fluid_in(k_7_23), .fluid_out(k_6_11), .air_in(c_7_1));
valve v_7_24 (.fluid_in(k_7_24), .fluid_out(k_6_12), .air_in(c_7_0));
valve v_7_25 (.fluid_in(k_7_25), .fluid_out(k_6_12), .air_in(c_7_1));
valve v_7_26 (.fluid_in(k_7_26), .fluid_out(k_6_13), .air_in(c_7_0));
valve v_7_27 (.fluid_in(k_7_27), .fluid_out(k_6_13), .air_in(c_7_1));
valve v_7_28 (.fluid_in(k_7_28), .fluid_out(k_6_14), .air_in(c_7_0));
valve v_7_29 (.fluid_in(k_7_29), .fluid_out(k_6_14), .air_in(c_7_1));
valve v_7_30 (.fluid_in(k_7_30), .fluid_out(k_6_15), .air_in(c_7_0));
valve v_7_31 (.fluid_in(k_7_31), .fluid_out(k_6_15), .air_in(c_7_1));
valve v_7_32 (.fluid_in(k_7_32), .fluid_out(k_6_16), .air_in(c_7_0));
valve v_7_33 (.fluid_in(k_7_33), .fluid_out(k_6_16), .air_in(c_7_1));
valve v_7_34 (.fluid_in(k_7_34), .fluid_out(k_6_17), .air_in(c_7_0));
valve v_7_35 (.fluid_in(k_7_35), .fluid_out(k_6_17), .air_in(c_7_1));
valve v_7_36 (.fluid_in(k_7_36), .fluid_out(k_6_18), .air_in(c_7_0));
valve v_7_37 (.fluid_in(k_7_37), .fluid_out(k_6_18), .air_in(c_7_1));
valve v_7_38 (.fluid_in(k_7_38), .fluid_out(k_6_19), .air_in(c_7_0));
valve v_7_39 (.fluid_in(k_7_39), .fluid_out(k_6_19), .air_in(c_7_1));
valve v_7_40 (.fluid_in(k_7_40), .fluid_out(k_6_20), .air_in(c_7_0));
valve v_7_41 (.fluid_in(k_7_41), .fluid_out(k_6_20), .air_in(c_7_1));
valve v_7_42 (.fluid_in(k_7_42), .fluid_out(k_6_21), .air_in(c_7_0));
valve v_7_43 (.fluid_in(k_7_43), .fluid_out(k_6_21), .air_in(c_7_1));
valve v_7_44 (.fluid_in(k_7_44), .fluid_out(k_6_22), .air_in(c_7_0));
valve v_7_45 (.fluid_in(k_7_45), .fluid_out(k_6_22), .air_in(c_7_1));
valve v_7_46 (.fluid_in(k_7_46), .fluid_out(k_6_23), .air_in(c_7_0));
valve v_7_47 (.fluid_in(k_7_47), .fluid_out(k_6_23), .air_in(c_7_1));
valve v_7_48 (.fluid_in(k_7_48), .fluid_out(k_6_24), .air_in(c_7_0));
valve v_7_49 (.fluid_in(k_7_49), .fluid_out(k_6_24), .air_in(c_7_1));
valve v_7_50 (.fluid_in(k_7_50), .fluid_out(k_6_25), .air_in(c_7_0));
valve v_7_51 (.fluid_in(k_7_51), .fluid_out(k_6_25), .air_in(c_7_1));
valve v_7_52 (.fluid_in(k_7_52), .fluid_out(k_6_26), .air_in(c_7_0));
valve v_7_53 (.fluid_in(k_7_53), .fluid_out(k_6_26), .air_in(c_7_1));
valve v_7_54 (.fluid_in(k_7_54), .fluid_out(k_6_27), .air_in(c_7_0));
valve v_7_55 (.fluid_in(k_7_55), .fluid_out(k_6_27), .air_in(c_7_1));
valve v_7_56 (.fluid_in(k_7_56), .fluid_out(k_6_28), .air_in(c_7_0));
valve v_7_57 (.fluid_in(k_7_57), .fluid_out(k_6_28), .air_in(c_7_1));
valve v_7_58 (.fluid_in(k_7_58), .fluid_out(k_6_29), .air_in(c_7_0));
valve v_7_59 (.fluid_in(k_7_59), .fluid_out(k_6_29), .air_in(c_7_1));
valve v_7_60 (.fluid_in(k_7_60), .fluid_out(k_6_30), .air_in(c_7_0));
valve v_7_61 (.fluid_in(k_7_61), .fluid_out(k_6_30), .air_in(c_7_1));
valve v_7_62 (.fluid_in(k_7_62), .fluid_out(k_6_31), .air_in(c_7_0));
valve v_7_63 (.fluid_in(k_7_63), .fluid_out(k_6_31), .air_in(c_7_1));
valve v_7_64 (.fluid_in(k_7_64), .fluid_out(k_6_32), .air_in(c_7_0));
valve v_7_65 (.fluid_in(k_7_65), .fluid_out(k_6_32), .air_in(c_7_1));
valve v_7_66 (.fluid_in(k_7_66), .fluid_out(k_6_33), .air_in(c_7_0));
valve v_7_67 (.fluid_in(k_7_67), .fluid_out(k_6_33), .air_in(c_7_1));
valve v_7_68 (.fluid_in(k_7_68), .fluid_out(k_6_34), .air_in(c_7_0));
valve v_7_69 (.fluid_in(k_7_69), .fluid_out(k_6_34), .air_in(c_7_1));
valve v_7_70 (.fluid_in(k_7_70), .fluid_out(k_6_35), .air_in(c_7_0));
valve v_7_71 (.fluid_in(k_7_71), .fluid_out(k_6_35), .air_in(c_7_1));
valve v_7_72 (.fluid_in(k_7_72), .fluid_out(k_6_36), .air_in(c_7_0));
valve v_7_73 (.fluid_in(k_7_73), .fluid_out(k_6_36), .air_in(c_7_1));
valve v_7_74 (.fluid_in(k_7_74), .fluid_out(k_6_37), .air_in(c_7_0));
valve v_7_75 (.fluid_in(k_7_75), .fluid_out(k_6_37), .air_in(c_7_1));
valve v_7_76 (.fluid_in(k_7_76), .fluid_out(k_6_38), .air_in(c_7_0));
valve v_7_77 (.fluid_in(k_7_77), .fluid_out(k_6_38), .air_in(c_7_1));
valve v_7_78 (.fluid_in(k_7_78), .fluid_out(k_6_39), .air_in(c_7_0));
valve v_7_79 (.fluid_in(k_7_79), .fluid_out(k_6_39), .air_in(c_7_1));
valve v_7_80 (.fluid_in(k_7_80), .fluid_out(k_6_40), .air_in(c_7_0));
valve v_7_81 (.fluid_in(k_7_81), .fluid_out(k_6_40), .air_in(c_7_1));
valve v_7_82 (.fluid_in(k_7_82), .fluid_out(k_6_41), .air_in(c_7_0));
valve v_7_83 (.fluid_in(k_7_83), .fluid_out(k_6_41), .air_in(c_7_1));
valve v_7_84 (.fluid_in(k_7_84), .fluid_out(k_6_42), .air_in(c_7_0));
valve v_7_85 (.fluid_in(k_7_85), .fluid_out(k_6_42), .air_in(c_7_1));
valve v_7_86 (.fluid_in(k_7_86), .fluid_out(k_6_43), .air_in(c_7_0));
valve v_7_87 (.fluid_in(k_7_87), .fluid_out(k_6_43), .air_in(c_7_1));
valve v_7_88 (.fluid_in(k_7_88), .fluid_out(k_6_44), .air_in(c_7_0));
valve v_7_89 (.fluid_in(k_7_89), .fluid_out(k_6_44), .air_in(c_7_1));
valve v_7_90 (.fluid_in(k_7_90), .fluid_out(k_6_45), .air_in(c_7_0));
valve v_7_91 (.fluid_in(k_7_91), .fluid_out(k_6_45), .air_in(c_7_1));
valve v_7_92 (.fluid_in(k_7_92), .fluid_out(k_6_46), .air_in(c_7_0));
valve v_7_93 (.fluid_in(k_7_93), .fluid_out(k_6_46), .air_in(c_7_1));
valve v_7_94 (.fluid_in(k_7_94), .fluid_out(k_6_47), .air_in(c_7_0));
valve v_7_95 (.fluid_in(k_7_95), .fluid_out(k_6_47), .air_in(c_7_1));
valve v_7_96 (.fluid_in(k_7_96), .fluid_out(k_6_48), .air_in(c_7_0));
valve v_7_97 (.fluid_in(k_7_97), .fluid_out(k_6_48), .air_in(c_7_1));
valve v_7_98 (.fluid_in(k_7_98), .fluid_out(k_6_49), .air_in(c_7_0));
valve v_7_99 (.fluid_in(k_7_99), .fluid_out(k_6_49), .air_in(c_7_1));
valve v_7_100 (.fluid_in(k_7_100), .fluid_out(k_6_50), .air_in(c_7_0));
valve v_7_101 (.fluid_in(k_7_101), .fluid_out(k_6_50), .air_in(c_7_1));
valve v_7_102 (.fluid_in(k_7_102), .fluid_out(k_6_51), .air_in(c_7_0));
valve v_7_103 (.fluid_in(k_7_103), .fluid_out(k_6_51), .air_in(c_7_1));
valve v_7_104 (.fluid_in(k_7_104), .fluid_out(k_6_52), .air_in(c_7_0));
valve v_7_105 (.fluid_in(k_7_105), .fluid_out(k_6_52), .air_in(c_7_1));
valve v_7_106 (.fluid_in(k_7_106), .fluid_out(k_6_53), .air_in(c_7_0));
valve v_7_107 (.fluid_in(k_7_107), .fluid_out(k_6_53), .air_in(c_7_1));
valve v_7_108 (.fluid_in(k_7_108), .fluid_out(k_6_54), .air_in(c_7_0));
valve v_7_109 (.fluid_in(k_7_109), .fluid_out(k_6_54), .air_in(c_7_1));
valve v_7_110 (.fluid_in(k_7_110), .fluid_out(k_6_55), .air_in(c_7_0));
valve v_7_111 (.fluid_in(k_7_111), .fluid_out(k_6_55), .air_in(c_7_1));
valve v_7_112 (.fluid_in(k_7_112), .fluid_out(k_6_56), .air_in(c_7_0));
valve v_7_113 (.fluid_in(k_7_113), .fluid_out(k_6_56), .air_in(c_7_1));
valve v_7_114 (.fluid_in(k_7_114), .fluid_out(k_6_57), .air_in(c_7_0));
valve v_7_115 (.fluid_in(k_7_115), .fluid_out(k_6_57), .air_in(c_7_1));
valve v_7_116 (.fluid_in(k_7_116), .fluid_out(k_6_58), .air_in(c_7_0));
valve v_7_117 (.fluid_in(k_7_117), .fluid_out(k_6_58), .air_in(c_7_1));
valve v_7_118 (.fluid_in(k_7_118), .fluid_out(k_6_59), .air_in(c_7_0));
valve v_7_119 (.fluid_in(k_7_119), .fluid_out(k_6_59), .air_in(c_7_1));
valve v_7_120 (.fluid_in(k_7_120), .fluid_out(k_6_60), .air_in(c_7_0));
valve v_7_121 (.fluid_in(k_7_121), .fluid_out(k_6_60), .air_in(c_7_1));
valve v_7_122 (.fluid_in(k_7_122), .fluid_out(k_6_61), .air_in(c_7_0));
valve v_7_123 (.fluid_in(k_7_123), .fluid_out(k_6_61), .air_in(c_7_1));
valve v_7_124 (.fluid_in(k_7_124), .fluid_out(k_6_62), .air_in(c_7_0));
valve v_7_125 (.fluid_in(k_7_125), .fluid_out(k_6_62), .air_in(c_7_1));
valve v_7_126 (.fluid_in(k_7_126), .fluid_out(k_6_63), .air_in(c_7_0));
valve v_7_127 (.fluid_in(k_7_127), .fluid_out(k_6_63), .air_in(c_7_1));
endmodule
