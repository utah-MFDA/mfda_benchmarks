module harries();
	mixer m_0(.a(e_0_1), .b(e_0_2), .y(e_0_3));
	mixer m_1(.a(e_0_1), .b(e_1_64), .y(e_1_67));
	mixer m_2(.a(e_0_2), .b(e_2_65), .y(e_2_66));
	mixer m_3(.a(e_0_3), .b(e_3_68), .y(e_3_69));
	mixer m_4(.a(e_4_10), .b(e_4_12), .y(e_4_16));
	mixer m_5(.a(e_5_11), .b(e_5_14), .y(e_5_15));
	mixer m_6(.a(e_6_9), .b(e_6_13), .y(e_6_17));
	mixer m_7(.a(e_7_8), .b(e_7_18), .y(e_7_19));
	mixer m_8(.a(e_7_8), .b(e_8_41), .y(e_8_43));
	mixer m_9(.a(e_6_9), .b(e_9_45), .y(e_9_46));
	mixer m_10(.a(e_4_10), .b(e_10_42), .y(e_10_47));
	mixer m_11(.a(e_5_11), .b(e_11_40), .y(e_11_44));
	mixer m_12(.a(e_4_12), .b(e_12_28), .y(e_12_32));
	mixer m_13(.a(e_6_13), .b(e_13_31), .y(e_13_33));
	mixer m_14(.a(e_5_14), .b(e_14_31), .y(e_14_35));
	mixer m_15(.a(e_5_15), .b(e_15_29), .y(e_15_37));
	mixer m_16(.a(e_4_16), .b(e_16_30), .y(e_16_34));
	mixer m_17(.a(e_6_17), .b(e_17_30), .y(e_17_36));
	mixer m_18(.a(e_7_18), .b(e_18_28), .y(e_18_39));
	mixer m_19(.a(e_7_19), .b(e_19_29), .y(e_19_38));
	mixer m_20(.a(e_20_32), .b(e_20_45), .y(e_20_50));
	mixer m_21(.a(e_21_34), .b(e_21_41), .y(e_21_48));
	mixer m_22(.a(e_22_37), .b(e_22_46), .y(e_22_48));
	mixer m_23(.a(e_23_33), .b(e_23_42), .y(e_23_49));
	mixer m_24(.a(e_24_35), .b(e_24_43), .y(e_24_50));
	mixer m_25(.a(e_25_38), .b(e_25_47), .y(e_25_51));
	mixer m_26(.a(e_26_36), .b(e_26_40), .y(e_26_51));
	mixer m_27(.a(e_27_39), .b(e_27_44), .y(e_27_49));
	mixer m_28(.a(e_12_28), .b(e_18_28), .y(e_28_62));
	mixer m_29(.a(e_15_29), .b(e_19_29), .y(e_29_63));
	mixer m_30(.a(e_16_30), .b(e_17_30), .y(e_30_63));
	mixer m_31(.a(e_13_31), .b(e_14_31), .y(e_31_62));
	mixer m_32(.a(e_12_32), .b(e_20_32), .y(e_32_54));
	mixer m_33(.a(e_13_33), .b(e_23_33), .y(e_33_55));
	mixer m_34(.a(e_16_34), .b(e_21_34), .y(e_34_58));
	mixer m_35(.a(e_14_35), .b(e_24_35), .y(e_35_59));
	mixer m_36(.a(e_17_36), .b(e_26_36), .y(e_36_56));
	mixer m_37(.a(e_15_37), .b(e_22_37), .y(e_37_57));
	mixer m_38(.a(e_19_38), .b(e_25_38), .y(e_38_61));
	mixer m_39(.a(e_18_39), .b(e_27_39), .y(e_39_60));
	mixer m_40(.a(e_11_40), .b(e_26_40), .y(e_40_54));
	mixer m_41(.a(e_8_41), .b(e_21_41), .y(e_41_55));
	mixer m_42(.a(e_10_42), .b(e_23_42), .y(e_42_57));
	mixer m_43(.a(e_8_43), .b(e_24_43), .y(e_43_56));
	mixer m_44(.a(e_11_44), .b(e_27_44), .y(e_44_58));
	mixer m_45(.a(e_9_45), .b(e_20_45), .y(e_45_61));
	mixer m_46(.a(e_9_46), .b(e_22_46), .y(e_46_60));
	mixer m_47(.a(e_10_47), .b(e_25_47), .y(e_47_59));
	mixer m_48(.a(e_21_48), .b(e_22_48), .y(e_48_52));
	mixer m_49(.a(e_23_49), .b(e_27_49), .y(e_49_53));
	mixer m_50(.a(e_20_50), .b(e_24_50), .y(e_50_53));
	mixer m_51(.a(e_25_51), .b(e_26_51), .y(e_51_52));
	mixer m_52(.a(e_48_52), .b(e_51_52), .y(e_52_69));
	mixer m_53(.a(e_49_53), .b(e_50_53), .y(e_53_68));
	mixer m_54(.a(e_32_54), .b(e_40_54), .y(e_54_64));
	mixer m_55(.a(e_33_55), .b(e_41_55), .y(e_55_64));
	mixer m_56(.a(e_36_56), .b(e_43_56), .y(e_56_65));
	mixer m_57(.a(e_37_57), .b(e_42_57), .y(e_57_65));
	mixer m_58(.a(e_34_58), .b(e_44_58), .y(e_58_66));
	mixer m_59(.a(e_35_59), .b(e_47_59), .y(e_59_67));
	mixer m_60(.a(e_39_60), .b(e_46_60), .y(e_60_67));
	mixer m_61(.a(e_38_61), .b(e_45_61), .y(e_61_66));
	mixer m_62(.a(e_28_62), .b(e_31_62), .y(e_62_69));
	mixer m_63(.a(e_29_63), .b(e_30_63), .y(e_63_68));
	mixer m_64(.a(e_1_64), .b(e_54_64), .y(e_55_64));
	mixer m_65(.a(e_2_65), .b(e_56_65), .y(e_57_65));
	mixer m_66(.a(e_2_66), .b(e_58_66), .y(e_61_66));
	mixer m_67(.a(e_1_67), .b(e_59_67), .y(e_60_67));
	mixer m_68(.a(e_3_68), .b(e_53_68), .y(e_63_68));
	mixer m_69(.a(e_3_69), .b(e_52_69), .y(e_62_69));
wire e_0_1,
	e_0_2,
	e_0_3,
	e_1_64,
	e_1_67,
	e_2_65,
	e_2_66,
	e_3_68,
	e_3_69,
	e_4_10,
	e_4_12,
	e_4_16,
	e_5_11,
	e_5_14,
	e_5_15,
	e_6_9,
	e_6_13,
	e_6_17,
	e_7_8,
	e_7_18,
	e_7_19,
	e_8_41,
	e_8_43,
	e_9_45,
	e_9_46,
	e_10_42,
	e_10_47,
	e_11_40,
	e_11_44,
	e_12_28,
	e_12_32,
	e_13_31,
	e_13_33,
	e_14_31,
	e_14_35,
	e_15_29,
	e_15_37,
	e_16_30,
	e_16_34,
	e_17_30,
	e_17_36,
	e_18_28,
	e_18_39,
	e_19_29,
	e_19_38,
	e_20_32,
	e_20_45,
	e_20_50,
	e_21_34,
	e_21_41,
	e_21_48,
	e_22_37,
	e_22_46,
	e_22_48,
	e_23_33,
	e_23_42,
	e_23_49,
	e_24_35,
	e_24_43,
	e_24_50,
	e_25_38,
	e_25_47,
	e_25_51,
	e_26_36,
	e_26_40,
	e_26_51,
	e_27_39,
	e_27_44,
	e_27_49,
	e_28_62,
	e_29_63,
	e_30_63,
	e_31_62,
	e_32_54,
	e_33_55,
	e_34_58,
	e_35_59,
	e_36_56,
	e_37_57,
	e_38_61,
	e_39_60,
	e_40_54,
	e_41_55,
	e_42_57,
	e_43_56,
	e_44_58,
	e_45_61,
	e_46_60,
	e_47_59,
	e_48_52,
	e_49_53,
	e_50_53,
	e_51_52,
	e_52_69,
	e_53_68,
	e_54_64,
	e_55_64,
	e_56_65,
	e_57_65,
	e_58_66,
	e_59_67,
	e_60_67,
	e_61_66,
	e_62_69,
	e_63_68;
endmodule
