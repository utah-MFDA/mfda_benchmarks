module fanout2_mesh_4_3 (
output output_0,output output_1,output output_2,output output_3,input input_0,input input_1,input input_2,input input_3
);
wire output_1_0, output_1_1, output_0_0;
diffmix_25px_0 gate_output_0_0(.a_fluid(output_1_0), .b_fluid(output_1_1), .out_fluid(output_0_0));
wire output_2_0, output_2_1, output_1_0;
diffmix_25px_0 gate_output_1_0(.a_fluid(output_2_0), .b_fluid(output_2_1), .out_fluid(output_1_0));
wire output_3_0, output_3_1, output_2_0;
diffmix_25px_0 gate_output_2_0(.a_fluid(output_3_0), .b_fluid(output_3_1), .out_fluid(output_2_0));
wire output_4_0, output_4_1, output_3_0;
diffmix_25px_0 gate_output_3_0(.a_fluid(output_4_0), .b_fluid(output_4_1), .out_fluid(output_3_0));
wire output_1_1, output_1_2, output_0_1;
diffmix_25px_0 gate_output_0_1(.a_fluid(output_1_1), .b_fluid(output_1_2), .out_fluid(output_0_1));
wire output_2_1, output_2_2, output_1_1;
diffmix_25px_0 gate_output_1_1(.a_fluid(output_2_1), .b_fluid(output_2_2), .out_fluid(output_1_1));
wire output_3_1, output_3_2, output_2_1;
diffmix_25px_0 gate_output_2_1(.a_fluid(output_3_1), .b_fluid(output_3_2), .out_fluid(output_2_1));
wire output_4_1, output_4_2, output_3_1;
diffmix_25px_0 gate_output_3_1(.a_fluid(output_4_1), .b_fluid(output_4_2), .out_fluid(output_3_1));
wire output_1_2, output_1_3, output_0_2;
diffmix_25px_0 gate_output_0_2(.a_fluid(output_1_2), .b_fluid(output_1_3), .out_fluid(output_0_2));
wire output_2_2, output_2_3, output_1_2;
diffmix_25px_0 gate_output_1_2(.a_fluid(output_2_2), .b_fluid(output_2_3), .out_fluid(output_1_2));
wire output_3_2, output_3_3, output_2_2;
diffmix_25px_0 gate_output_2_2(.a_fluid(output_3_2), .b_fluid(output_3_3), .out_fluid(output_2_2));
wire output_4_2, output_4_3, output_3_2;
diffmix_25px_0 gate_output_3_2(.a_fluid(output_4_2), .b_fluid(output_4_3), .out_fluid(output_3_2));
assign output_0 = output_0_0;
wire output_0_3;
assign output_0_3 = input_0;
assign output_1 = output_1_0;
wire output_1_3;
assign output_1_3 = input_1;
assign output_2 = output_2_0;
wire output_2_3;
assign output_2_3 = input_2;
assign output_3 = output_3_0;
wire output_3_3;
assign output_3_3 = input_3;
endmodule
