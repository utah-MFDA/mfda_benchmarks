module binary_tree_1_9 (
output out_0,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63,input input_64,input input_65,input input_66,input input_67,input input_68,input input_69,input input_70,input input_71,input input_72,input input_73,input input_74,input input_75,input input_76,input input_77,input input_78,input input_79,input input_80,input input_81,input input_82,input input_83,input input_84,input input_85,input input_86,input input_87,input input_88,input input_89,input input_90,input input_91,input input_92,input input_93,input input_94,input input_95,input input_96,input input_97,input input_98,input input_99,input input_100,input input_101,input input_102,input input_103,input input_104,input input_105,input input_106,input input_107,input input_108,input input_109,input input_110,input input_111,input input_112,input input_113,input input_114,input input_115,input input_116,input input_117,input input_118,input input_119,input input_120,input input_121,input input_122,input input_123,input input_124,input input_125,input input_126,input input_127,input input_128,input input_129,input input_130,input input_131,input input_132,input input_133,input input_134,input input_135,input input_136,input input_137,input input_138,input input_139,input input_140,input input_141,input input_142,input input_143,input input_144,input input_145,input input_146,input input_147,input input_148,input input_149,input input_150,input input_151,input input_152,input input_153,input input_154,input input_155,input input_156,input input_157,input input_158,input input_159,input input_160,input input_161,input input_162,input input_163,input input_164,input input_165,input input_166,input input_167,input input_168,input input_169,input input_170,input input_171,input input_172,input input_173,input input_174,input input_175,input input_176,input input_177,input input_178,input input_179,input input_180,input input_181,input input_182,input input_183,input input_184,input input_185,input input_186,input input_187,input input_188,input input_189,input input_190,input input_191,input input_192,input input_193,input input_194,input input_195,input input_196,input input_197,input input_198,input input_199,input input_200,input input_201,input input_202,input input_203,input input_204,input input_205,input input_206,input input_207,input input_208,input input_209,input input_210,input input_211,input input_212,input input_213,input input_214,input input_215,input input_216,input input_217,input input_218,input input_219,input input_220,input input_221,input input_222,input input_223,input input_224,input input_225,input input_226,input input_227,input input_228,input input_229,input input_230,input input_231,input input_232,input input_233,input input_234,input input_235,input input_236,input input_237,input input_238,input input_239,input input_240,input input_241,input input_242,input input_243,input input_244,input input_245,input input_246,input input_247,input input_248,input input_249,input input_250,input input_251,input input_252,input input_253,input input_254,input input_255,input input_256,input input_257,input input_258,input input_259,input input_260,input input_261,input input_262,input input_263,input input_264,input input_265,input input_266,input input_267,input input_268,input input_269,input input_270,input input_271,input input_272,input input_273,input input_274,input input_275,input input_276,input input_277,input input_278,input input_279,input input_280,input input_281,input input_282,input input_283,input input_284,input input_285,input input_286,input input_287,input input_288,input input_289,input input_290,input input_291,input input_292,input input_293,input input_294,input input_295,input input_296,input input_297,input input_298,input input_299,input input_300,input input_301,input input_302,input input_303,input input_304,input input_305,input input_306,input input_307,input input_308,input input_309,input input_310,input input_311,input input_312,input input_313,input input_314,input input_315,input input_316,input input_317,input input_318,input input_319,input input_320,input input_321,input input_322,input input_323,input input_324,input input_325,input input_326,input input_327,input input_328,input input_329,input input_330,input input_331,input input_332,input input_333,input input_334,input input_335,input input_336,input input_337,input input_338,input input_339,input input_340,input input_341,input input_342,input input_343,input input_344,input input_345,input input_346,input input_347,input input_348,input input_349,input input_350,input input_351,input input_352,input input_353,input input_354,input input_355,input input_356,input input_357,input input_358,input input_359,input input_360,input input_361,input input_362,input input_363,input input_364,input input_365,input input_366,input input_367,input input_368,input input_369,input input_370,input input_371,input input_372,input input_373,input input_374,input input_375,input input_376,input input_377,input input_378,input input_379,input input_380,input input_381,input input_382,input input_383,input input_384,input input_385,input input_386,input input_387,input input_388,input input_389,input input_390,input input_391,input input_392,input input_393,input input_394,input input_395,input input_396,input input_397,input input_398,input input_399,input input_400,input input_401,input input_402,input input_403,input input_404,input input_405,input input_406,input input_407,input input_408,input input_409,input input_410,input input_411,input input_412,input input_413,input input_414,input input_415,input input_416,input input_417,input input_418,input input_419,input input_420,input input_421,input input_422,input input_423,input input_424,input input_425,input input_426,input input_427,input input_428,input input_429,input input_430,input input_431,input input_432,input input_433,input input_434,input input_435,input input_436,input input_437,input input_438,input input_439,input input_440,input input_441,input input_442,input input_443,input input_444,input input_445,input input_446,input input_447,input input_448,input input_449,input input_450,input input_451,input input_452,input input_453,input input_454,input input_455,input input_456,input input_457,input input_458,input input_459,input input_460,input input_461,input input_462,input input_463,input input_464,input input_465,input input_466,input input_467,input input_468,input input_469,input input_470,input input_471,input input_472,input input_473,input input_474,input input_475,input input_476,input input_477,input input_478,input input_479,input input_480,input input_481,input input_482,input input_483,input input_484,input input_485,input input_486,input input_487,input input_488,input input_489,input input_490,input input_491,input input_492,input input_493,input input_494,input input_495,input input_496,input input_497,input input_498,input input_499,input input_500,input input_501,input input_502,input input_503,input input_504,input input_505,input input_506,input input_507,input input_508,input input_509,input input_510,input input_511
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_000000 (.a(t0_0000000), .b(t0_0000001), .y(t0_000000));
wire t0_0000000, t0_0000001;
mixer mix_t0_0000000 (.a(t0_00000000), .b(t0_00000001), .y(t0_0000000));
wire t0_00000000, t0_00000001;
mixer mix_t0_00000000 (.a(t0_000000000), .b(t0_000000001), .y(t0_00000000));
wire t0_000000000, t0_000000001;
mixer mix_t0_000000000 (.a(t0_0000000000), .b(t0_0000000001), .y(t0_000000000));
wire t0_0000000000, t0_0000000001;
mixer mix_t0_000000001 (.a(t0_0000000010), .b(t0_0000000011), .y(t0_000000001));
wire t0_0000000010, t0_0000000011;
mixer mix_t0_00000001 (.a(t0_000000010), .b(t0_000000011), .y(t0_00000001));
wire t0_000000010, t0_000000011;
mixer mix_t0_000000010 (.a(t0_0000000100), .b(t0_0000000101), .y(t0_000000010));
wire t0_0000000100, t0_0000000101;
mixer mix_t0_000000011 (.a(t0_0000000110), .b(t0_0000000111), .y(t0_000000011));
wire t0_0000000110, t0_0000000111;
mixer mix_t0_0000001 (.a(t0_00000010), .b(t0_00000011), .y(t0_0000001));
wire t0_00000010, t0_00000011;
mixer mix_t0_00000010 (.a(t0_000000100), .b(t0_000000101), .y(t0_00000010));
wire t0_000000100, t0_000000101;
mixer mix_t0_000000100 (.a(t0_0000001000), .b(t0_0000001001), .y(t0_000000100));
wire t0_0000001000, t0_0000001001;
mixer mix_t0_000000101 (.a(t0_0000001010), .b(t0_0000001011), .y(t0_000000101));
wire t0_0000001010, t0_0000001011;
mixer mix_t0_00000011 (.a(t0_000000110), .b(t0_000000111), .y(t0_00000011));
wire t0_000000110, t0_000000111;
mixer mix_t0_000000110 (.a(t0_0000001100), .b(t0_0000001101), .y(t0_000000110));
wire t0_0000001100, t0_0000001101;
mixer mix_t0_000000111 (.a(t0_0000001110), .b(t0_0000001111), .y(t0_000000111));
wire t0_0000001110, t0_0000001111;
mixer mix_t0_000001 (.a(t0_0000010), .b(t0_0000011), .y(t0_000001));
wire t0_0000010, t0_0000011;
mixer mix_t0_0000010 (.a(t0_00000100), .b(t0_00000101), .y(t0_0000010));
wire t0_00000100, t0_00000101;
mixer mix_t0_00000100 (.a(t0_000001000), .b(t0_000001001), .y(t0_00000100));
wire t0_000001000, t0_000001001;
mixer mix_t0_000001000 (.a(t0_0000010000), .b(t0_0000010001), .y(t0_000001000));
wire t0_0000010000, t0_0000010001;
mixer mix_t0_000001001 (.a(t0_0000010010), .b(t0_0000010011), .y(t0_000001001));
wire t0_0000010010, t0_0000010011;
mixer mix_t0_00000101 (.a(t0_000001010), .b(t0_000001011), .y(t0_00000101));
wire t0_000001010, t0_000001011;
mixer mix_t0_000001010 (.a(t0_0000010100), .b(t0_0000010101), .y(t0_000001010));
wire t0_0000010100, t0_0000010101;
mixer mix_t0_000001011 (.a(t0_0000010110), .b(t0_0000010111), .y(t0_000001011));
wire t0_0000010110, t0_0000010111;
mixer mix_t0_0000011 (.a(t0_00000110), .b(t0_00000111), .y(t0_0000011));
wire t0_00000110, t0_00000111;
mixer mix_t0_00000110 (.a(t0_000001100), .b(t0_000001101), .y(t0_00000110));
wire t0_000001100, t0_000001101;
mixer mix_t0_000001100 (.a(t0_0000011000), .b(t0_0000011001), .y(t0_000001100));
wire t0_0000011000, t0_0000011001;
mixer mix_t0_000001101 (.a(t0_0000011010), .b(t0_0000011011), .y(t0_000001101));
wire t0_0000011010, t0_0000011011;
mixer mix_t0_00000111 (.a(t0_000001110), .b(t0_000001111), .y(t0_00000111));
wire t0_000001110, t0_000001111;
mixer mix_t0_000001110 (.a(t0_0000011100), .b(t0_0000011101), .y(t0_000001110));
wire t0_0000011100, t0_0000011101;
mixer mix_t0_000001111 (.a(t0_0000011110), .b(t0_0000011111), .y(t0_000001111));
wire t0_0000011110, t0_0000011111;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_000010 (.a(t0_0000100), .b(t0_0000101), .y(t0_000010));
wire t0_0000100, t0_0000101;
mixer mix_t0_0000100 (.a(t0_00001000), .b(t0_00001001), .y(t0_0000100));
wire t0_00001000, t0_00001001;
mixer mix_t0_00001000 (.a(t0_000010000), .b(t0_000010001), .y(t0_00001000));
wire t0_000010000, t0_000010001;
mixer mix_t0_000010000 (.a(t0_0000100000), .b(t0_0000100001), .y(t0_000010000));
wire t0_0000100000, t0_0000100001;
mixer mix_t0_000010001 (.a(t0_0000100010), .b(t0_0000100011), .y(t0_000010001));
wire t0_0000100010, t0_0000100011;
mixer mix_t0_00001001 (.a(t0_000010010), .b(t0_000010011), .y(t0_00001001));
wire t0_000010010, t0_000010011;
mixer mix_t0_000010010 (.a(t0_0000100100), .b(t0_0000100101), .y(t0_000010010));
wire t0_0000100100, t0_0000100101;
mixer mix_t0_000010011 (.a(t0_0000100110), .b(t0_0000100111), .y(t0_000010011));
wire t0_0000100110, t0_0000100111;
mixer mix_t0_0000101 (.a(t0_00001010), .b(t0_00001011), .y(t0_0000101));
wire t0_00001010, t0_00001011;
mixer mix_t0_00001010 (.a(t0_000010100), .b(t0_000010101), .y(t0_00001010));
wire t0_000010100, t0_000010101;
mixer mix_t0_000010100 (.a(t0_0000101000), .b(t0_0000101001), .y(t0_000010100));
wire t0_0000101000, t0_0000101001;
mixer mix_t0_000010101 (.a(t0_0000101010), .b(t0_0000101011), .y(t0_000010101));
wire t0_0000101010, t0_0000101011;
mixer mix_t0_00001011 (.a(t0_000010110), .b(t0_000010111), .y(t0_00001011));
wire t0_000010110, t0_000010111;
mixer mix_t0_000010110 (.a(t0_0000101100), .b(t0_0000101101), .y(t0_000010110));
wire t0_0000101100, t0_0000101101;
mixer mix_t0_000010111 (.a(t0_0000101110), .b(t0_0000101111), .y(t0_000010111));
wire t0_0000101110, t0_0000101111;
mixer mix_t0_000011 (.a(t0_0000110), .b(t0_0000111), .y(t0_000011));
wire t0_0000110, t0_0000111;
mixer mix_t0_0000110 (.a(t0_00001100), .b(t0_00001101), .y(t0_0000110));
wire t0_00001100, t0_00001101;
mixer mix_t0_00001100 (.a(t0_000011000), .b(t0_000011001), .y(t0_00001100));
wire t0_000011000, t0_000011001;
mixer mix_t0_000011000 (.a(t0_0000110000), .b(t0_0000110001), .y(t0_000011000));
wire t0_0000110000, t0_0000110001;
mixer mix_t0_000011001 (.a(t0_0000110010), .b(t0_0000110011), .y(t0_000011001));
wire t0_0000110010, t0_0000110011;
mixer mix_t0_00001101 (.a(t0_000011010), .b(t0_000011011), .y(t0_00001101));
wire t0_000011010, t0_000011011;
mixer mix_t0_000011010 (.a(t0_0000110100), .b(t0_0000110101), .y(t0_000011010));
wire t0_0000110100, t0_0000110101;
mixer mix_t0_000011011 (.a(t0_0000110110), .b(t0_0000110111), .y(t0_000011011));
wire t0_0000110110, t0_0000110111;
mixer mix_t0_0000111 (.a(t0_00001110), .b(t0_00001111), .y(t0_0000111));
wire t0_00001110, t0_00001111;
mixer mix_t0_00001110 (.a(t0_000011100), .b(t0_000011101), .y(t0_00001110));
wire t0_000011100, t0_000011101;
mixer mix_t0_000011100 (.a(t0_0000111000), .b(t0_0000111001), .y(t0_000011100));
wire t0_0000111000, t0_0000111001;
mixer mix_t0_000011101 (.a(t0_0000111010), .b(t0_0000111011), .y(t0_000011101));
wire t0_0000111010, t0_0000111011;
mixer mix_t0_00001111 (.a(t0_000011110), .b(t0_000011111), .y(t0_00001111));
wire t0_000011110, t0_000011111;
mixer mix_t0_000011110 (.a(t0_0000111100), .b(t0_0000111101), .y(t0_000011110));
wire t0_0000111100, t0_0000111101;
mixer mix_t0_000011111 (.a(t0_0000111110), .b(t0_0000111111), .y(t0_000011111));
wire t0_0000111110, t0_0000111111;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_000100 (.a(t0_0001000), .b(t0_0001001), .y(t0_000100));
wire t0_0001000, t0_0001001;
mixer mix_t0_0001000 (.a(t0_00010000), .b(t0_00010001), .y(t0_0001000));
wire t0_00010000, t0_00010001;
mixer mix_t0_00010000 (.a(t0_000100000), .b(t0_000100001), .y(t0_00010000));
wire t0_000100000, t0_000100001;
mixer mix_t0_000100000 (.a(t0_0001000000), .b(t0_0001000001), .y(t0_000100000));
wire t0_0001000000, t0_0001000001;
mixer mix_t0_000100001 (.a(t0_0001000010), .b(t0_0001000011), .y(t0_000100001));
wire t0_0001000010, t0_0001000011;
mixer mix_t0_00010001 (.a(t0_000100010), .b(t0_000100011), .y(t0_00010001));
wire t0_000100010, t0_000100011;
mixer mix_t0_000100010 (.a(t0_0001000100), .b(t0_0001000101), .y(t0_000100010));
wire t0_0001000100, t0_0001000101;
mixer mix_t0_000100011 (.a(t0_0001000110), .b(t0_0001000111), .y(t0_000100011));
wire t0_0001000110, t0_0001000111;
mixer mix_t0_0001001 (.a(t0_00010010), .b(t0_00010011), .y(t0_0001001));
wire t0_00010010, t0_00010011;
mixer mix_t0_00010010 (.a(t0_000100100), .b(t0_000100101), .y(t0_00010010));
wire t0_000100100, t0_000100101;
mixer mix_t0_000100100 (.a(t0_0001001000), .b(t0_0001001001), .y(t0_000100100));
wire t0_0001001000, t0_0001001001;
mixer mix_t0_000100101 (.a(t0_0001001010), .b(t0_0001001011), .y(t0_000100101));
wire t0_0001001010, t0_0001001011;
mixer mix_t0_00010011 (.a(t0_000100110), .b(t0_000100111), .y(t0_00010011));
wire t0_000100110, t0_000100111;
mixer mix_t0_000100110 (.a(t0_0001001100), .b(t0_0001001101), .y(t0_000100110));
wire t0_0001001100, t0_0001001101;
mixer mix_t0_000100111 (.a(t0_0001001110), .b(t0_0001001111), .y(t0_000100111));
wire t0_0001001110, t0_0001001111;
mixer mix_t0_000101 (.a(t0_0001010), .b(t0_0001011), .y(t0_000101));
wire t0_0001010, t0_0001011;
mixer mix_t0_0001010 (.a(t0_00010100), .b(t0_00010101), .y(t0_0001010));
wire t0_00010100, t0_00010101;
mixer mix_t0_00010100 (.a(t0_000101000), .b(t0_000101001), .y(t0_00010100));
wire t0_000101000, t0_000101001;
mixer mix_t0_000101000 (.a(t0_0001010000), .b(t0_0001010001), .y(t0_000101000));
wire t0_0001010000, t0_0001010001;
mixer mix_t0_000101001 (.a(t0_0001010010), .b(t0_0001010011), .y(t0_000101001));
wire t0_0001010010, t0_0001010011;
mixer mix_t0_00010101 (.a(t0_000101010), .b(t0_000101011), .y(t0_00010101));
wire t0_000101010, t0_000101011;
mixer mix_t0_000101010 (.a(t0_0001010100), .b(t0_0001010101), .y(t0_000101010));
wire t0_0001010100, t0_0001010101;
mixer mix_t0_000101011 (.a(t0_0001010110), .b(t0_0001010111), .y(t0_000101011));
wire t0_0001010110, t0_0001010111;
mixer mix_t0_0001011 (.a(t0_00010110), .b(t0_00010111), .y(t0_0001011));
wire t0_00010110, t0_00010111;
mixer mix_t0_00010110 (.a(t0_000101100), .b(t0_000101101), .y(t0_00010110));
wire t0_000101100, t0_000101101;
mixer mix_t0_000101100 (.a(t0_0001011000), .b(t0_0001011001), .y(t0_000101100));
wire t0_0001011000, t0_0001011001;
mixer mix_t0_000101101 (.a(t0_0001011010), .b(t0_0001011011), .y(t0_000101101));
wire t0_0001011010, t0_0001011011;
mixer mix_t0_00010111 (.a(t0_000101110), .b(t0_000101111), .y(t0_00010111));
wire t0_000101110, t0_000101111;
mixer mix_t0_000101110 (.a(t0_0001011100), .b(t0_0001011101), .y(t0_000101110));
wire t0_0001011100, t0_0001011101;
mixer mix_t0_000101111 (.a(t0_0001011110), .b(t0_0001011111), .y(t0_000101111));
wire t0_0001011110, t0_0001011111;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_000110 (.a(t0_0001100), .b(t0_0001101), .y(t0_000110));
wire t0_0001100, t0_0001101;
mixer mix_t0_0001100 (.a(t0_00011000), .b(t0_00011001), .y(t0_0001100));
wire t0_00011000, t0_00011001;
mixer mix_t0_00011000 (.a(t0_000110000), .b(t0_000110001), .y(t0_00011000));
wire t0_000110000, t0_000110001;
mixer mix_t0_000110000 (.a(t0_0001100000), .b(t0_0001100001), .y(t0_000110000));
wire t0_0001100000, t0_0001100001;
mixer mix_t0_000110001 (.a(t0_0001100010), .b(t0_0001100011), .y(t0_000110001));
wire t0_0001100010, t0_0001100011;
mixer mix_t0_00011001 (.a(t0_000110010), .b(t0_000110011), .y(t0_00011001));
wire t0_000110010, t0_000110011;
mixer mix_t0_000110010 (.a(t0_0001100100), .b(t0_0001100101), .y(t0_000110010));
wire t0_0001100100, t0_0001100101;
mixer mix_t0_000110011 (.a(t0_0001100110), .b(t0_0001100111), .y(t0_000110011));
wire t0_0001100110, t0_0001100111;
mixer mix_t0_0001101 (.a(t0_00011010), .b(t0_00011011), .y(t0_0001101));
wire t0_00011010, t0_00011011;
mixer mix_t0_00011010 (.a(t0_000110100), .b(t0_000110101), .y(t0_00011010));
wire t0_000110100, t0_000110101;
mixer mix_t0_000110100 (.a(t0_0001101000), .b(t0_0001101001), .y(t0_000110100));
wire t0_0001101000, t0_0001101001;
mixer mix_t0_000110101 (.a(t0_0001101010), .b(t0_0001101011), .y(t0_000110101));
wire t0_0001101010, t0_0001101011;
mixer mix_t0_00011011 (.a(t0_000110110), .b(t0_000110111), .y(t0_00011011));
wire t0_000110110, t0_000110111;
mixer mix_t0_000110110 (.a(t0_0001101100), .b(t0_0001101101), .y(t0_000110110));
wire t0_0001101100, t0_0001101101;
mixer mix_t0_000110111 (.a(t0_0001101110), .b(t0_0001101111), .y(t0_000110111));
wire t0_0001101110, t0_0001101111;
mixer mix_t0_000111 (.a(t0_0001110), .b(t0_0001111), .y(t0_000111));
wire t0_0001110, t0_0001111;
mixer mix_t0_0001110 (.a(t0_00011100), .b(t0_00011101), .y(t0_0001110));
wire t0_00011100, t0_00011101;
mixer mix_t0_00011100 (.a(t0_000111000), .b(t0_000111001), .y(t0_00011100));
wire t0_000111000, t0_000111001;
mixer mix_t0_000111000 (.a(t0_0001110000), .b(t0_0001110001), .y(t0_000111000));
wire t0_0001110000, t0_0001110001;
mixer mix_t0_000111001 (.a(t0_0001110010), .b(t0_0001110011), .y(t0_000111001));
wire t0_0001110010, t0_0001110011;
mixer mix_t0_00011101 (.a(t0_000111010), .b(t0_000111011), .y(t0_00011101));
wire t0_000111010, t0_000111011;
mixer mix_t0_000111010 (.a(t0_0001110100), .b(t0_0001110101), .y(t0_000111010));
wire t0_0001110100, t0_0001110101;
mixer mix_t0_000111011 (.a(t0_0001110110), .b(t0_0001110111), .y(t0_000111011));
wire t0_0001110110, t0_0001110111;
mixer mix_t0_0001111 (.a(t0_00011110), .b(t0_00011111), .y(t0_0001111));
wire t0_00011110, t0_00011111;
mixer mix_t0_00011110 (.a(t0_000111100), .b(t0_000111101), .y(t0_00011110));
wire t0_000111100, t0_000111101;
mixer mix_t0_000111100 (.a(t0_0001111000), .b(t0_0001111001), .y(t0_000111100));
wire t0_0001111000, t0_0001111001;
mixer mix_t0_000111101 (.a(t0_0001111010), .b(t0_0001111011), .y(t0_000111101));
wire t0_0001111010, t0_0001111011;
mixer mix_t0_00011111 (.a(t0_000111110), .b(t0_000111111), .y(t0_00011111));
wire t0_000111110, t0_000111111;
mixer mix_t0_000111110 (.a(t0_0001111100), .b(t0_0001111101), .y(t0_000111110));
wire t0_0001111100, t0_0001111101;
mixer mix_t0_000111111 (.a(t0_0001111110), .b(t0_0001111111), .y(t0_000111111));
wire t0_0001111110, t0_0001111111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_001000 (.a(t0_0010000), .b(t0_0010001), .y(t0_001000));
wire t0_0010000, t0_0010001;
mixer mix_t0_0010000 (.a(t0_00100000), .b(t0_00100001), .y(t0_0010000));
wire t0_00100000, t0_00100001;
mixer mix_t0_00100000 (.a(t0_001000000), .b(t0_001000001), .y(t0_00100000));
wire t0_001000000, t0_001000001;
mixer mix_t0_001000000 (.a(t0_0010000000), .b(t0_0010000001), .y(t0_001000000));
wire t0_0010000000, t0_0010000001;
mixer mix_t0_001000001 (.a(t0_0010000010), .b(t0_0010000011), .y(t0_001000001));
wire t0_0010000010, t0_0010000011;
mixer mix_t0_00100001 (.a(t0_001000010), .b(t0_001000011), .y(t0_00100001));
wire t0_001000010, t0_001000011;
mixer mix_t0_001000010 (.a(t0_0010000100), .b(t0_0010000101), .y(t0_001000010));
wire t0_0010000100, t0_0010000101;
mixer mix_t0_001000011 (.a(t0_0010000110), .b(t0_0010000111), .y(t0_001000011));
wire t0_0010000110, t0_0010000111;
mixer mix_t0_0010001 (.a(t0_00100010), .b(t0_00100011), .y(t0_0010001));
wire t0_00100010, t0_00100011;
mixer mix_t0_00100010 (.a(t0_001000100), .b(t0_001000101), .y(t0_00100010));
wire t0_001000100, t0_001000101;
mixer mix_t0_001000100 (.a(t0_0010001000), .b(t0_0010001001), .y(t0_001000100));
wire t0_0010001000, t0_0010001001;
mixer mix_t0_001000101 (.a(t0_0010001010), .b(t0_0010001011), .y(t0_001000101));
wire t0_0010001010, t0_0010001011;
mixer mix_t0_00100011 (.a(t0_001000110), .b(t0_001000111), .y(t0_00100011));
wire t0_001000110, t0_001000111;
mixer mix_t0_001000110 (.a(t0_0010001100), .b(t0_0010001101), .y(t0_001000110));
wire t0_0010001100, t0_0010001101;
mixer mix_t0_001000111 (.a(t0_0010001110), .b(t0_0010001111), .y(t0_001000111));
wire t0_0010001110, t0_0010001111;
mixer mix_t0_001001 (.a(t0_0010010), .b(t0_0010011), .y(t0_001001));
wire t0_0010010, t0_0010011;
mixer mix_t0_0010010 (.a(t0_00100100), .b(t0_00100101), .y(t0_0010010));
wire t0_00100100, t0_00100101;
mixer mix_t0_00100100 (.a(t0_001001000), .b(t0_001001001), .y(t0_00100100));
wire t0_001001000, t0_001001001;
mixer mix_t0_001001000 (.a(t0_0010010000), .b(t0_0010010001), .y(t0_001001000));
wire t0_0010010000, t0_0010010001;
mixer mix_t0_001001001 (.a(t0_0010010010), .b(t0_0010010011), .y(t0_001001001));
wire t0_0010010010, t0_0010010011;
mixer mix_t0_00100101 (.a(t0_001001010), .b(t0_001001011), .y(t0_00100101));
wire t0_001001010, t0_001001011;
mixer mix_t0_001001010 (.a(t0_0010010100), .b(t0_0010010101), .y(t0_001001010));
wire t0_0010010100, t0_0010010101;
mixer mix_t0_001001011 (.a(t0_0010010110), .b(t0_0010010111), .y(t0_001001011));
wire t0_0010010110, t0_0010010111;
mixer mix_t0_0010011 (.a(t0_00100110), .b(t0_00100111), .y(t0_0010011));
wire t0_00100110, t0_00100111;
mixer mix_t0_00100110 (.a(t0_001001100), .b(t0_001001101), .y(t0_00100110));
wire t0_001001100, t0_001001101;
mixer mix_t0_001001100 (.a(t0_0010011000), .b(t0_0010011001), .y(t0_001001100));
wire t0_0010011000, t0_0010011001;
mixer mix_t0_001001101 (.a(t0_0010011010), .b(t0_0010011011), .y(t0_001001101));
wire t0_0010011010, t0_0010011011;
mixer mix_t0_00100111 (.a(t0_001001110), .b(t0_001001111), .y(t0_00100111));
wire t0_001001110, t0_001001111;
mixer mix_t0_001001110 (.a(t0_0010011100), .b(t0_0010011101), .y(t0_001001110));
wire t0_0010011100, t0_0010011101;
mixer mix_t0_001001111 (.a(t0_0010011110), .b(t0_0010011111), .y(t0_001001111));
wire t0_0010011110, t0_0010011111;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_001010 (.a(t0_0010100), .b(t0_0010101), .y(t0_001010));
wire t0_0010100, t0_0010101;
mixer mix_t0_0010100 (.a(t0_00101000), .b(t0_00101001), .y(t0_0010100));
wire t0_00101000, t0_00101001;
mixer mix_t0_00101000 (.a(t0_001010000), .b(t0_001010001), .y(t0_00101000));
wire t0_001010000, t0_001010001;
mixer mix_t0_001010000 (.a(t0_0010100000), .b(t0_0010100001), .y(t0_001010000));
wire t0_0010100000, t0_0010100001;
mixer mix_t0_001010001 (.a(t0_0010100010), .b(t0_0010100011), .y(t0_001010001));
wire t0_0010100010, t0_0010100011;
mixer mix_t0_00101001 (.a(t0_001010010), .b(t0_001010011), .y(t0_00101001));
wire t0_001010010, t0_001010011;
mixer mix_t0_001010010 (.a(t0_0010100100), .b(t0_0010100101), .y(t0_001010010));
wire t0_0010100100, t0_0010100101;
mixer mix_t0_001010011 (.a(t0_0010100110), .b(t0_0010100111), .y(t0_001010011));
wire t0_0010100110, t0_0010100111;
mixer mix_t0_0010101 (.a(t0_00101010), .b(t0_00101011), .y(t0_0010101));
wire t0_00101010, t0_00101011;
mixer mix_t0_00101010 (.a(t0_001010100), .b(t0_001010101), .y(t0_00101010));
wire t0_001010100, t0_001010101;
mixer mix_t0_001010100 (.a(t0_0010101000), .b(t0_0010101001), .y(t0_001010100));
wire t0_0010101000, t0_0010101001;
mixer mix_t0_001010101 (.a(t0_0010101010), .b(t0_0010101011), .y(t0_001010101));
wire t0_0010101010, t0_0010101011;
mixer mix_t0_00101011 (.a(t0_001010110), .b(t0_001010111), .y(t0_00101011));
wire t0_001010110, t0_001010111;
mixer mix_t0_001010110 (.a(t0_0010101100), .b(t0_0010101101), .y(t0_001010110));
wire t0_0010101100, t0_0010101101;
mixer mix_t0_001010111 (.a(t0_0010101110), .b(t0_0010101111), .y(t0_001010111));
wire t0_0010101110, t0_0010101111;
mixer mix_t0_001011 (.a(t0_0010110), .b(t0_0010111), .y(t0_001011));
wire t0_0010110, t0_0010111;
mixer mix_t0_0010110 (.a(t0_00101100), .b(t0_00101101), .y(t0_0010110));
wire t0_00101100, t0_00101101;
mixer mix_t0_00101100 (.a(t0_001011000), .b(t0_001011001), .y(t0_00101100));
wire t0_001011000, t0_001011001;
mixer mix_t0_001011000 (.a(t0_0010110000), .b(t0_0010110001), .y(t0_001011000));
wire t0_0010110000, t0_0010110001;
mixer mix_t0_001011001 (.a(t0_0010110010), .b(t0_0010110011), .y(t0_001011001));
wire t0_0010110010, t0_0010110011;
mixer mix_t0_00101101 (.a(t0_001011010), .b(t0_001011011), .y(t0_00101101));
wire t0_001011010, t0_001011011;
mixer mix_t0_001011010 (.a(t0_0010110100), .b(t0_0010110101), .y(t0_001011010));
wire t0_0010110100, t0_0010110101;
mixer mix_t0_001011011 (.a(t0_0010110110), .b(t0_0010110111), .y(t0_001011011));
wire t0_0010110110, t0_0010110111;
mixer mix_t0_0010111 (.a(t0_00101110), .b(t0_00101111), .y(t0_0010111));
wire t0_00101110, t0_00101111;
mixer mix_t0_00101110 (.a(t0_001011100), .b(t0_001011101), .y(t0_00101110));
wire t0_001011100, t0_001011101;
mixer mix_t0_001011100 (.a(t0_0010111000), .b(t0_0010111001), .y(t0_001011100));
wire t0_0010111000, t0_0010111001;
mixer mix_t0_001011101 (.a(t0_0010111010), .b(t0_0010111011), .y(t0_001011101));
wire t0_0010111010, t0_0010111011;
mixer mix_t0_00101111 (.a(t0_001011110), .b(t0_001011111), .y(t0_00101111));
wire t0_001011110, t0_001011111;
mixer mix_t0_001011110 (.a(t0_0010111100), .b(t0_0010111101), .y(t0_001011110));
wire t0_0010111100, t0_0010111101;
mixer mix_t0_001011111 (.a(t0_0010111110), .b(t0_0010111111), .y(t0_001011111));
wire t0_0010111110, t0_0010111111;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_001100 (.a(t0_0011000), .b(t0_0011001), .y(t0_001100));
wire t0_0011000, t0_0011001;
mixer mix_t0_0011000 (.a(t0_00110000), .b(t0_00110001), .y(t0_0011000));
wire t0_00110000, t0_00110001;
mixer mix_t0_00110000 (.a(t0_001100000), .b(t0_001100001), .y(t0_00110000));
wire t0_001100000, t0_001100001;
mixer mix_t0_001100000 (.a(t0_0011000000), .b(t0_0011000001), .y(t0_001100000));
wire t0_0011000000, t0_0011000001;
mixer mix_t0_001100001 (.a(t0_0011000010), .b(t0_0011000011), .y(t0_001100001));
wire t0_0011000010, t0_0011000011;
mixer mix_t0_00110001 (.a(t0_001100010), .b(t0_001100011), .y(t0_00110001));
wire t0_001100010, t0_001100011;
mixer mix_t0_001100010 (.a(t0_0011000100), .b(t0_0011000101), .y(t0_001100010));
wire t0_0011000100, t0_0011000101;
mixer mix_t0_001100011 (.a(t0_0011000110), .b(t0_0011000111), .y(t0_001100011));
wire t0_0011000110, t0_0011000111;
mixer mix_t0_0011001 (.a(t0_00110010), .b(t0_00110011), .y(t0_0011001));
wire t0_00110010, t0_00110011;
mixer mix_t0_00110010 (.a(t0_001100100), .b(t0_001100101), .y(t0_00110010));
wire t0_001100100, t0_001100101;
mixer mix_t0_001100100 (.a(t0_0011001000), .b(t0_0011001001), .y(t0_001100100));
wire t0_0011001000, t0_0011001001;
mixer mix_t0_001100101 (.a(t0_0011001010), .b(t0_0011001011), .y(t0_001100101));
wire t0_0011001010, t0_0011001011;
mixer mix_t0_00110011 (.a(t0_001100110), .b(t0_001100111), .y(t0_00110011));
wire t0_001100110, t0_001100111;
mixer mix_t0_001100110 (.a(t0_0011001100), .b(t0_0011001101), .y(t0_001100110));
wire t0_0011001100, t0_0011001101;
mixer mix_t0_001100111 (.a(t0_0011001110), .b(t0_0011001111), .y(t0_001100111));
wire t0_0011001110, t0_0011001111;
mixer mix_t0_001101 (.a(t0_0011010), .b(t0_0011011), .y(t0_001101));
wire t0_0011010, t0_0011011;
mixer mix_t0_0011010 (.a(t0_00110100), .b(t0_00110101), .y(t0_0011010));
wire t0_00110100, t0_00110101;
mixer mix_t0_00110100 (.a(t0_001101000), .b(t0_001101001), .y(t0_00110100));
wire t0_001101000, t0_001101001;
mixer mix_t0_001101000 (.a(t0_0011010000), .b(t0_0011010001), .y(t0_001101000));
wire t0_0011010000, t0_0011010001;
mixer mix_t0_001101001 (.a(t0_0011010010), .b(t0_0011010011), .y(t0_001101001));
wire t0_0011010010, t0_0011010011;
mixer mix_t0_00110101 (.a(t0_001101010), .b(t0_001101011), .y(t0_00110101));
wire t0_001101010, t0_001101011;
mixer mix_t0_001101010 (.a(t0_0011010100), .b(t0_0011010101), .y(t0_001101010));
wire t0_0011010100, t0_0011010101;
mixer mix_t0_001101011 (.a(t0_0011010110), .b(t0_0011010111), .y(t0_001101011));
wire t0_0011010110, t0_0011010111;
mixer mix_t0_0011011 (.a(t0_00110110), .b(t0_00110111), .y(t0_0011011));
wire t0_00110110, t0_00110111;
mixer mix_t0_00110110 (.a(t0_001101100), .b(t0_001101101), .y(t0_00110110));
wire t0_001101100, t0_001101101;
mixer mix_t0_001101100 (.a(t0_0011011000), .b(t0_0011011001), .y(t0_001101100));
wire t0_0011011000, t0_0011011001;
mixer mix_t0_001101101 (.a(t0_0011011010), .b(t0_0011011011), .y(t0_001101101));
wire t0_0011011010, t0_0011011011;
mixer mix_t0_00110111 (.a(t0_001101110), .b(t0_001101111), .y(t0_00110111));
wire t0_001101110, t0_001101111;
mixer mix_t0_001101110 (.a(t0_0011011100), .b(t0_0011011101), .y(t0_001101110));
wire t0_0011011100, t0_0011011101;
mixer mix_t0_001101111 (.a(t0_0011011110), .b(t0_0011011111), .y(t0_001101111));
wire t0_0011011110, t0_0011011111;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_001110 (.a(t0_0011100), .b(t0_0011101), .y(t0_001110));
wire t0_0011100, t0_0011101;
mixer mix_t0_0011100 (.a(t0_00111000), .b(t0_00111001), .y(t0_0011100));
wire t0_00111000, t0_00111001;
mixer mix_t0_00111000 (.a(t0_001110000), .b(t0_001110001), .y(t0_00111000));
wire t0_001110000, t0_001110001;
mixer mix_t0_001110000 (.a(t0_0011100000), .b(t0_0011100001), .y(t0_001110000));
wire t0_0011100000, t0_0011100001;
mixer mix_t0_001110001 (.a(t0_0011100010), .b(t0_0011100011), .y(t0_001110001));
wire t0_0011100010, t0_0011100011;
mixer mix_t0_00111001 (.a(t0_001110010), .b(t0_001110011), .y(t0_00111001));
wire t0_001110010, t0_001110011;
mixer mix_t0_001110010 (.a(t0_0011100100), .b(t0_0011100101), .y(t0_001110010));
wire t0_0011100100, t0_0011100101;
mixer mix_t0_001110011 (.a(t0_0011100110), .b(t0_0011100111), .y(t0_001110011));
wire t0_0011100110, t0_0011100111;
mixer mix_t0_0011101 (.a(t0_00111010), .b(t0_00111011), .y(t0_0011101));
wire t0_00111010, t0_00111011;
mixer mix_t0_00111010 (.a(t0_001110100), .b(t0_001110101), .y(t0_00111010));
wire t0_001110100, t0_001110101;
mixer mix_t0_001110100 (.a(t0_0011101000), .b(t0_0011101001), .y(t0_001110100));
wire t0_0011101000, t0_0011101001;
mixer mix_t0_001110101 (.a(t0_0011101010), .b(t0_0011101011), .y(t0_001110101));
wire t0_0011101010, t0_0011101011;
mixer mix_t0_00111011 (.a(t0_001110110), .b(t0_001110111), .y(t0_00111011));
wire t0_001110110, t0_001110111;
mixer mix_t0_001110110 (.a(t0_0011101100), .b(t0_0011101101), .y(t0_001110110));
wire t0_0011101100, t0_0011101101;
mixer mix_t0_001110111 (.a(t0_0011101110), .b(t0_0011101111), .y(t0_001110111));
wire t0_0011101110, t0_0011101111;
mixer mix_t0_001111 (.a(t0_0011110), .b(t0_0011111), .y(t0_001111));
wire t0_0011110, t0_0011111;
mixer mix_t0_0011110 (.a(t0_00111100), .b(t0_00111101), .y(t0_0011110));
wire t0_00111100, t0_00111101;
mixer mix_t0_00111100 (.a(t0_001111000), .b(t0_001111001), .y(t0_00111100));
wire t0_001111000, t0_001111001;
mixer mix_t0_001111000 (.a(t0_0011110000), .b(t0_0011110001), .y(t0_001111000));
wire t0_0011110000, t0_0011110001;
mixer mix_t0_001111001 (.a(t0_0011110010), .b(t0_0011110011), .y(t0_001111001));
wire t0_0011110010, t0_0011110011;
mixer mix_t0_00111101 (.a(t0_001111010), .b(t0_001111011), .y(t0_00111101));
wire t0_001111010, t0_001111011;
mixer mix_t0_001111010 (.a(t0_0011110100), .b(t0_0011110101), .y(t0_001111010));
wire t0_0011110100, t0_0011110101;
mixer mix_t0_001111011 (.a(t0_0011110110), .b(t0_0011110111), .y(t0_001111011));
wire t0_0011110110, t0_0011110111;
mixer mix_t0_0011111 (.a(t0_00111110), .b(t0_00111111), .y(t0_0011111));
wire t0_00111110, t0_00111111;
mixer mix_t0_00111110 (.a(t0_001111100), .b(t0_001111101), .y(t0_00111110));
wire t0_001111100, t0_001111101;
mixer mix_t0_001111100 (.a(t0_0011111000), .b(t0_0011111001), .y(t0_001111100));
wire t0_0011111000, t0_0011111001;
mixer mix_t0_001111101 (.a(t0_0011111010), .b(t0_0011111011), .y(t0_001111101));
wire t0_0011111010, t0_0011111011;
mixer mix_t0_00111111 (.a(t0_001111110), .b(t0_001111111), .y(t0_00111111));
wire t0_001111110, t0_001111111;
mixer mix_t0_001111110 (.a(t0_0011111100), .b(t0_0011111101), .y(t0_001111110));
wire t0_0011111100, t0_0011111101;
mixer mix_t0_001111111 (.a(t0_0011111110), .b(t0_0011111111), .y(t0_001111111));
wire t0_0011111110, t0_0011111111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_010000 (.a(t0_0100000), .b(t0_0100001), .y(t0_010000));
wire t0_0100000, t0_0100001;
mixer mix_t0_0100000 (.a(t0_01000000), .b(t0_01000001), .y(t0_0100000));
wire t0_01000000, t0_01000001;
mixer mix_t0_01000000 (.a(t0_010000000), .b(t0_010000001), .y(t0_01000000));
wire t0_010000000, t0_010000001;
mixer mix_t0_010000000 (.a(t0_0100000000), .b(t0_0100000001), .y(t0_010000000));
wire t0_0100000000, t0_0100000001;
mixer mix_t0_010000001 (.a(t0_0100000010), .b(t0_0100000011), .y(t0_010000001));
wire t0_0100000010, t0_0100000011;
mixer mix_t0_01000001 (.a(t0_010000010), .b(t0_010000011), .y(t0_01000001));
wire t0_010000010, t0_010000011;
mixer mix_t0_010000010 (.a(t0_0100000100), .b(t0_0100000101), .y(t0_010000010));
wire t0_0100000100, t0_0100000101;
mixer mix_t0_010000011 (.a(t0_0100000110), .b(t0_0100000111), .y(t0_010000011));
wire t0_0100000110, t0_0100000111;
mixer mix_t0_0100001 (.a(t0_01000010), .b(t0_01000011), .y(t0_0100001));
wire t0_01000010, t0_01000011;
mixer mix_t0_01000010 (.a(t0_010000100), .b(t0_010000101), .y(t0_01000010));
wire t0_010000100, t0_010000101;
mixer mix_t0_010000100 (.a(t0_0100001000), .b(t0_0100001001), .y(t0_010000100));
wire t0_0100001000, t0_0100001001;
mixer mix_t0_010000101 (.a(t0_0100001010), .b(t0_0100001011), .y(t0_010000101));
wire t0_0100001010, t0_0100001011;
mixer mix_t0_01000011 (.a(t0_010000110), .b(t0_010000111), .y(t0_01000011));
wire t0_010000110, t0_010000111;
mixer mix_t0_010000110 (.a(t0_0100001100), .b(t0_0100001101), .y(t0_010000110));
wire t0_0100001100, t0_0100001101;
mixer mix_t0_010000111 (.a(t0_0100001110), .b(t0_0100001111), .y(t0_010000111));
wire t0_0100001110, t0_0100001111;
mixer mix_t0_010001 (.a(t0_0100010), .b(t0_0100011), .y(t0_010001));
wire t0_0100010, t0_0100011;
mixer mix_t0_0100010 (.a(t0_01000100), .b(t0_01000101), .y(t0_0100010));
wire t0_01000100, t0_01000101;
mixer mix_t0_01000100 (.a(t0_010001000), .b(t0_010001001), .y(t0_01000100));
wire t0_010001000, t0_010001001;
mixer mix_t0_010001000 (.a(t0_0100010000), .b(t0_0100010001), .y(t0_010001000));
wire t0_0100010000, t0_0100010001;
mixer mix_t0_010001001 (.a(t0_0100010010), .b(t0_0100010011), .y(t0_010001001));
wire t0_0100010010, t0_0100010011;
mixer mix_t0_01000101 (.a(t0_010001010), .b(t0_010001011), .y(t0_01000101));
wire t0_010001010, t0_010001011;
mixer mix_t0_010001010 (.a(t0_0100010100), .b(t0_0100010101), .y(t0_010001010));
wire t0_0100010100, t0_0100010101;
mixer mix_t0_010001011 (.a(t0_0100010110), .b(t0_0100010111), .y(t0_010001011));
wire t0_0100010110, t0_0100010111;
mixer mix_t0_0100011 (.a(t0_01000110), .b(t0_01000111), .y(t0_0100011));
wire t0_01000110, t0_01000111;
mixer mix_t0_01000110 (.a(t0_010001100), .b(t0_010001101), .y(t0_01000110));
wire t0_010001100, t0_010001101;
mixer mix_t0_010001100 (.a(t0_0100011000), .b(t0_0100011001), .y(t0_010001100));
wire t0_0100011000, t0_0100011001;
mixer mix_t0_010001101 (.a(t0_0100011010), .b(t0_0100011011), .y(t0_010001101));
wire t0_0100011010, t0_0100011011;
mixer mix_t0_01000111 (.a(t0_010001110), .b(t0_010001111), .y(t0_01000111));
wire t0_010001110, t0_010001111;
mixer mix_t0_010001110 (.a(t0_0100011100), .b(t0_0100011101), .y(t0_010001110));
wire t0_0100011100, t0_0100011101;
mixer mix_t0_010001111 (.a(t0_0100011110), .b(t0_0100011111), .y(t0_010001111));
wire t0_0100011110, t0_0100011111;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_010010 (.a(t0_0100100), .b(t0_0100101), .y(t0_010010));
wire t0_0100100, t0_0100101;
mixer mix_t0_0100100 (.a(t0_01001000), .b(t0_01001001), .y(t0_0100100));
wire t0_01001000, t0_01001001;
mixer mix_t0_01001000 (.a(t0_010010000), .b(t0_010010001), .y(t0_01001000));
wire t0_010010000, t0_010010001;
mixer mix_t0_010010000 (.a(t0_0100100000), .b(t0_0100100001), .y(t0_010010000));
wire t0_0100100000, t0_0100100001;
mixer mix_t0_010010001 (.a(t0_0100100010), .b(t0_0100100011), .y(t0_010010001));
wire t0_0100100010, t0_0100100011;
mixer mix_t0_01001001 (.a(t0_010010010), .b(t0_010010011), .y(t0_01001001));
wire t0_010010010, t0_010010011;
mixer mix_t0_010010010 (.a(t0_0100100100), .b(t0_0100100101), .y(t0_010010010));
wire t0_0100100100, t0_0100100101;
mixer mix_t0_010010011 (.a(t0_0100100110), .b(t0_0100100111), .y(t0_010010011));
wire t0_0100100110, t0_0100100111;
mixer mix_t0_0100101 (.a(t0_01001010), .b(t0_01001011), .y(t0_0100101));
wire t0_01001010, t0_01001011;
mixer mix_t0_01001010 (.a(t0_010010100), .b(t0_010010101), .y(t0_01001010));
wire t0_010010100, t0_010010101;
mixer mix_t0_010010100 (.a(t0_0100101000), .b(t0_0100101001), .y(t0_010010100));
wire t0_0100101000, t0_0100101001;
mixer mix_t0_010010101 (.a(t0_0100101010), .b(t0_0100101011), .y(t0_010010101));
wire t0_0100101010, t0_0100101011;
mixer mix_t0_01001011 (.a(t0_010010110), .b(t0_010010111), .y(t0_01001011));
wire t0_010010110, t0_010010111;
mixer mix_t0_010010110 (.a(t0_0100101100), .b(t0_0100101101), .y(t0_010010110));
wire t0_0100101100, t0_0100101101;
mixer mix_t0_010010111 (.a(t0_0100101110), .b(t0_0100101111), .y(t0_010010111));
wire t0_0100101110, t0_0100101111;
mixer mix_t0_010011 (.a(t0_0100110), .b(t0_0100111), .y(t0_010011));
wire t0_0100110, t0_0100111;
mixer mix_t0_0100110 (.a(t0_01001100), .b(t0_01001101), .y(t0_0100110));
wire t0_01001100, t0_01001101;
mixer mix_t0_01001100 (.a(t0_010011000), .b(t0_010011001), .y(t0_01001100));
wire t0_010011000, t0_010011001;
mixer mix_t0_010011000 (.a(t0_0100110000), .b(t0_0100110001), .y(t0_010011000));
wire t0_0100110000, t0_0100110001;
mixer mix_t0_010011001 (.a(t0_0100110010), .b(t0_0100110011), .y(t0_010011001));
wire t0_0100110010, t0_0100110011;
mixer mix_t0_01001101 (.a(t0_010011010), .b(t0_010011011), .y(t0_01001101));
wire t0_010011010, t0_010011011;
mixer mix_t0_010011010 (.a(t0_0100110100), .b(t0_0100110101), .y(t0_010011010));
wire t0_0100110100, t0_0100110101;
mixer mix_t0_010011011 (.a(t0_0100110110), .b(t0_0100110111), .y(t0_010011011));
wire t0_0100110110, t0_0100110111;
mixer mix_t0_0100111 (.a(t0_01001110), .b(t0_01001111), .y(t0_0100111));
wire t0_01001110, t0_01001111;
mixer mix_t0_01001110 (.a(t0_010011100), .b(t0_010011101), .y(t0_01001110));
wire t0_010011100, t0_010011101;
mixer mix_t0_010011100 (.a(t0_0100111000), .b(t0_0100111001), .y(t0_010011100));
wire t0_0100111000, t0_0100111001;
mixer mix_t0_010011101 (.a(t0_0100111010), .b(t0_0100111011), .y(t0_010011101));
wire t0_0100111010, t0_0100111011;
mixer mix_t0_01001111 (.a(t0_010011110), .b(t0_010011111), .y(t0_01001111));
wire t0_010011110, t0_010011111;
mixer mix_t0_010011110 (.a(t0_0100111100), .b(t0_0100111101), .y(t0_010011110));
wire t0_0100111100, t0_0100111101;
mixer mix_t0_010011111 (.a(t0_0100111110), .b(t0_0100111111), .y(t0_010011111));
wire t0_0100111110, t0_0100111111;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_010100 (.a(t0_0101000), .b(t0_0101001), .y(t0_010100));
wire t0_0101000, t0_0101001;
mixer mix_t0_0101000 (.a(t0_01010000), .b(t0_01010001), .y(t0_0101000));
wire t0_01010000, t0_01010001;
mixer mix_t0_01010000 (.a(t0_010100000), .b(t0_010100001), .y(t0_01010000));
wire t0_010100000, t0_010100001;
mixer mix_t0_010100000 (.a(t0_0101000000), .b(t0_0101000001), .y(t0_010100000));
wire t0_0101000000, t0_0101000001;
mixer mix_t0_010100001 (.a(t0_0101000010), .b(t0_0101000011), .y(t0_010100001));
wire t0_0101000010, t0_0101000011;
mixer mix_t0_01010001 (.a(t0_010100010), .b(t0_010100011), .y(t0_01010001));
wire t0_010100010, t0_010100011;
mixer mix_t0_010100010 (.a(t0_0101000100), .b(t0_0101000101), .y(t0_010100010));
wire t0_0101000100, t0_0101000101;
mixer mix_t0_010100011 (.a(t0_0101000110), .b(t0_0101000111), .y(t0_010100011));
wire t0_0101000110, t0_0101000111;
mixer mix_t0_0101001 (.a(t0_01010010), .b(t0_01010011), .y(t0_0101001));
wire t0_01010010, t0_01010011;
mixer mix_t0_01010010 (.a(t0_010100100), .b(t0_010100101), .y(t0_01010010));
wire t0_010100100, t0_010100101;
mixer mix_t0_010100100 (.a(t0_0101001000), .b(t0_0101001001), .y(t0_010100100));
wire t0_0101001000, t0_0101001001;
mixer mix_t0_010100101 (.a(t0_0101001010), .b(t0_0101001011), .y(t0_010100101));
wire t0_0101001010, t0_0101001011;
mixer mix_t0_01010011 (.a(t0_010100110), .b(t0_010100111), .y(t0_01010011));
wire t0_010100110, t0_010100111;
mixer mix_t0_010100110 (.a(t0_0101001100), .b(t0_0101001101), .y(t0_010100110));
wire t0_0101001100, t0_0101001101;
mixer mix_t0_010100111 (.a(t0_0101001110), .b(t0_0101001111), .y(t0_010100111));
wire t0_0101001110, t0_0101001111;
mixer mix_t0_010101 (.a(t0_0101010), .b(t0_0101011), .y(t0_010101));
wire t0_0101010, t0_0101011;
mixer mix_t0_0101010 (.a(t0_01010100), .b(t0_01010101), .y(t0_0101010));
wire t0_01010100, t0_01010101;
mixer mix_t0_01010100 (.a(t0_010101000), .b(t0_010101001), .y(t0_01010100));
wire t0_010101000, t0_010101001;
mixer mix_t0_010101000 (.a(t0_0101010000), .b(t0_0101010001), .y(t0_010101000));
wire t0_0101010000, t0_0101010001;
mixer mix_t0_010101001 (.a(t0_0101010010), .b(t0_0101010011), .y(t0_010101001));
wire t0_0101010010, t0_0101010011;
mixer mix_t0_01010101 (.a(t0_010101010), .b(t0_010101011), .y(t0_01010101));
wire t0_010101010, t0_010101011;
mixer mix_t0_010101010 (.a(t0_0101010100), .b(t0_0101010101), .y(t0_010101010));
wire t0_0101010100, t0_0101010101;
mixer mix_t0_010101011 (.a(t0_0101010110), .b(t0_0101010111), .y(t0_010101011));
wire t0_0101010110, t0_0101010111;
mixer mix_t0_0101011 (.a(t0_01010110), .b(t0_01010111), .y(t0_0101011));
wire t0_01010110, t0_01010111;
mixer mix_t0_01010110 (.a(t0_010101100), .b(t0_010101101), .y(t0_01010110));
wire t0_010101100, t0_010101101;
mixer mix_t0_010101100 (.a(t0_0101011000), .b(t0_0101011001), .y(t0_010101100));
wire t0_0101011000, t0_0101011001;
mixer mix_t0_010101101 (.a(t0_0101011010), .b(t0_0101011011), .y(t0_010101101));
wire t0_0101011010, t0_0101011011;
mixer mix_t0_01010111 (.a(t0_010101110), .b(t0_010101111), .y(t0_01010111));
wire t0_010101110, t0_010101111;
mixer mix_t0_010101110 (.a(t0_0101011100), .b(t0_0101011101), .y(t0_010101110));
wire t0_0101011100, t0_0101011101;
mixer mix_t0_010101111 (.a(t0_0101011110), .b(t0_0101011111), .y(t0_010101111));
wire t0_0101011110, t0_0101011111;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_010110 (.a(t0_0101100), .b(t0_0101101), .y(t0_010110));
wire t0_0101100, t0_0101101;
mixer mix_t0_0101100 (.a(t0_01011000), .b(t0_01011001), .y(t0_0101100));
wire t0_01011000, t0_01011001;
mixer mix_t0_01011000 (.a(t0_010110000), .b(t0_010110001), .y(t0_01011000));
wire t0_010110000, t0_010110001;
mixer mix_t0_010110000 (.a(t0_0101100000), .b(t0_0101100001), .y(t0_010110000));
wire t0_0101100000, t0_0101100001;
mixer mix_t0_010110001 (.a(t0_0101100010), .b(t0_0101100011), .y(t0_010110001));
wire t0_0101100010, t0_0101100011;
mixer mix_t0_01011001 (.a(t0_010110010), .b(t0_010110011), .y(t0_01011001));
wire t0_010110010, t0_010110011;
mixer mix_t0_010110010 (.a(t0_0101100100), .b(t0_0101100101), .y(t0_010110010));
wire t0_0101100100, t0_0101100101;
mixer mix_t0_010110011 (.a(t0_0101100110), .b(t0_0101100111), .y(t0_010110011));
wire t0_0101100110, t0_0101100111;
mixer mix_t0_0101101 (.a(t0_01011010), .b(t0_01011011), .y(t0_0101101));
wire t0_01011010, t0_01011011;
mixer mix_t0_01011010 (.a(t0_010110100), .b(t0_010110101), .y(t0_01011010));
wire t0_010110100, t0_010110101;
mixer mix_t0_010110100 (.a(t0_0101101000), .b(t0_0101101001), .y(t0_010110100));
wire t0_0101101000, t0_0101101001;
mixer mix_t0_010110101 (.a(t0_0101101010), .b(t0_0101101011), .y(t0_010110101));
wire t0_0101101010, t0_0101101011;
mixer mix_t0_01011011 (.a(t0_010110110), .b(t0_010110111), .y(t0_01011011));
wire t0_010110110, t0_010110111;
mixer mix_t0_010110110 (.a(t0_0101101100), .b(t0_0101101101), .y(t0_010110110));
wire t0_0101101100, t0_0101101101;
mixer mix_t0_010110111 (.a(t0_0101101110), .b(t0_0101101111), .y(t0_010110111));
wire t0_0101101110, t0_0101101111;
mixer mix_t0_010111 (.a(t0_0101110), .b(t0_0101111), .y(t0_010111));
wire t0_0101110, t0_0101111;
mixer mix_t0_0101110 (.a(t0_01011100), .b(t0_01011101), .y(t0_0101110));
wire t0_01011100, t0_01011101;
mixer mix_t0_01011100 (.a(t0_010111000), .b(t0_010111001), .y(t0_01011100));
wire t0_010111000, t0_010111001;
mixer mix_t0_010111000 (.a(t0_0101110000), .b(t0_0101110001), .y(t0_010111000));
wire t0_0101110000, t0_0101110001;
mixer mix_t0_010111001 (.a(t0_0101110010), .b(t0_0101110011), .y(t0_010111001));
wire t0_0101110010, t0_0101110011;
mixer mix_t0_01011101 (.a(t0_010111010), .b(t0_010111011), .y(t0_01011101));
wire t0_010111010, t0_010111011;
mixer mix_t0_010111010 (.a(t0_0101110100), .b(t0_0101110101), .y(t0_010111010));
wire t0_0101110100, t0_0101110101;
mixer mix_t0_010111011 (.a(t0_0101110110), .b(t0_0101110111), .y(t0_010111011));
wire t0_0101110110, t0_0101110111;
mixer mix_t0_0101111 (.a(t0_01011110), .b(t0_01011111), .y(t0_0101111));
wire t0_01011110, t0_01011111;
mixer mix_t0_01011110 (.a(t0_010111100), .b(t0_010111101), .y(t0_01011110));
wire t0_010111100, t0_010111101;
mixer mix_t0_010111100 (.a(t0_0101111000), .b(t0_0101111001), .y(t0_010111100));
wire t0_0101111000, t0_0101111001;
mixer mix_t0_010111101 (.a(t0_0101111010), .b(t0_0101111011), .y(t0_010111101));
wire t0_0101111010, t0_0101111011;
mixer mix_t0_01011111 (.a(t0_010111110), .b(t0_010111111), .y(t0_01011111));
wire t0_010111110, t0_010111111;
mixer mix_t0_010111110 (.a(t0_0101111100), .b(t0_0101111101), .y(t0_010111110));
wire t0_0101111100, t0_0101111101;
mixer mix_t0_010111111 (.a(t0_0101111110), .b(t0_0101111111), .y(t0_010111111));
wire t0_0101111110, t0_0101111111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_011000 (.a(t0_0110000), .b(t0_0110001), .y(t0_011000));
wire t0_0110000, t0_0110001;
mixer mix_t0_0110000 (.a(t0_01100000), .b(t0_01100001), .y(t0_0110000));
wire t0_01100000, t0_01100001;
mixer mix_t0_01100000 (.a(t0_011000000), .b(t0_011000001), .y(t0_01100000));
wire t0_011000000, t0_011000001;
mixer mix_t0_011000000 (.a(t0_0110000000), .b(t0_0110000001), .y(t0_011000000));
wire t0_0110000000, t0_0110000001;
mixer mix_t0_011000001 (.a(t0_0110000010), .b(t0_0110000011), .y(t0_011000001));
wire t0_0110000010, t0_0110000011;
mixer mix_t0_01100001 (.a(t0_011000010), .b(t0_011000011), .y(t0_01100001));
wire t0_011000010, t0_011000011;
mixer mix_t0_011000010 (.a(t0_0110000100), .b(t0_0110000101), .y(t0_011000010));
wire t0_0110000100, t0_0110000101;
mixer mix_t0_011000011 (.a(t0_0110000110), .b(t0_0110000111), .y(t0_011000011));
wire t0_0110000110, t0_0110000111;
mixer mix_t0_0110001 (.a(t0_01100010), .b(t0_01100011), .y(t0_0110001));
wire t0_01100010, t0_01100011;
mixer mix_t0_01100010 (.a(t0_011000100), .b(t0_011000101), .y(t0_01100010));
wire t0_011000100, t0_011000101;
mixer mix_t0_011000100 (.a(t0_0110001000), .b(t0_0110001001), .y(t0_011000100));
wire t0_0110001000, t0_0110001001;
mixer mix_t0_011000101 (.a(t0_0110001010), .b(t0_0110001011), .y(t0_011000101));
wire t0_0110001010, t0_0110001011;
mixer mix_t0_01100011 (.a(t0_011000110), .b(t0_011000111), .y(t0_01100011));
wire t0_011000110, t0_011000111;
mixer mix_t0_011000110 (.a(t0_0110001100), .b(t0_0110001101), .y(t0_011000110));
wire t0_0110001100, t0_0110001101;
mixer mix_t0_011000111 (.a(t0_0110001110), .b(t0_0110001111), .y(t0_011000111));
wire t0_0110001110, t0_0110001111;
mixer mix_t0_011001 (.a(t0_0110010), .b(t0_0110011), .y(t0_011001));
wire t0_0110010, t0_0110011;
mixer mix_t0_0110010 (.a(t0_01100100), .b(t0_01100101), .y(t0_0110010));
wire t0_01100100, t0_01100101;
mixer mix_t0_01100100 (.a(t0_011001000), .b(t0_011001001), .y(t0_01100100));
wire t0_011001000, t0_011001001;
mixer mix_t0_011001000 (.a(t0_0110010000), .b(t0_0110010001), .y(t0_011001000));
wire t0_0110010000, t0_0110010001;
mixer mix_t0_011001001 (.a(t0_0110010010), .b(t0_0110010011), .y(t0_011001001));
wire t0_0110010010, t0_0110010011;
mixer mix_t0_01100101 (.a(t0_011001010), .b(t0_011001011), .y(t0_01100101));
wire t0_011001010, t0_011001011;
mixer mix_t0_011001010 (.a(t0_0110010100), .b(t0_0110010101), .y(t0_011001010));
wire t0_0110010100, t0_0110010101;
mixer mix_t0_011001011 (.a(t0_0110010110), .b(t0_0110010111), .y(t0_011001011));
wire t0_0110010110, t0_0110010111;
mixer mix_t0_0110011 (.a(t0_01100110), .b(t0_01100111), .y(t0_0110011));
wire t0_01100110, t0_01100111;
mixer mix_t0_01100110 (.a(t0_011001100), .b(t0_011001101), .y(t0_01100110));
wire t0_011001100, t0_011001101;
mixer mix_t0_011001100 (.a(t0_0110011000), .b(t0_0110011001), .y(t0_011001100));
wire t0_0110011000, t0_0110011001;
mixer mix_t0_011001101 (.a(t0_0110011010), .b(t0_0110011011), .y(t0_011001101));
wire t0_0110011010, t0_0110011011;
mixer mix_t0_01100111 (.a(t0_011001110), .b(t0_011001111), .y(t0_01100111));
wire t0_011001110, t0_011001111;
mixer mix_t0_011001110 (.a(t0_0110011100), .b(t0_0110011101), .y(t0_011001110));
wire t0_0110011100, t0_0110011101;
mixer mix_t0_011001111 (.a(t0_0110011110), .b(t0_0110011111), .y(t0_011001111));
wire t0_0110011110, t0_0110011111;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_011010 (.a(t0_0110100), .b(t0_0110101), .y(t0_011010));
wire t0_0110100, t0_0110101;
mixer mix_t0_0110100 (.a(t0_01101000), .b(t0_01101001), .y(t0_0110100));
wire t0_01101000, t0_01101001;
mixer mix_t0_01101000 (.a(t0_011010000), .b(t0_011010001), .y(t0_01101000));
wire t0_011010000, t0_011010001;
mixer mix_t0_011010000 (.a(t0_0110100000), .b(t0_0110100001), .y(t0_011010000));
wire t0_0110100000, t0_0110100001;
mixer mix_t0_011010001 (.a(t0_0110100010), .b(t0_0110100011), .y(t0_011010001));
wire t0_0110100010, t0_0110100011;
mixer mix_t0_01101001 (.a(t0_011010010), .b(t0_011010011), .y(t0_01101001));
wire t0_011010010, t0_011010011;
mixer mix_t0_011010010 (.a(t0_0110100100), .b(t0_0110100101), .y(t0_011010010));
wire t0_0110100100, t0_0110100101;
mixer mix_t0_011010011 (.a(t0_0110100110), .b(t0_0110100111), .y(t0_011010011));
wire t0_0110100110, t0_0110100111;
mixer mix_t0_0110101 (.a(t0_01101010), .b(t0_01101011), .y(t0_0110101));
wire t0_01101010, t0_01101011;
mixer mix_t0_01101010 (.a(t0_011010100), .b(t0_011010101), .y(t0_01101010));
wire t0_011010100, t0_011010101;
mixer mix_t0_011010100 (.a(t0_0110101000), .b(t0_0110101001), .y(t0_011010100));
wire t0_0110101000, t0_0110101001;
mixer mix_t0_011010101 (.a(t0_0110101010), .b(t0_0110101011), .y(t0_011010101));
wire t0_0110101010, t0_0110101011;
mixer mix_t0_01101011 (.a(t0_011010110), .b(t0_011010111), .y(t0_01101011));
wire t0_011010110, t0_011010111;
mixer mix_t0_011010110 (.a(t0_0110101100), .b(t0_0110101101), .y(t0_011010110));
wire t0_0110101100, t0_0110101101;
mixer mix_t0_011010111 (.a(t0_0110101110), .b(t0_0110101111), .y(t0_011010111));
wire t0_0110101110, t0_0110101111;
mixer mix_t0_011011 (.a(t0_0110110), .b(t0_0110111), .y(t0_011011));
wire t0_0110110, t0_0110111;
mixer mix_t0_0110110 (.a(t0_01101100), .b(t0_01101101), .y(t0_0110110));
wire t0_01101100, t0_01101101;
mixer mix_t0_01101100 (.a(t0_011011000), .b(t0_011011001), .y(t0_01101100));
wire t0_011011000, t0_011011001;
mixer mix_t0_011011000 (.a(t0_0110110000), .b(t0_0110110001), .y(t0_011011000));
wire t0_0110110000, t0_0110110001;
mixer mix_t0_011011001 (.a(t0_0110110010), .b(t0_0110110011), .y(t0_011011001));
wire t0_0110110010, t0_0110110011;
mixer mix_t0_01101101 (.a(t0_011011010), .b(t0_011011011), .y(t0_01101101));
wire t0_011011010, t0_011011011;
mixer mix_t0_011011010 (.a(t0_0110110100), .b(t0_0110110101), .y(t0_011011010));
wire t0_0110110100, t0_0110110101;
mixer mix_t0_011011011 (.a(t0_0110110110), .b(t0_0110110111), .y(t0_011011011));
wire t0_0110110110, t0_0110110111;
mixer mix_t0_0110111 (.a(t0_01101110), .b(t0_01101111), .y(t0_0110111));
wire t0_01101110, t0_01101111;
mixer mix_t0_01101110 (.a(t0_011011100), .b(t0_011011101), .y(t0_01101110));
wire t0_011011100, t0_011011101;
mixer mix_t0_011011100 (.a(t0_0110111000), .b(t0_0110111001), .y(t0_011011100));
wire t0_0110111000, t0_0110111001;
mixer mix_t0_011011101 (.a(t0_0110111010), .b(t0_0110111011), .y(t0_011011101));
wire t0_0110111010, t0_0110111011;
mixer mix_t0_01101111 (.a(t0_011011110), .b(t0_011011111), .y(t0_01101111));
wire t0_011011110, t0_011011111;
mixer mix_t0_011011110 (.a(t0_0110111100), .b(t0_0110111101), .y(t0_011011110));
wire t0_0110111100, t0_0110111101;
mixer mix_t0_011011111 (.a(t0_0110111110), .b(t0_0110111111), .y(t0_011011111));
wire t0_0110111110, t0_0110111111;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_011100 (.a(t0_0111000), .b(t0_0111001), .y(t0_011100));
wire t0_0111000, t0_0111001;
mixer mix_t0_0111000 (.a(t0_01110000), .b(t0_01110001), .y(t0_0111000));
wire t0_01110000, t0_01110001;
mixer mix_t0_01110000 (.a(t0_011100000), .b(t0_011100001), .y(t0_01110000));
wire t0_011100000, t0_011100001;
mixer mix_t0_011100000 (.a(t0_0111000000), .b(t0_0111000001), .y(t0_011100000));
wire t0_0111000000, t0_0111000001;
mixer mix_t0_011100001 (.a(t0_0111000010), .b(t0_0111000011), .y(t0_011100001));
wire t0_0111000010, t0_0111000011;
mixer mix_t0_01110001 (.a(t0_011100010), .b(t0_011100011), .y(t0_01110001));
wire t0_011100010, t0_011100011;
mixer mix_t0_011100010 (.a(t0_0111000100), .b(t0_0111000101), .y(t0_011100010));
wire t0_0111000100, t0_0111000101;
mixer mix_t0_011100011 (.a(t0_0111000110), .b(t0_0111000111), .y(t0_011100011));
wire t0_0111000110, t0_0111000111;
mixer mix_t0_0111001 (.a(t0_01110010), .b(t0_01110011), .y(t0_0111001));
wire t0_01110010, t0_01110011;
mixer mix_t0_01110010 (.a(t0_011100100), .b(t0_011100101), .y(t0_01110010));
wire t0_011100100, t0_011100101;
mixer mix_t0_011100100 (.a(t0_0111001000), .b(t0_0111001001), .y(t0_011100100));
wire t0_0111001000, t0_0111001001;
mixer mix_t0_011100101 (.a(t0_0111001010), .b(t0_0111001011), .y(t0_011100101));
wire t0_0111001010, t0_0111001011;
mixer mix_t0_01110011 (.a(t0_011100110), .b(t0_011100111), .y(t0_01110011));
wire t0_011100110, t0_011100111;
mixer mix_t0_011100110 (.a(t0_0111001100), .b(t0_0111001101), .y(t0_011100110));
wire t0_0111001100, t0_0111001101;
mixer mix_t0_011100111 (.a(t0_0111001110), .b(t0_0111001111), .y(t0_011100111));
wire t0_0111001110, t0_0111001111;
mixer mix_t0_011101 (.a(t0_0111010), .b(t0_0111011), .y(t0_011101));
wire t0_0111010, t0_0111011;
mixer mix_t0_0111010 (.a(t0_01110100), .b(t0_01110101), .y(t0_0111010));
wire t0_01110100, t0_01110101;
mixer mix_t0_01110100 (.a(t0_011101000), .b(t0_011101001), .y(t0_01110100));
wire t0_011101000, t0_011101001;
mixer mix_t0_011101000 (.a(t0_0111010000), .b(t0_0111010001), .y(t0_011101000));
wire t0_0111010000, t0_0111010001;
mixer mix_t0_011101001 (.a(t0_0111010010), .b(t0_0111010011), .y(t0_011101001));
wire t0_0111010010, t0_0111010011;
mixer mix_t0_01110101 (.a(t0_011101010), .b(t0_011101011), .y(t0_01110101));
wire t0_011101010, t0_011101011;
mixer mix_t0_011101010 (.a(t0_0111010100), .b(t0_0111010101), .y(t0_011101010));
wire t0_0111010100, t0_0111010101;
mixer mix_t0_011101011 (.a(t0_0111010110), .b(t0_0111010111), .y(t0_011101011));
wire t0_0111010110, t0_0111010111;
mixer mix_t0_0111011 (.a(t0_01110110), .b(t0_01110111), .y(t0_0111011));
wire t0_01110110, t0_01110111;
mixer mix_t0_01110110 (.a(t0_011101100), .b(t0_011101101), .y(t0_01110110));
wire t0_011101100, t0_011101101;
mixer mix_t0_011101100 (.a(t0_0111011000), .b(t0_0111011001), .y(t0_011101100));
wire t0_0111011000, t0_0111011001;
mixer mix_t0_011101101 (.a(t0_0111011010), .b(t0_0111011011), .y(t0_011101101));
wire t0_0111011010, t0_0111011011;
mixer mix_t0_01110111 (.a(t0_011101110), .b(t0_011101111), .y(t0_01110111));
wire t0_011101110, t0_011101111;
mixer mix_t0_011101110 (.a(t0_0111011100), .b(t0_0111011101), .y(t0_011101110));
wire t0_0111011100, t0_0111011101;
mixer mix_t0_011101111 (.a(t0_0111011110), .b(t0_0111011111), .y(t0_011101111));
wire t0_0111011110, t0_0111011111;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
mixer mix_t0_011110 (.a(t0_0111100), .b(t0_0111101), .y(t0_011110));
wire t0_0111100, t0_0111101;
mixer mix_t0_0111100 (.a(t0_01111000), .b(t0_01111001), .y(t0_0111100));
wire t0_01111000, t0_01111001;
mixer mix_t0_01111000 (.a(t0_011110000), .b(t0_011110001), .y(t0_01111000));
wire t0_011110000, t0_011110001;
mixer mix_t0_011110000 (.a(t0_0111100000), .b(t0_0111100001), .y(t0_011110000));
wire t0_0111100000, t0_0111100001;
mixer mix_t0_011110001 (.a(t0_0111100010), .b(t0_0111100011), .y(t0_011110001));
wire t0_0111100010, t0_0111100011;
mixer mix_t0_01111001 (.a(t0_011110010), .b(t0_011110011), .y(t0_01111001));
wire t0_011110010, t0_011110011;
mixer mix_t0_011110010 (.a(t0_0111100100), .b(t0_0111100101), .y(t0_011110010));
wire t0_0111100100, t0_0111100101;
mixer mix_t0_011110011 (.a(t0_0111100110), .b(t0_0111100111), .y(t0_011110011));
wire t0_0111100110, t0_0111100111;
mixer mix_t0_0111101 (.a(t0_01111010), .b(t0_01111011), .y(t0_0111101));
wire t0_01111010, t0_01111011;
mixer mix_t0_01111010 (.a(t0_011110100), .b(t0_011110101), .y(t0_01111010));
wire t0_011110100, t0_011110101;
mixer mix_t0_011110100 (.a(t0_0111101000), .b(t0_0111101001), .y(t0_011110100));
wire t0_0111101000, t0_0111101001;
mixer mix_t0_011110101 (.a(t0_0111101010), .b(t0_0111101011), .y(t0_011110101));
wire t0_0111101010, t0_0111101011;
mixer mix_t0_01111011 (.a(t0_011110110), .b(t0_011110111), .y(t0_01111011));
wire t0_011110110, t0_011110111;
mixer mix_t0_011110110 (.a(t0_0111101100), .b(t0_0111101101), .y(t0_011110110));
wire t0_0111101100, t0_0111101101;
mixer mix_t0_011110111 (.a(t0_0111101110), .b(t0_0111101111), .y(t0_011110111));
wire t0_0111101110, t0_0111101111;
mixer mix_t0_011111 (.a(t0_0111110), .b(t0_0111111), .y(t0_011111));
wire t0_0111110, t0_0111111;
mixer mix_t0_0111110 (.a(t0_01111100), .b(t0_01111101), .y(t0_0111110));
wire t0_01111100, t0_01111101;
mixer mix_t0_01111100 (.a(t0_011111000), .b(t0_011111001), .y(t0_01111100));
wire t0_011111000, t0_011111001;
mixer mix_t0_011111000 (.a(t0_0111110000), .b(t0_0111110001), .y(t0_011111000));
wire t0_0111110000, t0_0111110001;
mixer mix_t0_011111001 (.a(t0_0111110010), .b(t0_0111110011), .y(t0_011111001));
wire t0_0111110010, t0_0111110011;
mixer mix_t0_01111101 (.a(t0_011111010), .b(t0_011111011), .y(t0_01111101));
wire t0_011111010, t0_011111011;
mixer mix_t0_011111010 (.a(t0_0111110100), .b(t0_0111110101), .y(t0_011111010));
wire t0_0111110100, t0_0111110101;
mixer mix_t0_011111011 (.a(t0_0111110110), .b(t0_0111110111), .y(t0_011111011));
wire t0_0111110110, t0_0111110111;
mixer mix_t0_0111111 (.a(t0_01111110), .b(t0_01111111), .y(t0_0111111));
wire t0_01111110, t0_01111111;
mixer mix_t0_01111110 (.a(t0_011111100), .b(t0_011111101), .y(t0_01111110));
wire t0_011111100, t0_011111101;
mixer mix_t0_011111100 (.a(t0_0111111000), .b(t0_0111111001), .y(t0_011111100));
wire t0_0111111000, t0_0111111001;
mixer mix_t0_011111101 (.a(t0_0111111010), .b(t0_0111111011), .y(t0_011111101));
wire t0_0111111010, t0_0111111011;
mixer mix_t0_01111111 (.a(t0_011111110), .b(t0_011111111), .y(t0_01111111));
wire t0_011111110, t0_011111111;
mixer mix_t0_011111110 (.a(t0_0111111100), .b(t0_0111111101), .y(t0_011111110));
wire t0_0111111100, t0_0111111101;
mixer mix_t0_011111111 (.a(t0_0111111110), .b(t0_0111111111), .y(t0_011111111));
wire t0_0111111110, t0_0111111111;
wire t0_0;
assign out_0 = t0_0;
assign input_0 = t0_0000000000;
assign input_1 = t0_0000000001;
assign input_2 = t0_0000000010;
assign input_3 = t0_0000000011;
assign input_4 = t0_0000000100;
assign input_5 = t0_0000000101;
assign input_6 = t0_0000000110;
assign input_7 = t0_0000000111;
assign input_8 = t0_0000001000;
assign input_9 = t0_0000001001;
assign input_10 = t0_0000001010;
assign input_11 = t0_0000001011;
assign input_12 = t0_0000001100;
assign input_13 = t0_0000001101;
assign input_14 = t0_0000001110;
assign input_15 = t0_0000001111;
assign input_16 = t0_0000010000;
assign input_17 = t0_0000010001;
assign input_18 = t0_0000010010;
assign input_19 = t0_0000010011;
assign input_20 = t0_0000010100;
assign input_21 = t0_0000010101;
assign input_22 = t0_0000010110;
assign input_23 = t0_0000010111;
assign input_24 = t0_0000011000;
assign input_25 = t0_0000011001;
assign input_26 = t0_0000011010;
assign input_27 = t0_0000011011;
assign input_28 = t0_0000011100;
assign input_29 = t0_0000011101;
assign input_30 = t0_0000011110;
assign input_31 = t0_0000011111;
assign input_32 = t0_0000100000;
assign input_33 = t0_0000100001;
assign input_34 = t0_0000100010;
assign input_35 = t0_0000100011;
assign input_36 = t0_0000100100;
assign input_37 = t0_0000100101;
assign input_38 = t0_0000100110;
assign input_39 = t0_0000100111;
assign input_40 = t0_0000101000;
assign input_41 = t0_0000101001;
assign input_42 = t0_0000101010;
assign input_43 = t0_0000101011;
assign input_44 = t0_0000101100;
assign input_45 = t0_0000101101;
assign input_46 = t0_0000101110;
assign input_47 = t0_0000101111;
assign input_48 = t0_0000110000;
assign input_49 = t0_0000110001;
assign input_50 = t0_0000110010;
assign input_51 = t0_0000110011;
assign input_52 = t0_0000110100;
assign input_53 = t0_0000110101;
assign input_54 = t0_0000110110;
assign input_55 = t0_0000110111;
assign input_56 = t0_0000111000;
assign input_57 = t0_0000111001;
assign input_58 = t0_0000111010;
assign input_59 = t0_0000111011;
assign input_60 = t0_0000111100;
assign input_61 = t0_0000111101;
assign input_62 = t0_0000111110;
assign input_63 = t0_0000111111;
assign input_64 = t0_0001000000;
assign input_65 = t0_0001000001;
assign input_66 = t0_0001000010;
assign input_67 = t0_0001000011;
assign input_68 = t0_0001000100;
assign input_69 = t0_0001000101;
assign input_70 = t0_0001000110;
assign input_71 = t0_0001000111;
assign input_72 = t0_0001001000;
assign input_73 = t0_0001001001;
assign input_74 = t0_0001001010;
assign input_75 = t0_0001001011;
assign input_76 = t0_0001001100;
assign input_77 = t0_0001001101;
assign input_78 = t0_0001001110;
assign input_79 = t0_0001001111;
assign input_80 = t0_0001010000;
assign input_81 = t0_0001010001;
assign input_82 = t0_0001010010;
assign input_83 = t0_0001010011;
assign input_84 = t0_0001010100;
assign input_85 = t0_0001010101;
assign input_86 = t0_0001010110;
assign input_87 = t0_0001010111;
assign input_88 = t0_0001011000;
assign input_89 = t0_0001011001;
assign input_90 = t0_0001011010;
assign input_91 = t0_0001011011;
assign input_92 = t0_0001011100;
assign input_93 = t0_0001011101;
assign input_94 = t0_0001011110;
assign input_95 = t0_0001011111;
assign input_96 = t0_0001100000;
assign input_97 = t0_0001100001;
assign input_98 = t0_0001100010;
assign input_99 = t0_0001100011;
assign input_100 = t0_0001100100;
assign input_101 = t0_0001100101;
assign input_102 = t0_0001100110;
assign input_103 = t0_0001100111;
assign input_104 = t0_0001101000;
assign input_105 = t0_0001101001;
assign input_106 = t0_0001101010;
assign input_107 = t0_0001101011;
assign input_108 = t0_0001101100;
assign input_109 = t0_0001101101;
assign input_110 = t0_0001101110;
assign input_111 = t0_0001101111;
assign input_112 = t0_0001110000;
assign input_113 = t0_0001110001;
assign input_114 = t0_0001110010;
assign input_115 = t0_0001110011;
assign input_116 = t0_0001110100;
assign input_117 = t0_0001110101;
assign input_118 = t0_0001110110;
assign input_119 = t0_0001110111;
assign input_120 = t0_0001111000;
assign input_121 = t0_0001111001;
assign input_122 = t0_0001111010;
assign input_123 = t0_0001111011;
assign input_124 = t0_0001111100;
assign input_125 = t0_0001111101;
assign input_126 = t0_0001111110;
assign input_127 = t0_0001111111;
assign input_128 = t0_0010000000;
assign input_129 = t0_0010000001;
assign input_130 = t0_0010000010;
assign input_131 = t0_0010000011;
assign input_132 = t0_0010000100;
assign input_133 = t0_0010000101;
assign input_134 = t0_0010000110;
assign input_135 = t0_0010000111;
assign input_136 = t0_0010001000;
assign input_137 = t0_0010001001;
assign input_138 = t0_0010001010;
assign input_139 = t0_0010001011;
assign input_140 = t0_0010001100;
assign input_141 = t0_0010001101;
assign input_142 = t0_0010001110;
assign input_143 = t0_0010001111;
assign input_144 = t0_0010010000;
assign input_145 = t0_0010010001;
assign input_146 = t0_0010010010;
assign input_147 = t0_0010010011;
assign input_148 = t0_0010010100;
assign input_149 = t0_0010010101;
assign input_150 = t0_0010010110;
assign input_151 = t0_0010010111;
assign input_152 = t0_0010011000;
assign input_153 = t0_0010011001;
assign input_154 = t0_0010011010;
assign input_155 = t0_0010011011;
assign input_156 = t0_0010011100;
assign input_157 = t0_0010011101;
assign input_158 = t0_0010011110;
assign input_159 = t0_0010011111;
assign input_160 = t0_0010100000;
assign input_161 = t0_0010100001;
assign input_162 = t0_0010100010;
assign input_163 = t0_0010100011;
assign input_164 = t0_0010100100;
assign input_165 = t0_0010100101;
assign input_166 = t0_0010100110;
assign input_167 = t0_0010100111;
assign input_168 = t0_0010101000;
assign input_169 = t0_0010101001;
assign input_170 = t0_0010101010;
assign input_171 = t0_0010101011;
assign input_172 = t0_0010101100;
assign input_173 = t0_0010101101;
assign input_174 = t0_0010101110;
assign input_175 = t0_0010101111;
assign input_176 = t0_0010110000;
assign input_177 = t0_0010110001;
assign input_178 = t0_0010110010;
assign input_179 = t0_0010110011;
assign input_180 = t0_0010110100;
assign input_181 = t0_0010110101;
assign input_182 = t0_0010110110;
assign input_183 = t0_0010110111;
assign input_184 = t0_0010111000;
assign input_185 = t0_0010111001;
assign input_186 = t0_0010111010;
assign input_187 = t0_0010111011;
assign input_188 = t0_0010111100;
assign input_189 = t0_0010111101;
assign input_190 = t0_0010111110;
assign input_191 = t0_0010111111;
assign input_192 = t0_0011000000;
assign input_193 = t0_0011000001;
assign input_194 = t0_0011000010;
assign input_195 = t0_0011000011;
assign input_196 = t0_0011000100;
assign input_197 = t0_0011000101;
assign input_198 = t0_0011000110;
assign input_199 = t0_0011000111;
assign input_200 = t0_0011001000;
assign input_201 = t0_0011001001;
assign input_202 = t0_0011001010;
assign input_203 = t0_0011001011;
assign input_204 = t0_0011001100;
assign input_205 = t0_0011001101;
assign input_206 = t0_0011001110;
assign input_207 = t0_0011001111;
assign input_208 = t0_0011010000;
assign input_209 = t0_0011010001;
assign input_210 = t0_0011010010;
assign input_211 = t0_0011010011;
assign input_212 = t0_0011010100;
assign input_213 = t0_0011010101;
assign input_214 = t0_0011010110;
assign input_215 = t0_0011010111;
assign input_216 = t0_0011011000;
assign input_217 = t0_0011011001;
assign input_218 = t0_0011011010;
assign input_219 = t0_0011011011;
assign input_220 = t0_0011011100;
assign input_221 = t0_0011011101;
assign input_222 = t0_0011011110;
assign input_223 = t0_0011011111;
assign input_224 = t0_0011100000;
assign input_225 = t0_0011100001;
assign input_226 = t0_0011100010;
assign input_227 = t0_0011100011;
assign input_228 = t0_0011100100;
assign input_229 = t0_0011100101;
assign input_230 = t0_0011100110;
assign input_231 = t0_0011100111;
assign input_232 = t0_0011101000;
assign input_233 = t0_0011101001;
assign input_234 = t0_0011101010;
assign input_235 = t0_0011101011;
assign input_236 = t0_0011101100;
assign input_237 = t0_0011101101;
assign input_238 = t0_0011101110;
assign input_239 = t0_0011101111;
assign input_240 = t0_0011110000;
assign input_241 = t0_0011110001;
assign input_242 = t0_0011110010;
assign input_243 = t0_0011110011;
assign input_244 = t0_0011110100;
assign input_245 = t0_0011110101;
assign input_246 = t0_0011110110;
assign input_247 = t0_0011110111;
assign input_248 = t0_0011111000;
assign input_249 = t0_0011111001;
assign input_250 = t0_0011111010;
assign input_251 = t0_0011111011;
assign input_252 = t0_0011111100;
assign input_253 = t0_0011111101;
assign input_254 = t0_0011111110;
assign input_255 = t0_0011111111;
assign input_256 = t0_0100000000;
assign input_257 = t0_0100000001;
assign input_258 = t0_0100000010;
assign input_259 = t0_0100000011;
assign input_260 = t0_0100000100;
assign input_261 = t0_0100000101;
assign input_262 = t0_0100000110;
assign input_263 = t0_0100000111;
assign input_264 = t0_0100001000;
assign input_265 = t0_0100001001;
assign input_266 = t0_0100001010;
assign input_267 = t0_0100001011;
assign input_268 = t0_0100001100;
assign input_269 = t0_0100001101;
assign input_270 = t0_0100001110;
assign input_271 = t0_0100001111;
assign input_272 = t0_0100010000;
assign input_273 = t0_0100010001;
assign input_274 = t0_0100010010;
assign input_275 = t0_0100010011;
assign input_276 = t0_0100010100;
assign input_277 = t0_0100010101;
assign input_278 = t0_0100010110;
assign input_279 = t0_0100010111;
assign input_280 = t0_0100011000;
assign input_281 = t0_0100011001;
assign input_282 = t0_0100011010;
assign input_283 = t0_0100011011;
assign input_284 = t0_0100011100;
assign input_285 = t0_0100011101;
assign input_286 = t0_0100011110;
assign input_287 = t0_0100011111;
assign input_288 = t0_0100100000;
assign input_289 = t0_0100100001;
assign input_290 = t0_0100100010;
assign input_291 = t0_0100100011;
assign input_292 = t0_0100100100;
assign input_293 = t0_0100100101;
assign input_294 = t0_0100100110;
assign input_295 = t0_0100100111;
assign input_296 = t0_0100101000;
assign input_297 = t0_0100101001;
assign input_298 = t0_0100101010;
assign input_299 = t0_0100101011;
assign input_300 = t0_0100101100;
assign input_301 = t0_0100101101;
assign input_302 = t0_0100101110;
assign input_303 = t0_0100101111;
assign input_304 = t0_0100110000;
assign input_305 = t0_0100110001;
assign input_306 = t0_0100110010;
assign input_307 = t0_0100110011;
assign input_308 = t0_0100110100;
assign input_309 = t0_0100110101;
assign input_310 = t0_0100110110;
assign input_311 = t0_0100110111;
assign input_312 = t0_0100111000;
assign input_313 = t0_0100111001;
assign input_314 = t0_0100111010;
assign input_315 = t0_0100111011;
assign input_316 = t0_0100111100;
assign input_317 = t0_0100111101;
assign input_318 = t0_0100111110;
assign input_319 = t0_0100111111;
assign input_320 = t0_0101000000;
assign input_321 = t0_0101000001;
assign input_322 = t0_0101000010;
assign input_323 = t0_0101000011;
assign input_324 = t0_0101000100;
assign input_325 = t0_0101000101;
assign input_326 = t0_0101000110;
assign input_327 = t0_0101000111;
assign input_328 = t0_0101001000;
assign input_329 = t0_0101001001;
assign input_330 = t0_0101001010;
assign input_331 = t0_0101001011;
assign input_332 = t0_0101001100;
assign input_333 = t0_0101001101;
assign input_334 = t0_0101001110;
assign input_335 = t0_0101001111;
assign input_336 = t0_0101010000;
assign input_337 = t0_0101010001;
assign input_338 = t0_0101010010;
assign input_339 = t0_0101010011;
assign input_340 = t0_0101010100;
assign input_341 = t0_0101010101;
assign input_342 = t0_0101010110;
assign input_343 = t0_0101010111;
assign input_344 = t0_0101011000;
assign input_345 = t0_0101011001;
assign input_346 = t0_0101011010;
assign input_347 = t0_0101011011;
assign input_348 = t0_0101011100;
assign input_349 = t0_0101011101;
assign input_350 = t0_0101011110;
assign input_351 = t0_0101011111;
assign input_352 = t0_0101100000;
assign input_353 = t0_0101100001;
assign input_354 = t0_0101100010;
assign input_355 = t0_0101100011;
assign input_356 = t0_0101100100;
assign input_357 = t0_0101100101;
assign input_358 = t0_0101100110;
assign input_359 = t0_0101100111;
assign input_360 = t0_0101101000;
assign input_361 = t0_0101101001;
assign input_362 = t0_0101101010;
assign input_363 = t0_0101101011;
assign input_364 = t0_0101101100;
assign input_365 = t0_0101101101;
assign input_366 = t0_0101101110;
assign input_367 = t0_0101101111;
assign input_368 = t0_0101110000;
assign input_369 = t0_0101110001;
assign input_370 = t0_0101110010;
assign input_371 = t0_0101110011;
assign input_372 = t0_0101110100;
assign input_373 = t0_0101110101;
assign input_374 = t0_0101110110;
assign input_375 = t0_0101110111;
assign input_376 = t0_0101111000;
assign input_377 = t0_0101111001;
assign input_378 = t0_0101111010;
assign input_379 = t0_0101111011;
assign input_380 = t0_0101111100;
assign input_381 = t0_0101111101;
assign input_382 = t0_0101111110;
assign input_383 = t0_0101111111;
assign input_384 = t0_0110000000;
assign input_385 = t0_0110000001;
assign input_386 = t0_0110000010;
assign input_387 = t0_0110000011;
assign input_388 = t0_0110000100;
assign input_389 = t0_0110000101;
assign input_390 = t0_0110000110;
assign input_391 = t0_0110000111;
assign input_392 = t0_0110001000;
assign input_393 = t0_0110001001;
assign input_394 = t0_0110001010;
assign input_395 = t0_0110001011;
assign input_396 = t0_0110001100;
assign input_397 = t0_0110001101;
assign input_398 = t0_0110001110;
assign input_399 = t0_0110001111;
assign input_400 = t0_0110010000;
assign input_401 = t0_0110010001;
assign input_402 = t0_0110010010;
assign input_403 = t0_0110010011;
assign input_404 = t0_0110010100;
assign input_405 = t0_0110010101;
assign input_406 = t0_0110010110;
assign input_407 = t0_0110010111;
assign input_408 = t0_0110011000;
assign input_409 = t0_0110011001;
assign input_410 = t0_0110011010;
assign input_411 = t0_0110011011;
assign input_412 = t0_0110011100;
assign input_413 = t0_0110011101;
assign input_414 = t0_0110011110;
assign input_415 = t0_0110011111;
assign input_416 = t0_0110100000;
assign input_417 = t0_0110100001;
assign input_418 = t0_0110100010;
assign input_419 = t0_0110100011;
assign input_420 = t0_0110100100;
assign input_421 = t0_0110100101;
assign input_422 = t0_0110100110;
assign input_423 = t0_0110100111;
assign input_424 = t0_0110101000;
assign input_425 = t0_0110101001;
assign input_426 = t0_0110101010;
assign input_427 = t0_0110101011;
assign input_428 = t0_0110101100;
assign input_429 = t0_0110101101;
assign input_430 = t0_0110101110;
assign input_431 = t0_0110101111;
assign input_432 = t0_0110110000;
assign input_433 = t0_0110110001;
assign input_434 = t0_0110110010;
assign input_435 = t0_0110110011;
assign input_436 = t0_0110110100;
assign input_437 = t0_0110110101;
assign input_438 = t0_0110110110;
assign input_439 = t0_0110110111;
assign input_440 = t0_0110111000;
assign input_441 = t0_0110111001;
assign input_442 = t0_0110111010;
assign input_443 = t0_0110111011;
assign input_444 = t0_0110111100;
assign input_445 = t0_0110111101;
assign input_446 = t0_0110111110;
assign input_447 = t0_0110111111;
assign input_448 = t0_0111000000;
assign input_449 = t0_0111000001;
assign input_450 = t0_0111000010;
assign input_451 = t0_0111000011;
assign input_452 = t0_0111000100;
assign input_453 = t0_0111000101;
assign input_454 = t0_0111000110;
assign input_455 = t0_0111000111;
assign input_456 = t0_0111001000;
assign input_457 = t0_0111001001;
assign input_458 = t0_0111001010;
assign input_459 = t0_0111001011;
assign input_460 = t0_0111001100;
assign input_461 = t0_0111001101;
assign input_462 = t0_0111001110;
assign input_463 = t0_0111001111;
assign input_464 = t0_0111010000;
assign input_465 = t0_0111010001;
assign input_466 = t0_0111010010;
assign input_467 = t0_0111010011;
assign input_468 = t0_0111010100;
assign input_469 = t0_0111010101;
assign input_470 = t0_0111010110;
assign input_471 = t0_0111010111;
assign input_472 = t0_0111011000;
assign input_473 = t0_0111011001;
assign input_474 = t0_0111011010;
assign input_475 = t0_0111011011;
assign input_476 = t0_0111011100;
assign input_477 = t0_0111011101;
assign input_478 = t0_0111011110;
assign input_479 = t0_0111011111;
assign input_480 = t0_0111100000;
assign input_481 = t0_0111100001;
assign input_482 = t0_0111100010;
assign input_483 = t0_0111100011;
assign input_484 = t0_0111100100;
assign input_485 = t0_0111100101;
assign input_486 = t0_0111100110;
assign input_487 = t0_0111100111;
assign input_488 = t0_0111101000;
assign input_489 = t0_0111101001;
assign input_490 = t0_0111101010;
assign input_491 = t0_0111101011;
assign input_492 = t0_0111101100;
assign input_493 = t0_0111101101;
assign input_494 = t0_0111101110;
assign input_495 = t0_0111101111;
assign input_496 = t0_0111110000;
assign input_497 = t0_0111110001;
assign input_498 = t0_0111110010;
assign input_499 = t0_0111110011;
assign input_500 = t0_0111110100;
assign input_501 = t0_0111110101;
assign input_502 = t0_0111110110;
assign input_503 = t0_0111110111;
assign input_504 = t0_0111111000;
assign input_505 = t0_0111111001;
assign input_506 = t0_0111111010;
assign input_507 = t0_0111111011;
assign input_508 = t0_0111111100;
assign input_509 = t0_0111111101;
assign input_510 = t0_0111111110;
assign input_511 = t0_0111111111;
endmodule
