module chain_32 (
inout k0, k32
);
wire {wires};
chamber ch0 (.in(k0), .out(k1)
chamber ch1 (.in(k1), .out(k2)
chamber ch2 (.in(k2), .out(k3)
chamber ch3 (.in(k3), .out(k4)
chamber ch4 (.in(k4), .out(k5)
chamber ch5 (.in(k5), .out(k6)
chamber ch6 (.in(k6), .out(k7)
chamber ch7 (.in(k7), .out(k8)
chamber ch8 (.in(k8), .out(k9)
chamber ch9 (.in(k9), .out(k10)
chamber ch10 (.in(k10), .out(k11)
chamber ch11 (.in(k11), .out(k12)
chamber ch12 (.in(k12), .out(k13)
chamber ch13 (.in(k13), .out(k14)
chamber ch14 (.in(k14), .out(k15)
chamber ch15 (.in(k15), .out(k16)
chamber ch16 (.in(k16), .out(k17)
chamber ch17 (.in(k17), .out(k18)
chamber ch18 (.in(k18), .out(k19)
chamber ch19 (.in(k19), .out(k20)
chamber ch20 (.in(k20), .out(k21)
chamber ch21 (.in(k21), .out(k22)
chamber ch22 (.in(k22), .out(k23)
chamber ch23 (.in(k23), .out(k24)
chamber ch24 (.in(k24), .out(k25)
chamber ch25 (.in(k25), .out(k26)
chamber ch26 (.in(k26), .out(k27)
chamber ch27 (.in(k27), .out(k28)
chamber ch28 (.in(k28), .out(k29)
chamber ch29 (.in(k29), .out(k30)
chamber ch30 (.in(k30), .out(k31)
chamber ch31 (.in(k31), .out(k32)
endmodule
