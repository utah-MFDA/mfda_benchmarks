module complete_4 (
inout io_0,inout io_1,inout io_2,inout io_3
);
assign io_0 = input_0;
assign io_0 = input_1;
assign io_0 = input_2;
assign io_0 = input_3;
assign io_1 = input_1;
assign io_1 = input_2;
assign io_1 = input_3;
assign io_2 = input_2;
assign io_2 = input_3;
assign io_3 = input_3;
endmodule
