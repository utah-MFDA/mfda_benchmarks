module binary_tree_8_4 (
output out_0,output out_1,output out_2,output out_3,output out_4,output out_5,output out_6,output out_7,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63,input input_64,input input_65,input input_66,input input_67,input input_68,input input_69,input input_70,input input_71,input input_72,input input_73,input input_74,input input_75,input input_76,input input_77,input input_78,input input_79,input input_80,input input_81,input input_82,input input_83,input input_84,input input_85,input input_86,input input_87,input input_88,input input_89,input input_90,input input_91,input input_92,input input_93,input input_94,input input_95,input input_96,input input_97,input input_98,input input_99,input input_100,input input_101,input input_102,input input_103,input input_104,input input_105,input input_106,input input_107,input input_108,input input_109,input input_110,input input_111,input input_112,input input_113,input input_114,input input_115,input input_116,input input_117,input input_118,input input_119,input input_120,input input_121,input input_122,input input_123,input input_124,input input_125,input input_126,input input_127
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t1_0 (.a(t1_00), .b(t1_01), .y(t1_0));
wire t1_00, t1_01;
mixer mix_t1_00 (.a(t1_000), .b(t1_001), .y(t1_00));
wire t1_000, t1_001;
mixer mix_t1_000 (.a(t1_0000), .b(t1_0001), .y(t1_000));
wire t1_0000, t1_0001;
mixer mix_t1_0000 (.a(t1_00000), .b(t1_00001), .y(t1_0000));
wire t1_00000, t1_00001;
mixer mix_t1_0001 (.a(t1_00010), .b(t1_00011), .y(t1_0001));
wire t1_00010, t1_00011;
mixer mix_t1_001 (.a(t1_0010), .b(t1_0011), .y(t1_001));
wire t1_0010, t1_0011;
mixer mix_t1_0010 (.a(t1_00100), .b(t1_00101), .y(t1_0010));
wire t1_00100, t1_00101;
mixer mix_t1_0011 (.a(t1_00110), .b(t1_00111), .y(t1_0011));
wire t1_00110, t1_00111;
mixer mix_t1_01 (.a(t1_010), .b(t1_011), .y(t1_01));
wire t1_010, t1_011;
mixer mix_t1_010 (.a(t1_0100), .b(t1_0101), .y(t1_010));
wire t1_0100, t1_0101;
mixer mix_t1_0100 (.a(t1_01000), .b(t1_01001), .y(t1_0100));
wire t1_01000, t1_01001;
mixer mix_t1_0101 (.a(t1_01010), .b(t1_01011), .y(t1_0101));
wire t1_01010, t1_01011;
mixer mix_t1_011 (.a(t1_0110), .b(t1_0111), .y(t1_011));
wire t1_0110, t1_0111;
mixer mix_t1_0110 (.a(t1_01100), .b(t1_01101), .y(t1_0110));
wire t1_01100, t1_01101;
mixer mix_t1_0111 (.a(t1_01110), .b(t1_01111), .y(t1_0111));
wire t1_01110, t1_01111;
mixer mix_t2_0 (.a(t2_00), .b(t2_01), .y(t2_0));
wire t2_00, t2_01;
mixer mix_t2_00 (.a(t2_000), .b(t2_001), .y(t2_00));
wire t2_000, t2_001;
mixer mix_t2_000 (.a(t2_0000), .b(t2_0001), .y(t2_000));
wire t2_0000, t2_0001;
mixer mix_t2_0000 (.a(t2_00000), .b(t2_00001), .y(t2_0000));
wire t2_00000, t2_00001;
mixer mix_t2_0001 (.a(t2_00010), .b(t2_00011), .y(t2_0001));
wire t2_00010, t2_00011;
mixer mix_t2_001 (.a(t2_0010), .b(t2_0011), .y(t2_001));
wire t2_0010, t2_0011;
mixer mix_t2_0010 (.a(t2_00100), .b(t2_00101), .y(t2_0010));
wire t2_00100, t2_00101;
mixer mix_t2_0011 (.a(t2_00110), .b(t2_00111), .y(t2_0011));
wire t2_00110, t2_00111;
mixer mix_t2_01 (.a(t2_010), .b(t2_011), .y(t2_01));
wire t2_010, t2_011;
mixer mix_t2_010 (.a(t2_0100), .b(t2_0101), .y(t2_010));
wire t2_0100, t2_0101;
mixer mix_t2_0100 (.a(t2_01000), .b(t2_01001), .y(t2_0100));
wire t2_01000, t2_01001;
mixer mix_t2_0101 (.a(t2_01010), .b(t2_01011), .y(t2_0101));
wire t2_01010, t2_01011;
mixer mix_t2_011 (.a(t2_0110), .b(t2_0111), .y(t2_011));
wire t2_0110, t2_0111;
mixer mix_t2_0110 (.a(t2_01100), .b(t2_01101), .y(t2_0110));
wire t2_01100, t2_01101;
mixer mix_t2_0111 (.a(t2_01110), .b(t2_01111), .y(t2_0111));
wire t2_01110, t2_01111;
mixer mix_t3_0 (.a(t3_00), .b(t3_01), .y(t3_0));
wire t3_00, t3_01;
mixer mix_t3_00 (.a(t3_000), .b(t3_001), .y(t3_00));
wire t3_000, t3_001;
mixer mix_t3_000 (.a(t3_0000), .b(t3_0001), .y(t3_000));
wire t3_0000, t3_0001;
mixer mix_t3_0000 (.a(t3_00000), .b(t3_00001), .y(t3_0000));
wire t3_00000, t3_00001;
mixer mix_t3_0001 (.a(t3_00010), .b(t3_00011), .y(t3_0001));
wire t3_00010, t3_00011;
mixer mix_t3_001 (.a(t3_0010), .b(t3_0011), .y(t3_001));
wire t3_0010, t3_0011;
mixer mix_t3_0010 (.a(t3_00100), .b(t3_00101), .y(t3_0010));
wire t3_00100, t3_00101;
mixer mix_t3_0011 (.a(t3_00110), .b(t3_00111), .y(t3_0011));
wire t3_00110, t3_00111;
mixer mix_t3_01 (.a(t3_010), .b(t3_011), .y(t3_01));
wire t3_010, t3_011;
mixer mix_t3_010 (.a(t3_0100), .b(t3_0101), .y(t3_010));
wire t3_0100, t3_0101;
mixer mix_t3_0100 (.a(t3_01000), .b(t3_01001), .y(t3_0100));
wire t3_01000, t3_01001;
mixer mix_t3_0101 (.a(t3_01010), .b(t3_01011), .y(t3_0101));
wire t3_01010, t3_01011;
mixer mix_t3_011 (.a(t3_0110), .b(t3_0111), .y(t3_011));
wire t3_0110, t3_0111;
mixer mix_t3_0110 (.a(t3_01100), .b(t3_01101), .y(t3_0110));
wire t3_01100, t3_01101;
mixer mix_t3_0111 (.a(t3_01110), .b(t3_01111), .y(t3_0111));
wire t3_01110, t3_01111;
mixer mix_t4_0 (.a(t4_00), .b(t4_01), .y(t4_0));
wire t4_00, t4_01;
mixer mix_t4_00 (.a(t4_000), .b(t4_001), .y(t4_00));
wire t4_000, t4_001;
mixer mix_t4_000 (.a(t4_0000), .b(t4_0001), .y(t4_000));
wire t4_0000, t4_0001;
mixer mix_t4_0000 (.a(t4_00000), .b(t4_00001), .y(t4_0000));
wire t4_00000, t4_00001;
mixer mix_t4_0001 (.a(t4_00010), .b(t4_00011), .y(t4_0001));
wire t4_00010, t4_00011;
mixer mix_t4_001 (.a(t4_0010), .b(t4_0011), .y(t4_001));
wire t4_0010, t4_0011;
mixer mix_t4_0010 (.a(t4_00100), .b(t4_00101), .y(t4_0010));
wire t4_00100, t4_00101;
mixer mix_t4_0011 (.a(t4_00110), .b(t4_00111), .y(t4_0011));
wire t4_00110, t4_00111;
mixer mix_t4_01 (.a(t4_010), .b(t4_011), .y(t4_01));
wire t4_010, t4_011;
mixer mix_t4_010 (.a(t4_0100), .b(t4_0101), .y(t4_010));
wire t4_0100, t4_0101;
mixer mix_t4_0100 (.a(t4_01000), .b(t4_01001), .y(t4_0100));
wire t4_01000, t4_01001;
mixer mix_t4_0101 (.a(t4_01010), .b(t4_01011), .y(t4_0101));
wire t4_01010, t4_01011;
mixer mix_t4_011 (.a(t4_0110), .b(t4_0111), .y(t4_011));
wire t4_0110, t4_0111;
mixer mix_t4_0110 (.a(t4_01100), .b(t4_01101), .y(t4_0110));
wire t4_01100, t4_01101;
mixer mix_t4_0111 (.a(t4_01110), .b(t4_01111), .y(t4_0111));
wire t4_01110, t4_01111;
mixer mix_t5_0 (.a(t5_00), .b(t5_01), .y(t5_0));
wire t5_00, t5_01;
mixer mix_t5_00 (.a(t5_000), .b(t5_001), .y(t5_00));
wire t5_000, t5_001;
mixer mix_t5_000 (.a(t5_0000), .b(t5_0001), .y(t5_000));
wire t5_0000, t5_0001;
mixer mix_t5_0000 (.a(t5_00000), .b(t5_00001), .y(t5_0000));
wire t5_00000, t5_00001;
mixer mix_t5_0001 (.a(t5_00010), .b(t5_00011), .y(t5_0001));
wire t5_00010, t5_00011;
mixer mix_t5_001 (.a(t5_0010), .b(t5_0011), .y(t5_001));
wire t5_0010, t5_0011;
mixer mix_t5_0010 (.a(t5_00100), .b(t5_00101), .y(t5_0010));
wire t5_00100, t5_00101;
mixer mix_t5_0011 (.a(t5_00110), .b(t5_00111), .y(t5_0011));
wire t5_00110, t5_00111;
mixer mix_t5_01 (.a(t5_010), .b(t5_011), .y(t5_01));
wire t5_010, t5_011;
mixer mix_t5_010 (.a(t5_0100), .b(t5_0101), .y(t5_010));
wire t5_0100, t5_0101;
mixer mix_t5_0100 (.a(t5_01000), .b(t5_01001), .y(t5_0100));
wire t5_01000, t5_01001;
mixer mix_t5_0101 (.a(t5_01010), .b(t5_01011), .y(t5_0101));
wire t5_01010, t5_01011;
mixer mix_t5_011 (.a(t5_0110), .b(t5_0111), .y(t5_011));
wire t5_0110, t5_0111;
mixer mix_t5_0110 (.a(t5_01100), .b(t5_01101), .y(t5_0110));
wire t5_01100, t5_01101;
mixer mix_t5_0111 (.a(t5_01110), .b(t5_01111), .y(t5_0111));
wire t5_01110, t5_01111;
mixer mix_t6_0 (.a(t6_00), .b(t6_01), .y(t6_0));
wire t6_00, t6_01;
mixer mix_t6_00 (.a(t6_000), .b(t6_001), .y(t6_00));
wire t6_000, t6_001;
mixer mix_t6_000 (.a(t6_0000), .b(t6_0001), .y(t6_000));
wire t6_0000, t6_0001;
mixer mix_t6_0000 (.a(t6_00000), .b(t6_00001), .y(t6_0000));
wire t6_00000, t6_00001;
mixer mix_t6_0001 (.a(t6_00010), .b(t6_00011), .y(t6_0001));
wire t6_00010, t6_00011;
mixer mix_t6_001 (.a(t6_0010), .b(t6_0011), .y(t6_001));
wire t6_0010, t6_0011;
mixer mix_t6_0010 (.a(t6_00100), .b(t6_00101), .y(t6_0010));
wire t6_00100, t6_00101;
mixer mix_t6_0011 (.a(t6_00110), .b(t6_00111), .y(t6_0011));
wire t6_00110, t6_00111;
mixer mix_t6_01 (.a(t6_010), .b(t6_011), .y(t6_01));
wire t6_010, t6_011;
mixer mix_t6_010 (.a(t6_0100), .b(t6_0101), .y(t6_010));
wire t6_0100, t6_0101;
mixer mix_t6_0100 (.a(t6_01000), .b(t6_01001), .y(t6_0100));
wire t6_01000, t6_01001;
mixer mix_t6_0101 (.a(t6_01010), .b(t6_01011), .y(t6_0101));
wire t6_01010, t6_01011;
mixer mix_t6_011 (.a(t6_0110), .b(t6_0111), .y(t6_011));
wire t6_0110, t6_0111;
mixer mix_t6_0110 (.a(t6_01100), .b(t6_01101), .y(t6_0110));
wire t6_01100, t6_01101;
mixer mix_t6_0111 (.a(t6_01110), .b(t6_01111), .y(t6_0111));
wire t6_01110, t6_01111;
mixer mix_t7_0 (.a(t7_00), .b(t7_01), .y(t7_0));
wire t7_00, t7_01;
mixer mix_t7_00 (.a(t7_000), .b(t7_001), .y(t7_00));
wire t7_000, t7_001;
mixer mix_t7_000 (.a(t7_0000), .b(t7_0001), .y(t7_000));
wire t7_0000, t7_0001;
mixer mix_t7_0000 (.a(t7_00000), .b(t7_00001), .y(t7_0000));
wire t7_00000, t7_00001;
mixer mix_t7_0001 (.a(t7_00010), .b(t7_00011), .y(t7_0001));
wire t7_00010, t7_00011;
mixer mix_t7_001 (.a(t7_0010), .b(t7_0011), .y(t7_001));
wire t7_0010, t7_0011;
mixer mix_t7_0010 (.a(t7_00100), .b(t7_00101), .y(t7_0010));
wire t7_00100, t7_00101;
mixer mix_t7_0011 (.a(t7_00110), .b(t7_00111), .y(t7_0011));
wire t7_00110, t7_00111;
mixer mix_t7_01 (.a(t7_010), .b(t7_011), .y(t7_01));
wire t7_010, t7_011;
mixer mix_t7_010 (.a(t7_0100), .b(t7_0101), .y(t7_010));
wire t7_0100, t7_0101;
mixer mix_t7_0100 (.a(t7_01000), .b(t7_01001), .y(t7_0100));
wire t7_01000, t7_01001;
mixer mix_t7_0101 (.a(t7_01010), .b(t7_01011), .y(t7_0101));
wire t7_01010, t7_01011;
mixer mix_t7_011 (.a(t7_0110), .b(t7_0111), .y(t7_011));
wire t7_0110, t7_0111;
mixer mix_t7_0110 (.a(t7_01100), .b(t7_01101), .y(t7_0110));
wire t7_01100, t7_01101;
mixer mix_t7_0111 (.a(t7_01110), .b(t7_01111), .y(t7_0111));
wire t7_01110, t7_01111;
wire t0_0;
assign out_0 = t0_0;
wire t1_0;
assign out_1 = t1_0;
wire t2_0;
assign out_2 = t2_0;
wire t3_0;
assign out_3 = t3_0;
wire t4_0;
assign out_4 = t4_0;
wire t5_0;
assign out_5 = t5_0;
wire t6_0;
assign out_6 = t6_0;
wire t7_0;
assign out_7 = t7_0;
assign input_0 = t0_00000;
assign input_1 = t0_00001;
assign input_2 = t0_00010;
assign input_3 = t0_00011;
assign input_4 = t0_00100;
assign input_5 = t0_00101;
assign input_6 = t0_00110;
assign input_7 = t0_00111;
assign input_8 = t0_01000;
assign input_9 = t0_01001;
assign input_10 = t0_01010;
assign input_11 = t0_01011;
assign input_12 = t0_01100;
assign input_13 = t0_01101;
assign input_14 = t0_01110;
assign input_15 = t0_01111;
assign input_16 = t1_00000;
assign input_17 = t1_00001;
assign input_18 = t1_00010;
assign input_19 = t1_00011;
assign input_20 = t1_00100;
assign input_21 = t1_00101;
assign input_22 = t1_00110;
assign input_23 = t1_00111;
assign input_24 = t1_01000;
assign input_25 = t1_01001;
assign input_26 = t1_01010;
assign input_27 = t1_01011;
assign input_28 = t1_01100;
assign input_29 = t1_01101;
assign input_30 = t1_01110;
assign input_31 = t1_01111;
assign input_32 = t2_00000;
assign input_33 = t2_00001;
assign input_34 = t2_00010;
assign input_35 = t2_00011;
assign input_36 = t2_00100;
assign input_37 = t2_00101;
assign input_38 = t2_00110;
assign input_39 = t2_00111;
assign input_40 = t2_01000;
assign input_41 = t2_01001;
assign input_42 = t2_01010;
assign input_43 = t2_01011;
assign input_44 = t2_01100;
assign input_45 = t2_01101;
assign input_46 = t2_01110;
assign input_47 = t2_01111;
assign input_48 = t3_00000;
assign input_49 = t3_00001;
assign input_50 = t3_00010;
assign input_51 = t3_00011;
assign input_52 = t3_00100;
assign input_53 = t3_00101;
assign input_54 = t3_00110;
assign input_55 = t3_00111;
assign input_56 = t3_01000;
assign input_57 = t3_01001;
assign input_58 = t3_01010;
assign input_59 = t3_01011;
assign input_60 = t3_01100;
assign input_61 = t3_01101;
assign input_62 = t3_01110;
assign input_63 = t3_01111;
assign input_64 = t4_00000;
assign input_65 = t4_00001;
assign input_66 = t4_00010;
assign input_67 = t4_00011;
assign input_68 = t4_00100;
assign input_69 = t4_00101;
assign input_70 = t4_00110;
assign input_71 = t4_00111;
assign input_72 = t4_01000;
assign input_73 = t4_01001;
assign input_74 = t4_01010;
assign input_75 = t4_01011;
assign input_76 = t4_01100;
assign input_77 = t4_01101;
assign input_78 = t4_01110;
assign input_79 = t4_01111;
assign input_80 = t5_00000;
assign input_81 = t5_00001;
assign input_82 = t5_00010;
assign input_83 = t5_00011;
assign input_84 = t5_00100;
assign input_85 = t5_00101;
assign input_86 = t5_00110;
assign input_87 = t5_00111;
assign input_88 = t5_01000;
assign input_89 = t5_01001;
assign input_90 = t5_01010;
assign input_91 = t5_01011;
assign input_92 = t5_01100;
assign input_93 = t5_01101;
assign input_94 = t5_01110;
assign input_95 = t5_01111;
assign input_96 = t6_00000;
assign input_97 = t6_00001;
assign input_98 = t6_00010;
assign input_99 = t6_00011;
assign input_100 = t6_00100;
assign input_101 = t6_00101;
assign input_102 = t6_00110;
assign input_103 = t6_00111;
assign input_104 = t6_01000;
assign input_105 = t6_01001;
assign input_106 = t6_01010;
assign input_107 = t6_01011;
assign input_108 = t6_01100;
assign input_109 = t6_01101;
assign input_110 = t6_01110;
assign input_111 = t6_01111;
assign input_112 = t7_00000;
assign input_113 = t7_00001;
assign input_114 = t7_00010;
assign input_115 = t7_00011;
assign input_116 = t7_00100;
assign input_117 = t7_00101;
assign input_118 = t7_00110;
assign input_119 = t7_00111;
assign input_120 = t7_01000;
assign input_121 = t7_01001;
assign input_122 = t7_01010;
assign input_123 = t7_01011;
assign input_124 = t7_01100;
assign input_125 = t7_01101;
assign input_126 = t7_01110;
assign input_127 = t7_01111;
endmodule
