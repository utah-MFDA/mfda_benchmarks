module DROPLET_GENERATOR_FLOW_FOCUS(inout port0, port1, port2, port3);
endmodule

module DROPLET_GENERATOR_T()
module GRADIENT_GENERATOR()

module LONG_CELL_TRAP 2port
module MIXER 2port
module MUX 25, 5, 9, 15, ports
module NODE, 4, 2, 3,
module ROTARY_MIXER 7 ports
module SQUARE_CELL_TRAP 4 ports
module TREE 5, 3, 9 ports
module VALVE 3 ports
