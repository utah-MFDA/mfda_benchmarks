module fanout2_braid_3_512 (
output output_0,output output_1,output output_2,input input_0,input input_1,input input_2
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_1_2, output_1_0, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_0), .y(output_0_2));
wire output_2_2, output_2_0, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_0), .y(output_1_2));
wire output_3_2, output_3_0, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_0), .y(output_2_2));
wire output_1_3, output_1_1, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_1), .y(output_0_3));
wire output_2_3, output_2_1, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_1), .y(output_1_3));
wire output_3_3, output_3_1, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_1), .y(output_2_3));
wire output_1_4, output_1_2, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_2), .y(output_0_4));
wire output_2_4, output_2_2, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_2), .y(output_1_4));
wire output_3_4, output_3_2, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_2), .y(output_2_4));
wire output_1_5, output_1_0, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_0), .y(output_0_5));
wire output_2_5, output_2_0, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_0), .y(output_1_5));
wire output_3_5, output_3_0, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_0), .y(output_2_5));
wire output_1_6, output_1_1, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_1), .y(output_0_6));
wire output_2_6, output_2_1, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_1), .y(output_1_6));
wire output_3_6, output_3_1, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_1), .y(output_2_6));
wire output_1_7, output_1_2, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_2), .y(output_0_7));
wire output_2_7, output_2_2, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_2), .y(output_1_7));
wire output_3_7, output_3_2, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_2), .y(output_2_7));
wire output_1_8, output_1_0, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_0), .y(output_0_8));
wire output_2_8, output_2_0, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_0), .y(output_1_8));
wire output_3_8, output_3_0, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_0), .y(output_2_8));
wire output_1_9, output_1_1, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_1), .y(output_0_9));
wire output_2_9, output_2_1, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_1), .y(output_1_9));
wire output_3_9, output_3_1, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_1), .y(output_2_9));
wire output_1_10, output_1_2, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_2), .y(output_0_10));
wire output_2_10, output_2_2, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_2), .y(output_1_10));
wire output_3_10, output_3_2, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_2), .y(output_2_10));
wire output_1_11, output_1_0, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_0), .y(output_0_11));
wire output_2_11, output_2_0, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_0), .y(output_1_11));
wire output_3_11, output_3_0, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_0), .y(output_2_11));
wire output_1_12, output_1_1, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_1), .y(output_0_12));
wire output_2_12, output_2_1, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_1), .y(output_1_12));
wire output_3_12, output_3_1, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_1), .y(output_2_12));
wire output_1_13, output_1_2, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_2), .y(output_0_13));
wire output_2_13, output_2_2, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_2), .y(output_1_13));
wire output_3_13, output_3_2, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_2), .y(output_2_13));
wire output_1_14, output_1_0, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_0), .y(output_0_14));
wire output_2_14, output_2_0, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_0), .y(output_1_14));
wire output_3_14, output_3_0, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_0), .y(output_2_14));
wire output_1_15, output_1_1, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_1), .y(output_0_15));
wire output_2_15, output_2_1, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_1), .y(output_1_15));
wire output_3_15, output_3_1, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_1), .y(output_2_15));
wire output_1_16, output_1_2, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_2), .y(output_0_16));
wire output_2_16, output_2_2, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_2), .y(output_1_16));
wire output_3_16, output_3_2, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_2), .y(output_2_16));
wire output_1_17, output_1_0, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_0), .y(output_0_17));
wire output_2_17, output_2_0, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_0), .y(output_1_17));
wire output_3_17, output_3_0, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_0), .y(output_2_17));
wire output_1_18, output_1_1, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_1), .y(output_0_18));
wire output_2_18, output_2_1, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_1), .y(output_1_18));
wire output_3_18, output_3_1, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_1), .y(output_2_18));
wire output_1_19, output_1_2, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_2), .y(output_0_19));
wire output_2_19, output_2_2, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_2), .y(output_1_19));
wire output_3_19, output_3_2, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_2), .y(output_2_19));
wire output_1_20, output_1_0, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_0), .y(output_0_20));
wire output_2_20, output_2_0, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_0), .y(output_1_20));
wire output_3_20, output_3_0, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_0), .y(output_2_20));
wire output_1_21, output_1_1, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_1), .y(output_0_21));
wire output_2_21, output_2_1, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_1), .y(output_1_21));
wire output_3_21, output_3_1, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_1), .y(output_2_21));
wire output_1_22, output_1_2, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_2), .y(output_0_22));
wire output_2_22, output_2_2, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_2), .y(output_1_22));
wire output_3_22, output_3_2, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_2), .y(output_2_22));
wire output_1_23, output_1_0, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_0), .y(output_0_23));
wire output_2_23, output_2_0, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_0), .y(output_1_23));
wire output_3_23, output_3_0, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_0), .y(output_2_23));
wire output_1_24, output_1_1, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_1), .y(output_0_24));
wire output_2_24, output_2_1, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_1), .y(output_1_24));
wire output_3_24, output_3_1, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_1), .y(output_2_24));
wire output_1_25, output_1_2, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_2), .y(output_0_25));
wire output_2_25, output_2_2, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_2), .y(output_1_25));
wire output_3_25, output_3_2, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_2), .y(output_2_25));
wire output_1_26, output_1_0, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_0), .y(output_0_26));
wire output_2_26, output_2_0, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_0), .y(output_1_26));
wire output_3_26, output_3_0, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_0), .y(output_2_26));
wire output_1_27, output_1_1, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_1), .y(output_0_27));
wire output_2_27, output_2_1, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_1), .y(output_1_27));
wire output_3_27, output_3_1, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_1), .y(output_2_27));
wire output_1_28, output_1_2, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_2), .y(output_0_28));
wire output_2_28, output_2_2, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_2), .y(output_1_28));
wire output_3_28, output_3_2, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_2), .y(output_2_28));
wire output_1_29, output_1_0, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_0), .y(output_0_29));
wire output_2_29, output_2_0, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_0), .y(output_1_29));
wire output_3_29, output_3_0, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_0), .y(output_2_29));
wire output_1_30, output_1_1, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_1), .y(output_0_30));
wire output_2_30, output_2_1, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_1), .y(output_1_30));
wire output_3_30, output_3_1, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_1), .y(output_2_30));
wire output_1_31, output_1_2, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_2), .y(output_0_31));
wire output_2_31, output_2_2, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_2), .y(output_1_31));
wire output_3_31, output_3_2, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_2), .y(output_2_31));
wire output_1_32, output_1_0, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_0), .y(output_0_32));
wire output_2_32, output_2_0, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_0), .y(output_1_32));
wire output_3_32, output_3_0, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_0), .y(output_2_32));
wire output_1_33, output_1_1, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_1), .y(output_0_33));
wire output_2_33, output_2_1, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_1), .y(output_1_33));
wire output_3_33, output_3_1, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_1), .y(output_2_33));
wire output_1_34, output_1_2, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_2), .y(output_0_34));
wire output_2_34, output_2_2, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_2), .y(output_1_34));
wire output_3_34, output_3_2, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_2), .y(output_2_34));
wire output_1_35, output_1_0, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_0), .y(output_0_35));
wire output_2_35, output_2_0, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_0), .y(output_1_35));
wire output_3_35, output_3_0, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_0), .y(output_2_35));
wire output_1_36, output_1_1, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_1), .y(output_0_36));
wire output_2_36, output_2_1, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_1), .y(output_1_36));
wire output_3_36, output_3_1, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_1), .y(output_2_36));
wire output_1_37, output_1_2, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_2), .y(output_0_37));
wire output_2_37, output_2_2, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_2), .y(output_1_37));
wire output_3_37, output_3_2, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_2), .y(output_2_37));
wire output_1_38, output_1_0, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_0), .y(output_0_38));
wire output_2_38, output_2_0, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_0), .y(output_1_38));
wire output_3_38, output_3_0, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_0), .y(output_2_38));
wire output_1_39, output_1_1, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_1), .y(output_0_39));
wire output_2_39, output_2_1, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_1), .y(output_1_39));
wire output_3_39, output_3_1, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_1), .y(output_2_39));
wire output_1_40, output_1_2, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_2), .y(output_0_40));
wire output_2_40, output_2_2, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_2), .y(output_1_40));
wire output_3_40, output_3_2, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_2), .y(output_2_40));
wire output_1_41, output_1_0, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_0), .y(output_0_41));
wire output_2_41, output_2_0, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_0), .y(output_1_41));
wire output_3_41, output_3_0, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_0), .y(output_2_41));
wire output_1_42, output_1_1, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_1), .y(output_0_42));
wire output_2_42, output_2_1, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_1), .y(output_1_42));
wire output_3_42, output_3_1, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_1), .y(output_2_42));
wire output_1_43, output_1_2, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_2), .y(output_0_43));
wire output_2_43, output_2_2, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_2), .y(output_1_43));
wire output_3_43, output_3_2, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_2), .y(output_2_43));
wire output_1_44, output_1_0, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_0), .y(output_0_44));
wire output_2_44, output_2_0, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_0), .y(output_1_44));
wire output_3_44, output_3_0, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_0), .y(output_2_44));
wire output_1_45, output_1_1, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_1), .y(output_0_45));
wire output_2_45, output_2_1, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_1), .y(output_1_45));
wire output_3_45, output_3_1, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_1), .y(output_2_45));
wire output_1_46, output_1_2, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_2), .y(output_0_46));
wire output_2_46, output_2_2, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_2), .y(output_1_46));
wire output_3_46, output_3_2, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_2), .y(output_2_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_1_50, output_1_0, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_0), .y(output_0_50));
wire output_2_50, output_2_0, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_0), .y(output_1_50));
wire output_3_50, output_3_0, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_0), .y(output_2_50));
wire output_1_51, output_1_1, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_1), .y(output_0_51));
wire output_2_51, output_2_1, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_1), .y(output_1_51));
wire output_3_51, output_3_1, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_1), .y(output_2_51));
wire output_1_52, output_1_2, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_2), .y(output_0_52));
wire output_2_52, output_2_2, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_2), .y(output_1_52));
wire output_3_52, output_3_2, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_2), .y(output_2_52));
wire output_1_53, output_1_0, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_0), .y(output_0_53));
wire output_2_53, output_2_0, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_0), .y(output_1_53));
wire output_3_53, output_3_0, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_0), .y(output_2_53));
wire output_1_54, output_1_1, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_1), .y(output_0_54));
wire output_2_54, output_2_1, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_1), .y(output_1_54));
wire output_3_54, output_3_1, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_1), .y(output_2_54));
wire output_1_55, output_1_2, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_2), .y(output_0_55));
wire output_2_55, output_2_2, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_2), .y(output_1_55));
wire output_3_55, output_3_2, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_2), .y(output_2_55));
wire output_1_56, output_1_0, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_0), .y(output_0_56));
wire output_2_56, output_2_0, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_0), .y(output_1_56));
wire output_3_56, output_3_0, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_0), .y(output_2_56));
wire output_1_57, output_1_1, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_1), .y(output_0_57));
wire output_2_57, output_2_1, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_1), .y(output_1_57));
wire output_3_57, output_3_1, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_1), .y(output_2_57));
wire output_1_58, output_1_2, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_2), .y(output_0_58));
wire output_2_58, output_2_2, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_2), .y(output_1_58));
wire output_3_58, output_3_2, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_2), .y(output_2_58));
wire output_1_59, output_1_0, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_0), .y(output_0_59));
wire output_2_59, output_2_0, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_0), .y(output_1_59));
wire output_3_59, output_3_0, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_0), .y(output_2_59));
wire output_1_60, output_1_1, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_1), .y(output_0_60));
wire output_2_60, output_2_1, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_1), .y(output_1_60));
wire output_3_60, output_3_1, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_1), .y(output_2_60));
wire output_1_61, output_1_2, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_2), .y(output_0_61));
wire output_2_61, output_2_2, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_2), .y(output_1_61));
wire output_3_61, output_3_2, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_2), .y(output_2_61));
wire output_1_62, output_1_0, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_0), .y(output_0_62));
wire output_2_62, output_2_0, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_0), .y(output_1_62));
wire output_3_62, output_3_0, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_0), .y(output_2_62));
wire output_1_63, output_1_1, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_1), .y(output_0_63));
wire output_2_63, output_2_1, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_1), .y(output_1_63));
wire output_3_63, output_3_1, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_1), .y(output_2_63));
wire output_1_64, output_1_2, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_2), .y(output_0_64));
wire output_2_64, output_2_2, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_2), .y(output_1_64));
wire output_3_64, output_3_2, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_2), .y(output_2_64));
wire output_1_65, output_1_0, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_0), .y(output_0_65));
wire output_2_65, output_2_0, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_0), .y(output_1_65));
wire output_3_65, output_3_0, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_0), .y(output_2_65));
wire output_1_66, output_1_1, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_1), .y(output_0_66));
wire output_2_66, output_2_1, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_1), .y(output_1_66));
wire output_3_66, output_3_1, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_1), .y(output_2_66));
wire output_1_67, output_1_2, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_2), .y(output_0_67));
wire output_2_67, output_2_2, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_2), .y(output_1_67));
wire output_3_67, output_3_2, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_2), .y(output_2_67));
wire output_1_68, output_1_0, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_0), .y(output_0_68));
wire output_2_68, output_2_0, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_0), .y(output_1_68));
wire output_3_68, output_3_0, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_0), .y(output_2_68));
wire output_1_69, output_1_1, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_1), .y(output_0_69));
wire output_2_69, output_2_1, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_1), .y(output_1_69));
wire output_3_69, output_3_1, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_1), .y(output_2_69));
wire output_1_70, output_1_2, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_2), .y(output_0_70));
wire output_2_70, output_2_2, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_2), .y(output_1_70));
wire output_3_70, output_3_2, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_2), .y(output_2_70));
wire output_1_71, output_1_0, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_0), .y(output_0_71));
wire output_2_71, output_2_0, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_0), .y(output_1_71));
wire output_3_71, output_3_0, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_0), .y(output_2_71));
wire output_1_72, output_1_1, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_1), .y(output_0_72));
wire output_2_72, output_2_1, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_1), .y(output_1_72));
wire output_3_72, output_3_1, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_1), .y(output_2_72));
wire output_1_73, output_1_2, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_2), .y(output_0_73));
wire output_2_73, output_2_2, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_2), .y(output_1_73));
wire output_3_73, output_3_2, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_2), .y(output_2_73));
wire output_1_74, output_1_0, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_0), .y(output_0_74));
wire output_2_74, output_2_0, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_0), .y(output_1_74));
wire output_3_74, output_3_0, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_0), .y(output_2_74));
wire output_1_75, output_1_1, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_1), .y(output_0_75));
wire output_2_75, output_2_1, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_1), .y(output_1_75));
wire output_3_75, output_3_1, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_1), .y(output_2_75));
wire output_1_76, output_1_2, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_2), .y(output_0_76));
wire output_2_76, output_2_2, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_2), .y(output_1_76));
wire output_3_76, output_3_2, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_2), .y(output_2_76));
wire output_1_77, output_1_0, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_0), .y(output_0_77));
wire output_2_77, output_2_0, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_0), .y(output_1_77));
wire output_3_77, output_3_0, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_0), .y(output_2_77));
wire output_1_78, output_1_1, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_1), .y(output_0_78));
wire output_2_78, output_2_1, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_1), .y(output_1_78));
wire output_3_78, output_3_1, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_1), .y(output_2_78));
wire output_1_79, output_1_2, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_2), .y(output_0_79));
wire output_2_79, output_2_2, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_2), .y(output_1_79));
wire output_3_79, output_3_2, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_2), .y(output_2_79));
wire output_1_80, output_1_0, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_0), .y(output_0_80));
wire output_2_80, output_2_0, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_0), .y(output_1_80));
wire output_3_80, output_3_0, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_0), .y(output_2_80));
wire output_1_81, output_1_1, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_1), .y(output_0_81));
wire output_2_81, output_2_1, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_1), .y(output_1_81));
wire output_3_81, output_3_1, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_1), .y(output_2_81));
wire output_1_82, output_1_2, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_2), .y(output_0_82));
wire output_2_82, output_2_2, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_2), .y(output_1_82));
wire output_3_82, output_3_2, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_2), .y(output_2_82));
wire output_1_83, output_1_0, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_0), .y(output_0_83));
wire output_2_83, output_2_0, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_0), .y(output_1_83));
wire output_3_83, output_3_0, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_0), .y(output_2_83));
wire output_1_84, output_1_1, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_1), .y(output_0_84));
wire output_2_84, output_2_1, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_1), .y(output_1_84));
wire output_3_84, output_3_1, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_1), .y(output_2_84));
wire output_1_85, output_1_2, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_2), .y(output_0_85));
wire output_2_85, output_2_2, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_2), .y(output_1_85));
wire output_3_85, output_3_2, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_2), .y(output_2_85));
wire output_1_86, output_1_0, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_0), .y(output_0_86));
wire output_2_86, output_2_0, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_0), .y(output_1_86));
wire output_3_86, output_3_0, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_0), .y(output_2_86));
wire output_1_87, output_1_1, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_1), .y(output_0_87));
wire output_2_87, output_2_1, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_1), .y(output_1_87));
wire output_3_87, output_3_1, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_1), .y(output_2_87));
wire output_1_88, output_1_2, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_2), .y(output_0_88));
wire output_2_88, output_2_2, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_2), .y(output_1_88));
wire output_3_88, output_3_2, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_2), .y(output_2_88));
wire output_1_89, output_1_0, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_0), .y(output_0_89));
wire output_2_89, output_2_0, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_0), .y(output_1_89));
wire output_3_89, output_3_0, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_0), .y(output_2_89));
wire output_1_90, output_1_1, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_1), .y(output_0_90));
wire output_2_90, output_2_1, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_1), .y(output_1_90));
wire output_3_90, output_3_1, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_1), .y(output_2_90));
wire output_1_91, output_1_2, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_2), .y(output_0_91));
wire output_2_91, output_2_2, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_2), .y(output_1_91));
wire output_3_91, output_3_2, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_2), .y(output_2_91));
wire output_1_92, output_1_0, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_0), .y(output_0_92));
wire output_2_92, output_2_0, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_0), .y(output_1_92));
wire output_3_92, output_3_0, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_0), .y(output_2_92));
wire output_1_93, output_1_1, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_1), .y(output_0_93));
wire output_2_93, output_2_1, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_1), .y(output_1_93));
wire output_3_93, output_3_1, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_1), .y(output_2_93));
wire output_1_94, output_1_2, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_2), .y(output_0_94));
wire output_2_94, output_2_2, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_2), .y(output_1_94));
wire output_3_94, output_3_2, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_2), .y(output_2_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_1_96, output_1_1, output_0_96;
mixer gate_output_0_96(.a(output_1_96), .b(output_1_1), .y(output_0_96));
wire output_2_96, output_2_1, output_1_96;
mixer gate_output_1_96(.a(output_2_96), .b(output_2_1), .y(output_1_96));
wire output_3_96, output_3_1, output_2_96;
mixer gate_output_2_96(.a(output_3_96), .b(output_3_1), .y(output_2_96));
wire output_1_97, output_1_2, output_0_97;
mixer gate_output_0_97(.a(output_1_97), .b(output_1_2), .y(output_0_97));
wire output_2_97, output_2_2, output_1_97;
mixer gate_output_1_97(.a(output_2_97), .b(output_2_2), .y(output_1_97));
wire output_3_97, output_3_2, output_2_97;
mixer gate_output_2_97(.a(output_3_97), .b(output_3_2), .y(output_2_97));
wire output_1_98, output_1_0, output_0_98;
mixer gate_output_0_98(.a(output_1_98), .b(output_1_0), .y(output_0_98));
wire output_2_98, output_2_0, output_1_98;
mixer gate_output_1_98(.a(output_2_98), .b(output_2_0), .y(output_1_98));
wire output_3_98, output_3_0, output_2_98;
mixer gate_output_2_98(.a(output_3_98), .b(output_3_0), .y(output_2_98));
wire output_1_99, output_1_1, output_0_99;
mixer gate_output_0_99(.a(output_1_99), .b(output_1_1), .y(output_0_99));
wire output_2_99, output_2_1, output_1_99;
mixer gate_output_1_99(.a(output_2_99), .b(output_2_1), .y(output_1_99));
wire output_3_99, output_3_1, output_2_99;
mixer gate_output_2_99(.a(output_3_99), .b(output_3_1), .y(output_2_99));
wire output_1_100, output_1_2, output_0_100;
mixer gate_output_0_100(.a(output_1_100), .b(output_1_2), .y(output_0_100));
wire output_2_100, output_2_2, output_1_100;
mixer gate_output_1_100(.a(output_2_100), .b(output_2_2), .y(output_1_100));
wire output_3_100, output_3_2, output_2_100;
mixer gate_output_2_100(.a(output_3_100), .b(output_3_2), .y(output_2_100));
wire output_1_101, output_1_0, output_0_101;
mixer gate_output_0_101(.a(output_1_101), .b(output_1_0), .y(output_0_101));
wire output_2_101, output_2_0, output_1_101;
mixer gate_output_1_101(.a(output_2_101), .b(output_2_0), .y(output_1_101));
wire output_3_101, output_3_0, output_2_101;
mixer gate_output_2_101(.a(output_3_101), .b(output_3_0), .y(output_2_101));
wire output_1_102, output_1_1, output_0_102;
mixer gate_output_0_102(.a(output_1_102), .b(output_1_1), .y(output_0_102));
wire output_2_102, output_2_1, output_1_102;
mixer gate_output_1_102(.a(output_2_102), .b(output_2_1), .y(output_1_102));
wire output_3_102, output_3_1, output_2_102;
mixer gate_output_2_102(.a(output_3_102), .b(output_3_1), .y(output_2_102));
wire output_1_103, output_1_2, output_0_103;
mixer gate_output_0_103(.a(output_1_103), .b(output_1_2), .y(output_0_103));
wire output_2_103, output_2_2, output_1_103;
mixer gate_output_1_103(.a(output_2_103), .b(output_2_2), .y(output_1_103));
wire output_3_103, output_3_2, output_2_103;
mixer gate_output_2_103(.a(output_3_103), .b(output_3_2), .y(output_2_103));
wire output_1_104, output_1_0, output_0_104;
mixer gate_output_0_104(.a(output_1_104), .b(output_1_0), .y(output_0_104));
wire output_2_104, output_2_0, output_1_104;
mixer gate_output_1_104(.a(output_2_104), .b(output_2_0), .y(output_1_104));
wire output_3_104, output_3_0, output_2_104;
mixer gate_output_2_104(.a(output_3_104), .b(output_3_0), .y(output_2_104));
wire output_1_105, output_1_1, output_0_105;
mixer gate_output_0_105(.a(output_1_105), .b(output_1_1), .y(output_0_105));
wire output_2_105, output_2_1, output_1_105;
mixer gate_output_1_105(.a(output_2_105), .b(output_2_1), .y(output_1_105));
wire output_3_105, output_3_1, output_2_105;
mixer gate_output_2_105(.a(output_3_105), .b(output_3_1), .y(output_2_105));
wire output_1_106, output_1_2, output_0_106;
mixer gate_output_0_106(.a(output_1_106), .b(output_1_2), .y(output_0_106));
wire output_2_106, output_2_2, output_1_106;
mixer gate_output_1_106(.a(output_2_106), .b(output_2_2), .y(output_1_106));
wire output_3_106, output_3_2, output_2_106;
mixer gate_output_2_106(.a(output_3_106), .b(output_3_2), .y(output_2_106));
wire output_1_107, output_1_0, output_0_107;
mixer gate_output_0_107(.a(output_1_107), .b(output_1_0), .y(output_0_107));
wire output_2_107, output_2_0, output_1_107;
mixer gate_output_1_107(.a(output_2_107), .b(output_2_0), .y(output_1_107));
wire output_3_107, output_3_0, output_2_107;
mixer gate_output_2_107(.a(output_3_107), .b(output_3_0), .y(output_2_107));
wire output_1_108, output_1_1, output_0_108;
mixer gate_output_0_108(.a(output_1_108), .b(output_1_1), .y(output_0_108));
wire output_2_108, output_2_1, output_1_108;
mixer gate_output_1_108(.a(output_2_108), .b(output_2_1), .y(output_1_108));
wire output_3_108, output_3_1, output_2_108;
mixer gate_output_2_108(.a(output_3_108), .b(output_3_1), .y(output_2_108));
wire output_1_109, output_1_2, output_0_109;
mixer gate_output_0_109(.a(output_1_109), .b(output_1_2), .y(output_0_109));
wire output_2_109, output_2_2, output_1_109;
mixer gate_output_1_109(.a(output_2_109), .b(output_2_2), .y(output_1_109));
wire output_3_109, output_3_2, output_2_109;
mixer gate_output_2_109(.a(output_3_109), .b(output_3_2), .y(output_2_109));
wire output_1_110, output_1_0, output_0_110;
mixer gate_output_0_110(.a(output_1_110), .b(output_1_0), .y(output_0_110));
wire output_2_110, output_2_0, output_1_110;
mixer gate_output_1_110(.a(output_2_110), .b(output_2_0), .y(output_1_110));
wire output_3_110, output_3_0, output_2_110;
mixer gate_output_2_110(.a(output_3_110), .b(output_3_0), .y(output_2_110));
wire output_1_111, output_1_1, output_0_111;
mixer gate_output_0_111(.a(output_1_111), .b(output_1_1), .y(output_0_111));
wire output_2_111, output_2_1, output_1_111;
mixer gate_output_1_111(.a(output_2_111), .b(output_2_1), .y(output_1_111));
wire output_3_111, output_3_1, output_2_111;
mixer gate_output_2_111(.a(output_3_111), .b(output_3_1), .y(output_2_111));
wire output_1_112, output_1_2, output_0_112;
mixer gate_output_0_112(.a(output_1_112), .b(output_1_2), .y(output_0_112));
wire output_2_112, output_2_2, output_1_112;
mixer gate_output_1_112(.a(output_2_112), .b(output_2_2), .y(output_1_112));
wire output_3_112, output_3_2, output_2_112;
mixer gate_output_2_112(.a(output_3_112), .b(output_3_2), .y(output_2_112));
wire output_1_113, output_1_0, output_0_113;
mixer gate_output_0_113(.a(output_1_113), .b(output_1_0), .y(output_0_113));
wire output_2_113, output_2_0, output_1_113;
mixer gate_output_1_113(.a(output_2_113), .b(output_2_0), .y(output_1_113));
wire output_3_113, output_3_0, output_2_113;
mixer gate_output_2_113(.a(output_3_113), .b(output_3_0), .y(output_2_113));
wire output_1_114, output_1_1, output_0_114;
mixer gate_output_0_114(.a(output_1_114), .b(output_1_1), .y(output_0_114));
wire output_2_114, output_2_1, output_1_114;
mixer gate_output_1_114(.a(output_2_114), .b(output_2_1), .y(output_1_114));
wire output_3_114, output_3_1, output_2_114;
mixer gate_output_2_114(.a(output_3_114), .b(output_3_1), .y(output_2_114));
wire output_1_115, output_1_2, output_0_115;
mixer gate_output_0_115(.a(output_1_115), .b(output_1_2), .y(output_0_115));
wire output_2_115, output_2_2, output_1_115;
mixer gate_output_1_115(.a(output_2_115), .b(output_2_2), .y(output_1_115));
wire output_3_115, output_3_2, output_2_115;
mixer gate_output_2_115(.a(output_3_115), .b(output_3_2), .y(output_2_115));
wire output_1_116, output_1_0, output_0_116;
mixer gate_output_0_116(.a(output_1_116), .b(output_1_0), .y(output_0_116));
wire output_2_116, output_2_0, output_1_116;
mixer gate_output_1_116(.a(output_2_116), .b(output_2_0), .y(output_1_116));
wire output_3_116, output_3_0, output_2_116;
mixer gate_output_2_116(.a(output_3_116), .b(output_3_0), .y(output_2_116));
wire output_1_117, output_1_1, output_0_117;
mixer gate_output_0_117(.a(output_1_117), .b(output_1_1), .y(output_0_117));
wire output_2_117, output_2_1, output_1_117;
mixer gate_output_1_117(.a(output_2_117), .b(output_2_1), .y(output_1_117));
wire output_3_117, output_3_1, output_2_117;
mixer gate_output_2_117(.a(output_3_117), .b(output_3_1), .y(output_2_117));
wire output_1_118, output_1_2, output_0_118;
mixer gate_output_0_118(.a(output_1_118), .b(output_1_2), .y(output_0_118));
wire output_2_118, output_2_2, output_1_118;
mixer gate_output_1_118(.a(output_2_118), .b(output_2_2), .y(output_1_118));
wire output_3_118, output_3_2, output_2_118;
mixer gate_output_2_118(.a(output_3_118), .b(output_3_2), .y(output_2_118));
wire output_1_119, output_1_0, output_0_119;
mixer gate_output_0_119(.a(output_1_119), .b(output_1_0), .y(output_0_119));
wire output_2_119, output_2_0, output_1_119;
mixer gate_output_1_119(.a(output_2_119), .b(output_2_0), .y(output_1_119));
wire output_3_119, output_3_0, output_2_119;
mixer gate_output_2_119(.a(output_3_119), .b(output_3_0), .y(output_2_119));
wire output_1_120, output_1_1, output_0_120;
mixer gate_output_0_120(.a(output_1_120), .b(output_1_1), .y(output_0_120));
wire output_2_120, output_2_1, output_1_120;
mixer gate_output_1_120(.a(output_2_120), .b(output_2_1), .y(output_1_120));
wire output_3_120, output_3_1, output_2_120;
mixer gate_output_2_120(.a(output_3_120), .b(output_3_1), .y(output_2_120));
wire output_1_121, output_1_2, output_0_121;
mixer gate_output_0_121(.a(output_1_121), .b(output_1_2), .y(output_0_121));
wire output_2_121, output_2_2, output_1_121;
mixer gate_output_1_121(.a(output_2_121), .b(output_2_2), .y(output_1_121));
wire output_3_121, output_3_2, output_2_121;
mixer gate_output_2_121(.a(output_3_121), .b(output_3_2), .y(output_2_121));
wire output_1_122, output_1_0, output_0_122;
mixer gate_output_0_122(.a(output_1_122), .b(output_1_0), .y(output_0_122));
wire output_2_122, output_2_0, output_1_122;
mixer gate_output_1_122(.a(output_2_122), .b(output_2_0), .y(output_1_122));
wire output_3_122, output_3_0, output_2_122;
mixer gate_output_2_122(.a(output_3_122), .b(output_3_0), .y(output_2_122));
wire output_1_123, output_1_1, output_0_123;
mixer gate_output_0_123(.a(output_1_123), .b(output_1_1), .y(output_0_123));
wire output_2_123, output_2_1, output_1_123;
mixer gate_output_1_123(.a(output_2_123), .b(output_2_1), .y(output_1_123));
wire output_3_123, output_3_1, output_2_123;
mixer gate_output_2_123(.a(output_3_123), .b(output_3_1), .y(output_2_123));
wire output_1_124, output_1_2, output_0_124;
mixer gate_output_0_124(.a(output_1_124), .b(output_1_2), .y(output_0_124));
wire output_2_124, output_2_2, output_1_124;
mixer gate_output_1_124(.a(output_2_124), .b(output_2_2), .y(output_1_124));
wire output_3_124, output_3_2, output_2_124;
mixer gate_output_2_124(.a(output_3_124), .b(output_3_2), .y(output_2_124));
wire output_1_125, output_1_0, output_0_125;
mixer gate_output_0_125(.a(output_1_125), .b(output_1_0), .y(output_0_125));
wire output_2_125, output_2_0, output_1_125;
mixer gate_output_1_125(.a(output_2_125), .b(output_2_0), .y(output_1_125));
wire output_3_125, output_3_0, output_2_125;
mixer gate_output_2_125(.a(output_3_125), .b(output_3_0), .y(output_2_125));
wire output_1_126, output_1_1, output_0_126;
mixer gate_output_0_126(.a(output_1_126), .b(output_1_1), .y(output_0_126));
wire output_2_126, output_2_1, output_1_126;
mixer gate_output_1_126(.a(output_2_126), .b(output_2_1), .y(output_1_126));
wire output_3_126, output_3_1, output_2_126;
mixer gate_output_2_126(.a(output_3_126), .b(output_3_1), .y(output_2_126));
wire output_1_127, output_1_2, output_0_127;
mixer gate_output_0_127(.a(output_1_127), .b(output_1_2), .y(output_0_127));
wire output_2_127, output_2_2, output_1_127;
mixer gate_output_1_127(.a(output_2_127), .b(output_2_2), .y(output_1_127));
wire output_3_127, output_3_2, output_2_127;
mixer gate_output_2_127(.a(output_3_127), .b(output_3_2), .y(output_2_127));
wire output_1_128, output_1_0, output_0_128;
mixer gate_output_0_128(.a(output_1_128), .b(output_1_0), .y(output_0_128));
wire output_2_128, output_2_0, output_1_128;
mixer gate_output_1_128(.a(output_2_128), .b(output_2_0), .y(output_1_128));
wire output_3_128, output_3_0, output_2_128;
mixer gate_output_2_128(.a(output_3_128), .b(output_3_0), .y(output_2_128));
wire output_1_129, output_1_1, output_0_129;
mixer gate_output_0_129(.a(output_1_129), .b(output_1_1), .y(output_0_129));
wire output_2_129, output_2_1, output_1_129;
mixer gate_output_1_129(.a(output_2_129), .b(output_2_1), .y(output_1_129));
wire output_3_129, output_3_1, output_2_129;
mixer gate_output_2_129(.a(output_3_129), .b(output_3_1), .y(output_2_129));
wire output_1_130, output_1_2, output_0_130;
mixer gate_output_0_130(.a(output_1_130), .b(output_1_2), .y(output_0_130));
wire output_2_130, output_2_2, output_1_130;
mixer gate_output_1_130(.a(output_2_130), .b(output_2_2), .y(output_1_130));
wire output_3_130, output_3_2, output_2_130;
mixer gate_output_2_130(.a(output_3_130), .b(output_3_2), .y(output_2_130));
wire output_1_131, output_1_0, output_0_131;
mixer gate_output_0_131(.a(output_1_131), .b(output_1_0), .y(output_0_131));
wire output_2_131, output_2_0, output_1_131;
mixer gate_output_1_131(.a(output_2_131), .b(output_2_0), .y(output_1_131));
wire output_3_131, output_3_0, output_2_131;
mixer gate_output_2_131(.a(output_3_131), .b(output_3_0), .y(output_2_131));
wire output_1_132, output_1_1, output_0_132;
mixer gate_output_0_132(.a(output_1_132), .b(output_1_1), .y(output_0_132));
wire output_2_132, output_2_1, output_1_132;
mixer gate_output_1_132(.a(output_2_132), .b(output_2_1), .y(output_1_132));
wire output_3_132, output_3_1, output_2_132;
mixer gate_output_2_132(.a(output_3_132), .b(output_3_1), .y(output_2_132));
wire output_1_133, output_1_2, output_0_133;
mixer gate_output_0_133(.a(output_1_133), .b(output_1_2), .y(output_0_133));
wire output_2_133, output_2_2, output_1_133;
mixer gate_output_1_133(.a(output_2_133), .b(output_2_2), .y(output_1_133));
wire output_3_133, output_3_2, output_2_133;
mixer gate_output_2_133(.a(output_3_133), .b(output_3_2), .y(output_2_133));
wire output_1_134, output_1_0, output_0_134;
mixer gate_output_0_134(.a(output_1_134), .b(output_1_0), .y(output_0_134));
wire output_2_134, output_2_0, output_1_134;
mixer gate_output_1_134(.a(output_2_134), .b(output_2_0), .y(output_1_134));
wire output_3_134, output_3_0, output_2_134;
mixer gate_output_2_134(.a(output_3_134), .b(output_3_0), .y(output_2_134));
wire output_1_135, output_1_1, output_0_135;
mixer gate_output_0_135(.a(output_1_135), .b(output_1_1), .y(output_0_135));
wire output_2_135, output_2_1, output_1_135;
mixer gate_output_1_135(.a(output_2_135), .b(output_2_1), .y(output_1_135));
wire output_3_135, output_3_1, output_2_135;
mixer gate_output_2_135(.a(output_3_135), .b(output_3_1), .y(output_2_135));
wire output_1_136, output_1_2, output_0_136;
mixer gate_output_0_136(.a(output_1_136), .b(output_1_2), .y(output_0_136));
wire output_2_136, output_2_2, output_1_136;
mixer gate_output_1_136(.a(output_2_136), .b(output_2_2), .y(output_1_136));
wire output_3_136, output_3_2, output_2_136;
mixer gate_output_2_136(.a(output_3_136), .b(output_3_2), .y(output_2_136));
wire output_1_137, output_1_0, output_0_137;
mixer gate_output_0_137(.a(output_1_137), .b(output_1_0), .y(output_0_137));
wire output_2_137, output_2_0, output_1_137;
mixer gate_output_1_137(.a(output_2_137), .b(output_2_0), .y(output_1_137));
wire output_3_137, output_3_0, output_2_137;
mixer gate_output_2_137(.a(output_3_137), .b(output_3_0), .y(output_2_137));
wire output_1_138, output_1_1, output_0_138;
mixer gate_output_0_138(.a(output_1_138), .b(output_1_1), .y(output_0_138));
wire output_2_138, output_2_1, output_1_138;
mixer gate_output_1_138(.a(output_2_138), .b(output_2_1), .y(output_1_138));
wire output_3_138, output_3_1, output_2_138;
mixer gate_output_2_138(.a(output_3_138), .b(output_3_1), .y(output_2_138));
wire output_1_139, output_1_2, output_0_139;
mixer gate_output_0_139(.a(output_1_139), .b(output_1_2), .y(output_0_139));
wire output_2_139, output_2_2, output_1_139;
mixer gate_output_1_139(.a(output_2_139), .b(output_2_2), .y(output_1_139));
wire output_3_139, output_3_2, output_2_139;
mixer gate_output_2_139(.a(output_3_139), .b(output_3_2), .y(output_2_139));
wire output_1_140, output_1_0, output_0_140;
mixer gate_output_0_140(.a(output_1_140), .b(output_1_0), .y(output_0_140));
wire output_2_140, output_2_0, output_1_140;
mixer gate_output_1_140(.a(output_2_140), .b(output_2_0), .y(output_1_140));
wire output_3_140, output_3_0, output_2_140;
mixer gate_output_2_140(.a(output_3_140), .b(output_3_0), .y(output_2_140));
wire output_1_141, output_1_1, output_0_141;
mixer gate_output_0_141(.a(output_1_141), .b(output_1_1), .y(output_0_141));
wire output_2_141, output_2_1, output_1_141;
mixer gate_output_1_141(.a(output_2_141), .b(output_2_1), .y(output_1_141));
wire output_3_141, output_3_1, output_2_141;
mixer gate_output_2_141(.a(output_3_141), .b(output_3_1), .y(output_2_141));
wire output_1_142, output_1_2, output_0_142;
mixer gate_output_0_142(.a(output_1_142), .b(output_1_2), .y(output_0_142));
wire output_2_142, output_2_2, output_1_142;
mixer gate_output_1_142(.a(output_2_142), .b(output_2_2), .y(output_1_142));
wire output_3_142, output_3_2, output_2_142;
mixer gate_output_2_142(.a(output_3_142), .b(output_3_2), .y(output_2_142));
wire output_1_143, output_1_0, output_0_143;
mixer gate_output_0_143(.a(output_1_143), .b(output_1_0), .y(output_0_143));
wire output_2_143, output_2_0, output_1_143;
mixer gate_output_1_143(.a(output_2_143), .b(output_2_0), .y(output_1_143));
wire output_3_143, output_3_0, output_2_143;
mixer gate_output_2_143(.a(output_3_143), .b(output_3_0), .y(output_2_143));
wire output_1_144, output_1_1, output_0_144;
mixer gate_output_0_144(.a(output_1_144), .b(output_1_1), .y(output_0_144));
wire output_2_144, output_2_1, output_1_144;
mixer gate_output_1_144(.a(output_2_144), .b(output_2_1), .y(output_1_144));
wire output_3_144, output_3_1, output_2_144;
mixer gate_output_2_144(.a(output_3_144), .b(output_3_1), .y(output_2_144));
wire output_1_145, output_1_2, output_0_145;
mixer gate_output_0_145(.a(output_1_145), .b(output_1_2), .y(output_0_145));
wire output_2_145, output_2_2, output_1_145;
mixer gate_output_1_145(.a(output_2_145), .b(output_2_2), .y(output_1_145));
wire output_3_145, output_3_2, output_2_145;
mixer gate_output_2_145(.a(output_3_145), .b(output_3_2), .y(output_2_145));
wire output_1_146, output_1_0, output_0_146;
mixer gate_output_0_146(.a(output_1_146), .b(output_1_0), .y(output_0_146));
wire output_2_146, output_2_0, output_1_146;
mixer gate_output_1_146(.a(output_2_146), .b(output_2_0), .y(output_1_146));
wire output_3_146, output_3_0, output_2_146;
mixer gate_output_2_146(.a(output_3_146), .b(output_3_0), .y(output_2_146));
wire output_1_147, output_1_1, output_0_147;
mixer gate_output_0_147(.a(output_1_147), .b(output_1_1), .y(output_0_147));
wire output_2_147, output_2_1, output_1_147;
mixer gate_output_1_147(.a(output_2_147), .b(output_2_1), .y(output_1_147));
wire output_3_147, output_3_1, output_2_147;
mixer gate_output_2_147(.a(output_3_147), .b(output_3_1), .y(output_2_147));
wire output_1_148, output_1_2, output_0_148;
mixer gate_output_0_148(.a(output_1_148), .b(output_1_2), .y(output_0_148));
wire output_2_148, output_2_2, output_1_148;
mixer gate_output_1_148(.a(output_2_148), .b(output_2_2), .y(output_1_148));
wire output_3_148, output_3_2, output_2_148;
mixer gate_output_2_148(.a(output_3_148), .b(output_3_2), .y(output_2_148));
wire output_1_149, output_1_0, output_0_149;
mixer gate_output_0_149(.a(output_1_149), .b(output_1_0), .y(output_0_149));
wire output_2_149, output_2_0, output_1_149;
mixer gate_output_1_149(.a(output_2_149), .b(output_2_0), .y(output_1_149));
wire output_3_149, output_3_0, output_2_149;
mixer gate_output_2_149(.a(output_3_149), .b(output_3_0), .y(output_2_149));
wire output_1_150, output_1_1, output_0_150;
mixer gate_output_0_150(.a(output_1_150), .b(output_1_1), .y(output_0_150));
wire output_2_150, output_2_1, output_1_150;
mixer gate_output_1_150(.a(output_2_150), .b(output_2_1), .y(output_1_150));
wire output_3_150, output_3_1, output_2_150;
mixer gate_output_2_150(.a(output_3_150), .b(output_3_1), .y(output_2_150));
wire output_1_151, output_1_2, output_0_151;
mixer gate_output_0_151(.a(output_1_151), .b(output_1_2), .y(output_0_151));
wire output_2_151, output_2_2, output_1_151;
mixer gate_output_1_151(.a(output_2_151), .b(output_2_2), .y(output_1_151));
wire output_3_151, output_3_2, output_2_151;
mixer gate_output_2_151(.a(output_3_151), .b(output_3_2), .y(output_2_151));
wire output_1_152, output_1_0, output_0_152;
mixer gate_output_0_152(.a(output_1_152), .b(output_1_0), .y(output_0_152));
wire output_2_152, output_2_0, output_1_152;
mixer gate_output_1_152(.a(output_2_152), .b(output_2_0), .y(output_1_152));
wire output_3_152, output_3_0, output_2_152;
mixer gate_output_2_152(.a(output_3_152), .b(output_3_0), .y(output_2_152));
wire output_1_153, output_1_1, output_0_153;
mixer gate_output_0_153(.a(output_1_153), .b(output_1_1), .y(output_0_153));
wire output_2_153, output_2_1, output_1_153;
mixer gate_output_1_153(.a(output_2_153), .b(output_2_1), .y(output_1_153));
wire output_3_153, output_3_1, output_2_153;
mixer gate_output_2_153(.a(output_3_153), .b(output_3_1), .y(output_2_153));
wire output_1_154, output_1_2, output_0_154;
mixer gate_output_0_154(.a(output_1_154), .b(output_1_2), .y(output_0_154));
wire output_2_154, output_2_2, output_1_154;
mixer gate_output_1_154(.a(output_2_154), .b(output_2_2), .y(output_1_154));
wire output_3_154, output_3_2, output_2_154;
mixer gate_output_2_154(.a(output_3_154), .b(output_3_2), .y(output_2_154));
wire output_1_155, output_1_0, output_0_155;
mixer gate_output_0_155(.a(output_1_155), .b(output_1_0), .y(output_0_155));
wire output_2_155, output_2_0, output_1_155;
mixer gate_output_1_155(.a(output_2_155), .b(output_2_0), .y(output_1_155));
wire output_3_155, output_3_0, output_2_155;
mixer gate_output_2_155(.a(output_3_155), .b(output_3_0), .y(output_2_155));
wire output_1_156, output_1_1, output_0_156;
mixer gate_output_0_156(.a(output_1_156), .b(output_1_1), .y(output_0_156));
wire output_2_156, output_2_1, output_1_156;
mixer gate_output_1_156(.a(output_2_156), .b(output_2_1), .y(output_1_156));
wire output_3_156, output_3_1, output_2_156;
mixer gate_output_2_156(.a(output_3_156), .b(output_3_1), .y(output_2_156));
wire output_1_157, output_1_2, output_0_157;
mixer gate_output_0_157(.a(output_1_157), .b(output_1_2), .y(output_0_157));
wire output_2_157, output_2_2, output_1_157;
mixer gate_output_1_157(.a(output_2_157), .b(output_2_2), .y(output_1_157));
wire output_3_157, output_3_2, output_2_157;
mixer gate_output_2_157(.a(output_3_157), .b(output_3_2), .y(output_2_157));
wire output_1_158, output_1_0, output_0_158;
mixer gate_output_0_158(.a(output_1_158), .b(output_1_0), .y(output_0_158));
wire output_2_158, output_2_0, output_1_158;
mixer gate_output_1_158(.a(output_2_158), .b(output_2_0), .y(output_1_158));
wire output_3_158, output_3_0, output_2_158;
mixer gate_output_2_158(.a(output_3_158), .b(output_3_0), .y(output_2_158));
wire output_1_159, output_1_1, output_0_159;
mixer gate_output_0_159(.a(output_1_159), .b(output_1_1), .y(output_0_159));
wire output_2_159, output_2_1, output_1_159;
mixer gate_output_1_159(.a(output_2_159), .b(output_2_1), .y(output_1_159));
wire output_3_159, output_3_1, output_2_159;
mixer gate_output_2_159(.a(output_3_159), .b(output_3_1), .y(output_2_159));
wire output_1_160, output_1_2, output_0_160;
mixer gate_output_0_160(.a(output_1_160), .b(output_1_2), .y(output_0_160));
wire output_2_160, output_2_2, output_1_160;
mixer gate_output_1_160(.a(output_2_160), .b(output_2_2), .y(output_1_160));
wire output_3_160, output_3_2, output_2_160;
mixer gate_output_2_160(.a(output_3_160), .b(output_3_2), .y(output_2_160));
wire output_1_161, output_1_0, output_0_161;
mixer gate_output_0_161(.a(output_1_161), .b(output_1_0), .y(output_0_161));
wire output_2_161, output_2_0, output_1_161;
mixer gate_output_1_161(.a(output_2_161), .b(output_2_0), .y(output_1_161));
wire output_3_161, output_3_0, output_2_161;
mixer gate_output_2_161(.a(output_3_161), .b(output_3_0), .y(output_2_161));
wire output_1_162, output_1_1, output_0_162;
mixer gate_output_0_162(.a(output_1_162), .b(output_1_1), .y(output_0_162));
wire output_2_162, output_2_1, output_1_162;
mixer gate_output_1_162(.a(output_2_162), .b(output_2_1), .y(output_1_162));
wire output_3_162, output_3_1, output_2_162;
mixer gate_output_2_162(.a(output_3_162), .b(output_3_1), .y(output_2_162));
wire output_1_163, output_1_2, output_0_163;
mixer gate_output_0_163(.a(output_1_163), .b(output_1_2), .y(output_0_163));
wire output_2_163, output_2_2, output_1_163;
mixer gate_output_1_163(.a(output_2_163), .b(output_2_2), .y(output_1_163));
wire output_3_163, output_3_2, output_2_163;
mixer gate_output_2_163(.a(output_3_163), .b(output_3_2), .y(output_2_163));
wire output_1_164, output_1_0, output_0_164;
mixer gate_output_0_164(.a(output_1_164), .b(output_1_0), .y(output_0_164));
wire output_2_164, output_2_0, output_1_164;
mixer gate_output_1_164(.a(output_2_164), .b(output_2_0), .y(output_1_164));
wire output_3_164, output_3_0, output_2_164;
mixer gate_output_2_164(.a(output_3_164), .b(output_3_0), .y(output_2_164));
wire output_1_165, output_1_1, output_0_165;
mixer gate_output_0_165(.a(output_1_165), .b(output_1_1), .y(output_0_165));
wire output_2_165, output_2_1, output_1_165;
mixer gate_output_1_165(.a(output_2_165), .b(output_2_1), .y(output_1_165));
wire output_3_165, output_3_1, output_2_165;
mixer gate_output_2_165(.a(output_3_165), .b(output_3_1), .y(output_2_165));
wire output_1_166, output_1_2, output_0_166;
mixer gate_output_0_166(.a(output_1_166), .b(output_1_2), .y(output_0_166));
wire output_2_166, output_2_2, output_1_166;
mixer gate_output_1_166(.a(output_2_166), .b(output_2_2), .y(output_1_166));
wire output_3_166, output_3_2, output_2_166;
mixer gate_output_2_166(.a(output_3_166), .b(output_3_2), .y(output_2_166));
wire output_1_167, output_1_0, output_0_167;
mixer gate_output_0_167(.a(output_1_167), .b(output_1_0), .y(output_0_167));
wire output_2_167, output_2_0, output_1_167;
mixer gate_output_1_167(.a(output_2_167), .b(output_2_0), .y(output_1_167));
wire output_3_167, output_3_0, output_2_167;
mixer gate_output_2_167(.a(output_3_167), .b(output_3_0), .y(output_2_167));
wire output_1_168, output_1_1, output_0_168;
mixer gate_output_0_168(.a(output_1_168), .b(output_1_1), .y(output_0_168));
wire output_2_168, output_2_1, output_1_168;
mixer gate_output_1_168(.a(output_2_168), .b(output_2_1), .y(output_1_168));
wire output_3_168, output_3_1, output_2_168;
mixer gate_output_2_168(.a(output_3_168), .b(output_3_1), .y(output_2_168));
wire output_1_169, output_1_2, output_0_169;
mixer gate_output_0_169(.a(output_1_169), .b(output_1_2), .y(output_0_169));
wire output_2_169, output_2_2, output_1_169;
mixer gate_output_1_169(.a(output_2_169), .b(output_2_2), .y(output_1_169));
wire output_3_169, output_3_2, output_2_169;
mixer gate_output_2_169(.a(output_3_169), .b(output_3_2), .y(output_2_169));
wire output_1_170, output_1_0, output_0_170;
mixer gate_output_0_170(.a(output_1_170), .b(output_1_0), .y(output_0_170));
wire output_2_170, output_2_0, output_1_170;
mixer gate_output_1_170(.a(output_2_170), .b(output_2_0), .y(output_1_170));
wire output_3_170, output_3_0, output_2_170;
mixer gate_output_2_170(.a(output_3_170), .b(output_3_0), .y(output_2_170));
wire output_1_171, output_1_1, output_0_171;
mixer gate_output_0_171(.a(output_1_171), .b(output_1_1), .y(output_0_171));
wire output_2_171, output_2_1, output_1_171;
mixer gate_output_1_171(.a(output_2_171), .b(output_2_1), .y(output_1_171));
wire output_3_171, output_3_1, output_2_171;
mixer gate_output_2_171(.a(output_3_171), .b(output_3_1), .y(output_2_171));
wire output_1_172, output_1_2, output_0_172;
mixer gate_output_0_172(.a(output_1_172), .b(output_1_2), .y(output_0_172));
wire output_2_172, output_2_2, output_1_172;
mixer gate_output_1_172(.a(output_2_172), .b(output_2_2), .y(output_1_172));
wire output_3_172, output_3_2, output_2_172;
mixer gate_output_2_172(.a(output_3_172), .b(output_3_2), .y(output_2_172));
wire output_1_173, output_1_0, output_0_173;
mixer gate_output_0_173(.a(output_1_173), .b(output_1_0), .y(output_0_173));
wire output_2_173, output_2_0, output_1_173;
mixer gate_output_1_173(.a(output_2_173), .b(output_2_0), .y(output_1_173));
wire output_3_173, output_3_0, output_2_173;
mixer gate_output_2_173(.a(output_3_173), .b(output_3_0), .y(output_2_173));
wire output_1_174, output_1_1, output_0_174;
mixer gate_output_0_174(.a(output_1_174), .b(output_1_1), .y(output_0_174));
wire output_2_174, output_2_1, output_1_174;
mixer gate_output_1_174(.a(output_2_174), .b(output_2_1), .y(output_1_174));
wire output_3_174, output_3_1, output_2_174;
mixer gate_output_2_174(.a(output_3_174), .b(output_3_1), .y(output_2_174));
wire output_1_175, output_1_2, output_0_175;
mixer gate_output_0_175(.a(output_1_175), .b(output_1_2), .y(output_0_175));
wire output_2_175, output_2_2, output_1_175;
mixer gate_output_1_175(.a(output_2_175), .b(output_2_2), .y(output_1_175));
wire output_3_175, output_3_2, output_2_175;
mixer gate_output_2_175(.a(output_3_175), .b(output_3_2), .y(output_2_175));
wire output_1_176, output_1_0, output_0_176;
mixer gate_output_0_176(.a(output_1_176), .b(output_1_0), .y(output_0_176));
wire output_2_176, output_2_0, output_1_176;
mixer gate_output_1_176(.a(output_2_176), .b(output_2_0), .y(output_1_176));
wire output_3_176, output_3_0, output_2_176;
mixer gate_output_2_176(.a(output_3_176), .b(output_3_0), .y(output_2_176));
wire output_1_177, output_1_1, output_0_177;
mixer gate_output_0_177(.a(output_1_177), .b(output_1_1), .y(output_0_177));
wire output_2_177, output_2_1, output_1_177;
mixer gate_output_1_177(.a(output_2_177), .b(output_2_1), .y(output_1_177));
wire output_3_177, output_3_1, output_2_177;
mixer gate_output_2_177(.a(output_3_177), .b(output_3_1), .y(output_2_177));
wire output_1_178, output_1_2, output_0_178;
mixer gate_output_0_178(.a(output_1_178), .b(output_1_2), .y(output_0_178));
wire output_2_178, output_2_2, output_1_178;
mixer gate_output_1_178(.a(output_2_178), .b(output_2_2), .y(output_1_178));
wire output_3_178, output_3_2, output_2_178;
mixer gate_output_2_178(.a(output_3_178), .b(output_3_2), .y(output_2_178));
wire output_1_179, output_1_0, output_0_179;
mixer gate_output_0_179(.a(output_1_179), .b(output_1_0), .y(output_0_179));
wire output_2_179, output_2_0, output_1_179;
mixer gate_output_1_179(.a(output_2_179), .b(output_2_0), .y(output_1_179));
wire output_3_179, output_3_0, output_2_179;
mixer gate_output_2_179(.a(output_3_179), .b(output_3_0), .y(output_2_179));
wire output_1_180, output_1_1, output_0_180;
mixer gate_output_0_180(.a(output_1_180), .b(output_1_1), .y(output_0_180));
wire output_2_180, output_2_1, output_1_180;
mixer gate_output_1_180(.a(output_2_180), .b(output_2_1), .y(output_1_180));
wire output_3_180, output_3_1, output_2_180;
mixer gate_output_2_180(.a(output_3_180), .b(output_3_1), .y(output_2_180));
wire output_1_181, output_1_2, output_0_181;
mixer gate_output_0_181(.a(output_1_181), .b(output_1_2), .y(output_0_181));
wire output_2_181, output_2_2, output_1_181;
mixer gate_output_1_181(.a(output_2_181), .b(output_2_2), .y(output_1_181));
wire output_3_181, output_3_2, output_2_181;
mixer gate_output_2_181(.a(output_3_181), .b(output_3_2), .y(output_2_181));
wire output_1_182, output_1_0, output_0_182;
mixer gate_output_0_182(.a(output_1_182), .b(output_1_0), .y(output_0_182));
wire output_2_182, output_2_0, output_1_182;
mixer gate_output_1_182(.a(output_2_182), .b(output_2_0), .y(output_1_182));
wire output_3_182, output_3_0, output_2_182;
mixer gate_output_2_182(.a(output_3_182), .b(output_3_0), .y(output_2_182));
wire output_1_183, output_1_1, output_0_183;
mixer gate_output_0_183(.a(output_1_183), .b(output_1_1), .y(output_0_183));
wire output_2_183, output_2_1, output_1_183;
mixer gate_output_1_183(.a(output_2_183), .b(output_2_1), .y(output_1_183));
wire output_3_183, output_3_1, output_2_183;
mixer gate_output_2_183(.a(output_3_183), .b(output_3_1), .y(output_2_183));
wire output_1_184, output_1_2, output_0_184;
mixer gate_output_0_184(.a(output_1_184), .b(output_1_2), .y(output_0_184));
wire output_2_184, output_2_2, output_1_184;
mixer gate_output_1_184(.a(output_2_184), .b(output_2_2), .y(output_1_184));
wire output_3_184, output_3_2, output_2_184;
mixer gate_output_2_184(.a(output_3_184), .b(output_3_2), .y(output_2_184));
wire output_1_185, output_1_0, output_0_185;
mixer gate_output_0_185(.a(output_1_185), .b(output_1_0), .y(output_0_185));
wire output_2_185, output_2_0, output_1_185;
mixer gate_output_1_185(.a(output_2_185), .b(output_2_0), .y(output_1_185));
wire output_3_185, output_3_0, output_2_185;
mixer gate_output_2_185(.a(output_3_185), .b(output_3_0), .y(output_2_185));
wire output_1_186, output_1_1, output_0_186;
mixer gate_output_0_186(.a(output_1_186), .b(output_1_1), .y(output_0_186));
wire output_2_186, output_2_1, output_1_186;
mixer gate_output_1_186(.a(output_2_186), .b(output_2_1), .y(output_1_186));
wire output_3_186, output_3_1, output_2_186;
mixer gate_output_2_186(.a(output_3_186), .b(output_3_1), .y(output_2_186));
wire output_1_187, output_1_2, output_0_187;
mixer gate_output_0_187(.a(output_1_187), .b(output_1_2), .y(output_0_187));
wire output_2_187, output_2_2, output_1_187;
mixer gate_output_1_187(.a(output_2_187), .b(output_2_2), .y(output_1_187));
wire output_3_187, output_3_2, output_2_187;
mixer gate_output_2_187(.a(output_3_187), .b(output_3_2), .y(output_2_187));
wire output_1_188, output_1_0, output_0_188;
mixer gate_output_0_188(.a(output_1_188), .b(output_1_0), .y(output_0_188));
wire output_2_188, output_2_0, output_1_188;
mixer gate_output_1_188(.a(output_2_188), .b(output_2_0), .y(output_1_188));
wire output_3_188, output_3_0, output_2_188;
mixer gate_output_2_188(.a(output_3_188), .b(output_3_0), .y(output_2_188));
wire output_1_189, output_1_1, output_0_189;
mixer gate_output_0_189(.a(output_1_189), .b(output_1_1), .y(output_0_189));
wire output_2_189, output_2_1, output_1_189;
mixer gate_output_1_189(.a(output_2_189), .b(output_2_1), .y(output_1_189));
wire output_3_189, output_3_1, output_2_189;
mixer gate_output_2_189(.a(output_3_189), .b(output_3_1), .y(output_2_189));
wire output_1_190, output_1_2, output_0_190;
mixer gate_output_0_190(.a(output_1_190), .b(output_1_2), .y(output_0_190));
wire output_2_190, output_2_2, output_1_190;
mixer gate_output_1_190(.a(output_2_190), .b(output_2_2), .y(output_1_190));
wire output_3_190, output_3_2, output_2_190;
mixer gate_output_2_190(.a(output_3_190), .b(output_3_2), .y(output_2_190));
wire output_1_191, output_1_0, output_0_191;
mixer gate_output_0_191(.a(output_1_191), .b(output_1_0), .y(output_0_191));
wire output_2_191, output_2_0, output_1_191;
mixer gate_output_1_191(.a(output_2_191), .b(output_2_0), .y(output_1_191));
wire output_3_191, output_3_0, output_2_191;
mixer gate_output_2_191(.a(output_3_191), .b(output_3_0), .y(output_2_191));
wire output_1_192, output_1_1, output_0_192;
mixer gate_output_0_192(.a(output_1_192), .b(output_1_1), .y(output_0_192));
wire output_2_192, output_2_1, output_1_192;
mixer gate_output_1_192(.a(output_2_192), .b(output_2_1), .y(output_1_192));
wire output_3_192, output_3_1, output_2_192;
mixer gate_output_2_192(.a(output_3_192), .b(output_3_1), .y(output_2_192));
wire output_1_193, output_1_2, output_0_193;
mixer gate_output_0_193(.a(output_1_193), .b(output_1_2), .y(output_0_193));
wire output_2_193, output_2_2, output_1_193;
mixer gate_output_1_193(.a(output_2_193), .b(output_2_2), .y(output_1_193));
wire output_3_193, output_3_2, output_2_193;
mixer gate_output_2_193(.a(output_3_193), .b(output_3_2), .y(output_2_193));
wire output_1_194, output_1_0, output_0_194;
mixer gate_output_0_194(.a(output_1_194), .b(output_1_0), .y(output_0_194));
wire output_2_194, output_2_0, output_1_194;
mixer gate_output_1_194(.a(output_2_194), .b(output_2_0), .y(output_1_194));
wire output_3_194, output_3_0, output_2_194;
mixer gate_output_2_194(.a(output_3_194), .b(output_3_0), .y(output_2_194));
wire output_1_195, output_1_1, output_0_195;
mixer gate_output_0_195(.a(output_1_195), .b(output_1_1), .y(output_0_195));
wire output_2_195, output_2_1, output_1_195;
mixer gate_output_1_195(.a(output_2_195), .b(output_2_1), .y(output_1_195));
wire output_3_195, output_3_1, output_2_195;
mixer gate_output_2_195(.a(output_3_195), .b(output_3_1), .y(output_2_195));
wire output_1_196, output_1_2, output_0_196;
mixer gate_output_0_196(.a(output_1_196), .b(output_1_2), .y(output_0_196));
wire output_2_196, output_2_2, output_1_196;
mixer gate_output_1_196(.a(output_2_196), .b(output_2_2), .y(output_1_196));
wire output_3_196, output_3_2, output_2_196;
mixer gate_output_2_196(.a(output_3_196), .b(output_3_2), .y(output_2_196));
wire output_1_197, output_1_0, output_0_197;
mixer gate_output_0_197(.a(output_1_197), .b(output_1_0), .y(output_0_197));
wire output_2_197, output_2_0, output_1_197;
mixer gate_output_1_197(.a(output_2_197), .b(output_2_0), .y(output_1_197));
wire output_3_197, output_3_0, output_2_197;
mixer gate_output_2_197(.a(output_3_197), .b(output_3_0), .y(output_2_197));
wire output_1_198, output_1_1, output_0_198;
mixer gate_output_0_198(.a(output_1_198), .b(output_1_1), .y(output_0_198));
wire output_2_198, output_2_1, output_1_198;
mixer gate_output_1_198(.a(output_2_198), .b(output_2_1), .y(output_1_198));
wire output_3_198, output_3_1, output_2_198;
mixer gate_output_2_198(.a(output_3_198), .b(output_3_1), .y(output_2_198));
wire output_1_199, output_1_2, output_0_199;
mixer gate_output_0_199(.a(output_1_199), .b(output_1_2), .y(output_0_199));
wire output_2_199, output_2_2, output_1_199;
mixer gate_output_1_199(.a(output_2_199), .b(output_2_2), .y(output_1_199));
wire output_3_199, output_3_2, output_2_199;
mixer gate_output_2_199(.a(output_3_199), .b(output_3_2), .y(output_2_199));
wire output_1_200, output_1_0, output_0_200;
mixer gate_output_0_200(.a(output_1_200), .b(output_1_0), .y(output_0_200));
wire output_2_200, output_2_0, output_1_200;
mixer gate_output_1_200(.a(output_2_200), .b(output_2_0), .y(output_1_200));
wire output_3_200, output_3_0, output_2_200;
mixer gate_output_2_200(.a(output_3_200), .b(output_3_0), .y(output_2_200));
wire output_1_201, output_1_1, output_0_201;
mixer gate_output_0_201(.a(output_1_201), .b(output_1_1), .y(output_0_201));
wire output_2_201, output_2_1, output_1_201;
mixer gate_output_1_201(.a(output_2_201), .b(output_2_1), .y(output_1_201));
wire output_3_201, output_3_1, output_2_201;
mixer gate_output_2_201(.a(output_3_201), .b(output_3_1), .y(output_2_201));
wire output_1_202, output_1_2, output_0_202;
mixer gate_output_0_202(.a(output_1_202), .b(output_1_2), .y(output_0_202));
wire output_2_202, output_2_2, output_1_202;
mixer gate_output_1_202(.a(output_2_202), .b(output_2_2), .y(output_1_202));
wire output_3_202, output_3_2, output_2_202;
mixer gate_output_2_202(.a(output_3_202), .b(output_3_2), .y(output_2_202));
wire output_1_203, output_1_0, output_0_203;
mixer gate_output_0_203(.a(output_1_203), .b(output_1_0), .y(output_0_203));
wire output_2_203, output_2_0, output_1_203;
mixer gate_output_1_203(.a(output_2_203), .b(output_2_0), .y(output_1_203));
wire output_3_203, output_3_0, output_2_203;
mixer gate_output_2_203(.a(output_3_203), .b(output_3_0), .y(output_2_203));
wire output_1_204, output_1_1, output_0_204;
mixer gate_output_0_204(.a(output_1_204), .b(output_1_1), .y(output_0_204));
wire output_2_204, output_2_1, output_1_204;
mixer gate_output_1_204(.a(output_2_204), .b(output_2_1), .y(output_1_204));
wire output_3_204, output_3_1, output_2_204;
mixer gate_output_2_204(.a(output_3_204), .b(output_3_1), .y(output_2_204));
wire output_1_205, output_1_2, output_0_205;
mixer gate_output_0_205(.a(output_1_205), .b(output_1_2), .y(output_0_205));
wire output_2_205, output_2_2, output_1_205;
mixer gate_output_1_205(.a(output_2_205), .b(output_2_2), .y(output_1_205));
wire output_3_205, output_3_2, output_2_205;
mixer gate_output_2_205(.a(output_3_205), .b(output_3_2), .y(output_2_205));
wire output_1_206, output_1_0, output_0_206;
mixer gate_output_0_206(.a(output_1_206), .b(output_1_0), .y(output_0_206));
wire output_2_206, output_2_0, output_1_206;
mixer gate_output_1_206(.a(output_2_206), .b(output_2_0), .y(output_1_206));
wire output_3_206, output_3_0, output_2_206;
mixer gate_output_2_206(.a(output_3_206), .b(output_3_0), .y(output_2_206));
wire output_1_207, output_1_1, output_0_207;
mixer gate_output_0_207(.a(output_1_207), .b(output_1_1), .y(output_0_207));
wire output_2_207, output_2_1, output_1_207;
mixer gate_output_1_207(.a(output_2_207), .b(output_2_1), .y(output_1_207));
wire output_3_207, output_3_1, output_2_207;
mixer gate_output_2_207(.a(output_3_207), .b(output_3_1), .y(output_2_207));
wire output_1_208, output_1_2, output_0_208;
mixer gate_output_0_208(.a(output_1_208), .b(output_1_2), .y(output_0_208));
wire output_2_208, output_2_2, output_1_208;
mixer gate_output_1_208(.a(output_2_208), .b(output_2_2), .y(output_1_208));
wire output_3_208, output_3_2, output_2_208;
mixer gate_output_2_208(.a(output_3_208), .b(output_3_2), .y(output_2_208));
wire output_1_209, output_1_0, output_0_209;
mixer gate_output_0_209(.a(output_1_209), .b(output_1_0), .y(output_0_209));
wire output_2_209, output_2_0, output_1_209;
mixer gate_output_1_209(.a(output_2_209), .b(output_2_0), .y(output_1_209));
wire output_3_209, output_3_0, output_2_209;
mixer gate_output_2_209(.a(output_3_209), .b(output_3_0), .y(output_2_209));
wire output_1_210, output_1_1, output_0_210;
mixer gate_output_0_210(.a(output_1_210), .b(output_1_1), .y(output_0_210));
wire output_2_210, output_2_1, output_1_210;
mixer gate_output_1_210(.a(output_2_210), .b(output_2_1), .y(output_1_210));
wire output_3_210, output_3_1, output_2_210;
mixer gate_output_2_210(.a(output_3_210), .b(output_3_1), .y(output_2_210));
wire output_1_211, output_1_2, output_0_211;
mixer gate_output_0_211(.a(output_1_211), .b(output_1_2), .y(output_0_211));
wire output_2_211, output_2_2, output_1_211;
mixer gate_output_1_211(.a(output_2_211), .b(output_2_2), .y(output_1_211));
wire output_3_211, output_3_2, output_2_211;
mixer gate_output_2_211(.a(output_3_211), .b(output_3_2), .y(output_2_211));
wire output_1_212, output_1_0, output_0_212;
mixer gate_output_0_212(.a(output_1_212), .b(output_1_0), .y(output_0_212));
wire output_2_212, output_2_0, output_1_212;
mixer gate_output_1_212(.a(output_2_212), .b(output_2_0), .y(output_1_212));
wire output_3_212, output_3_0, output_2_212;
mixer gate_output_2_212(.a(output_3_212), .b(output_3_0), .y(output_2_212));
wire output_1_213, output_1_1, output_0_213;
mixer gate_output_0_213(.a(output_1_213), .b(output_1_1), .y(output_0_213));
wire output_2_213, output_2_1, output_1_213;
mixer gate_output_1_213(.a(output_2_213), .b(output_2_1), .y(output_1_213));
wire output_3_213, output_3_1, output_2_213;
mixer gate_output_2_213(.a(output_3_213), .b(output_3_1), .y(output_2_213));
wire output_1_214, output_1_2, output_0_214;
mixer gate_output_0_214(.a(output_1_214), .b(output_1_2), .y(output_0_214));
wire output_2_214, output_2_2, output_1_214;
mixer gate_output_1_214(.a(output_2_214), .b(output_2_2), .y(output_1_214));
wire output_3_214, output_3_2, output_2_214;
mixer gate_output_2_214(.a(output_3_214), .b(output_3_2), .y(output_2_214));
wire output_1_215, output_1_0, output_0_215;
mixer gate_output_0_215(.a(output_1_215), .b(output_1_0), .y(output_0_215));
wire output_2_215, output_2_0, output_1_215;
mixer gate_output_1_215(.a(output_2_215), .b(output_2_0), .y(output_1_215));
wire output_3_215, output_3_0, output_2_215;
mixer gate_output_2_215(.a(output_3_215), .b(output_3_0), .y(output_2_215));
wire output_1_216, output_1_1, output_0_216;
mixer gate_output_0_216(.a(output_1_216), .b(output_1_1), .y(output_0_216));
wire output_2_216, output_2_1, output_1_216;
mixer gate_output_1_216(.a(output_2_216), .b(output_2_1), .y(output_1_216));
wire output_3_216, output_3_1, output_2_216;
mixer gate_output_2_216(.a(output_3_216), .b(output_3_1), .y(output_2_216));
wire output_1_217, output_1_2, output_0_217;
mixer gate_output_0_217(.a(output_1_217), .b(output_1_2), .y(output_0_217));
wire output_2_217, output_2_2, output_1_217;
mixer gate_output_1_217(.a(output_2_217), .b(output_2_2), .y(output_1_217));
wire output_3_217, output_3_2, output_2_217;
mixer gate_output_2_217(.a(output_3_217), .b(output_3_2), .y(output_2_217));
wire output_1_218, output_1_0, output_0_218;
mixer gate_output_0_218(.a(output_1_218), .b(output_1_0), .y(output_0_218));
wire output_2_218, output_2_0, output_1_218;
mixer gate_output_1_218(.a(output_2_218), .b(output_2_0), .y(output_1_218));
wire output_3_218, output_3_0, output_2_218;
mixer gate_output_2_218(.a(output_3_218), .b(output_3_0), .y(output_2_218));
wire output_1_219, output_1_1, output_0_219;
mixer gate_output_0_219(.a(output_1_219), .b(output_1_1), .y(output_0_219));
wire output_2_219, output_2_1, output_1_219;
mixer gate_output_1_219(.a(output_2_219), .b(output_2_1), .y(output_1_219));
wire output_3_219, output_3_1, output_2_219;
mixer gate_output_2_219(.a(output_3_219), .b(output_3_1), .y(output_2_219));
wire output_1_220, output_1_2, output_0_220;
mixer gate_output_0_220(.a(output_1_220), .b(output_1_2), .y(output_0_220));
wire output_2_220, output_2_2, output_1_220;
mixer gate_output_1_220(.a(output_2_220), .b(output_2_2), .y(output_1_220));
wire output_3_220, output_3_2, output_2_220;
mixer gate_output_2_220(.a(output_3_220), .b(output_3_2), .y(output_2_220));
wire output_1_221, output_1_0, output_0_221;
mixer gate_output_0_221(.a(output_1_221), .b(output_1_0), .y(output_0_221));
wire output_2_221, output_2_0, output_1_221;
mixer gate_output_1_221(.a(output_2_221), .b(output_2_0), .y(output_1_221));
wire output_3_221, output_3_0, output_2_221;
mixer gate_output_2_221(.a(output_3_221), .b(output_3_0), .y(output_2_221));
wire output_1_222, output_1_1, output_0_222;
mixer gate_output_0_222(.a(output_1_222), .b(output_1_1), .y(output_0_222));
wire output_2_222, output_2_1, output_1_222;
mixer gate_output_1_222(.a(output_2_222), .b(output_2_1), .y(output_1_222));
wire output_3_222, output_3_1, output_2_222;
mixer gate_output_2_222(.a(output_3_222), .b(output_3_1), .y(output_2_222));
wire output_1_223, output_1_2, output_0_223;
mixer gate_output_0_223(.a(output_1_223), .b(output_1_2), .y(output_0_223));
wire output_2_223, output_2_2, output_1_223;
mixer gate_output_1_223(.a(output_2_223), .b(output_2_2), .y(output_1_223));
wire output_3_223, output_3_2, output_2_223;
mixer gate_output_2_223(.a(output_3_223), .b(output_3_2), .y(output_2_223));
wire output_1_224, output_1_0, output_0_224;
mixer gate_output_0_224(.a(output_1_224), .b(output_1_0), .y(output_0_224));
wire output_2_224, output_2_0, output_1_224;
mixer gate_output_1_224(.a(output_2_224), .b(output_2_0), .y(output_1_224));
wire output_3_224, output_3_0, output_2_224;
mixer gate_output_2_224(.a(output_3_224), .b(output_3_0), .y(output_2_224));
wire output_1_225, output_1_1, output_0_225;
mixer gate_output_0_225(.a(output_1_225), .b(output_1_1), .y(output_0_225));
wire output_2_225, output_2_1, output_1_225;
mixer gate_output_1_225(.a(output_2_225), .b(output_2_1), .y(output_1_225));
wire output_3_225, output_3_1, output_2_225;
mixer gate_output_2_225(.a(output_3_225), .b(output_3_1), .y(output_2_225));
wire output_1_226, output_1_2, output_0_226;
mixer gate_output_0_226(.a(output_1_226), .b(output_1_2), .y(output_0_226));
wire output_2_226, output_2_2, output_1_226;
mixer gate_output_1_226(.a(output_2_226), .b(output_2_2), .y(output_1_226));
wire output_3_226, output_3_2, output_2_226;
mixer gate_output_2_226(.a(output_3_226), .b(output_3_2), .y(output_2_226));
wire output_1_227, output_1_0, output_0_227;
mixer gate_output_0_227(.a(output_1_227), .b(output_1_0), .y(output_0_227));
wire output_2_227, output_2_0, output_1_227;
mixer gate_output_1_227(.a(output_2_227), .b(output_2_0), .y(output_1_227));
wire output_3_227, output_3_0, output_2_227;
mixer gate_output_2_227(.a(output_3_227), .b(output_3_0), .y(output_2_227));
wire output_1_228, output_1_1, output_0_228;
mixer gate_output_0_228(.a(output_1_228), .b(output_1_1), .y(output_0_228));
wire output_2_228, output_2_1, output_1_228;
mixer gate_output_1_228(.a(output_2_228), .b(output_2_1), .y(output_1_228));
wire output_3_228, output_3_1, output_2_228;
mixer gate_output_2_228(.a(output_3_228), .b(output_3_1), .y(output_2_228));
wire output_1_229, output_1_2, output_0_229;
mixer gate_output_0_229(.a(output_1_229), .b(output_1_2), .y(output_0_229));
wire output_2_229, output_2_2, output_1_229;
mixer gate_output_1_229(.a(output_2_229), .b(output_2_2), .y(output_1_229));
wire output_3_229, output_3_2, output_2_229;
mixer gate_output_2_229(.a(output_3_229), .b(output_3_2), .y(output_2_229));
wire output_1_230, output_1_0, output_0_230;
mixer gate_output_0_230(.a(output_1_230), .b(output_1_0), .y(output_0_230));
wire output_2_230, output_2_0, output_1_230;
mixer gate_output_1_230(.a(output_2_230), .b(output_2_0), .y(output_1_230));
wire output_3_230, output_3_0, output_2_230;
mixer gate_output_2_230(.a(output_3_230), .b(output_3_0), .y(output_2_230));
wire output_1_231, output_1_1, output_0_231;
mixer gate_output_0_231(.a(output_1_231), .b(output_1_1), .y(output_0_231));
wire output_2_231, output_2_1, output_1_231;
mixer gate_output_1_231(.a(output_2_231), .b(output_2_1), .y(output_1_231));
wire output_3_231, output_3_1, output_2_231;
mixer gate_output_2_231(.a(output_3_231), .b(output_3_1), .y(output_2_231));
wire output_1_232, output_1_2, output_0_232;
mixer gate_output_0_232(.a(output_1_232), .b(output_1_2), .y(output_0_232));
wire output_2_232, output_2_2, output_1_232;
mixer gate_output_1_232(.a(output_2_232), .b(output_2_2), .y(output_1_232));
wire output_3_232, output_3_2, output_2_232;
mixer gate_output_2_232(.a(output_3_232), .b(output_3_2), .y(output_2_232));
wire output_1_233, output_1_0, output_0_233;
mixer gate_output_0_233(.a(output_1_233), .b(output_1_0), .y(output_0_233));
wire output_2_233, output_2_0, output_1_233;
mixer gate_output_1_233(.a(output_2_233), .b(output_2_0), .y(output_1_233));
wire output_3_233, output_3_0, output_2_233;
mixer gate_output_2_233(.a(output_3_233), .b(output_3_0), .y(output_2_233));
wire output_1_234, output_1_1, output_0_234;
mixer gate_output_0_234(.a(output_1_234), .b(output_1_1), .y(output_0_234));
wire output_2_234, output_2_1, output_1_234;
mixer gate_output_1_234(.a(output_2_234), .b(output_2_1), .y(output_1_234));
wire output_3_234, output_3_1, output_2_234;
mixer gate_output_2_234(.a(output_3_234), .b(output_3_1), .y(output_2_234));
wire output_1_235, output_1_2, output_0_235;
mixer gate_output_0_235(.a(output_1_235), .b(output_1_2), .y(output_0_235));
wire output_2_235, output_2_2, output_1_235;
mixer gate_output_1_235(.a(output_2_235), .b(output_2_2), .y(output_1_235));
wire output_3_235, output_3_2, output_2_235;
mixer gate_output_2_235(.a(output_3_235), .b(output_3_2), .y(output_2_235));
wire output_1_236, output_1_0, output_0_236;
mixer gate_output_0_236(.a(output_1_236), .b(output_1_0), .y(output_0_236));
wire output_2_236, output_2_0, output_1_236;
mixer gate_output_1_236(.a(output_2_236), .b(output_2_0), .y(output_1_236));
wire output_3_236, output_3_0, output_2_236;
mixer gate_output_2_236(.a(output_3_236), .b(output_3_0), .y(output_2_236));
wire output_1_237, output_1_1, output_0_237;
mixer gate_output_0_237(.a(output_1_237), .b(output_1_1), .y(output_0_237));
wire output_2_237, output_2_1, output_1_237;
mixer gate_output_1_237(.a(output_2_237), .b(output_2_1), .y(output_1_237));
wire output_3_237, output_3_1, output_2_237;
mixer gate_output_2_237(.a(output_3_237), .b(output_3_1), .y(output_2_237));
wire output_1_238, output_1_2, output_0_238;
mixer gate_output_0_238(.a(output_1_238), .b(output_1_2), .y(output_0_238));
wire output_2_238, output_2_2, output_1_238;
mixer gate_output_1_238(.a(output_2_238), .b(output_2_2), .y(output_1_238));
wire output_3_238, output_3_2, output_2_238;
mixer gate_output_2_238(.a(output_3_238), .b(output_3_2), .y(output_2_238));
wire output_1_239, output_1_0, output_0_239;
mixer gate_output_0_239(.a(output_1_239), .b(output_1_0), .y(output_0_239));
wire output_2_239, output_2_0, output_1_239;
mixer gate_output_1_239(.a(output_2_239), .b(output_2_0), .y(output_1_239));
wire output_3_239, output_3_0, output_2_239;
mixer gate_output_2_239(.a(output_3_239), .b(output_3_0), .y(output_2_239));
wire output_1_240, output_1_1, output_0_240;
mixer gate_output_0_240(.a(output_1_240), .b(output_1_1), .y(output_0_240));
wire output_2_240, output_2_1, output_1_240;
mixer gate_output_1_240(.a(output_2_240), .b(output_2_1), .y(output_1_240));
wire output_3_240, output_3_1, output_2_240;
mixer gate_output_2_240(.a(output_3_240), .b(output_3_1), .y(output_2_240));
wire output_1_241, output_1_2, output_0_241;
mixer gate_output_0_241(.a(output_1_241), .b(output_1_2), .y(output_0_241));
wire output_2_241, output_2_2, output_1_241;
mixer gate_output_1_241(.a(output_2_241), .b(output_2_2), .y(output_1_241));
wire output_3_241, output_3_2, output_2_241;
mixer gate_output_2_241(.a(output_3_241), .b(output_3_2), .y(output_2_241));
wire output_1_242, output_1_0, output_0_242;
mixer gate_output_0_242(.a(output_1_242), .b(output_1_0), .y(output_0_242));
wire output_2_242, output_2_0, output_1_242;
mixer gate_output_1_242(.a(output_2_242), .b(output_2_0), .y(output_1_242));
wire output_3_242, output_3_0, output_2_242;
mixer gate_output_2_242(.a(output_3_242), .b(output_3_0), .y(output_2_242));
wire output_1_243, output_1_1, output_0_243;
mixer gate_output_0_243(.a(output_1_243), .b(output_1_1), .y(output_0_243));
wire output_2_243, output_2_1, output_1_243;
mixer gate_output_1_243(.a(output_2_243), .b(output_2_1), .y(output_1_243));
wire output_3_243, output_3_1, output_2_243;
mixer gate_output_2_243(.a(output_3_243), .b(output_3_1), .y(output_2_243));
wire output_1_244, output_1_2, output_0_244;
mixer gate_output_0_244(.a(output_1_244), .b(output_1_2), .y(output_0_244));
wire output_2_244, output_2_2, output_1_244;
mixer gate_output_1_244(.a(output_2_244), .b(output_2_2), .y(output_1_244));
wire output_3_244, output_3_2, output_2_244;
mixer gate_output_2_244(.a(output_3_244), .b(output_3_2), .y(output_2_244));
wire output_1_245, output_1_0, output_0_245;
mixer gate_output_0_245(.a(output_1_245), .b(output_1_0), .y(output_0_245));
wire output_2_245, output_2_0, output_1_245;
mixer gate_output_1_245(.a(output_2_245), .b(output_2_0), .y(output_1_245));
wire output_3_245, output_3_0, output_2_245;
mixer gate_output_2_245(.a(output_3_245), .b(output_3_0), .y(output_2_245));
wire output_1_246, output_1_1, output_0_246;
mixer gate_output_0_246(.a(output_1_246), .b(output_1_1), .y(output_0_246));
wire output_2_246, output_2_1, output_1_246;
mixer gate_output_1_246(.a(output_2_246), .b(output_2_1), .y(output_1_246));
wire output_3_246, output_3_1, output_2_246;
mixer gate_output_2_246(.a(output_3_246), .b(output_3_1), .y(output_2_246));
wire output_1_247, output_1_2, output_0_247;
mixer gate_output_0_247(.a(output_1_247), .b(output_1_2), .y(output_0_247));
wire output_2_247, output_2_2, output_1_247;
mixer gate_output_1_247(.a(output_2_247), .b(output_2_2), .y(output_1_247));
wire output_3_247, output_3_2, output_2_247;
mixer gate_output_2_247(.a(output_3_247), .b(output_3_2), .y(output_2_247));
wire output_1_248, output_1_0, output_0_248;
mixer gate_output_0_248(.a(output_1_248), .b(output_1_0), .y(output_0_248));
wire output_2_248, output_2_0, output_1_248;
mixer gate_output_1_248(.a(output_2_248), .b(output_2_0), .y(output_1_248));
wire output_3_248, output_3_0, output_2_248;
mixer gate_output_2_248(.a(output_3_248), .b(output_3_0), .y(output_2_248));
wire output_1_249, output_1_1, output_0_249;
mixer gate_output_0_249(.a(output_1_249), .b(output_1_1), .y(output_0_249));
wire output_2_249, output_2_1, output_1_249;
mixer gate_output_1_249(.a(output_2_249), .b(output_2_1), .y(output_1_249));
wire output_3_249, output_3_1, output_2_249;
mixer gate_output_2_249(.a(output_3_249), .b(output_3_1), .y(output_2_249));
wire output_1_250, output_1_2, output_0_250;
mixer gate_output_0_250(.a(output_1_250), .b(output_1_2), .y(output_0_250));
wire output_2_250, output_2_2, output_1_250;
mixer gate_output_1_250(.a(output_2_250), .b(output_2_2), .y(output_1_250));
wire output_3_250, output_3_2, output_2_250;
mixer gate_output_2_250(.a(output_3_250), .b(output_3_2), .y(output_2_250));
wire output_1_251, output_1_0, output_0_251;
mixer gate_output_0_251(.a(output_1_251), .b(output_1_0), .y(output_0_251));
wire output_2_251, output_2_0, output_1_251;
mixer gate_output_1_251(.a(output_2_251), .b(output_2_0), .y(output_1_251));
wire output_3_251, output_3_0, output_2_251;
mixer gate_output_2_251(.a(output_3_251), .b(output_3_0), .y(output_2_251));
wire output_1_252, output_1_1, output_0_252;
mixer gate_output_0_252(.a(output_1_252), .b(output_1_1), .y(output_0_252));
wire output_2_252, output_2_1, output_1_252;
mixer gate_output_1_252(.a(output_2_252), .b(output_2_1), .y(output_1_252));
wire output_3_252, output_3_1, output_2_252;
mixer gate_output_2_252(.a(output_3_252), .b(output_3_1), .y(output_2_252));
wire output_1_253, output_1_2, output_0_253;
mixer gate_output_0_253(.a(output_1_253), .b(output_1_2), .y(output_0_253));
wire output_2_253, output_2_2, output_1_253;
mixer gate_output_1_253(.a(output_2_253), .b(output_2_2), .y(output_1_253));
wire output_3_253, output_3_2, output_2_253;
mixer gate_output_2_253(.a(output_3_253), .b(output_3_2), .y(output_2_253));
wire output_1_254, output_1_0, output_0_254;
mixer gate_output_0_254(.a(output_1_254), .b(output_1_0), .y(output_0_254));
wire output_2_254, output_2_0, output_1_254;
mixer gate_output_1_254(.a(output_2_254), .b(output_2_0), .y(output_1_254));
wire output_3_254, output_3_0, output_2_254;
mixer gate_output_2_254(.a(output_3_254), .b(output_3_0), .y(output_2_254));
wire output_1_255, output_1_1, output_0_255;
mixer gate_output_0_255(.a(output_1_255), .b(output_1_1), .y(output_0_255));
wire output_2_255, output_2_1, output_1_255;
mixer gate_output_1_255(.a(output_2_255), .b(output_2_1), .y(output_1_255));
wire output_3_255, output_3_1, output_2_255;
mixer gate_output_2_255(.a(output_3_255), .b(output_3_1), .y(output_2_255));
wire output_1_256, output_1_2, output_0_256;
mixer gate_output_0_256(.a(output_1_256), .b(output_1_2), .y(output_0_256));
wire output_2_256, output_2_2, output_1_256;
mixer gate_output_1_256(.a(output_2_256), .b(output_2_2), .y(output_1_256));
wire output_3_256, output_3_2, output_2_256;
mixer gate_output_2_256(.a(output_3_256), .b(output_3_2), .y(output_2_256));
wire output_1_257, output_1_0, output_0_257;
mixer gate_output_0_257(.a(output_1_257), .b(output_1_0), .y(output_0_257));
wire output_2_257, output_2_0, output_1_257;
mixer gate_output_1_257(.a(output_2_257), .b(output_2_0), .y(output_1_257));
wire output_3_257, output_3_0, output_2_257;
mixer gate_output_2_257(.a(output_3_257), .b(output_3_0), .y(output_2_257));
wire output_1_258, output_1_1, output_0_258;
mixer gate_output_0_258(.a(output_1_258), .b(output_1_1), .y(output_0_258));
wire output_2_258, output_2_1, output_1_258;
mixer gate_output_1_258(.a(output_2_258), .b(output_2_1), .y(output_1_258));
wire output_3_258, output_3_1, output_2_258;
mixer gate_output_2_258(.a(output_3_258), .b(output_3_1), .y(output_2_258));
wire output_1_259, output_1_2, output_0_259;
mixer gate_output_0_259(.a(output_1_259), .b(output_1_2), .y(output_0_259));
wire output_2_259, output_2_2, output_1_259;
mixer gate_output_1_259(.a(output_2_259), .b(output_2_2), .y(output_1_259));
wire output_3_259, output_3_2, output_2_259;
mixer gate_output_2_259(.a(output_3_259), .b(output_3_2), .y(output_2_259));
wire output_1_260, output_1_0, output_0_260;
mixer gate_output_0_260(.a(output_1_260), .b(output_1_0), .y(output_0_260));
wire output_2_260, output_2_0, output_1_260;
mixer gate_output_1_260(.a(output_2_260), .b(output_2_0), .y(output_1_260));
wire output_3_260, output_3_0, output_2_260;
mixer gate_output_2_260(.a(output_3_260), .b(output_3_0), .y(output_2_260));
wire output_1_261, output_1_1, output_0_261;
mixer gate_output_0_261(.a(output_1_261), .b(output_1_1), .y(output_0_261));
wire output_2_261, output_2_1, output_1_261;
mixer gate_output_1_261(.a(output_2_261), .b(output_2_1), .y(output_1_261));
wire output_3_261, output_3_1, output_2_261;
mixer gate_output_2_261(.a(output_3_261), .b(output_3_1), .y(output_2_261));
wire output_1_262, output_1_2, output_0_262;
mixer gate_output_0_262(.a(output_1_262), .b(output_1_2), .y(output_0_262));
wire output_2_262, output_2_2, output_1_262;
mixer gate_output_1_262(.a(output_2_262), .b(output_2_2), .y(output_1_262));
wire output_3_262, output_3_2, output_2_262;
mixer gate_output_2_262(.a(output_3_262), .b(output_3_2), .y(output_2_262));
wire output_1_263, output_1_0, output_0_263;
mixer gate_output_0_263(.a(output_1_263), .b(output_1_0), .y(output_0_263));
wire output_2_263, output_2_0, output_1_263;
mixer gate_output_1_263(.a(output_2_263), .b(output_2_0), .y(output_1_263));
wire output_3_263, output_3_0, output_2_263;
mixer gate_output_2_263(.a(output_3_263), .b(output_3_0), .y(output_2_263));
wire output_1_264, output_1_1, output_0_264;
mixer gate_output_0_264(.a(output_1_264), .b(output_1_1), .y(output_0_264));
wire output_2_264, output_2_1, output_1_264;
mixer gate_output_1_264(.a(output_2_264), .b(output_2_1), .y(output_1_264));
wire output_3_264, output_3_1, output_2_264;
mixer gate_output_2_264(.a(output_3_264), .b(output_3_1), .y(output_2_264));
wire output_1_265, output_1_2, output_0_265;
mixer gate_output_0_265(.a(output_1_265), .b(output_1_2), .y(output_0_265));
wire output_2_265, output_2_2, output_1_265;
mixer gate_output_1_265(.a(output_2_265), .b(output_2_2), .y(output_1_265));
wire output_3_265, output_3_2, output_2_265;
mixer gate_output_2_265(.a(output_3_265), .b(output_3_2), .y(output_2_265));
wire output_1_266, output_1_0, output_0_266;
mixer gate_output_0_266(.a(output_1_266), .b(output_1_0), .y(output_0_266));
wire output_2_266, output_2_0, output_1_266;
mixer gate_output_1_266(.a(output_2_266), .b(output_2_0), .y(output_1_266));
wire output_3_266, output_3_0, output_2_266;
mixer gate_output_2_266(.a(output_3_266), .b(output_3_0), .y(output_2_266));
wire output_1_267, output_1_1, output_0_267;
mixer gate_output_0_267(.a(output_1_267), .b(output_1_1), .y(output_0_267));
wire output_2_267, output_2_1, output_1_267;
mixer gate_output_1_267(.a(output_2_267), .b(output_2_1), .y(output_1_267));
wire output_3_267, output_3_1, output_2_267;
mixer gate_output_2_267(.a(output_3_267), .b(output_3_1), .y(output_2_267));
wire output_1_268, output_1_2, output_0_268;
mixer gate_output_0_268(.a(output_1_268), .b(output_1_2), .y(output_0_268));
wire output_2_268, output_2_2, output_1_268;
mixer gate_output_1_268(.a(output_2_268), .b(output_2_2), .y(output_1_268));
wire output_3_268, output_3_2, output_2_268;
mixer gate_output_2_268(.a(output_3_268), .b(output_3_2), .y(output_2_268));
wire output_1_269, output_1_0, output_0_269;
mixer gate_output_0_269(.a(output_1_269), .b(output_1_0), .y(output_0_269));
wire output_2_269, output_2_0, output_1_269;
mixer gate_output_1_269(.a(output_2_269), .b(output_2_0), .y(output_1_269));
wire output_3_269, output_3_0, output_2_269;
mixer gate_output_2_269(.a(output_3_269), .b(output_3_0), .y(output_2_269));
wire output_1_270, output_1_1, output_0_270;
mixer gate_output_0_270(.a(output_1_270), .b(output_1_1), .y(output_0_270));
wire output_2_270, output_2_1, output_1_270;
mixer gate_output_1_270(.a(output_2_270), .b(output_2_1), .y(output_1_270));
wire output_3_270, output_3_1, output_2_270;
mixer gate_output_2_270(.a(output_3_270), .b(output_3_1), .y(output_2_270));
wire output_1_271, output_1_2, output_0_271;
mixer gate_output_0_271(.a(output_1_271), .b(output_1_2), .y(output_0_271));
wire output_2_271, output_2_2, output_1_271;
mixer gate_output_1_271(.a(output_2_271), .b(output_2_2), .y(output_1_271));
wire output_3_271, output_3_2, output_2_271;
mixer gate_output_2_271(.a(output_3_271), .b(output_3_2), .y(output_2_271));
wire output_1_272, output_1_0, output_0_272;
mixer gate_output_0_272(.a(output_1_272), .b(output_1_0), .y(output_0_272));
wire output_2_272, output_2_0, output_1_272;
mixer gate_output_1_272(.a(output_2_272), .b(output_2_0), .y(output_1_272));
wire output_3_272, output_3_0, output_2_272;
mixer gate_output_2_272(.a(output_3_272), .b(output_3_0), .y(output_2_272));
wire output_1_273, output_1_1, output_0_273;
mixer gate_output_0_273(.a(output_1_273), .b(output_1_1), .y(output_0_273));
wire output_2_273, output_2_1, output_1_273;
mixer gate_output_1_273(.a(output_2_273), .b(output_2_1), .y(output_1_273));
wire output_3_273, output_3_1, output_2_273;
mixer gate_output_2_273(.a(output_3_273), .b(output_3_1), .y(output_2_273));
wire output_1_274, output_1_2, output_0_274;
mixer gate_output_0_274(.a(output_1_274), .b(output_1_2), .y(output_0_274));
wire output_2_274, output_2_2, output_1_274;
mixer gate_output_1_274(.a(output_2_274), .b(output_2_2), .y(output_1_274));
wire output_3_274, output_3_2, output_2_274;
mixer gate_output_2_274(.a(output_3_274), .b(output_3_2), .y(output_2_274));
wire output_1_275, output_1_0, output_0_275;
mixer gate_output_0_275(.a(output_1_275), .b(output_1_0), .y(output_0_275));
wire output_2_275, output_2_0, output_1_275;
mixer gate_output_1_275(.a(output_2_275), .b(output_2_0), .y(output_1_275));
wire output_3_275, output_3_0, output_2_275;
mixer gate_output_2_275(.a(output_3_275), .b(output_3_0), .y(output_2_275));
wire output_1_276, output_1_1, output_0_276;
mixer gate_output_0_276(.a(output_1_276), .b(output_1_1), .y(output_0_276));
wire output_2_276, output_2_1, output_1_276;
mixer gate_output_1_276(.a(output_2_276), .b(output_2_1), .y(output_1_276));
wire output_3_276, output_3_1, output_2_276;
mixer gate_output_2_276(.a(output_3_276), .b(output_3_1), .y(output_2_276));
wire output_1_277, output_1_2, output_0_277;
mixer gate_output_0_277(.a(output_1_277), .b(output_1_2), .y(output_0_277));
wire output_2_277, output_2_2, output_1_277;
mixer gate_output_1_277(.a(output_2_277), .b(output_2_2), .y(output_1_277));
wire output_3_277, output_3_2, output_2_277;
mixer gate_output_2_277(.a(output_3_277), .b(output_3_2), .y(output_2_277));
wire output_1_278, output_1_0, output_0_278;
mixer gate_output_0_278(.a(output_1_278), .b(output_1_0), .y(output_0_278));
wire output_2_278, output_2_0, output_1_278;
mixer gate_output_1_278(.a(output_2_278), .b(output_2_0), .y(output_1_278));
wire output_3_278, output_3_0, output_2_278;
mixer gate_output_2_278(.a(output_3_278), .b(output_3_0), .y(output_2_278));
wire output_1_279, output_1_1, output_0_279;
mixer gate_output_0_279(.a(output_1_279), .b(output_1_1), .y(output_0_279));
wire output_2_279, output_2_1, output_1_279;
mixer gate_output_1_279(.a(output_2_279), .b(output_2_1), .y(output_1_279));
wire output_3_279, output_3_1, output_2_279;
mixer gate_output_2_279(.a(output_3_279), .b(output_3_1), .y(output_2_279));
wire output_1_280, output_1_2, output_0_280;
mixer gate_output_0_280(.a(output_1_280), .b(output_1_2), .y(output_0_280));
wire output_2_280, output_2_2, output_1_280;
mixer gate_output_1_280(.a(output_2_280), .b(output_2_2), .y(output_1_280));
wire output_3_280, output_3_2, output_2_280;
mixer gate_output_2_280(.a(output_3_280), .b(output_3_2), .y(output_2_280));
wire output_1_281, output_1_0, output_0_281;
mixer gate_output_0_281(.a(output_1_281), .b(output_1_0), .y(output_0_281));
wire output_2_281, output_2_0, output_1_281;
mixer gate_output_1_281(.a(output_2_281), .b(output_2_0), .y(output_1_281));
wire output_3_281, output_3_0, output_2_281;
mixer gate_output_2_281(.a(output_3_281), .b(output_3_0), .y(output_2_281));
wire output_1_282, output_1_1, output_0_282;
mixer gate_output_0_282(.a(output_1_282), .b(output_1_1), .y(output_0_282));
wire output_2_282, output_2_1, output_1_282;
mixer gate_output_1_282(.a(output_2_282), .b(output_2_1), .y(output_1_282));
wire output_3_282, output_3_1, output_2_282;
mixer gate_output_2_282(.a(output_3_282), .b(output_3_1), .y(output_2_282));
wire output_1_283, output_1_2, output_0_283;
mixer gate_output_0_283(.a(output_1_283), .b(output_1_2), .y(output_0_283));
wire output_2_283, output_2_2, output_1_283;
mixer gate_output_1_283(.a(output_2_283), .b(output_2_2), .y(output_1_283));
wire output_3_283, output_3_2, output_2_283;
mixer gate_output_2_283(.a(output_3_283), .b(output_3_2), .y(output_2_283));
wire output_1_284, output_1_0, output_0_284;
mixer gate_output_0_284(.a(output_1_284), .b(output_1_0), .y(output_0_284));
wire output_2_284, output_2_0, output_1_284;
mixer gate_output_1_284(.a(output_2_284), .b(output_2_0), .y(output_1_284));
wire output_3_284, output_3_0, output_2_284;
mixer gate_output_2_284(.a(output_3_284), .b(output_3_0), .y(output_2_284));
wire output_1_285, output_1_1, output_0_285;
mixer gate_output_0_285(.a(output_1_285), .b(output_1_1), .y(output_0_285));
wire output_2_285, output_2_1, output_1_285;
mixer gate_output_1_285(.a(output_2_285), .b(output_2_1), .y(output_1_285));
wire output_3_285, output_3_1, output_2_285;
mixer gate_output_2_285(.a(output_3_285), .b(output_3_1), .y(output_2_285));
wire output_1_286, output_1_2, output_0_286;
mixer gate_output_0_286(.a(output_1_286), .b(output_1_2), .y(output_0_286));
wire output_2_286, output_2_2, output_1_286;
mixer gate_output_1_286(.a(output_2_286), .b(output_2_2), .y(output_1_286));
wire output_3_286, output_3_2, output_2_286;
mixer gate_output_2_286(.a(output_3_286), .b(output_3_2), .y(output_2_286));
wire output_1_287, output_1_0, output_0_287;
mixer gate_output_0_287(.a(output_1_287), .b(output_1_0), .y(output_0_287));
wire output_2_287, output_2_0, output_1_287;
mixer gate_output_1_287(.a(output_2_287), .b(output_2_0), .y(output_1_287));
wire output_3_287, output_3_0, output_2_287;
mixer gate_output_2_287(.a(output_3_287), .b(output_3_0), .y(output_2_287));
wire output_1_288, output_1_1, output_0_288;
mixer gate_output_0_288(.a(output_1_288), .b(output_1_1), .y(output_0_288));
wire output_2_288, output_2_1, output_1_288;
mixer gate_output_1_288(.a(output_2_288), .b(output_2_1), .y(output_1_288));
wire output_3_288, output_3_1, output_2_288;
mixer gate_output_2_288(.a(output_3_288), .b(output_3_1), .y(output_2_288));
wire output_1_289, output_1_2, output_0_289;
mixer gate_output_0_289(.a(output_1_289), .b(output_1_2), .y(output_0_289));
wire output_2_289, output_2_2, output_1_289;
mixer gate_output_1_289(.a(output_2_289), .b(output_2_2), .y(output_1_289));
wire output_3_289, output_3_2, output_2_289;
mixer gate_output_2_289(.a(output_3_289), .b(output_3_2), .y(output_2_289));
wire output_1_290, output_1_0, output_0_290;
mixer gate_output_0_290(.a(output_1_290), .b(output_1_0), .y(output_0_290));
wire output_2_290, output_2_0, output_1_290;
mixer gate_output_1_290(.a(output_2_290), .b(output_2_0), .y(output_1_290));
wire output_3_290, output_3_0, output_2_290;
mixer gate_output_2_290(.a(output_3_290), .b(output_3_0), .y(output_2_290));
wire output_1_291, output_1_1, output_0_291;
mixer gate_output_0_291(.a(output_1_291), .b(output_1_1), .y(output_0_291));
wire output_2_291, output_2_1, output_1_291;
mixer gate_output_1_291(.a(output_2_291), .b(output_2_1), .y(output_1_291));
wire output_3_291, output_3_1, output_2_291;
mixer gate_output_2_291(.a(output_3_291), .b(output_3_1), .y(output_2_291));
wire output_1_292, output_1_2, output_0_292;
mixer gate_output_0_292(.a(output_1_292), .b(output_1_2), .y(output_0_292));
wire output_2_292, output_2_2, output_1_292;
mixer gate_output_1_292(.a(output_2_292), .b(output_2_2), .y(output_1_292));
wire output_3_292, output_3_2, output_2_292;
mixer gate_output_2_292(.a(output_3_292), .b(output_3_2), .y(output_2_292));
wire output_1_293, output_1_0, output_0_293;
mixer gate_output_0_293(.a(output_1_293), .b(output_1_0), .y(output_0_293));
wire output_2_293, output_2_0, output_1_293;
mixer gate_output_1_293(.a(output_2_293), .b(output_2_0), .y(output_1_293));
wire output_3_293, output_3_0, output_2_293;
mixer gate_output_2_293(.a(output_3_293), .b(output_3_0), .y(output_2_293));
wire output_1_294, output_1_1, output_0_294;
mixer gate_output_0_294(.a(output_1_294), .b(output_1_1), .y(output_0_294));
wire output_2_294, output_2_1, output_1_294;
mixer gate_output_1_294(.a(output_2_294), .b(output_2_1), .y(output_1_294));
wire output_3_294, output_3_1, output_2_294;
mixer gate_output_2_294(.a(output_3_294), .b(output_3_1), .y(output_2_294));
wire output_1_295, output_1_2, output_0_295;
mixer gate_output_0_295(.a(output_1_295), .b(output_1_2), .y(output_0_295));
wire output_2_295, output_2_2, output_1_295;
mixer gate_output_1_295(.a(output_2_295), .b(output_2_2), .y(output_1_295));
wire output_3_295, output_3_2, output_2_295;
mixer gate_output_2_295(.a(output_3_295), .b(output_3_2), .y(output_2_295));
wire output_1_296, output_1_0, output_0_296;
mixer gate_output_0_296(.a(output_1_296), .b(output_1_0), .y(output_0_296));
wire output_2_296, output_2_0, output_1_296;
mixer gate_output_1_296(.a(output_2_296), .b(output_2_0), .y(output_1_296));
wire output_3_296, output_3_0, output_2_296;
mixer gate_output_2_296(.a(output_3_296), .b(output_3_0), .y(output_2_296));
wire output_1_297, output_1_1, output_0_297;
mixer gate_output_0_297(.a(output_1_297), .b(output_1_1), .y(output_0_297));
wire output_2_297, output_2_1, output_1_297;
mixer gate_output_1_297(.a(output_2_297), .b(output_2_1), .y(output_1_297));
wire output_3_297, output_3_1, output_2_297;
mixer gate_output_2_297(.a(output_3_297), .b(output_3_1), .y(output_2_297));
wire output_1_298, output_1_2, output_0_298;
mixer gate_output_0_298(.a(output_1_298), .b(output_1_2), .y(output_0_298));
wire output_2_298, output_2_2, output_1_298;
mixer gate_output_1_298(.a(output_2_298), .b(output_2_2), .y(output_1_298));
wire output_3_298, output_3_2, output_2_298;
mixer gate_output_2_298(.a(output_3_298), .b(output_3_2), .y(output_2_298));
wire output_1_299, output_1_0, output_0_299;
mixer gate_output_0_299(.a(output_1_299), .b(output_1_0), .y(output_0_299));
wire output_2_299, output_2_0, output_1_299;
mixer gate_output_1_299(.a(output_2_299), .b(output_2_0), .y(output_1_299));
wire output_3_299, output_3_0, output_2_299;
mixer gate_output_2_299(.a(output_3_299), .b(output_3_0), .y(output_2_299));
wire output_1_300, output_1_1, output_0_300;
mixer gate_output_0_300(.a(output_1_300), .b(output_1_1), .y(output_0_300));
wire output_2_300, output_2_1, output_1_300;
mixer gate_output_1_300(.a(output_2_300), .b(output_2_1), .y(output_1_300));
wire output_3_300, output_3_1, output_2_300;
mixer gate_output_2_300(.a(output_3_300), .b(output_3_1), .y(output_2_300));
wire output_1_301, output_1_2, output_0_301;
mixer gate_output_0_301(.a(output_1_301), .b(output_1_2), .y(output_0_301));
wire output_2_301, output_2_2, output_1_301;
mixer gate_output_1_301(.a(output_2_301), .b(output_2_2), .y(output_1_301));
wire output_3_301, output_3_2, output_2_301;
mixer gate_output_2_301(.a(output_3_301), .b(output_3_2), .y(output_2_301));
wire output_1_302, output_1_0, output_0_302;
mixer gate_output_0_302(.a(output_1_302), .b(output_1_0), .y(output_0_302));
wire output_2_302, output_2_0, output_1_302;
mixer gate_output_1_302(.a(output_2_302), .b(output_2_0), .y(output_1_302));
wire output_3_302, output_3_0, output_2_302;
mixer gate_output_2_302(.a(output_3_302), .b(output_3_0), .y(output_2_302));
wire output_1_303, output_1_1, output_0_303;
mixer gate_output_0_303(.a(output_1_303), .b(output_1_1), .y(output_0_303));
wire output_2_303, output_2_1, output_1_303;
mixer gate_output_1_303(.a(output_2_303), .b(output_2_1), .y(output_1_303));
wire output_3_303, output_3_1, output_2_303;
mixer gate_output_2_303(.a(output_3_303), .b(output_3_1), .y(output_2_303));
wire output_1_304, output_1_2, output_0_304;
mixer gate_output_0_304(.a(output_1_304), .b(output_1_2), .y(output_0_304));
wire output_2_304, output_2_2, output_1_304;
mixer gate_output_1_304(.a(output_2_304), .b(output_2_2), .y(output_1_304));
wire output_3_304, output_3_2, output_2_304;
mixer gate_output_2_304(.a(output_3_304), .b(output_3_2), .y(output_2_304));
wire output_1_305, output_1_0, output_0_305;
mixer gate_output_0_305(.a(output_1_305), .b(output_1_0), .y(output_0_305));
wire output_2_305, output_2_0, output_1_305;
mixer gate_output_1_305(.a(output_2_305), .b(output_2_0), .y(output_1_305));
wire output_3_305, output_3_0, output_2_305;
mixer gate_output_2_305(.a(output_3_305), .b(output_3_0), .y(output_2_305));
wire output_1_306, output_1_1, output_0_306;
mixer gate_output_0_306(.a(output_1_306), .b(output_1_1), .y(output_0_306));
wire output_2_306, output_2_1, output_1_306;
mixer gate_output_1_306(.a(output_2_306), .b(output_2_1), .y(output_1_306));
wire output_3_306, output_3_1, output_2_306;
mixer gate_output_2_306(.a(output_3_306), .b(output_3_1), .y(output_2_306));
wire output_1_307, output_1_2, output_0_307;
mixer gate_output_0_307(.a(output_1_307), .b(output_1_2), .y(output_0_307));
wire output_2_307, output_2_2, output_1_307;
mixer gate_output_1_307(.a(output_2_307), .b(output_2_2), .y(output_1_307));
wire output_3_307, output_3_2, output_2_307;
mixer gate_output_2_307(.a(output_3_307), .b(output_3_2), .y(output_2_307));
wire output_1_308, output_1_0, output_0_308;
mixer gate_output_0_308(.a(output_1_308), .b(output_1_0), .y(output_0_308));
wire output_2_308, output_2_0, output_1_308;
mixer gate_output_1_308(.a(output_2_308), .b(output_2_0), .y(output_1_308));
wire output_3_308, output_3_0, output_2_308;
mixer gate_output_2_308(.a(output_3_308), .b(output_3_0), .y(output_2_308));
wire output_1_309, output_1_1, output_0_309;
mixer gate_output_0_309(.a(output_1_309), .b(output_1_1), .y(output_0_309));
wire output_2_309, output_2_1, output_1_309;
mixer gate_output_1_309(.a(output_2_309), .b(output_2_1), .y(output_1_309));
wire output_3_309, output_3_1, output_2_309;
mixer gate_output_2_309(.a(output_3_309), .b(output_3_1), .y(output_2_309));
wire output_1_310, output_1_2, output_0_310;
mixer gate_output_0_310(.a(output_1_310), .b(output_1_2), .y(output_0_310));
wire output_2_310, output_2_2, output_1_310;
mixer gate_output_1_310(.a(output_2_310), .b(output_2_2), .y(output_1_310));
wire output_3_310, output_3_2, output_2_310;
mixer gate_output_2_310(.a(output_3_310), .b(output_3_2), .y(output_2_310));
wire output_1_311, output_1_0, output_0_311;
mixer gate_output_0_311(.a(output_1_311), .b(output_1_0), .y(output_0_311));
wire output_2_311, output_2_0, output_1_311;
mixer gate_output_1_311(.a(output_2_311), .b(output_2_0), .y(output_1_311));
wire output_3_311, output_3_0, output_2_311;
mixer gate_output_2_311(.a(output_3_311), .b(output_3_0), .y(output_2_311));
wire output_1_312, output_1_1, output_0_312;
mixer gate_output_0_312(.a(output_1_312), .b(output_1_1), .y(output_0_312));
wire output_2_312, output_2_1, output_1_312;
mixer gate_output_1_312(.a(output_2_312), .b(output_2_1), .y(output_1_312));
wire output_3_312, output_3_1, output_2_312;
mixer gate_output_2_312(.a(output_3_312), .b(output_3_1), .y(output_2_312));
wire output_1_313, output_1_2, output_0_313;
mixer gate_output_0_313(.a(output_1_313), .b(output_1_2), .y(output_0_313));
wire output_2_313, output_2_2, output_1_313;
mixer gate_output_1_313(.a(output_2_313), .b(output_2_2), .y(output_1_313));
wire output_3_313, output_3_2, output_2_313;
mixer gate_output_2_313(.a(output_3_313), .b(output_3_2), .y(output_2_313));
wire output_1_314, output_1_0, output_0_314;
mixer gate_output_0_314(.a(output_1_314), .b(output_1_0), .y(output_0_314));
wire output_2_314, output_2_0, output_1_314;
mixer gate_output_1_314(.a(output_2_314), .b(output_2_0), .y(output_1_314));
wire output_3_314, output_3_0, output_2_314;
mixer gate_output_2_314(.a(output_3_314), .b(output_3_0), .y(output_2_314));
wire output_1_315, output_1_1, output_0_315;
mixer gate_output_0_315(.a(output_1_315), .b(output_1_1), .y(output_0_315));
wire output_2_315, output_2_1, output_1_315;
mixer gate_output_1_315(.a(output_2_315), .b(output_2_1), .y(output_1_315));
wire output_3_315, output_3_1, output_2_315;
mixer gate_output_2_315(.a(output_3_315), .b(output_3_1), .y(output_2_315));
wire output_1_316, output_1_2, output_0_316;
mixer gate_output_0_316(.a(output_1_316), .b(output_1_2), .y(output_0_316));
wire output_2_316, output_2_2, output_1_316;
mixer gate_output_1_316(.a(output_2_316), .b(output_2_2), .y(output_1_316));
wire output_3_316, output_3_2, output_2_316;
mixer gate_output_2_316(.a(output_3_316), .b(output_3_2), .y(output_2_316));
wire output_1_317, output_1_0, output_0_317;
mixer gate_output_0_317(.a(output_1_317), .b(output_1_0), .y(output_0_317));
wire output_2_317, output_2_0, output_1_317;
mixer gate_output_1_317(.a(output_2_317), .b(output_2_0), .y(output_1_317));
wire output_3_317, output_3_0, output_2_317;
mixer gate_output_2_317(.a(output_3_317), .b(output_3_0), .y(output_2_317));
wire output_1_318, output_1_1, output_0_318;
mixer gate_output_0_318(.a(output_1_318), .b(output_1_1), .y(output_0_318));
wire output_2_318, output_2_1, output_1_318;
mixer gate_output_1_318(.a(output_2_318), .b(output_2_1), .y(output_1_318));
wire output_3_318, output_3_1, output_2_318;
mixer gate_output_2_318(.a(output_3_318), .b(output_3_1), .y(output_2_318));
wire output_1_319, output_1_2, output_0_319;
mixer gate_output_0_319(.a(output_1_319), .b(output_1_2), .y(output_0_319));
wire output_2_319, output_2_2, output_1_319;
mixer gate_output_1_319(.a(output_2_319), .b(output_2_2), .y(output_1_319));
wire output_3_319, output_3_2, output_2_319;
mixer gate_output_2_319(.a(output_3_319), .b(output_3_2), .y(output_2_319));
wire output_1_320, output_1_0, output_0_320;
mixer gate_output_0_320(.a(output_1_320), .b(output_1_0), .y(output_0_320));
wire output_2_320, output_2_0, output_1_320;
mixer gate_output_1_320(.a(output_2_320), .b(output_2_0), .y(output_1_320));
wire output_3_320, output_3_0, output_2_320;
mixer gate_output_2_320(.a(output_3_320), .b(output_3_0), .y(output_2_320));
wire output_1_321, output_1_1, output_0_321;
mixer gate_output_0_321(.a(output_1_321), .b(output_1_1), .y(output_0_321));
wire output_2_321, output_2_1, output_1_321;
mixer gate_output_1_321(.a(output_2_321), .b(output_2_1), .y(output_1_321));
wire output_3_321, output_3_1, output_2_321;
mixer gate_output_2_321(.a(output_3_321), .b(output_3_1), .y(output_2_321));
wire output_1_322, output_1_2, output_0_322;
mixer gate_output_0_322(.a(output_1_322), .b(output_1_2), .y(output_0_322));
wire output_2_322, output_2_2, output_1_322;
mixer gate_output_1_322(.a(output_2_322), .b(output_2_2), .y(output_1_322));
wire output_3_322, output_3_2, output_2_322;
mixer gate_output_2_322(.a(output_3_322), .b(output_3_2), .y(output_2_322));
wire output_1_323, output_1_0, output_0_323;
mixer gate_output_0_323(.a(output_1_323), .b(output_1_0), .y(output_0_323));
wire output_2_323, output_2_0, output_1_323;
mixer gate_output_1_323(.a(output_2_323), .b(output_2_0), .y(output_1_323));
wire output_3_323, output_3_0, output_2_323;
mixer gate_output_2_323(.a(output_3_323), .b(output_3_0), .y(output_2_323));
wire output_1_324, output_1_1, output_0_324;
mixer gate_output_0_324(.a(output_1_324), .b(output_1_1), .y(output_0_324));
wire output_2_324, output_2_1, output_1_324;
mixer gate_output_1_324(.a(output_2_324), .b(output_2_1), .y(output_1_324));
wire output_3_324, output_3_1, output_2_324;
mixer gate_output_2_324(.a(output_3_324), .b(output_3_1), .y(output_2_324));
wire output_1_325, output_1_2, output_0_325;
mixer gate_output_0_325(.a(output_1_325), .b(output_1_2), .y(output_0_325));
wire output_2_325, output_2_2, output_1_325;
mixer gate_output_1_325(.a(output_2_325), .b(output_2_2), .y(output_1_325));
wire output_3_325, output_3_2, output_2_325;
mixer gate_output_2_325(.a(output_3_325), .b(output_3_2), .y(output_2_325));
wire output_1_326, output_1_0, output_0_326;
mixer gate_output_0_326(.a(output_1_326), .b(output_1_0), .y(output_0_326));
wire output_2_326, output_2_0, output_1_326;
mixer gate_output_1_326(.a(output_2_326), .b(output_2_0), .y(output_1_326));
wire output_3_326, output_3_0, output_2_326;
mixer gate_output_2_326(.a(output_3_326), .b(output_3_0), .y(output_2_326));
wire output_1_327, output_1_1, output_0_327;
mixer gate_output_0_327(.a(output_1_327), .b(output_1_1), .y(output_0_327));
wire output_2_327, output_2_1, output_1_327;
mixer gate_output_1_327(.a(output_2_327), .b(output_2_1), .y(output_1_327));
wire output_3_327, output_3_1, output_2_327;
mixer gate_output_2_327(.a(output_3_327), .b(output_3_1), .y(output_2_327));
wire output_1_328, output_1_2, output_0_328;
mixer gate_output_0_328(.a(output_1_328), .b(output_1_2), .y(output_0_328));
wire output_2_328, output_2_2, output_1_328;
mixer gate_output_1_328(.a(output_2_328), .b(output_2_2), .y(output_1_328));
wire output_3_328, output_3_2, output_2_328;
mixer gate_output_2_328(.a(output_3_328), .b(output_3_2), .y(output_2_328));
wire output_1_329, output_1_0, output_0_329;
mixer gate_output_0_329(.a(output_1_329), .b(output_1_0), .y(output_0_329));
wire output_2_329, output_2_0, output_1_329;
mixer gate_output_1_329(.a(output_2_329), .b(output_2_0), .y(output_1_329));
wire output_3_329, output_3_0, output_2_329;
mixer gate_output_2_329(.a(output_3_329), .b(output_3_0), .y(output_2_329));
wire output_1_330, output_1_1, output_0_330;
mixer gate_output_0_330(.a(output_1_330), .b(output_1_1), .y(output_0_330));
wire output_2_330, output_2_1, output_1_330;
mixer gate_output_1_330(.a(output_2_330), .b(output_2_1), .y(output_1_330));
wire output_3_330, output_3_1, output_2_330;
mixer gate_output_2_330(.a(output_3_330), .b(output_3_1), .y(output_2_330));
wire output_1_331, output_1_2, output_0_331;
mixer gate_output_0_331(.a(output_1_331), .b(output_1_2), .y(output_0_331));
wire output_2_331, output_2_2, output_1_331;
mixer gate_output_1_331(.a(output_2_331), .b(output_2_2), .y(output_1_331));
wire output_3_331, output_3_2, output_2_331;
mixer gate_output_2_331(.a(output_3_331), .b(output_3_2), .y(output_2_331));
wire output_1_332, output_1_0, output_0_332;
mixer gate_output_0_332(.a(output_1_332), .b(output_1_0), .y(output_0_332));
wire output_2_332, output_2_0, output_1_332;
mixer gate_output_1_332(.a(output_2_332), .b(output_2_0), .y(output_1_332));
wire output_3_332, output_3_0, output_2_332;
mixer gate_output_2_332(.a(output_3_332), .b(output_3_0), .y(output_2_332));
wire output_1_333, output_1_1, output_0_333;
mixer gate_output_0_333(.a(output_1_333), .b(output_1_1), .y(output_0_333));
wire output_2_333, output_2_1, output_1_333;
mixer gate_output_1_333(.a(output_2_333), .b(output_2_1), .y(output_1_333));
wire output_3_333, output_3_1, output_2_333;
mixer gate_output_2_333(.a(output_3_333), .b(output_3_1), .y(output_2_333));
wire output_1_334, output_1_2, output_0_334;
mixer gate_output_0_334(.a(output_1_334), .b(output_1_2), .y(output_0_334));
wire output_2_334, output_2_2, output_1_334;
mixer gate_output_1_334(.a(output_2_334), .b(output_2_2), .y(output_1_334));
wire output_3_334, output_3_2, output_2_334;
mixer gate_output_2_334(.a(output_3_334), .b(output_3_2), .y(output_2_334));
wire output_1_335, output_1_0, output_0_335;
mixer gate_output_0_335(.a(output_1_335), .b(output_1_0), .y(output_0_335));
wire output_2_335, output_2_0, output_1_335;
mixer gate_output_1_335(.a(output_2_335), .b(output_2_0), .y(output_1_335));
wire output_3_335, output_3_0, output_2_335;
mixer gate_output_2_335(.a(output_3_335), .b(output_3_0), .y(output_2_335));
wire output_1_336, output_1_1, output_0_336;
mixer gate_output_0_336(.a(output_1_336), .b(output_1_1), .y(output_0_336));
wire output_2_336, output_2_1, output_1_336;
mixer gate_output_1_336(.a(output_2_336), .b(output_2_1), .y(output_1_336));
wire output_3_336, output_3_1, output_2_336;
mixer gate_output_2_336(.a(output_3_336), .b(output_3_1), .y(output_2_336));
wire output_1_337, output_1_2, output_0_337;
mixer gate_output_0_337(.a(output_1_337), .b(output_1_2), .y(output_0_337));
wire output_2_337, output_2_2, output_1_337;
mixer gate_output_1_337(.a(output_2_337), .b(output_2_2), .y(output_1_337));
wire output_3_337, output_3_2, output_2_337;
mixer gate_output_2_337(.a(output_3_337), .b(output_3_2), .y(output_2_337));
wire output_1_338, output_1_0, output_0_338;
mixer gate_output_0_338(.a(output_1_338), .b(output_1_0), .y(output_0_338));
wire output_2_338, output_2_0, output_1_338;
mixer gate_output_1_338(.a(output_2_338), .b(output_2_0), .y(output_1_338));
wire output_3_338, output_3_0, output_2_338;
mixer gate_output_2_338(.a(output_3_338), .b(output_3_0), .y(output_2_338));
wire output_1_339, output_1_1, output_0_339;
mixer gate_output_0_339(.a(output_1_339), .b(output_1_1), .y(output_0_339));
wire output_2_339, output_2_1, output_1_339;
mixer gate_output_1_339(.a(output_2_339), .b(output_2_1), .y(output_1_339));
wire output_3_339, output_3_1, output_2_339;
mixer gate_output_2_339(.a(output_3_339), .b(output_3_1), .y(output_2_339));
wire output_1_340, output_1_2, output_0_340;
mixer gate_output_0_340(.a(output_1_340), .b(output_1_2), .y(output_0_340));
wire output_2_340, output_2_2, output_1_340;
mixer gate_output_1_340(.a(output_2_340), .b(output_2_2), .y(output_1_340));
wire output_3_340, output_3_2, output_2_340;
mixer gate_output_2_340(.a(output_3_340), .b(output_3_2), .y(output_2_340));
wire output_1_341, output_1_0, output_0_341;
mixer gate_output_0_341(.a(output_1_341), .b(output_1_0), .y(output_0_341));
wire output_2_341, output_2_0, output_1_341;
mixer gate_output_1_341(.a(output_2_341), .b(output_2_0), .y(output_1_341));
wire output_3_341, output_3_0, output_2_341;
mixer gate_output_2_341(.a(output_3_341), .b(output_3_0), .y(output_2_341));
wire output_1_342, output_1_1, output_0_342;
mixer gate_output_0_342(.a(output_1_342), .b(output_1_1), .y(output_0_342));
wire output_2_342, output_2_1, output_1_342;
mixer gate_output_1_342(.a(output_2_342), .b(output_2_1), .y(output_1_342));
wire output_3_342, output_3_1, output_2_342;
mixer gate_output_2_342(.a(output_3_342), .b(output_3_1), .y(output_2_342));
wire output_1_343, output_1_2, output_0_343;
mixer gate_output_0_343(.a(output_1_343), .b(output_1_2), .y(output_0_343));
wire output_2_343, output_2_2, output_1_343;
mixer gate_output_1_343(.a(output_2_343), .b(output_2_2), .y(output_1_343));
wire output_3_343, output_3_2, output_2_343;
mixer gate_output_2_343(.a(output_3_343), .b(output_3_2), .y(output_2_343));
wire output_1_344, output_1_0, output_0_344;
mixer gate_output_0_344(.a(output_1_344), .b(output_1_0), .y(output_0_344));
wire output_2_344, output_2_0, output_1_344;
mixer gate_output_1_344(.a(output_2_344), .b(output_2_0), .y(output_1_344));
wire output_3_344, output_3_0, output_2_344;
mixer gate_output_2_344(.a(output_3_344), .b(output_3_0), .y(output_2_344));
wire output_1_345, output_1_1, output_0_345;
mixer gate_output_0_345(.a(output_1_345), .b(output_1_1), .y(output_0_345));
wire output_2_345, output_2_1, output_1_345;
mixer gate_output_1_345(.a(output_2_345), .b(output_2_1), .y(output_1_345));
wire output_3_345, output_3_1, output_2_345;
mixer gate_output_2_345(.a(output_3_345), .b(output_3_1), .y(output_2_345));
wire output_1_346, output_1_2, output_0_346;
mixer gate_output_0_346(.a(output_1_346), .b(output_1_2), .y(output_0_346));
wire output_2_346, output_2_2, output_1_346;
mixer gate_output_1_346(.a(output_2_346), .b(output_2_2), .y(output_1_346));
wire output_3_346, output_3_2, output_2_346;
mixer gate_output_2_346(.a(output_3_346), .b(output_3_2), .y(output_2_346));
wire output_1_347, output_1_0, output_0_347;
mixer gate_output_0_347(.a(output_1_347), .b(output_1_0), .y(output_0_347));
wire output_2_347, output_2_0, output_1_347;
mixer gate_output_1_347(.a(output_2_347), .b(output_2_0), .y(output_1_347));
wire output_3_347, output_3_0, output_2_347;
mixer gate_output_2_347(.a(output_3_347), .b(output_3_0), .y(output_2_347));
wire output_1_348, output_1_1, output_0_348;
mixer gate_output_0_348(.a(output_1_348), .b(output_1_1), .y(output_0_348));
wire output_2_348, output_2_1, output_1_348;
mixer gate_output_1_348(.a(output_2_348), .b(output_2_1), .y(output_1_348));
wire output_3_348, output_3_1, output_2_348;
mixer gate_output_2_348(.a(output_3_348), .b(output_3_1), .y(output_2_348));
wire output_1_349, output_1_2, output_0_349;
mixer gate_output_0_349(.a(output_1_349), .b(output_1_2), .y(output_0_349));
wire output_2_349, output_2_2, output_1_349;
mixer gate_output_1_349(.a(output_2_349), .b(output_2_2), .y(output_1_349));
wire output_3_349, output_3_2, output_2_349;
mixer gate_output_2_349(.a(output_3_349), .b(output_3_2), .y(output_2_349));
wire output_1_350, output_1_0, output_0_350;
mixer gate_output_0_350(.a(output_1_350), .b(output_1_0), .y(output_0_350));
wire output_2_350, output_2_0, output_1_350;
mixer gate_output_1_350(.a(output_2_350), .b(output_2_0), .y(output_1_350));
wire output_3_350, output_3_0, output_2_350;
mixer gate_output_2_350(.a(output_3_350), .b(output_3_0), .y(output_2_350));
wire output_1_351, output_1_1, output_0_351;
mixer gate_output_0_351(.a(output_1_351), .b(output_1_1), .y(output_0_351));
wire output_2_351, output_2_1, output_1_351;
mixer gate_output_1_351(.a(output_2_351), .b(output_2_1), .y(output_1_351));
wire output_3_351, output_3_1, output_2_351;
mixer gate_output_2_351(.a(output_3_351), .b(output_3_1), .y(output_2_351));
wire output_1_352, output_1_2, output_0_352;
mixer gate_output_0_352(.a(output_1_352), .b(output_1_2), .y(output_0_352));
wire output_2_352, output_2_2, output_1_352;
mixer gate_output_1_352(.a(output_2_352), .b(output_2_2), .y(output_1_352));
wire output_3_352, output_3_2, output_2_352;
mixer gate_output_2_352(.a(output_3_352), .b(output_3_2), .y(output_2_352));
wire output_1_353, output_1_0, output_0_353;
mixer gate_output_0_353(.a(output_1_353), .b(output_1_0), .y(output_0_353));
wire output_2_353, output_2_0, output_1_353;
mixer gate_output_1_353(.a(output_2_353), .b(output_2_0), .y(output_1_353));
wire output_3_353, output_3_0, output_2_353;
mixer gate_output_2_353(.a(output_3_353), .b(output_3_0), .y(output_2_353));
wire output_1_354, output_1_1, output_0_354;
mixer gate_output_0_354(.a(output_1_354), .b(output_1_1), .y(output_0_354));
wire output_2_354, output_2_1, output_1_354;
mixer gate_output_1_354(.a(output_2_354), .b(output_2_1), .y(output_1_354));
wire output_3_354, output_3_1, output_2_354;
mixer gate_output_2_354(.a(output_3_354), .b(output_3_1), .y(output_2_354));
wire output_1_355, output_1_2, output_0_355;
mixer gate_output_0_355(.a(output_1_355), .b(output_1_2), .y(output_0_355));
wire output_2_355, output_2_2, output_1_355;
mixer gate_output_1_355(.a(output_2_355), .b(output_2_2), .y(output_1_355));
wire output_3_355, output_3_2, output_2_355;
mixer gate_output_2_355(.a(output_3_355), .b(output_3_2), .y(output_2_355));
wire output_1_356, output_1_0, output_0_356;
mixer gate_output_0_356(.a(output_1_356), .b(output_1_0), .y(output_0_356));
wire output_2_356, output_2_0, output_1_356;
mixer gate_output_1_356(.a(output_2_356), .b(output_2_0), .y(output_1_356));
wire output_3_356, output_3_0, output_2_356;
mixer gate_output_2_356(.a(output_3_356), .b(output_3_0), .y(output_2_356));
wire output_1_357, output_1_1, output_0_357;
mixer gate_output_0_357(.a(output_1_357), .b(output_1_1), .y(output_0_357));
wire output_2_357, output_2_1, output_1_357;
mixer gate_output_1_357(.a(output_2_357), .b(output_2_1), .y(output_1_357));
wire output_3_357, output_3_1, output_2_357;
mixer gate_output_2_357(.a(output_3_357), .b(output_3_1), .y(output_2_357));
wire output_1_358, output_1_2, output_0_358;
mixer gate_output_0_358(.a(output_1_358), .b(output_1_2), .y(output_0_358));
wire output_2_358, output_2_2, output_1_358;
mixer gate_output_1_358(.a(output_2_358), .b(output_2_2), .y(output_1_358));
wire output_3_358, output_3_2, output_2_358;
mixer gate_output_2_358(.a(output_3_358), .b(output_3_2), .y(output_2_358));
wire output_1_359, output_1_0, output_0_359;
mixer gate_output_0_359(.a(output_1_359), .b(output_1_0), .y(output_0_359));
wire output_2_359, output_2_0, output_1_359;
mixer gate_output_1_359(.a(output_2_359), .b(output_2_0), .y(output_1_359));
wire output_3_359, output_3_0, output_2_359;
mixer gate_output_2_359(.a(output_3_359), .b(output_3_0), .y(output_2_359));
wire output_1_360, output_1_1, output_0_360;
mixer gate_output_0_360(.a(output_1_360), .b(output_1_1), .y(output_0_360));
wire output_2_360, output_2_1, output_1_360;
mixer gate_output_1_360(.a(output_2_360), .b(output_2_1), .y(output_1_360));
wire output_3_360, output_3_1, output_2_360;
mixer gate_output_2_360(.a(output_3_360), .b(output_3_1), .y(output_2_360));
wire output_1_361, output_1_2, output_0_361;
mixer gate_output_0_361(.a(output_1_361), .b(output_1_2), .y(output_0_361));
wire output_2_361, output_2_2, output_1_361;
mixer gate_output_1_361(.a(output_2_361), .b(output_2_2), .y(output_1_361));
wire output_3_361, output_3_2, output_2_361;
mixer gate_output_2_361(.a(output_3_361), .b(output_3_2), .y(output_2_361));
wire output_1_362, output_1_0, output_0_362;
mixer gate_output_0_362(.a(output_1_362), .b(output_1_0), .y(output_0_362));
wire output_2_362, output_2_0, output_1_362;
mixer gate_output_1_362(.a(output_2_362), .b(output_2_0), .y(output_1_362));
wire output_3_362, output_3_0, output_2_362;
mixer gate_output_2_362(.a(output_3_362), .b(output_3_0), .y(output_2_362));
wire output_1_363, output_1_1, output_0_363;
mixer gate_output_0_363(.a(output_1_363), .b(output_1_1), .y(output_0_363));
wire output_2_363, output_2_1, output_1_363;
mixer gate_output_1_363(.a(output_2_363), .b(output_2_1), .y(output_1_363));
wire output_3_363, output_3_1, output_2_363;
mixer gate_output_2_363(.a(output_3_363), .b(output_3_1), .y(output_2_363));
wire output_1_364, output_1_2, output_0_364;
mixer gate_output_0_364(.a(output_1_364), .b(output_1_2), .y(output_0_364));
wire output_2_364, output_2_2, output_1_364;
mixer gate_output_1_364(.a(output_2_364), .b(output_2_2), .y(output_1_364));
wire output_3_364, output_3_2, output_2_364;
mixer gate_output_2_364(.a(output_3_364), .b(output_3_2), .y(output_2_364));
wire output_1_365, output_1_0, output_0_365;
mixer gate_output_0_365(.a(output_1_365), .b(output_1_0), .y(output_0_365));
wire output_2_365, output_2_0, output_1_365;
mixer gate_output_1_365(.a(output_2_365), .b(output_2_0), .y(output_1_365));
wire output_3_365, output_3_0, output_2_365;
mixer gate_output_2_365(.a(output_3_365), .b(output_3_0), .y(output_2_365));
wire output_1_366, output_1_1, output_0_366;
mixer gate_output_0_366(.a(output_1_366), .b(output_1_1), .y(output_0_366));
wire output_2_366, output_2_1, output_1_366;
mixer gate_output_1_366(.a(output_2_366), .b(output_2_1), .y(output_1_366));
wire output_3_366, output_3_1, output_2_366;
mixer gate_output_2_366(.a(output_3_366), .b(output_3_1), .y(output_2_366));
wire output_1_367, output_1_2, output_0_367;
mixer gate_output_0_367(.a(output_1_367), .b(output_1_2), .y(output_0_367));
wire output_2_367, output_2_2, output_1_367;
mixer gate_output_1_367(.a(output_2_367), .b(output_2_2), .y(output_1_367));
wire output_3_367, output_3_2, output_2_367;
mixer gate_output_2_367(.a(output_3_367), .b(output_3_2), .y(output_2_367));
wire output_1_368, output_1_0, output_0_368;
mixer gate_output_0_368(.a(output_1_368), .b(output_1_0), .y(output_0_368));
wire output_2_368, output_2_0, output_1_368;
mixer gate_output_1_368(.a(output_2_368), .b(output_2_0), .y(output_1_368));
wire output_3_368, output_3_0, output_2_368;
mixer gate_output_2_368(.a(output_3_368), .b(output_3_0), .y(output_2_368));
wire output_1_369, output_1_1, output_0_369;
mixer gate_output_0_369(.a(output_1_369), .b(output_1_1), .y(output_0_369));
wire output_2_369, output_2_1, output_1_369;
mixer gate_output_1_369(.a(output_2_369), .b(output_2_1), .y(output_1_369));
wire output_3_369, output_3_1, output_2_369;
mixer gate_output_2_369(.a(output_3_369), .b(output_3_1), .y(output_2_369));
wire output_1_370, output_1_2, output_0_370;
mixer gate_output_0_370(.a(output_1_370), .b(output_1_2), .y(output_0_370));
wire output_2_370, output_2_2, output_1_370;
mixer gate_output_1_370(.a(output_2_370), .b(output_2_2), .y(output_1_370));
wire output_3_370, output_3_2, output_2_370;
mixer gate_output_2_370(.a(output_3_370), .b(output_3_2), .y(output_2_370));
wire output_1_371, output_1_0, output_0_371;
mixer gate_output_0_371(.a(output_1_371), .b(output_1_0), .y(output_0_371));
wire output_2_371, output_2_0, output_1_371;
mixer gate_output_1_371(.a(output_2_371), .b(output_2_0), .y(output_1_371));
wire output_3_371, output_3_0, output_2_371;
mixer gate_output_2_371(.a(output_3_371), .b(output_3_0), .y(output_2_371));
wire output_1_372, output_1_1, output_0_372;
mixer gate_output_0_372(.a(output_1_372), .b(output_1_1), .y(output_0_372));
wire output_2_372, output_2_1, output_1_372;
mixer gate_output_1_372(.a(output_2_372), .b(output_2_1), .y(output_1_372));
wire output_3_372, output_3_1, output_2_372;
mixer gate_output_2_372(.a(output_3_372), .b(output_3_1), .y(output_2_372));
wire output_1_373, output_1_2, output_0_373;
mixer gate_output_0_373(.a(output_1_373), .b(output_1_2), .y(output_0_373));
wire output_2_373, output_2_2, output_1_373;
mixer gate_output_1_373(.a(output_2_373), .b(output_2_2), .y(output_1_373));
wire output_3_373, output_3_2, output_2_373;
mixer gate_output_2_373(.a(output_3_373), .b(output_3_2), .y(output_2_373));
wire output_1_374, output_1_0, output_0_374;
mixer gate_output_0_374(.a(output_1_374), .b(output_1_0), .y(output_0_374));
wire output_2_374, output_2_0, output_1_374;
mixer gate_output_1_374(.a(output_2_374), .b(output_2_0), .y(output_1_374));
wire output_3_374, output_3_0, output_2_374;
mixer gate_output_2_374(.a(output_3_374), .b(output_3_0), .y(output_2_374));
wire output_1_375, output_1_1, output_0_375;
mixer gate_output_0_375(.a(output_1_375), .b(output_1_1), .y(output_0_375));
wire output_2_375, output_2_1, output_1_375;
mixer gate_output_1_375(.a(output_2_375), .b(output_2_1), .y(output_1_375));
wire output_3_375, output_3_1, output_2_375;
mixer gate_output_2_375(.a(output_3_375), .b(output_3_1), .y(output_2_375));
wire output_1_376, output_1_2, output_0_376;
mixer gate_output_0_376(.a(output_1_376), .b(output_1_2), .y(output_0_376));
wire output_2_376, output_2_2, output_1_376;
mixer gate_output_1_376(.a(output_2_376), .b(output_2_2), .y(output_1_376));
wire output_3_376, output_3_2, output_2_376;
mixer gate_output_2_376(.a(output_3_376), .b(output_3_2), .y(output_2_376));
wire output_1_377, output_1_0, output_0_377;
mixer gate_output_0_377(.a(output_1_377), .b(output_1_0), .y(output_0_377));
wire output_2_377, output_2_0, output_1_377;
mixer gate_output_1_377(.a(output_2_377), .b(output_2_0), .y(output_1_377));
wire output_3_377, output_3_0, output_2_377;
mixer gate_output_2_377(.a(output_3_377), .b(output_3_0), .y(output_2_377));
wire output_1_378, output_1_1, output_0_378;
mixer gate_output_0_378(.a(output_1_378), .b(output_1_1), .y(output_0_378));
wire output_2_378, output_2_1, output_1_378;
mixer gate_output_1_378(.a(output_2_378), .b(output_2_1), .y(output_1_378));
wire output_3_378, output_3_1, output_2_378;
mixer gate_output_2_378(.a(output_3_378), .b(output_3_1), .y(output_2_378));
wire output_1_379, output_1_2, output_0_379;
mixer gate_output_0_379(.a(output_1_379), .b(output_1_2), .y(output_0_379));
wire output_2_379, output_2_2, output_1_379;
mixer gate_output_1_379(.a(output_2_379), .b(output_2_2), .y(output_1_379));
wire output_3_379, output_3_2, output_2_379;
mixer gate_output_2_379(.a(output_3_379), .b(output_3_2), .y(output_2_379));
wire output_1_380, output_1_0, output_0_380;
mixer gate_output_0_380(.a(output_1_380), .b(output_1_0), .y(output_0_380));
wire output_2_380, output_2_0, output_1_380;
mixer gate_output_1_380(.a(output_2_380), .b(output_2_0), .y(output_1_380));
wire output_3_380, output_3_0, output_2_380;
mixer gate_output_2_380(.a(output_3_380), .b(output_3_0), .y(output_2_380));
wire output_1_381, output_1_1, output_0_381;
mixer gate_output_0_381(.a(output_1_381), .b(output_1_1), .y(output_0_381));
wire output_2_381, output_2_1, output_1_381;
mixer gate_output_1_381(.a(output_2_381), .b(output_2_1), .y(output_1_381));
wire output_3_381, output_3_1, output_2_381;
mixer gate_output_2_381(.a(output_3_381), .b(output_3_1), .y(output_2_381));
wire output_1_382, output_1_2, output_0_382;
mixer gate_output_0_382(.a(output_1_382), .b(output_1_2), .y(output_0_382));
wire output_2_382, output_2_2, output_1_382;
mixer gate_output_1_382(.a(output_2_382), .b(output_2_2), .y(output_1_382));
wire output_3_382, output_3_2, output_2_382;
mixer gate_output_2_382(.a(output_3_382), .b(output_3_2), .y(output_2_382));
wire output_1_383, output_1_0, output_0_383;
mixer gate_output_0_383(.a(output_1_383), .b(output_1_0), .y(output_0_383));
wire output_2_383, output_2_0, output_1_383;
mixer gate_output_1_383(.a(output_2_383), .b(output_2_0), .y(output_1_383));
wire output_3_383, output_3_0, output_2_383;
mixer gate_output_2_383(.a(output_3_383), .b(output_3_0), .y(output_2_383));
wire output_1_384, output_1_1, output_0_384;
mixer gate_output_0_384(.a(output_1_384), .b(output_1_1), .y(output_0_384));
wire output_2_384, output_2_1, output_1_384;
mixer gate_output_1_384(.a(output_2_384), .b(output_2_1), .y(output_1_384));
wire output_3_384, output_3_1, output_2_384;
mixer gate_output_2_384(.a(output_3_384), .b(output_3_1), .y(output_2_384));
wire output_1_385, output_1_2, output_0_385;
mixer gate_output_0_385(.a(output_1_385), .b(output_1_2), .y(output_0_385));
wire output_2_385, output_2_2, output_1_385;
mixer gate_output_1_385(.a(output_2_385), .b(output_2_2), .y(output_1_385));
wire output_3_385, output_3_2, output_2_385;
mixer gate_output_2_385(.a(output_3_385), .b(output_3_2), .y(output_2_385));
wire output_1_386, output_1_0, output_0_386;
mixer gate_output_0_386(.a(output_1_386), .b(output_1_0), .y(output_0_386));
wire output_2_386, output_2_0, output_1_386;
mixer gate_output_1_386(.a(output_2_386), .b(output_2_0), .y(output_1_386));
wire output_3_386, output_3_0, output_2_386;
mixer gate_output_2_386(.a(output_3_386), .b(output_3_0), .y(output_2_386));
wire output_1_387, output_1_1, output_0_387;
mixer gate_output_0_387(.a(output_1_387), .b(output_1_1), .y(output_0_387));
wire output_2_387, output_2_1, output_1_387;
mixer gate_output_1_387(.a(output_2_387), .b(output_2_1), .y(output_1_387));
wire output_3_387, output_3_1, output_2_387;
mixer gate_output_2_387(.a(output_3_387), .b(output_3_1), .y(output_2_387));
wire output_1_388, output_1_2, output_0_388;
mixer gate_output_0_388(.a(output_1_388), .b(output_1_2), .y(output_0_388));
wire output_2_388, output_2_2, output_1_388;
mixer gate_output_1_388(.a(output_2_388), .b(output_2_2), .y(output_1_388));
wire output_3_388, output_3_2, output_2_388;
mixer gate_output_2_388(.a(output_3_388), .b(output_3_2), .y(output_2_388));
wire output_1_389, output_1_0, output_0_389;
mixer gate_output_0_389(.a(output_1_389), .b(output_1_0), .y(output_0_389));
wire output_2_389, output_2_0, output_1_389;
mixer gate_output_1_389(.a(output_2_389), .b(output_2_0), .y(output_1_389));
wire output_3_389, output_3_0, output_2_389;
mixer gate_output_2_389(.a(output_3_389), .b(output_3_0), .y(output_2_389));
wire output_1_390, output_1_1, output_0_390;
mixer gate_output_0_390(.a(output_1_390), .b(output_1_1), .y(output_0_390));
wire output_2_390, output_2_1, output_1_390;
mixer gate_output_1_390(.a(output_2_390), .b(output_2_1), .y(output_1_390));
wire output_3_390, output_3_1, output_2_390;
mixer gate_output_2_390(.a(output_3_390), .b(output_3_1), .y(output_2_390));
wire output_1_391, output_1_2, output_0_391;
mixer gate_output_0_391(.a(output_1_391), .b(output_1_2), .y(output_0_391));
wire output_2_391, output_2_2, output_1_391;
mixer gate_output_1_391(.a(output_2_391), .b(output_2_2), .y(output_1_391));
wire output_3_391, output_3_2, output_2_391;
mixer gate_output_2_391(.a(output_3_391), .b(output_3_2), .y(output_2_391));
wire output_1_392, output_1_0, output_0_392;
mixer gate_output_0_392(.a(output_1_392), .b(output_1_0), .y(output_0_392));
wire output_2_392, output_2_0, output_1_392;
mixer gate_output_1_392(.a(output_2_392), .b(output_2_0), .y(output_1_392));
wire output_3_392, output_3_0, output_2_392;
mixer gate_output_2_392(.a(output_3_392), .b(output_3_0), .y(output_2_392));
wire output_1_393, output_1_1, output_0_393;
mixer gate_output_0_393(.a(output_1_393), .b(output_1_1), .y(output_0_393));
wire output_2_393, output_2_1, output_1_393;
mixer gate_output_1_393(.a(output_2_393), .b(output_2_1), .y(output_1_393));
wire output_3_393, output_3_1, output_2_393;
mixer gate_output_2_393(.a(output_3_393), .b(output_3_1), .y(output_2_393));
wire output_1_394, output_1_2, output_0_394;
mixer gate_output_0_394(.a(output_1_394), .b(output_1_2), .y(output_0_394));
wire output_2_394, output_2_2, output_1_394;
mixer gate_output_1_394(.a(output_2_394), .b(output_2_2), .y(output_1_394));
wire output_3_394, output_3_2, output_2_394;
mixer gate_output_2_394(.a(output_3_394), .b(output_3_2), .y(output_2_394));
wire output_1_395, output_1_0, output_0_395;
mixer gate_output_0_395(.a(output_1_395), .b(output_1_0), .y(output_0_395));
wire output_2_395, output_2_0, output_1_395;
mixer gate_output_1_395(.a(output_2_395), .b(output_2_0), .y(output_1_395));
wire output_3_395, output_3_0, output_2_395;
mixer gate_output_2_395(.a(output_3_395), .b(output_3_0), .y(output_2_395));
wire output_1_396, output_1_1, output_0_396;
mixer gate_output_0_396(.a(output_1_396), .b(output_1_1), .y(output_0_396));
wire output_2_396, output_2_1, output_1_396;
mixer gate_output_1_396(.a(output_2_396), .b(output_2_1), .y(output_1_396));
wire output_3_396, output_3_1, output_2_396;
mixer gate_output_2_396(.a(output_3_396), .b(output_3_1), .y(output_2_396));
wire output_1_397, output_1_2, output_0_397;
mixer gate_output_0_397(.a(output_1_397), .b(output_1_2), .y(output_0_397));
wire output_2_397, output_2_2, output_1_397;
mixer gate_output_1_397(.a(output_2_397), .b(output_2_2), .y(output_1_397));
wire output_3_397, output_3_2, output_2_397;
mixer gate_output_2_397(.a(output_3_397), .b(output_3_2), .y(output_2_397));
wire output_1_398, output_1_0, output_0_398;
mixer gate_output_0_398(.a(output_1_398), .b(output_1_0), .y(output_0_398));
wire output_2_398, output_2_0, output_1_398;
mixer gate_output_1_398(.a(output_2_398), .b(output_2_0), .y(output_1_398));
wire output_3_398, output_3_0, output_2_398;
mixer gate_output_2_398(.a(output_3_398), .b(output_3_0), .y(output_2_398));
wire output_1_399, output_1_1, output_0_399;
mixer gate_output_0_399(.a(output_1_399), .b(output_1_1), .y(output_0_399));
wire output_2_399, output_2_1, output_1_399;
mixer gate_output_1_399(.a(output_2_399), .b(output_2_1), .y(output_1_399));
wire output_3_399, output_3_1, output_2_399;
mixer gate_output_2_399(.a(output_3_399), .b(output_3_1), .y(output_2_399));
wire output_1_400, output_1_2, output_0_400;
mixer gate_output_0_400(.a(output_1_400), .b(output_1_2), .y(output_0_400));
wire output_2_400, output_2_2, output_1_400;
mixer gate_output_1_400(.a(output_2_400), .b(output_2_2), .y(output_1_400));
wire output_3_400, output_3_2, output_2_400;
mixer gate_output_2_400(.a(output_3_400), .b(output_3_2), .y(output_2_400));
wire output_1_401, output_1_0, output_0_401;
mixer gate_output_0_401(.a(output_1_401), .b(output_1_0), .y(output_0_401));
wire output_2_401, output_2_0, output_1_401;
mixer gate_output_1_401(.a(output_2_401), .b(output_2_0), .y(output_1_401));
wire output_3_401, output_3_0, output_2_401;
mixer gate_output_2_401(.a(output_3_401), .b(output_3_0), .y(output_2_401));
wire output_1_402, output_1_1, output_0_402;
mixer gate_output_0_402(.a(output_1_402), .b(output_1_1), .y(output_0_402));
wire output_2_402, output_2_1, output_1_402;
mixer gate_output_1_402(.a(output_2_402), .b(output_2_1), .y(output_1_402));
wire output_3_402, output_3_1, output_2_402;
mixer gate_output_2_402(.a(output_3_402), .b(output_3_1), .y(output_2_402));
wire output_1_403, output_1_2, output_0_403;
mixer gate_output_0_403(.a(output_1_403), .b(output_1_2), .y(output_0_403));
wire output_2_403, output_2_2, output_1_403;
mixer gate_output_1_403(.a(output_2_403), .b(output_2_2), .y(output_1_403));
wire output_3_403, output_3_2, output_2_403;
mixer gate_output_2_403(.a(output_3_403), .b(output_3_2), .y(output_2_403));
wire output_1_404, output_1_0, output_0_404;
mixer gate_output_0_404(.a(output_1_404), .b(output_1_0), .y(output_0_404));
wire output_2_404, output_2_0, output_1_404;
mixer gate_output_1_404(.a(output_2_404), .b(output_2_0), .y(output_1_404));
wire output_3_404, output_3_0, output_2_404;
mixer gate_output_2_404(.a(output_3_404), .b(output_3_0), .y(output_2_404));
wire output_1_405, output_1_1, output_0_405;
mixer gate_output_0_405(.a(output_1_405), .b(output_1_1), .y(output_0_405));
wire output_2_405, output_2_1, output_1_405;
mixer gate_output_1_405(.a(output_2_405), .b(output_2_1), .y(output_1_405));
wire output_3_405, output_3_1, output_2_405;
mixer gate_output_2_405(.a(output_3_405), .b(output_3_1), .y(output_2_405));
wire output_1_406, output_1_2, output_0_406;
mixer gate_output_0_406(.a(output_1_406), .b(output_1_2), .y(output_0_406));
wire output_2_406, output_2_2, output_1_406;
mixer gate_output_1_406(.a(output_2_406), .b(output_2_2), .y(output_1_406));
wire output_3_406, output_3_2, output_2_406;
mixer gate_output_2_406(.a(output_3_406), .b(output_3_2), .y(output_2_406));
wire output_1_407, output_1_0, output_0_407;
mixer gate_output_0_407(.a(output_1_407), .b(output_1_0), .y(output_0_407));
wire output_2_407, output_2_0, output_1_407;
mixer gate_output_1_407(.a(output_2_407), .b(output_2_0), .y(output_1_407));
wire output_3_407, output_3_0, output_2_407;
mixer gate_output_2_407(.a(output_3_407), .b(output_3_0), .y(output_2_407));
wire output_1_408, output_1_1, output_0_408;
mixer gate_output_0_408(.a(output_1_408), .b(output_1_1), .y(output_0_408));
wire output_2_408, output_2_1, output_1_408;
mixer gate_output_1_408(.a(output_2_408), .b(output_2_1), .y(output_1_408));
wire output_3_408, output_3_1, output_2_408;
mixer gate_output_2_408(.a(output_3_408), .b(output_3_1), .y(output_2_408));
wire output_1_409, output_1_2, output_0_409;
mixer gate_output_0_409(.a(output_1_409), .b(output_1_2), .y(output_0_409));
wire output_2_409, output_2_2, output_1_409;
mixer gate_output_1_409(.a(output_2_409), .b(output_2_2), .y(output_1_409));
wire output_3_409, output_3_2, output_2_409;
mixer gate_output_2_409(.a(output_3_409), .b(output_3_2), .y(output_2_409));
wire output_1_410, output_1_0, output_0_410;
mixer gate_output_0_410(.a(output_1_410), .b(output_1_0), .y(output_0_410));
wire output_2_410, output_2_0, output_1_410;
mixer gate_output_1_410(.a(output_2_410), .b(output_2_0), .y(output_1_410));
wire output_3_410, output_3_0, output_2_410;
mixer gate_output_2_410(.a(output_3_410), .b(output_3_0), .y(output_2_410));
wire output_1_411, output_1_1, output_0_411;
mixer gate_output_0_411(.a(output_1_411), .b(output_1_1), .y(output_0_411));
wire output_2_411, output_2_1, output_1_411;
mixer gate_output_1_411(.a(output_2_411), .b(output_2_1), .y(output_1_411));
wire output_3_411, output_3_1, output_2_411;
mixer gate_output_2_411(.a(output_3_411), .b(output_3_1), .y(output_2_411));
wire output_1_412, output_1_2, output_0_412;
mixer gate_output_0_412(.a(output_1_412), .b(output_1_2), .y(output_0_412));
wire output_2_412, output_2_2, output_1_412;
mixer gate_output_1_412(.a(output_2_412), .b(output_2_2), .y(output_1_412));
wire output_3_412, output_3_2, output_2_412;
mixer gate_output_2_412(.a(output_3_412), .b(output_3_2), .y(output_2_412));
wire output_1_413, output_1_0, output_0_413;
mixer gate_output_0_413(.a(output_1_413), .b(output_1_0), .y(output_0_413));
wire output_2_413, output_2_0, output_1_413;
mixer gate_output_1_413(.a(output_2_413), .b(output_2_0), .y(output_1_413));
wire output_3_413, output_3_0, output_2_413;
mixer gate_output_2_413(.a(output_3_413), .b(output_3_0), .y(output_2_413));
wire output_1_414, output_1_1, output_0_414;
mixer gate_output_0_414(.a(output_1_414), .b(output_1_1), .y(output_0_414));
wire output_2_414, output_2_1, output_1_414;
mixer gate_output_1_414(.a(output_2_414), .b(output_2_1), .y(output_1_414));
wire output_3_414, output_3_1, output_2_414;
mixer gate_output_2_414(.a(output_3_414), .b(output_3_1), .y(output_2_414));
wire output_1_415, output_1_2, output_0_415;
mixer gate_output_0_415(.a(output_1_415), .b(output_1_2), .y(output_0_415));
wire output_2_415, output_2_2, output_1_415;
mixer gate_output_1_415(.a(output_2_415), .b(output_2_2), .y(output_1_415));
wire output_3_415, output_3_2, output_2_415;
mixer gate_output_2_415(.a(output_3_415), .b(output_3_2), .y(output_2_415));
wire output_1_416, output_1_0, output_0_416;
mixer gate_output_0_416(.a(output_1_416), .b(output_1_0), .y(output_0_416));
wire output_2_416, output_2_0, output_1_416;
mixer gate_output_1_416(.a(output_2_416), .b(output_2_0), .y(output_1_416));
wire output_3_416, output_3_0, output_2_416;
mixer gate_output_2_416(.a(output_3_416), .b(output_3_0), .y(output_2_416));
wire output_1_417, output_1_1, output_0_417;
mixer gate_output_0_417(.a(output_1_417), .b(output_1_1), .y(output_0_417));
wire output_2_417, output_2_1, output_1_417;
mixer gate_output_1_417(.a(output_2_417), .b(output_2_1), .y(output_1_417));
wire output_3_417, output_3_1, output_2_417;
mixer gate_output_2_417(.a(output_3_417), .b(output_3_1), .y(output_2_417));
wire output_1_418, output_1_2, output_0_418;
mixer gate_output_0_418(.a(output_1_418), .b(output_1_2), .y(output_0_418));
wire output_2_418, output_2_2, output_1_418;
mixer gate_output_1_418(.a(output_2_418), .b(output_2_2), .y(output_1_418));
wire output_3_418, output_3_2, output_2_418;
mixer gate_output_2_418(.a(output_3_418), .b(output_3_2), .y(output_2_418));
wire output_1_419, output_1_0, output_0_419;
mixer gate_output_0_419(.a(output_1_419), .b(output_1_0), .y(output_0_419));
wire output_2_419, output_2_0, output_1_419;
mixer gate_output_1_419(.a(output_2_419), .b(output_2_0), .y(output_1_419));
wire output_3_419, output_3_0, output_2_419;
mixer gate_output_2_419(.a(output_3_419), .b(output_3_0), .y(output_2_419));
wire output_1_420, output_1_1, output_0_420;
mixer gate_output_0_420(.a(output_1_420), .b(output_1_1), .y(output_0_420));
wire output_2_420, output_2_1, output_1_420;
mixer gate_output_1_420(.a(output_2_420), .b(output_2_1), .y(output_1_420));
wire output_3_420, output_3_1, output_2_420;
mixer gate_output_2_420(.a(output_3_420), .b(output_3_1), .y(output_2_420));
wire output_1_421, output_1_2, output_0_421;
mixer gate_output_0_421(.a(output_1_421), .b(output_1_2), .y(output_0_421));
wire output_2_421, output_2_2, output_1_421;
mixer gate_output_1_421(.a(output_2_421), .b(output_2_2), .y(output_1_421));
wire output_3_421, output_3_2, output_2_421;
mixer gate_output_2_421(.a(output_3_421), .b(output_3_2), .y(output_2_421));
wire output_1_422, output_1_0, output_0_422;
mixer gate_output_0_422(.a(output_1_422), .b(output_1_0), .y(output_0_422));
wire output_2_422, output_2_0, output_1_422;
mixer gate_output_1_422(.a(output_2_422), .b(output_2_0), .y(output_1_422));
wire output_3_422, output_3_0, output_2_422;
mixer gate_output_2_422(.a(output_3_422), .b(output_3_0), .y(output_2_422));
wire output_1_423, output_1_1, output_0_423;
mixer gate_output_0_423(.a(output_1_423), .b(output_1_1), .y(output_0_423));
wire output_2_423, output_2_1, output_1_423;
mixer gate_output_1_423(.a(output_2_423), .b(output_2_1), .y(output_1_423));
wire output_3_423, output_3_1, output_2_423;
mixer gate_output_2_423(.a(output_3_423), .b(output_3_1), .y(output_2_423));
wire output_1_424, output_1_2, output_0_424;
mixer gate_output_0_424(.a(output_1_424), .b(output_1_2), .y(output_0_424));
wire output_2_424, output_2_2, output_1_424;
mixer gate_output_1_424(.a(output_2_424), .b(output_2_2), .y(output_1_424));
wire output_3_424, output_3_2, output_2_424;
mixer gate_output_2_424(.a(output_3_424), .b(output_3_2), .y(output_2_424));
wire output_1_425, output_1_0, output_0_425;
mixer gate_output_0_425(.a(output_1_425), .b(output_1_0), .y(output_0_425));
wire output_2_425, output_2_0, output_1_425;
mixer gate_output_1_425(.a(output_2_425), .b(output_2_0), .y(output_1_425));
wire output_3_425, output_3_0, output_2_425;
mixer gate_output_2_425(.a(output_3_425), .b(output_3_0), .y(output_2_425));
wire output_1_426, output_1_1, output_0_426;
mixer gate_output_0_426(.a(output_1_426), .b(output_1_1), .y(output_0_426));
wire output_2_426, output_2_1, output_1_426;
mixer gate_output_1_426(.a(output_2_426), .b(output_2_1), .y(output_1_426));
wire output_3_426, output_3_1, output_2_426;
mixer gate_output_2_426(.a(output_3_426), .b(output_3_1), .y(output_2_426));
wire output_1_427, output_1_2, output_0_427;
mixer gate_output_0_427(.a(output_1_427), .b(output_1_2), .y(output_0_427));
wire output_2_427, output_2_2, output_1_427;
mixer gate_output_1_427(.a(output_2_427), .b(output_2_2), .y(output_1_427));
wire output_3_427, output_3_2, output_2_427;
mixer gate_output_2_427(.a(output_3_427), .b(output_3_2), .y(output_2_427));
wire output_1_428, output_1_0, output_0_428;
mixer gate_output_0_428(.a(output_1_428), .b(output_1_0), .y(output_0_428));
wire output_2_428, output_2_0, output_1_428;
mixer gate_output_1_428(.a(output_2_428), .b(output_2_0), .y(output_1_428));
wire output_3_428, output_3_0, output_2_428;
mixer gate_output_2_428(.a(output_3_428), .b(output_3_0), .y(output_2_428));
wire output_1_429, output_1_1, output_0_429;
mixer gate_output_0_429(.a(output_1_429), .b(output_1_1), .y(output_0_429));
wire output_2_429, output_2_1, output_1_429;
mixer gate_output_1_429(.a(output_2_429), .b(output_2_1), .y(output_1_429));
wire output_3_429, output_3_1, output_2_429;
mixer gate_output_2_429(.a(output_3_429), .b(output_3_1), .y(output_2_429));
wire output_1_430, output_1_2, output_0_430;
mixer gate_output_0_430(.a(output_1_430), .b(output_1_2), .y(output_0_430));
wire output_2_430, output_2_2, output_1_430;
mixer gate_output_1_430(.a(output_2_430), .b(output_2_2), .y(output_1_430));
wire output_3_430, output_3_2, output_2_430;
mixer gate_output_2_430(.a(output_3_430), .b(output_3_2), .y(output_2_430));
wire output_1_431, output_1_0, output_0_431;
mixer gate_output_0_431(.a(output_1_431), .b(output_1_0), .y(output_0_431));
wire output_2_431, output_2_0, output_1_431;
mixer gate_output_1_431(.a(output_2_431), .b(output_2_0), .y(output_1_431));
wire output_3_431, output_3_0, output_2_431;
mixer gate_output_2_431(.a(output_3_431), .b(output_3_0), .y(output_2_431));
wire output_1_432, output_1_1, output_0_432;
mixer gate_output_0_432(.a(output_1_432), .b(output_1_1), .y(output_0_432));
wire output_2_432, output_2_1, output_1_432;
mixer gate_output_1_432(.a(output_2_432), .b(output_2_1), .y(output_1_432));
wire output_3_432, output_3_1, output_2_432;
mixer gate_output_2_432(.a(output_3_432), .b(output_3_1), .y(output_2_432));
wire output_1_433, output_1_2, output_0_433;
mixer gate_output_0_433(.a(output_1_433), .b(output_1_2), .y(output_0_433));
wire output_2_433, output_2_2, output_1_433;
mixer gate_output_1_433(.a(output_2_433), .b(output_2_2), .y(output_1_433));
wire output_3_433, output_3_2, output_2_433;
mixer gate_output_2_433(.a(output_3_433), .b(output_3_2), .y(output_2_433));
wire output_1_434, output_1_0, output_0_434;
mixer gate_output_0_434(.a(output_1_434), .b(output_1_0), .y(output_0_434));
wire output_2_434, output_2_0, output_1_434;
mixer gate_output_1_434(.a(output_2_434), .b(output_2_0), .y(output_1_434));
wire output_3_434, output_3_0, output_2_434;
mixer gate_output_2_434(.a(output_3_434), .b(output_3_0), .y(output_2_434));
wire output_1_435, output_1_1, output_0_435;
mixer gate_output_0_435(.a(output_1_435), .b(output_1_1), .y(output_0_435));
wire output_2_435, output_2_1, output_1_435;
mixer gate_output_1_435(.a(output_2_435), .b(output_2_1), .y(output_1_435));
wire output_3_435, output_3_1, output_2_435;
mixer gate_output_2_435(.a(output_3_435), .b(output_3_1), .y(output_2_435));
wire output_1_436, output_1_2, output_0_436;
mixer gate_output_0_436(.a(output_1_436), .b(output_1_2), .y(output_0_436));
wire output_2_436, output_2_2, output_1_436;
mixer gate_output_1_436(.a(output_2_436), .b(output_2_2), .y(output_1_436));
wire output_3_436, output_3_2, output_2_436;
mixer gate_output_2_436(.a(output_3_436), .b(output_3_2), .y(output_2_436));
wire output_1_437, output_1_0, output_0_437;
mixer gate_output_0_437(.a(output_1_437), .b(output_1_0), .y(output_0_437));
wire output_2_437, output_2_0, output_1_437;
mixer gate_output_1_437(.a(output_2_437), .b(output_2_0), .y(output_1_437));
wire output_3_437, output_3_0, output_2_437;
mixer gate_output_2_437(.a(output_3_437), .b(output_3_0), .y(output_2_437));
wire output_1_438, output_1_1, output_0_438;
mixer gate_output_0_438(.a(output_1_438), .b(output_1_1), .y(output_0_438));
wire output_2_438, output_2_1, output_1_438;
mixer gate_output_1_438(.a(output_2_438), .b(output_2_1), .y(output_1_438));
wire output_3_438, output_3_1, output_2_438;
mixer gate_output_2_438(.a(output_3_438), .b(output_3_1), .y(output_2_438));
wire output_1_439, output_1_2, output_0_439;
mixer gate_output_0_439(.a(output_1_439), .b(output_1_2), .y(output_0_439));
wire output_2_439, output_2_2, output_1_439;
mixer gate_output_1_439(.a(output_2_439), .b(output_2_2), .y(output_1_439));
wire output_3_439, output_3_2, output_2_439;
mixer gate_output_2_439(.a(output_3_439), .b(output_3_2), .y(output_2_439));
wire output_1_440, output_1_0, output_0_440;
mixer gate_output_0_440(.a(output_1_440), .b(output_1_0), .y(output_0_440));
wire output_2_440, output_2_0, output_1_440;
mixer gate_output_1_440(.a(output_2_440), .b(output_2_0), .y(output_1_440));
wire output_3_440, output_3_0, output_2_440;
mixer gate_output_2_440(.a(output_3_440), .b(output_3_0), .y(output_2_440));
wire output_1_441, output_1_1, output_0_441;
mixer gate_output_0_441(.a(output_1_441), .b(output_1_1), .y(output_0_441));
wire output_2_441, output_2_1, output_1_441;
mixer gate_output_1_441(.a(output_2_441), .b(output_2_1), .y(output_1_441));
wire output_3_441, output_3_1, output_2_441;
mixer gate_output_2_441(.a(output_3_441), .b(output_3_1), .y(output_2_441));
wire output_1_442, output_1_2, output_0_442;
mixer gate_output_0_442(.a(output_1_442), .b(output_1_2), .y(output_0_442));
wire output_2_442, output_2_2, output_1_442;
mixer gate_output_1_442(.a(output_2_442), .b(output_2_2), .y(output_1_442));
wire output_3_442, output_3_2, output_2_442;
mixer gate_output_2_442(.a(output_3_442), .b(output_3_2), .y(output_2_442));
wire output_1_443, output_1_0, output_0_443;
mixer gate_output_0_443(.a(output_1_443), .b(output_1_0), .y(output_0_443));
wire output_2_443, output_2_0, output_1_443;
mixer gate_output_1_443(.a(output_2_443), .b(output_2_0), .y(output_1_443));
wire output_3_443, output_3_0, output_2_443;
mixer gate_output_2_443(.a(output_3_443), .b(output_3_0), .y(output_2_443));
wire output_1_444, output_1_1, output_0_444;
mixer gate_output_0_444(.a(output_1_444), .b(output_1_1), .y(output_0_444));
wire output_2_444, output_2_1, output_1_444;
mixer gate_output_1_444(.a(output_2_444), .b(output_2_1), .y(output_1_444));
wire output_3_444, output_3_1, output_2_444;
mixer gate_output_2_444(.a(output_3_444), .b(output_3_1), .y(output_2_444));
wire output_1_445, output_1_2, output_0_445;
mixer gate_output_0_445(.a(output_1_445), .b(output_1_2), .y(output_0_445));
wire output_2_445, output_2_2, output_1_445;
mixer gate_output_1_445(.a(output_2_445), .b(output_2_2), .y(output_1_445));
wire output_3_445, output_3_2, output_2_445;
mixer gate_output_2_445(.a(output_3_445), .b(output_3_2), .y(output_2_445));
wire output_1_446, output_1_0, output_0_446;
mixer gate_output_0_446(.a(output_1_446), .b(output_1_0), .y(output_0_446));
wire output_2_446, output_2_0, output_1_446;
mixer gate_output_1_446(.a(output_2_446), .b(output_2_0), .y(output_1_446));
wire output_3_446, output_3_0, output_2_446;
mixer gate_output_2_446(.a(output_3_446), .b(output_3_0), .y(output_2_446));
wire output_1_447, output_1_1, output_0_447;
mixer gate_output_0_447(.a(output_1_447), .b(output_1_1), .y(output_0_447));
wire output_2_447, output_2_1, output_1_447;
mixer gate_output_1_447(.a(output_2_447), .b(output_2_1), .y(output_1_447));
wire output_3_447, output_3_1, output_2_447;
mixer gate_output_2_447(.a(output_3_447), .b(output_3_1), .y(output_2_447));
wire output_1_448, output_1_2, output_0_448;
mixer gate_output_0_448(.a(output_1_448), .b(output_1_2), .y(output_0_448));
wire output_2_448, output_2_2, output_1_448;
mixer gate_output_1_448(.a(output_2_448), .b(output_2_2), .y(output_1_448));
wire output_3_448, output_3_2, output_2_448;
mixer gate_output_2_448(.a(output_3_448), .b(output_3_2), .y(output_2_448));
wire output_1_449, output_1_0, output_0_449;
mixer gate_output_0_449(.a(output_1_449), .b(output_1_0), .y(output_0_449));
wire output_2_449, output_2_0, output_1_449;
mixer gate_output_1_449(.a(output_2_449), .b(output_2_0), .y(output_1_449));
wire output_3_449, output_3_0, output_2_449;
mixer gate_output_2_449(.a(output_3_449), .b(output_3_0), .y(output_2_449));
wire output_1_450, output_1_1, output_0_450;
mixer gate_output_0_450(.a(output_1_450), .b(output_1_1), .y(output_0_450));
wire output_2_450, output_2_1, output_1_450;
mixer gate_output_1_450(.a(output_2_450), .b(output_2_1), .y(output_1_450));
wire output_3_450, output_3_1, output_2_450;
mixer gate_output_2_450(.a(output_3_450), .b(output_3_1), .y(output_2_450));
wire output_1_451, output_1_2, output_0_451;
mixer gate_output_0_451(.a(output_1_451), .b(output_1_2), .y(output_0_451));
wire output_2_451, output_2_2, output_1_451;
mixer gate_output_1_451(.a(output_2_451), .b(output_2_2), .y(output_1_451));
wire output_3_451, output_3_2, output_2_451;
mixer gate_output_2_451(.a(output_3_451), .b(output_3_2), .y(output_2_451));
wire output_1_452, output_1_0, output_0_452;
mixer gate_output_0_452(.a(output_1_452), .b(output_1_0), .y(output_0_452));
wire output_2_452, output_2_0, output_1_452;
mixer gate_output_1_452(.a(output_2_452), .b(output_2_0), .y(output_1_452));
wire output_3_452, output_3_0, output_2_452;
mixer gate_output_2_452(.a(output_3_452), .b(output_3_0), .y(output_2_452));
wire output_1_453, output_1_1, output_0_453;
mixer gate_output_0_453(.a(output_1_453), .b(output_1_1), .y(output_0_453));
wire output_2_453, output_2_1, output_1_453;
mixer gate_output_1_453(.a(output_2_453), .b(output_2_1), .y(output_1_453));
wire output_3_453, output_3_1, output_2_453;
mixer gate_output_2_453(.a(output_3_453), .b(output_3_1), .y(output_2_453));
wire output_1_454, output_1_2, output_0_454;
mixer gate_output_0_454(.a(output_1_454), .b(output_1_2), .y(output_0_454));
wire output_2_454, output_2_2, output_1_454;
mixer gate_output_1_454(.a(output_2_454), .b(output_2_2), .y(output_1_454));
wire output_3_454, output_3_2, output_2_454;
mixer gate_output_2_454(.a(output_3_454), .b(output_3_2), .y(output_2_454));
wire output_1_455, output_1_0, output_0_455;
mixer gate_output_0_455(.a(output_1_455), .b(output_1_0), .y(output_0_455));
wire output_2_455, output_2_0, output_1_455;
mixer gate_output_1_455(.a(output_2_455), .b(output_2_0), .y(output_1_455));
wire output_3_455, output_3_0, output_2_455;
mixer gate_output_2_455(.a(output_3_455), .b(output_3_0), .y(output_2_455));
wire output_1_456, output_1_1, output_0_456;
mixer gate_output_0_456(.a(output_1_456), .b(output_1_1), .y(output_0_456));
wire output_2_456, output_2_1, output_1_456;
mixer gate_output_1_456(.a(output_2_456), .b(output_2_1), .y(output_1_456));
wire output_3_456, output_3_1, output_2_456;
mixer gate_output_2_456(.a(output_3_456), .b(output_3_1), .y(output_2_456));
wire output_1_457, output_1_2, output_0_457;
mixer gate_output_0_457(.a(output_1_457), .b(output_1_2), .y(output_0_457));
wire output_2_457, output_2_2, output_1_457;
mixer gate_output_1_457(.a(output_2_457), .b(output_2_2), .y(output_1_457));
wire output_3_457, output_3_2, output_2_457;
mixer gate_output_2_457(.a(output_3_457), .b(output_3_2), .y(output_2_457));
wire output_1_458, output_1_0, output_0_458;
mixer gate_output_0_458(.a(output_1_458), .b(output_1_0), .y(output_0_458));
wire output_2_458, output_2_0, output_1_458;
mixer gate_output_1_458(.a(output_2_458), .b(output_2_0), .y(output_1_458));
wire output_3_458, output_3_0, output_2_458;
mixer gate_output_2_458(.a(output_3_458), .b(output_3_0), .y(output_2_458));
wire output_1_459, output_1_1, output_0_459;
mixer gate_output_0_459(.a(output_1_459), .b(output_1_1), .y(output_0_459));
wire output_2_459, output_2_1, output_1_459;
mixer gate_output_1_459(.a(output_2_459), .b(output_2_1), .y(output_1_459));
wire output_3_459, output_3_1, output_2_459;
mixer gate_output_2_459(.a(output_3_459), .b(output_3_1), .y(output_2_459));
wire output_1_460, output_1_2, output_0_460;
mixer gate_output_0_460(.a(output_1_460), .b(output_1_2), .y(output_0_460));
wire output_2_460, output_2_2, output_1_460;
mixer gate_output_1_460(.a(output_2_460), .b(output_2_2), .y(output_1_460));
wire output_3_460, output_3_2, output_2_460;
mixer gate_output_2_460(.a(output_3_460), .b(output_3_2), .y(output_2_460));
wire output_1_461, output_1_0, output_0_461;
mixer gate_output_0_461(.a(output_1_461), .b(output_1_0), .y(output_0_461));
wire output_2_461, output_2_0, output_1_461;
mixer gate_output_1_461(.a(output_2_461), .b(output_2_0), .y(output_1_461));
wire output_3_461, output_3_0, output_2_461;
mixer gate_output_2_461(.a(output_3_461), .b(output_3_0), .y(output_2_461));
wire output_1_462, output_1_1, output_0_462;
mixer gate_output_0_462(.a(output_1_462), .b(output_1_1), .y(output_0_462));
wire output_2_462, output_2_1, output_1_462;
mixer gate_output_1_462(.a(output_2_462), .b(output_2_1), .y(output_1_462));
wire output_3_462, output_3_1, output_2_462;
mixer gate_output_2_462(.a(output_3_462), .b(output_3_1), .y(output_2_462));
wire output_1_463, output_1_2, output_0_463;
mixer gate_output_0_463(.a(output_1_463), .b(output_1_2), .y(output_0_463));
wire output_2_463, output_2_2, output_1_463;
mixer gate_output_1_463(.a(output_2_463), .b(output_2_2), .y(output_1_463));
wire output_3_463, output_3_2, output_2_463;
mixer gate_output_2_463(.a(output_3_463), .b(output_3_2), .y(output_2_463));
wire output_1_464, output_1_0, output_0_464;
mixer gate_output_0_464(.a(output_1_464), .b(output_1_0), .y(output_0_464));
wire output_2_464, output_2_0, output_1_464;
mixer gate_output_1_464(.a(output_2_464), .b(output_2_0), .y(output_1_464));
wire output_3_464, output_3_0, output_2_464;
mixer gate_output_2_464(.a(output_3_464), .b(output_3_0), .y(output_2_464));
wire output_1_465, output_1_1, output_0_465;
mixer gate_output_0_465(.a(output_1_465), .b(output_1_1), .y(output_0_465));
wire output_2_465, output_2_1, output_1_465;
mixer gate_output_1_465(.a(output_2_465), .b(output_2_1), .y(output_1_465));
wire output_3_465, output_3_1, output_2_465;
mixer gate_output_2_465(.a(output_3_465), .b(output_3_1), .y(output_2_465));
wire output_1_466, output_1_2, output_0_466;
mixer gate_output_0_466(.a(output_1_466), .b(output_1_2), .y(output_0_466));
wire output_2_466, output_2_2, output_1_466;
mixer gate_output_1_466(.a(output_2_466), .b(output_2_2), .y(output_1_466));
wire output_3_466, output_3_2, output_2_466;
mixer gate_output_2_466(.a(output_3_466), .b(output_3_2), .y(output_2_466));
wire output_1_467, output_1_0, output_0_467;
mixer gate_output_0_467(.a(output_1_467), .b(output_1_0), .y(output_0_467));
wire output_2_467, output_2_0, output_1_467;
mixer gate_output_1_467(.a(output_2_467), .b(output_2_0), .y(output_1_467));
wire output_3_467, output_3_0, output_2_467;
mixer gate_output_2_467(.a(output_3_467), .b(output_3_0), .y(output_2_467));
wire output_1_468, output_1_1, output_0_468;
mixer gate_output_0_468(.a(output_1_468), .b(output_1_1), .y(output_0_468));
wire output_2_468, output_2_1, output_1_468;
mixer gate_output_1_468(.a(output_2_468), .b(output_2_1), .y(output_1_468));
wire output_3_468, output_3_1, output_2_468;
mixer gate_output_2_468(.a(output_3_468), .b(output_3_1), .y(output_2_468));
wire output_1_469, output_1_2, output_0_469;
mixer gate_output_0_469(.a(output_1_469), .b(output_1_2), .y(output_0_469));
wire output_2_469, output_2_2, output_1_469;
mixer gate_output_1_469(.a(output_2_469), .b(output_2_2), .y(output_1_469));
wire output_3_469, output_3_2, output_2_469;
mixer gate_output_2_469(.a(output_3_469), .b(output_3_2), .y(output_2_469));
wire output_1_470, output_1_0, output_0_470;
mixer gate_output_0_470(.a(output_1_470), .b(output_1_0), .y(output_0_470));
wire output_2_470, output_2_0, output_1_470;
mixer gate_output_1_470(.a(output_2_470), .b(output_2_0), .y(output_1_470));
wire output_3_470, output_3_0, output_2_470;
mixer gate_output_2_470(.a(output_3_470), .b(output_3_0), .y(output_2_470));
wire output_1_471, output_1_1, output_0_471;
mixer gate_output_0_471(.a(output_1_471), .b(output_1_1), .y(output_0_471));
wire output_2_471, output_2_1, output_1_471;
mixer gate_output_1_471(.a(output_2_471), .b(output_2_1), .y(output_1_471));
wire output_3_471, output_3_1, output_2_471;
mixer gate_output_2_471(.a(output_3_471), .b(output_3_1), .y(output_2_471));
wire output_1_472, output_1_2, output_0_472;
mixer gate_output_0_472(.a(output_1_472), .b(output_1_2), .y(output_0_472));
wire output_2_472, output_2_2, output_1_472;
mixer gate_output_1_472(.a(output_2_472), .b(output_2_2), .y(output_1_472));
wire output_3_472, output_3_2, output_2_472;
mixer gate_output_2_472(.a(output_3_472), .b(output_3_2), .y(output_2_472));
wire output_1_473, output_1_0, output_0_473;
mixer gate_output_0_473(.a(output_1_473), .b(output_1_0), .y(output_0_473));
wire output_2_473, output_2_0, output_1_473;
mixer gate_output_1_473(.a(output_2_473), .b(output_2_0), .y(output_1_473));
wire output_3_473, output_3_0, output_2_473;
mixer gate_output_2_473(.a(output_3_473), .b(output_3_0), .y(output_2_473));
wire output_1_474, output_1_1, output_0_474;
mixer gate_output_0_474(.a(output_1_474), .b(output_1_1), .y(output_0_474));
wire output_2_474, output_2_1, output_1_474;
mixer gate_output_1_474(.a(output_2_474), .b(output_2_1), .y(output_1_474));
wire output_3_474, output_3_1, output_2_474;
mixer gate_output_2_474(.a(output_3_474), .b(output_3_1), .y(output_2_474));
wire output_1_475, output_1_2, output_0_475;
mixer gate_output_0_475(.a(output_1_475), .b(output_1_2), .y(output_0_475));
wire output_2_475, output_2_2, output_1_475;
mixer gate_output_1_475(.a(output_2_475), .b(output_2_2), .y(output_1_475));
wire output_3_475, output_3_2, output_2_475;
mixer gate_output_2_475(.a(output_3_475), .b(output_3_2), .y(output_2_475));
wire output_1_476, output_1_0, output_0_476;
mixer gate_output_0_476(.a(output_1_476), .b(output_1_0), .y(output_0_476));
wire output_2_476, output_2_0, output_1_476;
mixer gate_output_1_476(.a(output_2_476), .b(output_2_0), .y(output_1_476));
wire output_3_476, output_3_0, output_2_476;
mixer gate_output_2_476(.a(output_3_476), .b(output_3_0), .y(output_2_476));
wire output_1_477, output_1_1, output_0_477;
mixer gate_output_0_477(.a(output_1_477), .b(output_1_1), .y(output_0_477));
wire output_2_477, output_2_1, output_1_477;
mixer gate_output_1_477(.a(output_2_477), .b(output_2_1), .y(output_1_477));
wire output_3_477, output_3_1, output_2_477;
mixer gate_output_2_477(.a(output_3_477), .b(output_3_1), .y(output_2_477));
wire output_1_478, output_1_2, output_0_478;
mixer gate_output_0_478(.a(output_1_478), .b(output_1_2), .y(output_0_478));
wire output_2_478, output_2_2, output_1_478;
mixer gate_output_1_478(.a(output_2_478), .b(output_2_2), .y(output_1_478));
wire output_3_478, output_3_2, output_2_478;
mixer gate_output_2_478(.a(output_3_478), .b(output_3_2), .y(output_2_478));
wire output_1_479, output_1_0, output_0_479;
mixer gate_output_0_479(.a(output_1_479), .b(output_1_0), .y(output_0_479));
wire output_2_479, output_2_0, output_1_479;
mixer gate_output_1_479(.a(output_2_479), .b(output_2_0), .y(output_1_479));
wire output_3_479, output_3_0, output_2_479;
mixer gate_output_2_479(.a(output_3_479), .b(output_3_0), .y(output_2_479));
wire output_1_480, output_1_1, output_0_480;
mixer gate_output_0_480(.a(output_1_480), .b(output_1_1), .y(output_0_480));
wire output_2_480, output_2_1, output_1_480;
mixer gate_output_1_480(.a(output_2_480), .b(output_2_1), .y(output_1_480));
wire output_3_480, output_3_1, output_2_480;
mixer gate_output_2_480(.a(output_3_480), .b(output_3_1), .y(output_2_480));
wire output_1_481, output_1_2, output_0_481;
mixer gate_output_0_481(.a(output_1_481), .b(output_1_2), .y(output_0_481));
wire output_2_481, output_2_2, output_1_481;
mixer gate_output_1_481(.a(output_2_481), .b(output_2_2), .y(output_1_481));
wire output_3_481, output_3_2, output_2_481;
mixer gate_output_2_481(.a(output_3_481), .b(output_3_2), .y(output_2_481));
wire output_1_482, output_1_0, output_0_482;
mixer gate_output_0_482(.a(output_1_482), .b(output_1_0), .y(output_0_482));
wire output_2_482, output_2_0, output_1_482;
mixer gate_output_1_482(.a(output_2_482), .b(output_2_0), .y(output_1_482));
wire output_3_482, output_3_0, output_2_482;
mixer gate_output_2_482(.a(output_3_482), .b(output_3_0), .y(output_2_482));
wire output_1_483, output_1_1, output_0_483;
mixer gate_output_0_483(.a(output_1_483), .b(output_1_1), .y(output_0_483));
wire output_2_483, output_2_1, output_1_483;
mixer gate_output_1_483(.a(output_2_483), .b(output_2_1), .y(output_1_483));
wire output_3_483, output_3_1, output_2_483;
mixer gate_output_2_483(.a(output_3_483), .b(output_3_1), .y(output_2_483));
wire output_1_484, output_1_2, output_0_484;
mixer gate_output_0_484(.a(output_1_484), .b(output_1_2), .y(output_0_484));
wire output_2_484, output_2_2, output_1_484;
mixer gate_output_1_484(.a(output_2_484), .b(output_2_2), .y(output_1_484));
wire output_3_484, output_3_2, output_2_484;
mixer gate_output_2_484(.a(output_3_484), .b(output_3_2), .y(output_2_484));
wire output_1_485, output_1_0, output_0_485;
mixer gate_output_0_485(.a(output_1_485), .b(output_1_0), .y(output_0_485));
wire output_2_485, output_2_0, output_1_485;
mixer gate_output_1_485(.a(output_2_485), .b(output_2_0), .y(output_1_485));
wire output_3_485, output_3_0, output_2_485;
mixer gate_output_2_485(.a(output_3_485), .b(output_3_0), .y(output_2_485));
wire output_1_486, output_1_1, output_0_486;
mixer gate_output_0_486(.a(output_1_486), .b(output_1_1), .y(output_0_486));
wire output_2_486, output_2_1, output_1_486;
mixer gate_output_1_486(.a(output_2_486), .b(output_2_1), .y(output_1_486));
wire output_3_486, output_3_1, output_2_486;
mixer gate_output_2_486(.a(output_3_486), .b(output_3_1), .y(output_2_486));
wire output_1_487, output_1_2, output_0_487;
mixer gate_output_0_487(.a(output_1_487), .b(output_1_2), .y(output_0_487));
wire output_2_487, output_2_2, output_1_487;
mixer gate_output_1_487(.a(output_2_487), .b(output_2_2), .y(output_1_487));
wire output_3_487, output_3_2, output_2_487;
mixer gate_output_2_487(.a(output_3_487), .b(output_3_2), .y(output_2_487));
wire output_1_488, output_1_0, output_0_488;
mixer gate_output_0_488(.a(output_1_488), .b(output_1_0), .y(output_0_488));
wire output_2_488, output_2_0, output_1_488;
mixer gate_output_1_488(.a(output_2_488), .b(output_2_0), .y(output_1_488));
wire output_3_488, output_3_0, output_2_488;
mixer gate_output_2_488(.a(output_3_488), .b(output_3_0), .y(output_2_488));
wire output_1_489, output_1_1, output_0_489;
mixer gate_output_0_489(.a(output_1_489), .b(output_1_1), .y(output_0_489));
wire output_2_489, output_2_1, output_1_489;
mixer gate_output_1_489(.a(output_2_489), .b(output_2_1), .y(output_1_489));
wire output_3_489, output_3_1, output_2_489;
mixer gate_output_2_489(.a(output_3_489), .b(output_3_1), .y(output_2_489));
wire output_1_490, output_1_2, output_0_490;
mixer gate_output_0_490(.a(output_1_490), .b(output_1_2), .y(output_0_490));
wire output_2_490, output_2_2, output_1_490;
mixer gate_output_1_490(.a(output_2_490), .b(output_2_2), .y(output_1_490));
wire output_3_490, output_3_2, output_2_490;
mixer gate_output_2_490(.a(output_3_490), .b(output_3_2), .y(output_2_490));
wire output_1_491, output_1_0, output_0_491;
mixer gate_output_0_491(.a(output_1_491), .b(output_1_0), .y(output_0_491));
wire output_2_491, output_2_0, output_1_491;
mixer gate_output_1_491(.a(output_2_491), .b(output_2_0), .y(output_1_491));
wire output_3_491, output_3_0, output_2_491;
mixer gate_output_2_491(.a(output_3_491), .b(output_3_0), .y(output_2_491));
wire output_1_492, output_1_1, output_0_492;
mixer gate_output_0_492(.a(output_1_492), .b(output_1_1), .y(output_0_492));
wire output_2_492, output_2_1, output_1_492;
mixer gate_output_1_492(.a(output_2_492), .b(output_2_1), .y(output_1_492));
wire output_3_492, output_3_1, output_2_492;
mixer gate_output_2_492(.a(output_3_492), .b(output_3_1), .y(output_2_492));
wire output_1_493, output_1_2, output_0_493;
mixer gate_output_0_493(.a(output_1_493), .b(output_1_2), .y(output_0_493));
wire output_2_493, output_2_2, output_1_493;
mixer gate_output_1_493(.a(output_2_493), .b(output_2_2), .y(output_1_493));
wire output_3_493, output_3_2, output_2_493;
mixer gate_output_2_493(.a(output_3_493), .b(output_3_2), .y(output_2_493));
wire output_1_494, output_1_0, output_0_494;
mixer gate_output_0_494(.a(output_1_494), .b(output_1_0), .y(output_0_494));
wire output_2_494, output_2_0, output_1_494;
mixer gate_output_1_494(.a(output_2_494), .b(output_2_0), .y(output_1_494));
wire output_3_494, output_3_0, output_2_494;
mixer gate_output_2_494(.a(output_3_494), .b(output_3_0), .y(output_2_494));
wire output_1_495, output_1_1, output_0_495;
mixer gate_output_0_495(.a(output_1_495), .b(output_1_1), .y(output_0_495));
wire output_2_495, output_2_1, output_1_495;
mixer gate_output_1_495(.a(output_2_495), .b(output_2_1), .y(output_1_495));
wire output_3_495, output_3_1, output_2_495;
mixer gate_output_2_495(.a(output_3_495), .b(output_3_1), .y(output_2_495));
wire output_1_496, output_1_2, output_0_496;
mixer gate_output_0_496(.a(output_1_496), .b(output_1_2), .y(output_0_496));
wire output_2_496, output_2_2, output_1_496;
mixer gate_output_1_496(.a(output_2_496), .b(output_2_2), .y(output_1_496));
wire output_3_496, output_3_2, output_2_496;
mixer gate_output_2_496(.a(output_3_496), .b(output_3_2), .y(output_2_496));
wire output_1_497, output_1_0, output_0_497;
mixer gate_output_0_497(.a(output_1_497), .b(output_1_0), .y(output_0_497));
wire output_2_497, output_2_0, output_1_497;
mixer gate_output_1_497(.a(output_2_497), .b(output_2_0), .y(output_1_497));
wire output_3_497, output_3_0, output_2_497;
mixer gate_output_2_497(.a(output_3_497), .b(output_3_0), .y(output_2_497));
wire output_1_498, output_1_1, output_0_498;
mixer gate_output_0_498(.a(output_1_498), .b(output_1_1), .y(output_0_498));
wire output_2_498, output_2_1, output_1_498;
mixer gate_output_1_498(.a(output_2_498), .b(output_2_1), .y(output_1_498));
wire output_3_498, output_3_1, output_2_498;
mixer gate_output_2_498(.a(output_3_498), .b(output_3_1), .y(output_2_498));
wire output_1_499, output_1_2, output_0_499;
mixer gate_output_0_499(.a(output_1_499), .b(output_1_2), .y(output_0_499));
wire output_2_499, output_2_2, output_1_499;
mixer gate_output_1_499(.a(output_2_499), .b(output_2_2), .y(output_1_499));
wire output_3_499, output_3_2, output_2_499;
mixer gate_output_2_499(.a(output_3_499), .b(output_3_2), .y(output_2_499));
wire output_1_500, output_1_0, output_0_500;
mixer gate_output_0_500(.a(output_1_500), .b(output_1_0), .y(output_0_500));
wire output_2_500, output_2_0, output_1_500;
mixer gate_output_1_500(.a(output_2_500), .b(output_2_0), .y(output_1_500));
wire output_3_500, output_3_0, output_2_500;
mixer gate_output_2_500(.a(output_3_500), .b(output_3_0), .y(output_2_500));
wire output_1_501, output_1_1, output_0_501;
mixer gate_output_0_501(.a(output_1_501), .b(output_1_1), .y(output_0_501));
wire output_2_501, output_2_1, output_1_501;
mixer gate_output_1_501(.a(output_2_501), .b(output_2_1), .y(output_1_501));
wire output_3_501, output_3_1, output_2_501;
mixer gate_output_2_501(.a(output_3_501), .b(output_3_1), .y(output_2_501));
wire output_1_502, output_1_2, output_0_502;
mixer gate_output_0_502(.a(output_1_502), .b(output_1_2), .y(output_0_502));
wire output_2_502, output_2_2, output_1_502;
mixer gate_output_1_502(.a(output_2_502), .b(output_2_2), .y(output_1_502));
wire output_3_502, output_3_2, output_2_502;
mixer gate_output_2_502(.a(output_3_502), .b(output_3_2), .y(output_2_502));
wire output_1_503, output_1_0, output_0_503;
mixer gate_output_0_503(.a(output_1_503), .b(output_1_0), .y(output_0_503));
wire output_2_503, output_2_0, output_1_503;
mixer gate_output_1_503(.a(output_2_503), .b(output_2_0), .y(output_1_503));
wire output_3_503, output_3_0, output_2_503;
mixer gate_output_2_503(.a(output_3_503), .b(output_3_0), .y(output_2_503));
wire output_1_504, output_1_1, output_0_504;
mixer gate_output_0_504(.a(output_1_504), .b(output_1_1), .y(output_0_504));
wire output_2_504, output_2_1, output_1_504;
mixer gate_output_1_504(.a(output_2_504), .b(output_2_1), .y(output_1_504));
wire output_3_504, output_3_1, output_2_504;
mixer gate_output_2_504(.a(output_3_504), .b(output_3_1), .y(output_2_504));
wire output_1_505, output_1_2, output_0_505;
mixer gate_output_0_505(.a(output_1_505), .b(output_1_2), .y(output_0_505));
wire output_2_505, output_2_2, output_1_505;
mixer gate_output_1_505(.a(output_2_505), .b(output_2_2), .y(output_1_505));
wire output_3_505, output_3_2, output_2_505;
mixer gate_output_2_505(.a(output_3_505), .b(output_3_2), .y(output_2_505));
wire output_1_506, output_1_0, output_0_506;
mixer gate_output_0_506(.a(output_1_506), .b(output_1_0), .y(output_0_506));
wire output_2_506, output_2_0, output_1_506;
mixer gate_output_1_506(.a(output_2_506), .b(output_2_0), .y(output_1_506));
wire output_3_506, output_3_0, output_2_506;
mixer gate_output_2_506(.a(output_3_506), .b(output_3_0), .y(output_2_506));
wire output_1_507, output_1_1, output_0_507;
mixer gate_output_0_507(.a(output_1_507), .b(output_1_1), .y(output_0_507));
wire output_2_507, output_2_1, output_1_507;
mixer gate_output_1_507(.a(output_2_507), .b(output_2_1), .y(output_1_507));
wire output_3_507, output_3_1, output_2_507;
mixer gate_output_2_507(.a(output_3_507), .b(output_3_1), .y(output_2_507));
wire output_1_508, output_1_2, output_0_508;
mixer gate_output_0_508(.a(output_1_508), .b(output_1_2), .y(output_0_508));
wire output_2_508, output_2_2, output_1_508;
mixer gate_output_1_508(.a(output_2_508), .b(output_2_2), .y(output_1_508));
wire output_3_508, output_3_2, output_2_508;
mixer gate_output_2_508(.a(output_3_508), .b(output_3_2), .y(output_2_508));
wire output_1_509, output_1_0, output_0_509;
mixer gate_output_0_509(.a(output_1_509), .b(output_1_0), .y(output_0_509));
wire output_2_509, output_2_0, output_1_509;
mixer gate_output_1_509(.a(output_2_509), .b(output_2_0), .y(output_1_509));
wire output_3_509, output_3_0, output_2_509;
mixer gate_output_2_509(.a(output_3_509), .b(output_3_0), .y(output_2_509));
wire output_1_510, output_1_1, output_0_510;
mixer gate_output_0_510(.a(output_1_510), .b(output_1_1), .y(output_0_510));
wire output_2_510, output_2_1, output_1_510;
mixer gate_output_1_510(.a(output_2_510), .b(output_2_1), .y(output_1_510));
wire output_3_510, output_3_1, output_2_510;
mixer gate_output_2_510(.a(output_3_510), .b(output_3_1), .y(output_2_510));
wire output_1_511, output_1_2, output_0_511;
mixer gate_output_0_511(.a(output_1_511), .b(output_1_2), .y(output_0_511));
wire output_2_511, output_2_2, output_1_511;
mixer gate_output_1_511(.a(output_2_511), .b(output_2_2), .y(output_1_511));
wire output_3_511, output_3_2, output_2_511;
mixer gate_output_2_511(.a(output_3_511), .b(output_3_2), .y(output_2_511));
assign output_0 = output_0_0;
wire output_0_512;
assign output_0_512 = input_0;
assign output_1 = output_1_0;
wire output_1_512;
assign output_1_512 = input_1;
assign output_2 = output_2_0;
wire output_2_512;
assign output_2_512 = input_2;
endmodule
