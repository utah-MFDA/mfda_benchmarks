module complete_16 (
inout io_0,inout io_1,inout io_2,inout io_3,inout io_4,inout io_5,inout io_6,inout io_7,inout io_8,inout io_9,inout io_10,inout io_11,inout io_12,inout io_13,inout io_14,inout io_15
);
assign io_0 = input_0;
assign io_0 = input_1;
assign io_0 = input_2;
assign io_0 = input_3;
assign io_0 = input_4;
assign io_0 = input_5;
assign io_0 = input_6;
assign io_0 = input_7;
assign io_0 = input_8;
assign io_0 = input_9;
assign io_0 = input_10;
assign io_0 = input_11;
assign io_0 = input_12;
assign io_0 = input_13;
assign io_0 = input_14;
assign io_0 = input_15;
assign io_1 = input_1;
assign io_1 = input_2;
assign io_1 = input_3;
assign io_1 = input_4;
assign io_1 = input_5;
assign io_1 = input_6;
assign io_1 = input_7;
assign io_1 = input_8;
assign io_1 = input_9;
assign io_1 = input_10;
assign io_1 = input_11;
assign io_1 = input_12;
assign io_1 = input_13;
assign io_1 = input_14;
assign io_1 = input_15;
assign io_2 = input_2;
assign io_2 = input_3;
assign io_2 = input_4;
assign io_2 = input_5;
assign io_2 = input_6;
assign io_2 = input_7;
assign io_2 = input_8;
assign io_2 = input_9;
assign io_2 = input_10;
assign io_2 = input_11;
assign io_2 = input_12;
assign io_2 = input_13;
assign io_2 = input_14;
assign io_2 = input_15;
assign io_3 = input_3;
assign io_3 = input_4;
assign io_3 = input_5;
assign io_3 = input_6;
assign io_3 = input_7;
assign io_3 = input_8;
assign io_3 = input_9;
assign io_3 = input_10;
assign io_3 = input_11;
assign io_3 = input_12;
assign io_3 = input_13;
assign io_3 = input_14;
assign io_3 = input_15;
assign io_4 = input_4;
assign io_4 = input_5;
assign io_4 = input_6;
assign io_4 = input_7;
assign io_4 = input_8;
assign io_4 = input_9;
assign io_4 = input_10;
assign io_4 = input_11;
assign io_4 = input_12;
assign io_4 = input_13;
assign io_4 = input_14;
assign io_4 = input_15;
assign io_5 = input_5;
assign io_5 = input_6;
assign io_5 = input_7;
assign io_5 = input_8;
assign io_5 = input_9;
assign io_5 = input_10;
assign io_5 = input_11;
assign io_5 = input_12;
assign io_5 = input_13;
assign io_5 = input_14;
assign io_5 = input_15;
assign io_6 = input_6;
assign io_6 = input_7;
assign io_6 = input_8;
assign io_6 = input_9;
assign io_6 = input_10;
assign io_6 = input_11;
assign io_6 = input_12;
assign io_6 = input_13;
assign io_6 = input_14;
assign io_6 = input_15;
assign io_7 = input_7;
assign io_7 = input_8;
assign io_7 = input_9;
assign io_7 = input_10;
assign io_7 = input_11;
assign io_7 = input_12;
assign io_7 = input_13;
assign io_7 = input_14;
assign io_7 = input_15;
assign io_8 = input_8;
assign io_8 = input_9;
assign io_8 = input_10;
assign io_8 = input_11;
assign io_8 = input_12;
assign io_8 = input_13;
assign io_8 = input_14;
assign io_8 = input_15;
assign io_9 = input_9;
assign io_9 = input_10;
assign io_9 = input_11;
assign io_9 = input_12;
assign io_9 = input_13;
assign io_9 = input_14;
assign io_9 = input_15;
assign io_10 = input_10;
assign io_10 = input_11;
assign io_10 = input_12;
assign io_10 = input_13;
assign io_10 = input_14;
assign io_10 = input_15;
assign io_11 = input_11;
assign io_11 = input_12;
assign io_11 = input_13;
assign io_11 = input_14;
assign io_11 = input_15;
assign io_12 = input_12;
assign io_12 = input_13;
assign io_12 = input_14;
assign io_12 = input_15;
assign io_13 = input_13;
assign io_13 = input_14;
assign io_13 = input_15;
assign io_14 = input_14;
assign io_14 = input_15;
assign io_15 = input_15;
endmodule
