module complete_32 (
inout io_0,inout io_1,inout io_2,inout io_3,inout io_4,inout io_5,inout io_6,inout io_7,inout io_8,inout io_9,inout io_10,inout io_11,inout io_12,inout io_13,inout io_14,inout io_15,inout io_16,inout io_17,inout io_18,inout io_19,inout io_20,inout io_21,inout io_22,inout io_23,inout io_24,inout io_25,inout io_26,inout io_27,inout io_28,inout io_29,inout io_30,inout io_31
);
assign io_0 = input_0;
assign io_0 = input_1;
assign io_0 = input_2;
assign io_0 = input_3;
assign io_0 = input_4;
assign io_0 = input_5;
assign io_0 = input_6;
assign io_0 = input_7;
assign io_0 = input_8;
assign io_0 = input_9;
assign io_0 = input_10;
assign io_0 = input_11;
assign io_0 = input_12;
assign io_0 = input_13;
assign io_0 = input_14;
assign io_0 = input_15;
assign io_0 = input_16;
assign io_0 = input_17;
assign io_0 = input_18;
assign io_0 = input_19;
assign io_0 = input_20;
assign io_0 = input_21;
assign io_0 = input_22;
assign io_0 = input_23;
assign io_0 = input_24;
assign io_0 = input_25;
assign io_0 = input_26;
assign io_0 = input_27;
assign io_0 = input_28;
assign io_0 = input_29;
assign io_0 = input_30;
assign io_0 = input_31;
assign io_1 = input_1;
assign io_1 = input_2;
assign io_1 = input_3;
assign io_1 = input_4;
assign io_1 = input_5;
assign io_1 = input_6;
assign io_1 = input_7;
assign io_1 = input_8;
assign io_1 = input_9;
assign io_1 = input_10;
assign io_1 = input_11;
assign io_1 = input_12;
assign io_1 = input_13;
assign io_1 = input_14;
assign io_1 = input_15;
assign io_1 = input_16;
assign io_1 = input_17;
assign io_1 = input_18;
assign io_1 = input_19;
assign io_1 = input_20;
assign io_1 = input_21;
assign io_1 = input_22;
assign io_1 = input_23;
assign io_1 = input_24;
assign io_1 = input_25;
assign io_1 = input_26;
assign io_1 = input_27;
assign io_1 = input_28;
assign io_1 = input_29;
assign io_1 = input_30;
assign io_1 = input_31;
assign io_2 = input_2;
assign io_2 = input_3;
assign io_2 = input_4;
assign io_2 = input_5;
assign io_2 = input_6;
assign io_2 = input_7;
assign io_2 = input_8;
assign io_2 = input_9;
assign io_2 = input_10;
assign io_2 = input_11;
assign io_2 = input_12;
assign io_2 = input_13;
assign io_2 = input_14;
assign io_2 = input_15;
assign io_2 = input_16;
assign io_2 = input_17;
assign io_2 = input_18;
assign io_2 = input_19;
assign io_2 = input_20;
assign io_2 = input_21;
assign io_2 = input_22;
assign io_2 = input_23;
assign io_2 = input_24;
assign io_2 = input_25;
assign io_2 = input_26;
assign io_2 = input_27;
assign io_2 = input_28;
assign io_2 = input_29;
assign io_2 = input_30;
assign io_2 = input_31;
assign io_3 = input_3;
assign io_3 = input_4;
assign io_3 = input_5;
assign io_3 = input_6;
assign io_3 = input_7;
assign io_3 = input_8;
assign io_3 = input_9;
assign io_3 = input_10;
assign io_3 = input_11;
assign io_3 = input_12;
assign io_3 = input_13;
assign io_3 = input_14;
assign io_3 = input_15;
assign io_3 = input_16;
assign io_3 = input_17;
assign io_3 = input_18;
assign io_3 = input_19;
assign io_3 = input_20;
assign io_3 = input_21;
assign io_3 = input_22;
assign io_3 = input_23;
assign io_3 = input_24;
assign io_3 = input_25;
assign io_3 = input_26;
assign io_3 = input_27;
assign io_3 = input_28;
assign io_3 = input_29;
assign io_3 = input_30;
assign io_3 = input_31;
assign io_4 = input_4;
assign io_4 = input_5;
assign io_4 = input_6;
assign io_4 = input_7;
assign io_4 = input_8;
assign io_4 = input_9;
assign io_4 = input_10;
assign io_4 = input_11;
assign io_4 = input_12;
assign io_4 = input_13;
assign io_4 = input_14;
assign io_4 = input_15;
assign io_4 = input_16;
assign io_4 = input_17;
assign io_4 = input_18;
assign io_4 = input_19;
assign io_4 = input_20;
assign io_4 = input_21;
assign io_4 = input_22;
assign io_4 = input_23;
assign io_4 = input_24;
assign io_4 = input_25;
assign io_4 = input_26;
assign io_4 = input_27;
assign io_4 = input_28;
assign io_4 = input_29;
assign io_4 = input_30;
assign io_4 = input_31;
assign io_5 = input_5;
assign io_5 = input_6;
assign io_5 = input_7;
assign io_5 = input_8;
assign io_5 = input_9;
assign io_5 = input_10;
assign io_5 = input_11;
assign io_5 = input_12;
assign io_5 = input_13;
assign io_5 = input_14;
assign io_5 = input_15;
assign io_5 = input_16;
assign io_5 = input_17;
assign io_5 = input_18;
assign io_5 = input_19;
assign io_5 = input_20;
assign io_5 = input_21;
assign io_5 = input_22;
assign io_5 = input_23;
assign io_5 = input_24;
assign io_5 = input_25;
assign io_5 = input_26;
assign io_5 = input_27;
assign io_5 = input_28;
assign io_5 = input_29;
assign io_5 = input_30;
assign io_5 = input_31;
assign io_6 = input_6;
assign io_6 = input_7;
assign io_6 = input_8;
assign io_6 = input_9;
assign io_6 = input_10;
assign io_6 = input_11;
assign io_6 = input_12;
assign io_6 = input_13;
assign io_6 = input_14;
assign io_6 = input_15;
assign io_6 = input_16;
assign io_6 = input_17;
assign io_6 = input_18;
assign io_6 = input_19;
assign io_6 = input_20;
assign io_6 = input_21;
assign io_6 = input_22;
assign io_6 = input_23;
assign io_6 = input_24;
assign io_6 = input_25;
assign io_6 = input_26;
assign io_6 = input_27;
assign io_6 = input_28;
assign io_6 = input_29;
assign io_6 = input_30;
assign io_6 = input_31;
assign io_7 = input_7;
assign io_7 = input_8;
assign io_7 = input_9;
assign io_7 = input_10;
assign io_7 = input_11;
assign io_7 = input_12;
assign io_7 = input_13;
assign io_7 = input_14;
assign io_7 = input_15;
assign io_7 = input_16;
assign io_7 = input_17;
assign io_7 = input_18;
assign io_7 = input_19;
assign io_7 = input_20;
assign io_7 = input_21;
assign io_7 = input_22;
assign io_7 = input_23;
assign io_7 = input_24;
assign io_7 = input_25;
assign io_7 = input_26;
assign io_7 = input_27;
assign io_7 = input_28;
assign io_7 = input_29;
assign io_7 = input_30;
assign io_7 = input_31;
assign io_8 = input_8;
assign io_8 = input_9;
assign io_8 = input_10;
assign io_8 = input_11;
assign io_8 = input_12;
assign io_8 = input_13;
assign io_8 = input_14;
assign io_8 = input_15;
assign io_8 = input_16;
assign io_8 = input_17;
assign io_8 = input_18;
assign io_8 = input_19;
assign io_8 = input_20;
assign io_8 = input_21;
assign io_8 = input_22;
assign io_8 = input_23;
assign io_8 = input_24;
assign io_8 = input_25;
assign io_8 = input_26;
assign io_8 = input_27;
assign io_8 = input_28;
assign io_8 = input_29;
assign io_8 = input_30;
assign io_8 = input_31;
assign io_9 = input_9;
assign io_9 = input_10;
assign io_9 = input_11;
assign io_9 = input_12;
assign io_9 = input_13;
assign io_9 = input_14;
assign io_9 = input_15;
assign io_9 = input_16;
assign io_9 = input_17;
assign io_9 = input_18;
assign io_9 = input_19;
assign io_9 = input_20;
assign io_9 = input_21;
assign io_9 = input_22;
assign io_9 = input_23;
assign io_9 = input_24;
assign io_9 = input_25;
assign io_9 = input_26;
assign io_9 = input_27;
assign io_9 = input_28;
assign io_9 = input_29;
assign io_9 = input_30;
assign io_9 = input_31;
assign io_10 = input_10;
assign io_10 = input_11;
assign io_10 = input_12;
assign io_10 = input_13;
assign io_10 = input_14;
assign io_10 = input_15;
assign io_10 = input_16;
assign io_10 = input_17;
assign io_10 = input_18;
assign io_10 = input_19;
assign io_10 = input_20;
assign io_10 = input_21;
assign io_10 = input_22;
assign io_10 = input_23;
assign io_10 = input_24;
assign io_10 = input_25;
assign io_10 = input_26;
assign io_10 = input_27;
assign io_10 = input_28;
assign io_10 = input_29;
assign io_10 = input_30;
assign io_10 = input_31;
assign io_11 = input_11;
assign io_11 = input_12;
assign io_11 = input_13;
assign io_11 = input_14;
assign io_11 = input_15;
assign io_11 = input_16;
assign io_11 = input_17;
assign io_11 = input_18;
assign io_11 = input_19;
assign io_11 = input_20;
assign io_11 = input_21;
assign io_11 = input_22;
assign io_11 = input_23;
assign io_11 = input_24;
assign io_11 = input_25;
assign io_11 = input_26;
assign io_11 = input_27;
assign io_11 = input_28;
assign io_11 = input_29;
assign io_11 = input_30;
assign io_11 = input_31;
assign io_12 = input_12;
assign io_12 = input_13;
assign io_12 = input_14;
assign io_12 = input_15;
assign io_12 = input_16;
assign io_12 = input_17;
assign io_12 = input_18;
assign io_12 = input_19;
assign io_12 = input_20;
assign io_12 = input_21;
assign io_12 = input_22;
assign io_12 = input_23;
assign io_12 = input_24;
assign io_12 = input_25;
assign io_12 = input_26;
assign io_12 = input_27;
assign io_12 = input_28;
assign io_12 = input_29;
assign io_12 = input_30;
assign io_12 = input_31;
assign io_13 = input_13;
assign io_13 = input_14;
assign io_13 = input_15;
assign io_13 = input_16;
assign io_13 = input_17;
assign io_13 = input_18;
assign io_13 = input_19;
assign io_13 = input_20;
assign io_13 = input_21;
assign io_13 = input_22;
assign io_13 = input_23;
assign io_13 = input_24;
assign io_13 = input_25;
assign io_13 = input_26;
assign io_13 = input_27;
assign io_13 = input_28;
assign io_13 = input_29;
assign io_13 = input_30;
assign io_13 = input_31;
assign io_14 = input_14;
assign io_14 = input_15;
assign io_14 = input_16;
assign io_14 = input_17;
assign io_14 = input_18;
assign io_14 = input_19;
assign io_14 = input_20;
assign io_14 = input_21;
assign io_14 = input_22;
assign io_14 = input_23;
assign io_14 = input_24;
assign io_14 = input_25;
assign io_14 = input_26;
assign io_14 = input_27;
assign io_14 = input_28;
assign io_14 = input_29;
assign io_14 = input_30;
assign io_14 = input_31;
assign io_15 = input_15;
assign io_15 = input_16;
assign io_15 = input_17;
assign io_15 = input_18;
assign io_15 = input_19;
assign io_15 = input_20;
assign io_15 = input_21;
assign io_15 = input_22;
assign io_15 = input_23;
assign io_15 = input_24;
assign io_15 = input_25;
assign io_15 = input_26;
assign io_15 = input_27;
assign io_15 = input_28;
assign io_15 = input_29;
assign io_15 = input_30;
assign io_15 = input_31;
assign io_16 = input_16;
assign io_16 = input_17;
assign io_16 = input_18;
assign io_16 = input_19;
assign io_16 = input_20;
assign io_16 = input_21;
assign io_16 = input_22;
assign io_16 = input_23;
assign io_16 = input_24;
assign io_16 = input_25;
assign io_16 = input_26;
assign io_16 = input_27;
assign io_16 = input_28;
assign io_16 = input_29;
assign io_16 = input_30;
assign io_16 = input_31;
assign io_17 = input_17;
assign io_17 = input_18;
assign io_17 = input_19;
assign io_17 = input_20;
assign io_17 = input_21;
assign io_17 = input_22;
assign io_17 = input_23;
assign io_17 = input_24;
assign io_17 = input_25;
assign io_17 = input_26;
assign io_17 = input_27;
assign io_17 = input_28;
assign io_17 = input_29;
assign io_17 = input_30;
assign io_17 = input_31;
assign io_18 = input_18;
assign io_18 = input_19;
assign io_18 = input_20;
assign io_18 = input_21;
assign io_18 = input_22;
assign io_18 = input_23;
assign io_18 = input_24;
assign io_18 = input_25;
assign io_18 = input_26;
assign io_18 = input_27;
assign io_18 = input_28;
assign io_18 = input_29;
assign io_18 = input_30;
assign io_18 = input_31;
assign io_19 = input_19;
assign io_19 = input_20;
assign io_19 = input_21;
assign io_19 = input_22;
assign io_19 = input_23;
assign io_19 = input_24;
assign io_19 = input_25;
assign io_19 = input_26;
assign io_19 = input_27;
assign io_19 = input_28;
assign io_19 = input_29;
assign io_19 = input_30;
assign io_19 = input_31;
assign io_20 = input_20;
assign io_20 = input_21;
assign io_20 = input_22;
assign io_20 = input_23;
assign io_20 = input_24;
assign io_20 = input_25;
assign io_20 = input_26;
assign io_20 = input_27;
assign io_20 = input_28;
assign io_20 = input_29;
assign io_20 = input_30;
assign io_20 = input_31;
assign io_21 = input_21;
assign io_21 = input_22;
assign io_21 = input_23;
assign io_21 = input_24;
assign io_21 = input_25;
assign io_21 = input_26;
assign io_21 = input_27;
assign io_21 = input_28;
assign io_21 = input_29;
assign io_21 = input_30;
assign io_21 = input_31;
assign io_22 = input_22;
assign io_22 = input_23;
assign io_22 = input_24;
assign io_22 = input_25;
assign io_22 = input_26;
assign io_22 = input_27;
assign io_22 = input_28;
assign io_22 = input_29;
assign io_22 = input_30;
assign io_22 = input_31;
assign io_23 = input_23;
assign io_23 = input_24;
assign io_23 = input_25;
assign io_23 = input_26;
assign io_23 = input_27;
assign io_23 = input_28;
assign io_23 = input_29;
assign io_23 = input_30;
assign io_23 = input_31;
assign io_24 = input_24;
assign io_24 = input_25;
assign io_24 = input_26;
assign io_24 = input_27;
assign io_24 = input_28;
assign io_24 = input_29;
assign io_24 = input_30;
assign io_24 = input_31;
assign io_25 = input_25;
assign io_25 = input_26;
assign io_25 = input_27;
assign io_25 = input_28;
assign io_25 = input_29;
assign io_25 = input_30;
assign io_25 = input_31;
assign io_26 = input_26;
assign io_26 = input_27;
assign io_26 = input_28;
assign io_26 = input_29;
assign io_26 = input_30;
assign io_26 = input_31;
assign io_27 = input_27;
assign io_27 = input_28;
assign io_27 = input_29;
assign io_27 = input_30;
assign io_27 = input_31;
assign io_28 = input_28;
assign io_28 = input_29;
assign io_28 = input_30;
assign io_28 = input_31;
assign io_29 = input_29;
assign io_29 = input_30;
assign io_29 = input_31;
assign io_30 = input_30;
assign io_30 = input_31;
assign io_31 = input_31;
endmodule
