module complete_bipartite_16_16 (
inout input_0,inout input_1,inout input_2,inout input_3,inout input_4,inout input_5,inout input_6,inout input_7,inout input_8,inout input_9,inout input_10,inout input_11,inout input_12,inout input_13,inout input_14,inout input_15,inout output_0,inout output_1,inout output_2,inout output_3,inout output_4,inout output_5,inout output_6,inout output_7,inout output_8,inout output_9,inout output_10,inout output_11,inout output_12,inout output_13,inout output_14,inout output_15
);
assign output_0 = input_0;
assign output_1 = input_0;
assign output_2 = input_0;
assign output_3 = input_0;
assign output_4 = input_0;
assign output_5 = input_0;
assign output_6 = input_0;
assign output_7 = input_0;
assign output_8 = input_0;
assign output_9 = input_0;
assign output_10 = input_0;
assign output_11 = input_0;
assign output_12 = input_0;
assign output_13 = input_0;
assign output_14 = input_0;
assign output_15 = input_0;
assign output_0 = input_1;
assign output_1 = input_1;
assign output_2 = input_1;
assign output_3 = input_1;
assign output_4 = input_1;
assign output_5 = input_1;
assign output_6 = input_1;
assign output_7 = input_1;
assign output_8 = input_1;
assign output_9 = input_1;
assign output_10 = input_1;
assign output_11 = input_1;
assign output_12 = input_1;
assign output_13 = input_1;
assign output_14 = input_1;
assign output_15 = input_1;
assign output_0 = input_2;
assign output_1 = input_2;
assign output_2 = input_2;
assign output_3 = input_2;
assign output_4 = input_2;
assign output_5 = input_2;
assign output_6 = input_2;
assign output_7 = input_2;
assign output_8 = input_2;
assign output_9 = input_2;
assign output_10 = input_2;
assign output_11 = input_2;
assign output_12 = input_2;
assign output_13 = input_2;
assign output_14 = input_2;
assign output_15 = input_2;
assign output_0 = input_3;
assign output_1 = input_3;
assign output_2 = input_3;
assign output_3 = input_3;
assign output_4 = input_3;
assign output_5 = input_3;
assign output_6 = input_3;
assign output_7 = input_3;
assign output_8 = input_3;
assign output_9 = input_3;
assign output_10 = input_3;
assign output_11 = input_3;
assign output_12 = input_3;
assign output_13 = input_3;
assign output_14 = input_3;
assign output_15 = input_3;
assign output_0 = input_4;
assign output_1 = input_4;
assign output_2 = input_4;
assign output_3 = input_4;
assign output_4 = input_4;
assign output_5 = input_4;
assign output_6 = input_4;
assign output_7 = input_4;
assign output_8 = input_4;
assign output_9 = input_4;
assign output_10 = input_4;
assign output_11 = input_4;
assign output_12 = input_4;
assign output_13 = input_4;
assign output_14 = input_4;
assign output_15 = input_4;
assign output_0 = input_5;
assign output_1 = input_5;
assign output_2 = input_5;
assign output_3 = input_5;
assign output_4 = input_5;
assign output_5 = input_5;
assign output_6 = input_5;
assign output_7 = input_5;
assign output_8 = input_5;
assign output_9 = input_5;
assign output_10 = input_5;
assign output_11 = input_5;
assign output_12 = input_5;
assign output_13 = input_5;
assign output_14 = input_5;
assign output_15 = input_5;
assign output_0 = input_6;
assign output_1 = input_6;
assign output_2 = input_6;
assign output_3 = input_6;
assign output_4 = input_6;
assign output_5 = input_6;
assign output_6 = input_6;
assign output_7 = input_6;
assign output_8 = input_6;
assign output_9 = input_6;
assign output_10 = input_6;
assign output_11 = input_6;
assign output_12 = input_6;
assign output_13 = input_6;
assign output_14 = input_6;
assign output_15 = input_6;
assign output_0 = input_7;
assign output_1 = input_7;
assign output_2 = input_7;
assign output_3 = input_7;
assign output_4 = input_7;
assign output_5 = input_7;
assign output_6 = input_7;
assign output_7 = input_7;
assign output_8 = input_7;
assign output_9 = input_7;
assign output_10 = input_7;
assign output_11 = input_7;
assign output_12 = input_7;
assign output_13 = input_7;
assign output_14 = input_7;
assign output_15 = input_7;
assign output_0 = input_8;
assign output_1 = input_8;
assign output_2 = input_8;
assign output_3 = input_8;
assign output_4 = input_8;
assign output_5 = input_8;
assign output_6 = input_8;
assign output_7 = input_8;
assign output_8 = input_8;
assign output_9 = input_8;
assign output_10 = input_8;
assign output_11 = input_8;
assign output_12 = input_8;
assign output_13 = input_8;
assign output_14 = input_8;
assign output_15 = input_8;
assign output_0 = input_9;
assign output_1 = input_9;
assign output_2 = input_9;
assign output_3 = input_9;
assign output_4 = input_9;
assign output_5 = input_9;
assign output_6 = input_9;
assign output_7 = input_9;
assign output_8 = input_9;
assign output_9 = input_9;
assign output_10 = input_9;
assign output_11 = input_9;
assign output_12 = input_9;
assign output_13 = input_9;
assign output_14 = input_9;
assign output_15 = input_9;
assign output_0 = input_10;
assign output_1 = input_10;
assign output_2 = input_10;
assign output_3 = input_10;
assign output_4 = input_10;
assign output_5 = input_10;
assign output_6 = input_10;
assign output_7 = input_10;
assign output_8 = input_10;
assign output_9 = input_10;
assign output_10 = input_10;
assign output_11 = input_10;
assign output_12 = input_10;
assign output_13 = input_10;
assign output_14 = input_10;
assign output_15 = input_10;
assign output_0 = input_11;
assign output_1 = input_11;
assign output_2 = input_11;
assign output_3 = input_11;
assign output_4 = input_11;
assign output_5 = input_11;
assign output_6 = input_11;
assign output_7 = input_11;
assign output_8 = input_11;
assign output_9 = input_11;
assign output_10 = input_11;
assign output_11 = input_11;
assign output_12 = input_11;
assign output_13 = input_11;
assign output_14 = input_11;
assign output_15 = input_11;
assign output_0 = input_12;
assign output_1 = input_12;
assign output_2 = input_12;
assign output_3 = input_12;
assign output_4 = input_12;
assign output_5 = input_12;
assign output_6 = input_12;
assign output_7 = input_12;
assign output_8 = input_12;
assign output_9 = input_12;
assign output_10 = input_12;
assign output_11 = input_12;
assign output_12 = input_12;
assign output_13 = input_12;
assign output_14 = input_12;
assign output_15 = input_12;
assign output_0 = input_13;
assign output_1 = input_13;
assign output_2 = input_13;
assign output_3 = input_13;
assign output_4 = input_13;
assign output_5 = input_13;
assign output_6 = input_13;
assign output_7 = input_13;
assign output_8 = input_13;
assign output_9 = input_13;
assign output_10 = input_13;
assign output_11 = input_13;
assign output_12 = input_13;
assign output_13 = input_13;
assign output_14 = input_13;
assign output_15 = input_13;
assign output_0 = input_14;
assign output_1 = input_14;
assign output_2 = input_14;
assign output_3 = input_14;
assign output_4 = input_14;
assign output_5 = input_14;
assign output_6 = input_14;
assign output_7 = input_14;
assign output_8 = input_14;
assign output_9 = input_14;
assign output_10 = input_14;
assign output_11 = input_14;
assign output_12 = input_14;
assign output_13 = input_14;
assign output_14 = input_14;
assign output_15 = input_14;
assign output_0 = input_15;
assign output_1 = input_15;
assign output_2 = input_15;
assign output_3 = input_15;
assign output_4 = input_15;
assign output_5 = input_15;
assign output_6 = input_15;
assign output_7 = input_15;
assign output_8 = input_15;
assign output_9 = input_15;
assign output_10 = input_15;
assign output_11 = input_15;
assign output_12 = input_15;
assign output_13 = input_15;
assign output_14 = input_15;
assign output_15 = input_15;
endmodule
