module biggs_smith();
	mixer m_0(.a(e_0_1), .b(e_0_2), .y(e_0_3));
	mixer m_1(.a(e_0_1), .b(e_1_96), .y(e_1_97));
	mixer m_2(.a(e_0_2), .b(e_2_98), .y(e_2_101));
	mixer m_3(.a(e_0_3), .b(e_3_99), .y(e_3_100));
	mixer m_4(.a(e_4_12), .b(e_4_14), .y(e_4_15));
	mixer m_5(.a(e_5_13), .b(e_5_16), .y(e_5_17));
	mixer m_6(.a(e_6_18), .b(e_6_19), .y(e_6_33));
	mixer m_7(.a(e_7_21), .b(e_7_23), .y(e_7_34));
	mixer m_8(.a(e_8_20), .b(e_8_25), .y(e_8_32));
	mixer m_9(.a(e_9_22), .b(e_9_24), .y(e_9_26));
	mixer m_10(.a(e_10_27), .b(e_10_31), .y(e_10_35));
	mixer m_11(.a(e_11_28), .b(e_11_29), .y(e_11_30));
	mixer m_12(.a(e_4_12), .b(e_12_13), .y(e_12_36));
	mixer m_13(.a(e_5_13), .b(e_12_13), .y(e_13_38));
	mixer m_14(.a(e_4_14), .b(e_14_35), .y(e_14_59));
	mixer m_15(.a(e_4_15), .b(e_15_34), .y(e_15_58));
	mixer m_16(.a(e_5_16), .b(e_16_33), .y(e_16_57));
	mixer m_17(.a(e_5_17), .b(e_17_32), .y(e_17_41));
	mixer m_18(.a(e_6_18), .b(e_18_31), .y(e_18_37));
	mixer m_19(.a(e_6_19), .b(e_19_30), .y(e_19_46));
	mixer m_20(.a(e_8_20), .b(e_20_21), .y(e_20_49));
	mixer m_21(.a(e_7_21), .b(e_20_21), .y(e_21_39));
	mixer m_22(.a(e_9_22), .b(e_22_23), .y(e_22_51));
	mixer m_23(.a(e_7_23), .b(e_22_23), .y(e_23_45));
	mixer m_24(.a(e_9_24), .b(e_24_27), .y(e_24_52));
	mixer m_25(.a(e_8_25), .b(e_25_29), .y(e_25_44));
	mixer m_26(.a(e_9_26), .b(e_26_28), .y(e_26_40));
	mixer m_27(.a(e_10_27), .b(e_24_27), .y(e_27_53));
	mixer m_28(.a(e_11_28), .b(e_26_28), .y(e_28_54));
	mixer m_29(.a(e_11_29), .b(e_25_29), .y(e_29_47));
	mixer m_30(.a(e_11_30), .b(e_19_30), .y(e_30_56));
	mixer m_31(.a(e_10_31), .b(e_18_31), .y(e_31_55));
	mixer m_32(.a(e_8_32), .b(e_17_32), .y(e_32_48));
	mixer m_33(.a(e_6_33), .b(e_16_33), .y(e_33_43));
	mixer m_34(.a(e_7_34), .b(e_15_34), .y(e_34_50));
	mixer m_35(.a(e_10_35), .b(e_14_35), .y(e_35_42));
	mixer m_36(.a(e_12_36), .b(e_36_37), .y(e_36_60));
	mixer m_37(.a(e_18_37), .b(e_36_37), .y(e_37_79));
	mixer m_38(.a(e_13_38), .b(e_38_39), .y(e_38_63));
	mixer m_39(.a(e_21_39), .b(e_38_39), .y(e_39_80));
	mixer m_40(.a(e_26_40), .b(e_40_49), .y(e_40_64));
	mixer m_41(.a(e_17_41), .b(e_41_56), .y(e_41_65));
	mixer m_42(.a(e_35_42), .b(e_42_57), .y(e_42_76));
	mixer m_43(.a(e_33_43), .b(e_43_44), .y(e_43_71));
	mixer m_44(.a(e_25_44), .b(e_43_44), .y(e_44_77));
	mixer m_45(.a(e_23_45), .b(e_45_47), .y(e_45_72));
	mixer m_46(.a(e_19_46), .b(e_46_52), .y(e_46_73));
	mixer m_47(.a(e_29_47), .b(e_45_47), .y(e_47_75));
	mixer m_48(.a(e_32_48), .b(e_48_58), .y(e_48_67));
	mixer m_49(.a(e_20_49), .b(e_40_49), .y(e_49_78));
	mixer m_50(.a(e_34_50), .b(e_50_53), .y(e_50_81));
	mixer m_51(.a(e_22_51), .b(e_51_59), .y(e_51_70));
	mixer m_52(.a(e_24_52), .b(e_46_52), .y(e_52_66));
	mixer m_53(.a(e_27_53), .b(e_50_53), .y(e_53_68));
	mixer m_54(.a(e_28_54), .b(e_54_55), .y(e_54_62));
	mixer m_55(.a(e_31_55), .b(e_54_55), .y(e_55_82));
	mixer m_56(.a(e_30_56), .b(e_41_56), .y(e_56_61));
	mixer m_57(.a(e_16_57), .b(e_42_57), .y(e_57_69));
	mixer m_58(.a(e_15_58), .b(e_48_58), .y(e_58_74));
	mixer m_59(.a(e_14_59), .b(e_51_59), .y(e_59_83));
	mixer m_60(.a(e_36_60), .b(e_60_61), .y(e_60_84));
	mixer m_61(.a(e_56_61), .b(e_60_61), .y(e_61_91));
	mixer m_62(.a(e_54_62), .b(e_62_83), .y(e_62_84));
	mixer m_63(.a(e_38_63), .b(e_63_70), .y(e_63_85));
	mixer m_64(.a(e_40_64), .b(e_64_65), .y(e_64_85));
	mixer m_65(.a(e_41_65), .b(e_64_65), .y(e_65_88));
	mixer m_66(.a(e_52_66), .b(e_66_69), .y(e_66_88));
	mixer m_67(.a(e_48_67), .b(e_67_76), .y(e_67_89));
	mixer m_68(.a(e_53_68), .b(e_68_78), .y(e_68_89));
	mixer m_69(.a(e_57_69), .b(e_66_69), .y(e_69_92));
	mixer m_70(.a(e_51_70), .b(e_63_70), .y(e_70_92));
	mixer m_71(.a(e_43_71), .b(e_71_80), .y(e_71_95));
	mixer m_72(.a(e_45_72), .b(e_72_73), .y(e_72_95));
	mixer m_73(.a(e_46_73), .b(e_72_73), .y(e_73_90));
	mixer m_74(.a(e_58_74), .b(e_74_75), .y(e_74_91));
	mixer m_75(.a(e_47_75), .b(e_74_75), .y(e_75_93));
	mixer m_76(.a(e_42_76), .b(e_67_76), .y(e_76_94));
	mixer m_77(.a(e_44_77), .b(e_77_82), .y(e_77_94));
	mixer m_78(.a(e_49_78), .b(e_68_78), .y(e_78_86));
	mixer m_79(.a(e_37_79), .b(e_79_81), .y(e_79_87));
	mixer m_80(.a(e_39_80), .b(e_71_80), .y(e_80_87));
	mixer m_81(.a(e_50_81), .b(e_79_81), .y(e_81_90));
	mixer m_82(.a(e_55_82), .b(e_77_82), .y(e_82_86));
	mixer m_83(.a(e_59_83), .b(e_62_83), .y(e_83_93));
	mixer m_84(.a(e_60_84), .b(e_62_84), .y(e_84_96));
	mixer m_85(.a(e_63_85), .b(e_64_85), .y(e_85_96));
	mixer m_86(.a(e_78_86), .b(e_82_86), .y(e_86_97));
	mixer m_87(.a(e_79_87), .b(e_80_87), .y(e_87_97));
	mixer m_88(.a(e_65_88), .b(e_66_88), .y(e_88_98));
	mixer m_89(.a(e_67_89), .b(e_68_89), .y(e_89_98));
	mixer m_90(.a(e_73_90), .b(e_81_90), .y(e_90_101));
	mixer m_91(.a(e_61_91), .b(e_74_91), .y(e_91_101));
	mixer m_92(.a(e_69_92), .b(e_70_92), .y(e_92_99));
	mixer m_93(.a(e_75_93), .b(e_83_93), .y(e_93_100));
	mixer m_94(.a(e_76_94), .b(e_77_94), .y(e_94_100));
	mixer m_95(.a(e_71_95), .b(e_72_95), .y(e_95_99));
	mixer m_96(.a(e_1_96), .b(e_84_96), .y(e_85_96));
	mixer m_97(.a(e_1_97), .b(e_86_97), .y(e_87_97));
	mixer m_98(.a(e_2_98), .b(e_88_98), .y(e_89_98));
	mixer m_99(.a(e_3_99), .b(e_92_99), .y(e_95_99));
	mixer m_100(.a(e_3_100), .b(e_93_100), .y(e_94_100));
	mixer m_101(.a(e_2_101), .b(e_90_101), .y(e_91_101));
wire e_0_1,
	e_0_2,
	e_0_3,
	e_1_96,
	e_1_97,
	e_2_98,
	e_2_101,
	e_3_99,
	e_3_100,
	e_4_12,
	e_4_14,
	e_4_15,
	e_5_13,
	e_5_16,
	e_5_17,
	e_6_18,
	e_6_19,
	e_6_33,
	e_7_21,
	e_7_23,
	e_7_34,
	e_8_20,
	e_8_25,
	e_8_32,
	e_9_22,
	e_9_24,
	e_9_26,
	e_10_27,
	e_10_31,
	e_10_35,
	e_11_28,
	e_11_29,
	e_11_30,
	e_12_13,
	e_12_36,
	e_13_38,
	e_14_35,
	e_14_59,
	e_15_34,
	e_15_58,
	e_16_33,
	e_16_57,
	e_17_32,
	e_17_41,
	e_18_31,
	e_18_37,
	e_19_30,
	e_19_46,
	e_20_21,
	e_20_49,
	e_21_39,
	e_22_23,
	e_22_51,
	e_23_45,
	e_24_27,
	e_24_52,
	e_25_29,
	e_25_44,
	e_26_28,
	e_26_40,
	e_27_53,
	e_28_54,
	e_29_47,
	e_30_56,
	e_31_55,
	e_32_48,
	e_33_43,
	e_34_50,
	e_35_42,
	e_36_37,
	e_36_60,
	e_37_79,
	e_38_39,
	e_38_63,
	e_39_80,
	e_40_49,
	e_40_64,
	e_41_56,
	e_41_65,
	e_42_57,
	e_42_76,
	e_43_44,
	e_43_71,
	e_44_77,
	e_45_47,
	e_45_72,
	e_46_52,
	e_46_73,
	e_47_75,
	e_48_58,
	e_48_67,
	e_49_78,
	e_50_53,
	e_50_81,
	e_51_59,
	e_51_70,
	e_52_66,
	e_53_68,
	e_54_55,
	e_54_62,
	e_55_82,
	e_56_61,
	e_57_69,
	e_58_74,
	e_59_83,
	e_60_61,
	e_60_84,
	e_61_91,
	e_62_83,
	e_62_84,
	e_63_70,
	e_63_85,
	e_64_65,
	e_64_85,
	e_65_88,
	e_66_69,
	e_66_88,
	e_67_76,
	e_67_89,
	e_68_78,
	e_68_89,
	e_69_92,
	e_70_92,
	e_71_80,
	e_71_95,
	e_72_73,
	e_72_95,
	e_73_90,
	e_74_75,
	e_74_91,
	e_75_93,
	e_76_94,
	e_77_82,
	e_77_94,
	e_78_86,
	e_79_81,
	e_79_87,
	e_80_87,
	e_81_90,
	e_82_86,
	e_83_93,
	e_84_96,
	e_85_96,
	e_86_97,
	e_87_97,
	e_88_98,
	e_89_98,
	e_90_101,
	e_91_101,
	e_92_99,
	e_93_100,
	e_94_100,
	e_95_99;
endmodule
