module fanout2_braid_8_512 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_1_7, output_1_0, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_0), .y(output_0_7));
wire output_2_7, output_2_0, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_0), .y(output_1_7));
wire output_3_7, output_3_0, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_0), .y(output_2_7));
wire output_4_7, output_4_0, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_0), .y(output_3_7));
wire output_5_7, output_5_0, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_0), .y(output_4_7));
wire output_6_7, output_6_0, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_0), .y(output_5_7));
wire output_7_7, output_7_0, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_0), .y(output_6_7));
wire output_8_7, output_8_0, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_0), .y(output_7_7));
wire output_1_8, output_1_1, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_1), .y(output_0_8));
wire output_2_8, output_2_1, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_1), .y(output_1_8));
wire output_3_8, output_3_1, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_1), .y(output_2_8));
wire output_4_8, output_4_1, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_1), .y(output_3_8));
wire output_5_8, output_5_1, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_1), .y(output_4_8));
wire output_6_8, output_6_1, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_1), .y(output_5_8));
wire output_7_8, output_7_1, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_1), .y(output_6_8));
wire output_8_8, output_8_1, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_1), .y(output_7_8));
wire output_1_9, output_1_2, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_2), .y(output_0_9));
wire output_2_9, output_2_2, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_2), .y(output_1_9));
wire output_3_9, output_3_2, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_2), .y(output_2_9));
wire output_4_9, output_4_2, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_2), .y(output_3_9));
wire output_5_9, output_5_2, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_2), .y(output_4_9));
wire output_6_9, output_6_2, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_2), .y(output_5_9));
wire output_7_9, output_7_2, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_2), .y(output_6_9));
wire output_8_9, output_8_2, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_2), .y(output_7_9));
wire output_1_10, output_1_3, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_3), .y(output_0_10));
wire output_2_10, output_2_3, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_3), .y(output_1_10));
wire output_3_10, output_3_3, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_3), .y(output_2_10));
wire output_4_10, output_4_3, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_3), .y(output_3_10));
wire output_5_10, output_5_3, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_3), .y(output_4_10));
wire output_6_10, output_6_3, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_3), .y(output_5_10));
wire output_7_10, output_7_3, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_3), .y(output_6_10));
wire output_8_10, output_8_3, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_3), .y(output_7_10));
wire output_1_11, output_1_4, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_4), .y(output_0_11));
wire output_2_11, output_2_4, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_4), .y(output_1_11));
wire output_3_11, output_3_4, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_4), .y(output_2_11));
wire output_4_11, output_4_4, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_4), .y(output_3_11));
wire output_5_11, output_5_4, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_4), .y(output_4_11));
wire output_6_11, output_6_4, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_4), .y(output_5_11));
wire output_7_11, output_7_4, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_4), .y(output_6_11));
wire output_8_11, output_8_4, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_4), .y(output_7_11));
wire output_1_12, output_1_5, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_5), .y(output_0_12));
wire output_2_12, output_2_5, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_5), .y(output_1_12));
wire output_3_12, output_3_5, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_5), .y(output_2_12));
wire output_4_12, output_4_5, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_5), .y(output_3_12));
wire output_5_12, output_5_5, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_5), .y(output_4_12));
wire output_6_12, output_6_5, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_5), .y(output_5_12));
wire output_7_12, output_7_5, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_5), .y(output_6_12));
wire output_8_12, output_8_5, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_5), .y(output_7_12));
wire output_1_13, output_1_6, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_6), .y(output_0_13));
wire output_2_13, output_2_6, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_6), .y(output_1_13));
wire output_3_13, output_3_6, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_6), .y(output_2_13));
wire output_4_13, output_4_6, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_6), .y(output_3_13));
wire output_5_13, output_5_6, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_6), .y(output_4_13));
wire output_6_13, output_6_6, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_6), .y(output_5_13));
wire output_7_13, output_7_6, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_6), .y(output_6_13));
wire output_8_13, output_8_6, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_6), .y(output_7_13));
wire output_1_14, output_1_7, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_7), .y(output_0_14));
wire output_2_14, output_2_7, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_7), .y(output_1_14));
wire output_3_14, output_3_7, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_7), .y(output_2_14));
wire output_4_14, output_4_7, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_7), .y(output_3_14));
wire output_5_14, output_5_7, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_7), .y(output_4_14));
wire output_6_14, output_6_7, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_7), .y(output_5_14));
wire output_7_14, output_7_7, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_7), .y(output_6_14));
wire output_8_14, output_8_7, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_7), .y(output_7_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
wire output_1_16, output_1_1, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_1), .y(output_0_16));
wire output_2_16, output_2_1, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_1), .y(output_1_16));
wire output_3_16, output_3_1, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_1), .y(output_2_16));
wire output_4_16, output_4_1, output_3_16;
mixer gate_output_3_16(.a(output_4_16), .b(output_4_1), .y(output_3_16));
wire output_5_16, output_5_1, output_4_16;
mixer gate_output_4_16(.a(output_5_16), .b(output_5_1), .y(output_4_16));
wire output_6_16, output_6_1, output_5_16;
mixer gate_output_5_16(.a(output_6_16), .b(output_6_1), .y(output_5_16));
wire output_7_16, output_7_1, output_6_16;
mixer gate_output_6_16(.a(output_7_16), .b(output_7_1), .y(output_6_16));
wire output_8_16, output_8_1, output_7_16;
mixer gate_output_7_16(.a(output_8_16), .b(output_8_1), .y(output_7_16));
wire output_1_17, output_1_2, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_2), .y(output_0_17));
wire output_2_17, output_2_2, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_2), .y(output_1_17));
wire output_3_17, output_3_2, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_2), .y(output_2_17));
wire output_4_17, output_4_2, output_3_17;
mixer gate_output_3_17(.a(output_4_17), .b(output_4_2), .y(output_3_17));
wire output_5_17, output_5_2, output_4_17;
mixer gate_output_4_17(.a(output_5_17), .b(output_5_2), .y(output_4_17));
wire output_6_17, output_6_2, output_5_17;
mixer gate_output_5_17(.a(output_6_17), .b(output_6_2), .y(output_5_17));
wire output_7_17, output_7_2, output_6_17;
mixer gate_output_6_17(.a(output_7_17), .b(output_7_2), .y(output_6_17));
wire output_8_17, output_8_2, output_7_17;
mixer gate_output_7_17(.a(output_8_17), .b(output_8_2), .y(output_7_17));
wire output_1_18, output_1_3, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_3), .y(output_0_18));
wire output_2_18, output_2_3, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_3), .y(output_1_18));
wire output_3_18, output_3_3, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_3), .y(output_2_18));
wire output_4_18, output_4_3, output_3_18;
mixer gate_output_3_18(.a(output_4_18), .b(output_4_3), .y(output_3_18));
wire output_5_18, output_5_3, output_4_18;
mixer gate_output_4_18(.a(output_5_18), .b(output_5_3), .y(output_4_18));
wire output_6_18, output_6_3, output_5_18;
mixer gate_output_5_18(.a(output_6_18), .b(output_6_3), .y(output_5_18));
wire output_7_18, output_7_3, output_6_18;
mixer gate_output_6_18(.a(output_7_18), .b(output_7_3), .y(output_6_18));
wire output_8_18, output_8_3, output_7_18;
mixer gate_output_7_18(.a(output_8_18), .b(output_8_3), .y(output_7_18));
wire output_1_19, output_1_4, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_4), .y(output_0_19));
wire output_2_19, output_2_4, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_4), .y(output_1_19));
wire output_3_19, output_3_4, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_4), .y(output_2_19));
wire output_4_19, output_4_4, output_3_19;
mixer gate_output_3_19(.a(output_4_19), .b(output_4_4), .y(output_3_19));
wire output_5_19, output_5_4, output_4_19;
mixer gate_output_4_19(.a(output_5_19), .b(output_5_4), .y(output_4_19));
wire output_6_19, output_6_4, output_5_19;
mixer gate_output_5_19(.a(output_6_19), .b(output_6_4), .y(output_5_19));
wire output_7_19, output_7_4, output_6_19;
mixer gate_output_6_19(.a(output_7_19), .b(output_7_4), .y(output_6_19));
wire output_8_19, output_8_4, output_7_19;
mixer gate_output_7_19(.a(output_8_19), .b(output_8_4), .y(output_7_19));
wire output_1_20, output_1_5, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_5), .y(output_0_20));
wire output_2_20, output_2_5, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_5), .y(output_1_20));
wire output_3_20, output_3_5, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_5), .y(output_2_20));
wire output_4_20, output_4_5, output_3_20;
mixer gate_output_3_20(.a(output_4_20), .b(output_4_5), .y(output_3_20));
wire output_5_20, output_5_5, output_4_20;
mixer gate_output_4_20(.a(output_5_20), .b(output_5_5), .y(output_4_20));
wire output_6_20, output_6_5, output_5_20;
mixer gate_output_5_20(.a(output_6_20), .b(output_6_5), .y(output_5_20));
wire output_7_20, output_7_5, output_6_20;
mixer gate_output_6_20(.a(output_7_20), .b(output_7_5), .y(output_6_20));
wire output_8_20, output_8_5, output_7_20;
mixer gate_output_7_20(.a(output_8_20), .b(output_8_5), .y(output_7_20));
wire output_1_21, output_1_6, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_6), .y(output_0_21));
wire output_2_21, output_2_6, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_6), .y(output_1_21));
wire output_3_21, output_3_6, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_6), .y(output_2_21));
wire output_4_21, output_4_6, output_3_21;
mixer gate_output_3_21(.a(output_4_21), .b(output_4_6), .y(output_3_21));
wire output_5_21, output_5_6, output_4_21;
mixer gate_output_4_21(.a(output_5_21), .b(output_5_6), .y(output_4_21));
wire output_6_21, output_6_6, output_5_21;
mixer gate_output_5_21(.a(output_6_21), .b(output_6_6), .y(output_5_21));
wire output_7_21, output_7_6, output_6_21;
mixer gate_output_6_21(.a(output_7_21), .b(output_7_6), .y(output_6_21));
wire output_8_21, output_8_6, output_7_21;
mixer gate_output_7_21(.a(output_8_21), .b(output_8_6), .y(output_7_21));
wire output_1_22, output_1_7, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_7), .y(output_0_22));
wire output_2_22, output_2_7, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_7), .y(output_1_22));
wire output_3_22, output_3_7, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_7), .y(output_2_22));
wire output_4_22, output_4_7, output_3_22;
mixer gate_output_3_22(.a(output_4_22), .b(output_4_7), .y(output_3_22));
wire output_5_22, output_5_7, output_4_22;
mixer gate_output_4_22(.a(output_5_22), .b(output_5_7), .y(output_4_22));
wire output_6_22, output_6_7, output_5_22;
mixer gate_output_5_22(.a(output_6_22), .b(output_6_7), .y(output_5_22));
wire output_7_22, output_7_7, output_6_22;
mixer gate_output_6_22(.a(output_7_22), .b(output_7_7), .y(output_6_22));
wire output_8_22, output_8_7, output_7_22;
mixer gate_output_7_22(.a(output_8_22), .b(output_8_7), .y(output_7_22));
wire output_1_23, output_1_0, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_0), .y(output_0_23));
wire output_2_23, output_2_0, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_0), .y(output_1_23));
wire output_3_23, output_3_0, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_0), .y(output_2_23));
wire output_4_23, output_4_0, output_3_23;
mixer gate_output_3_23(.a(output_4_23), .b(output_4_0), .y(output_3_23));
wire output_5_23, output_5_0, output_4_23;
mixer gate_output_4_23(.a(output_5_23), .b(output_5_0), .y(output_4_23));
wire output_6_23, output_6_0, output_5_23;
mixer gate_output_5_23(.a(output_6_23), .b(output_6_0), .y(output_5_23));
wire output_7_23, output_7_0, output_6_23;
mixer gate_output_6_23(.a(output_7_23), .b(output_7_0), .y(output_6_23));
wire output_8_23, output_8_0, output_7_23;
mixer gate_output_7_23(.a(output_8_23), .b(output_8_0), .y(output_7_23));
wire output_1_24, output_1_1, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_1), .y(output_0_24));
wire output_2_24, output_2_1, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_1), .y(output_1_24));
wire output_3_24, output_3_1, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_1), .y(output_2_24));
wire output_4_24, output_4_1, output_3_24;
mixer gate_output_3_24(.a(output_4_24), .b(output_4_1), .y(output_3_24));
wire output_5_24, output_5_1, output_4_24;
mixer gate_output_4_24(.a(output_5_24), .b(output_5_1), .y(output_4_24));
wire output_6_24, output_6_1, output_5_24;
mixer gate_output_5_24(.a(output_6_24), .b(output_6_1), .y(output_5_24));
wire output_7_24, output_7_1, output_6_24;
mixer gate_output_6_24(.a(output_7_24), .b(output_7_1), .y(output_6_24));
wire output_8_24, output_8_1, output_7_24;
mixer gate_output_7_24(.a(output_8_24), .b(output_8_1), .y(output_7_24));
wire output_1_25, output_1_2, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_2), .y(output_0_25));
wire output_2_25, output_2_2, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_2), .y(output_1_25));
wire output_3_25, output_3_2, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_2), .y(output_2_25));
wire output_4_25, output_4_2, output_3_25;
mixer gate_output_3_25(.a(output_4_25), .b(output_4_2), .y(output_3_25));
wire output_5_25, output_5_2, output_4_25;
mixer gate_output_4_25(.a(output_5_25), .b(output_5_2), .y(output_4_25));
wire output_6_25, output_6_2, output_5_25;
mixer gate_output_5_25(.a(output_6_25), .b(output_6_2), .y(output_5_25));
wire output_7_25, output_7_2, output_6_25;
mixer gate_output_6_25(.a(output_7_25), .b(output_7_2), .y(output_6_25));
wire output_8_25, output_8_2, output_7_25;
mixer gate_output_7_25(.a(output_8_25), .b(output_8_2), .y(output_7_25));
wire output_1_26, output_1_3, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_3), .y(output_0_26));
wire output_2_26, output_2_3, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_3), .y(output_1_26));
wire output_3_26, output_3_3, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_3), .y(output_2_26));
wire output_4_26, output_4_3, output_3_26;
mixer gate_output_3_26(.a(output_4_26), .b(output_4_3), .y(output_3_26));
wire output_5_26, output_5_3, output_4_26;
mixer gate_output_4_26(.a(output_5_26), .b(output_5_3), .y(output_4_26));
wire output_6_26, output_6_3, output_5_26;
mixer gate_output_5_26(.a(output_6_26), .b(output_6_3), .y(output_5_26));
wire output_7_26, output_7_3, output_6_26;
mixer gate_output_6_26(.a(output_7_26), .b(output_7_3), .y(output_6_26));
wire output_8_26, output_8_3, output_7_26;
mixer gate_output_7_26(.a(output_8_26), .b(output_8_3), .y(output_7_26));
wire output_1_27, output_1_4, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_4), .y(output_0_27));
wire output_2_27, output_2_4, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_4), .y(output_1_27));
wire output_3_27, output_3_4, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_4), .y(output_2_27));
wire output_4_27, output_4_4, output_3_27;
mixer gate_output_3_27(.a(output_4_27), .b(output_4_4), .y(output_3_27));
wire output_5_27, output_5_4, output_4_27;
mixer gate_output_4_27(.a(output_5_27), .b(output_5_4), .y(output_4_27));
wire output_6_27, output_6_4, output_5_27;
mixer gate_output_5_27(.a(output_6_27), .b(output_6_4), .y(output_5_27));
wire output_7_27, output_7_4, output_6_27;
mixer gate_output_6_27(.a(output_7_27), .b(output_7_4), .y(output_6_27));
wire output_8_27, output_8_4, output_7_27;
mixer gate_output_7_27(.a(output_8_27), .b(output_8_4), .y(output_7_27));
wire output_1_28, output_1_5, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_5), .y(output_0_28));
wire output_2_28, output_2_5, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_5), .y(output_1_28));
wire output_3_28, output_3_5, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_5), .y(output_2_28));
wire output_4_28, output_4_5, output_3_28;
mixer gate_output_3_28(.a(output_4_28), .b(output_4_5), .y(output_3_28));
wire output_5_28, output_5_5, output_4_28;
mixer gate_output_4_28(.a(output_5_28), .b(output_5_5), .y(output_4_28));
wire output_6_28, output_6_5, output_5_28;
mixer gate_output_5_28(.a(output_6_28), .b(output_6_5), .y(output_5_28));
wire output_7_28, output_7_5, output_6_28;
mixer gate_output_6_28(.a(output_7_28), .b(output_7_5), .y(output_6_28));
wire output_8_28, output_8_5, output_7_28;
mixer gate_output_7_28(.a(output_8_28), .b(output_8_5), .y(output_7_28));
wire output_1_29, output_1_6, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_6), .y(output_0_29));
wire output_2_29, output_2_6, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_6), .y(output_1_29));
wire output_3_29, output_3_6, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_6), .y(output_2_29));
wire output_4_29, output_4_6, output_3_29;
mixer gate_output_3_29(.a(output_4_29), .b(output_4_6), .y(output_3_29));
wire output_5_29, output_5_6, output_4_29;
mixer gate_output_4_29(.a(output_5_29), .b(output_5_6), .y(output_4_29));
wire output_6_29, output_6_6, output_5_29;
mixer gate_output_5_29(.a(output_6_29), .b(output_6_6), .y(output_5_29));
wire output_7_29, output_7_6, output_6_29;
mixer gate_output_6_29(.a(output_7_29), .b(output_7_6), .y(output_6_29));
wire output_8_29, output_8_6, output_7_29;
mixer gate_output_7_29(.a(output_8_29), .b(output_8_6), .y(output_7_29));
wire output_1_30, output_1_7, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_7), .y(output_0_30));
wire output_2_30, output_2_7, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_7), .y(output_1_30));
wire output_3_30, output_3_7, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_7), .y(output_2_30));
wire output_4_30, output_4_7, output_3_30;
mixer gate_output_3_30(.a(output_4_30), .b(output_4_7), .y(output_3_30));
wire output_5_30, output_5_7, output_4_30;
mixer gate_output_4_30(.a(output_5_30), .b(output_5_7), .y(output_4_30));
wire output_6_30, output_6_7, output_5_30;
mixer gate_output_5_30(.a(output_6_30), .b(output_6_7), .y(output_5_30));
wire output_7_30, output_7_7, output_6_30;
mixer gate_output_6_30(.a(output_7_30), .b(output_7_7), .y(output_6_30));
wire output_8_30, output_8_7, output_7_30;
mixer gate_output_7_30(.a(output_8_30), .b(output_8_7), .y(output_7_30));
wire output_1_31, output_1_0, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_0), .y(output_0_31));
wire output_2_31, output_2_0, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_0), .y(output_1_31));
wire output_3_31, output_3_0, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_0), .y(output_2_31));
wire output_4_31, output_4_0, output_3_31;
mixer gate_output_3_31(.a(output_4_31), .b(output_4_0), .y(output_3_31));
wire output_5_31, output_5_0, output_4_31;
mixer gate_output_4_31(.a(output_5_31), .b(output_5_0), .y(output_4_31));
wire output_6_31, output_6_0, output_5_31;
mixer gate_output_5_31(.a(output_6_31), .b(output_6_0), .y(output_5_31));
wire output_7_31, output_7_0, output_6_31;
mixer gate_output_6_31(.a(output_7_31), .b(output_7_0), .y(output_6_31));
wire output_8_31, output_8_0, output_7_31;
mixer gate_output_7_31(.a(output_8_31), .b(output_8_0), .y(output_7_31));
wire output_1_32, output_1_1, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_1), .y(output_0_32));
wire output_2_32, output_2_1, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_1), .y(output_1_32));
wire output_3_32, output_3_1, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_1), .y(output_2_32));
wire output_4_32, output_4_1, output_3_32;
mixer gate_output_3_32(.a(output_4_32), .b(output_4_1), .y(output_3_32));
wire output_5_32, output_5_1, output_4_32;
mixer gate_output_4_32(.a(output_5_32), .b(output_5_1), .y(output_4_32));
wire output_6_32, output_6_1, output_5_32;
mixer gate_output_5_32(.a(output_6_32), .b(output_6_1), .y(output_5_32));
wire output_7_32, output_7_1, output_6_32;
mixer gate_output_6_32(.a(output_7_32), .b(output_7_1), .y(output_6_32));
wire output_8_32, output_8_1, output_7_32;
mixer gate_output_7_32(.a(output_8_32), .b(output_8_1), .y(output_7_32));
wire output_1_33, output_1_2, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_2), .y(output_0_33));
wire output_2_33, output_2_2, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_2), .y(output_1_33));
wire output_3_33, output_3_2, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_2), .y(output_2_33));
wire output_4_33, output_4_2, output_3_33;
mixer gate_output_3_33(.a(output_4_33), .b(output_4_2), .y(output_3_33));
wire output_5_33, output_5_2, output_4_33;
mixer gate_output_4_33(.a(output_5_33), .b(output_5_2), .y(output_4_33));
wire output_6_33, output_6_2, output_5_33;
mixer gate_output_5_33(.a(output_6_33), .b(output_6_2), .y(output_5_33));
wire output_7_33, output_7_2, output_6_33;
mixer gate_output_6_33(.a(output_7_33), .b(output_7_2), .y(output_6_33));
wire output_8_33, output_8_2, output_7_33;
mixer gate_output_7_33(.a(output_8_33), .b(output_8_2), .y(output_7_33));
wire output_1_34, output_1_3, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_3), .y(output_0_34));
wire output_2_34, output_2_3, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_3), .y(output_1_34));
wire output_3_34, output_3_3, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_3), .y(output_2_34));
wire output_4_34, output_4_3, output_3_34;
mixer gate_output_3_34(.a(output_4_34), .b(output_4_3), .y(output_3_34));
wire output_5_34, output_5_3, output_4_34;
mixer gate_output_4_34(.a(output_5_34), .b(output_5_3), .y(output_4_34));
wire output_6_34, output_6_3, output_5_34;
mixer gate_output_5_34(.a(output_6_34), .b(output_6_3), .y(output_5_34));
wire output_7_34, output_7_3, output_6_34;
mixer gate_output_6_34(.a(output_7_34), .b(output_7_3), .y(output_6_34));
wire output_8_34, output_8_3, output_7_34;
mixer gate_output_7_34(.a(output_8_34), .b(output_8_3), .y(output_7_34));
wire output_1_35, output_1_4, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_4), .y(output_0_35));
wire output_2_35, output_2_4, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_4), .y(output_1_35));
wire output_3_35, output_3_4, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_4), .y(output_2_35));
wire output_4_35, output_4_4, output_3_35;
mixer gate_output_3_35(.a(output_4_35), .b(output_4_4), .y(output_3_35));
wire output_5_35, output_5_4, output_4_35;
mixer gate_output_4_35(.a(output_5_35), .b(output_5_4), .y(output_4_35));
wire output_6_35, output_6_4, output_5_35;
mixer gate_output_5_35(.a(output_6_35), .b(output_6_4), .y(output_5_35));
wire output_7_35, output_7_4, output_6_35;
mixer gate_output_6_35(.a(output_7_35), .b(output_7_4), .y(output_6_35));
wire output_8_35, output_8_4, output_7_35;
mixer gate_output_7_35(.a(output_8_35), .b(output_8_4), .y(output_7_35));
wire output_1_36, output_1_5, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_5), .y(output_0_36));
wire output_2_36, output_2_5, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_5), .y(output_1_36));
wire output_3_36, output_3_5, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_5), .y(output_2_36));
wire output_4_36, output_4_5, output_3_36;
mixer gate_output_3_36(.a(output_4_36), .b(output_4_5), .y(output_3_36));
wire output_5_36, output_5_5, output_4_36;
mixer gate_output_4_36(.a(output_5_36), .b(output_5_5), .y(output_4_36));
wire output_6_36, output_6_5, output_5_36;
mixer gate_output_5_36(.a(output_6_36), .b(output_6_5), .y(output_5_36));
wire output_7_36, output_7_5, output_6_36;
mixer gate_output_6_36(.a(output_7_36), .b(output_7_5), .y(output_6_36));
wire output_8_36, output_8_5, output_7_36;
mixer gate_output_7_36(.a(output_8_36), .b(output_8_5), .y(output_7_36));
wire output_1_37, output_1_6, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_6), .y(output_0_37));
wire output_2_37, output_2_6, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_6), .y(output_1_37));
wire output_3_37, output_3_6, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_6), .y(output_2_37));
wire output_4_37, output_4_6, output_3_37;
mixer gate_output_3_37(.a(output_4_37), .b(output_4_6), .y(output_3_37));
wire output_5_37, output_5_6, output_4_37;
mixer gate_output_4_37(.a(output_5_37), .b(output_5_6), .y(output_4_37));
wire output_6_37, output_6_6, output_5_37;
mixer gate_output_5_37(.a(output_6_37), .b(output_6_6), .y(output_5_37));
wire output_7_37, output_7_6, output_6_37;
mixer gate_output_6_37(.a(output_7_37), .b(output_7_6), .y(output_6_37));
wire output_8_37, output_8_6, output_7_37;
mixer gate_output_7_37(.a(output_8_37), .b(output_8_6), .y(output_7_37));
wire output_1_38, output_1_7, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_7), .y(output_0_38));
wire output_2_38, output_2_7, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_7), .y(output_1_38));
wire output_3_38, output_3_7, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_7), .y(output_2_38));
wire output_4_38, output_4_7, output_3_38;
mixer gate_output_3_38(.a(output_4_38), .b(output_4_7), .y(output_3_38));
wire output_5_38, output_5_7, output_4_38;
mixer gate_output_4_38(.a(output_5_38), .b(output_5_7), .y(output_4_38));
wire output_6_38, output_6_7, output_5_38;
mixer gate_output_5_38(.a(output_6_38), .b(output_6_7), .y(output_5_38));
wire output_7_38, output_7_7, output_6_38;
mixer gate_output_6_38(.a(output_7_38), .b(output_7_7), .y(output_6_38));
wire output_8_38, output_8_7, output_7_38;
mixer gate_output_7_38(.a(output_8_38), .b(output_8_7), .y(output_7_38));
wire output_1_39, output_1_0, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_0), .y(output_0_39));
wire output_2_39, output_2_0, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_0), .y(output_1_39));
wire output_3_39, output_3_0, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_0), .y(output_2_39));
wire output_4_39, output_4_0, output_3_39;
mixer gate_output_3_39(.a(output_4_39), .b(output_4_0), .y(output_3_39));
wire output_5_39, output_5_0, output_4_39;
mixer gate_output_4_39(.a(output_5_39), .b(output_5_0), .y(output_4_39));
wire output_6_39, output_6_0, output_5_39;
mixer gate_output_5_39(.a(output_6_39), .b(output_6_0), .y(output_5_39));
wire output_7_39, output_7_0, output_6_39;
mixer gate_output_6_39(.a(output_7_39), .b(output_7_0), .y(output_6_39));
wire output_8_39, output_8_0, output_7_39;
mixer gate_output_7_39(.a(output_8_39), .b(output_8_0), .y(output_7_39));
wire output_1_40, output_1_1, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_1), .y(output_0_40));
wire output_2_40, output_2_1, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_1), .y(output_1_40));
wire output_3_40, output_3_1, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_1), .y(output_2_40));
wire output_4_40, output_4_1, output_3_40;
mixer gate_output_3_40(.a(output_4_40), .b(output_4_1), .y(output_3_40));
wire output_5_40, output_5_1, output_4_40;
mixer gate_output_4_40(.a(output_5_40), .b(output_5_1), .y(output_4_40));
wire output_6_40, output_6_1, output_5_40;
mixer gate_output_5_40(.a(output_6_40), .b(output_6_1), .y(output_5_40));
wire output_7_40, output_7_1, output_6_40;
mixer gate_output_6_40(.a(output_7_40), .b(output_7_1), .y(output_6_40));
wire output_8_40, output_8_1, output_7_40;
mixer gate_output_7_40(.a(output_8_40), .b(output_8_1), .y(output_7_40));
wire output_1_41, output_1_2, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_2), .y(output_0_41));
wire output_2_41, output_2_2, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_2), .y(output_1_41));
wire output_3_41, output_3_2, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_2), .y(output_2_41));
wire output_4_41, output_4_2, output_3_41;
mixer gate_output_3_41(.a(output_4_41), .b(output_4_2), .y(output_3_41));
wire output_5_41, output_5_2, output_4_41;
mixer gate_output_4_41(.a(output_5_41), .b(output_5_2), .y(output_4_41));
wire output_6_41, output_6_2, output_5_41;
mixer gate_output_5_41(.a(output_6_41), .b(output_6_2), .y(output_5_41));
wire output_7_41, output_7_2, output_6_41;
mixer gate_output_6_41(.a(output_7_41), .b(output_7_2), .y(output_6_41));
wire output_8_41, output_8_2, output_7_41;
mixer gate_output_7_41(.a(output_8_41), .b(output_8_2), .y(output_7_41));
wire output_1_42, output_1_3, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_3), .y(output_0_42));
wire output_2_42, output_2_3, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_3), .y(output_1_42));
wire output_3_42, output_3_3, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_3), .y(output_2_42));
wire output_4_42, output_4_3, output_3_42;
mixer gate_output_3_42(.a(output_4_42), .b(output_4_3), .y(output_3_42));
wire output_5_42, output_5_3, output_4_42;
mixer gate_output_4_42(.a(output_5_42), .b(output_5_3), .y(output_4_42));
wire output_6_42, output_6_3, output_5_42;
mixer gate_output_5_42(.a(output_6_42), .b(output_6_3), .y(output_5_42));
wire output_7_42, output_7_3, output_6_42;
mixer gate_output_6_42(.a(output_7_42), .b(output_7_3), .y(output_6_42));
wire output_8_42, output_8_3, output_7_42;
mixer gate_output_7_42(.a(output_8_42), .b(output_8_3), .y(output_7_42));
wire output_1_43, output_1_4, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_4), .y(output_0_43));
wire output_2_43, output_2_4, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_4), .y(output_1_43));
wire output_3_43, output_3_4, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_4), .y(output_2_43));
wire output_4_43, output_4_4, output_3_43;
mixer gate_output_3_43(.a(output_4_43), .b(output_4_4), .y(output_3_43));
wire output_5_43, output_5_4, output_4_43;
mixer gate_output_4_43(.a(output_5_43), .b(output_5_4), .y(output_4_43));
wire output_6_43, output_6_4, output_5_43;
mixer gate_output_5_43(.a(output_6_43), .b(output_6_4), .y(output_5_43));
wire output_7_43, output_7_4, output_6_43;
mixer gate_output_6_43(.a(output_7_43), .b(output_7_4), .y(output_6_43));
wire output_8_43, output_8_4, output_7_43;
mixer gate_output_7_43(.a(output_8_43), .b(output_8_4), .y(output_7_43));
wire output_1_44, output_1_5, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_5), .y(output_0_44));
wire output_2_44, output_2_5, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_5), .y(output_1_44));
wire output_3_44, output_3_5, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_5), .y(output_2_44));
wire output_4_44, output_4_5, output_3_44;
mixer gate_output_3_44(.a(output_4_44), .b(output_4_5), .y(output_3_44));
wire output_5_44, output_5_5, output_4_44;
mixer gate_output_4_44(.a(output_5_44), .b(output_5_5), .y(output_4_44));
wire output_6_44, output_6_5, output_5_44;
mixer gate_output_5_44(.a(output_6_44), .b(output_6_5), .y(output_5_44));
wire output_7_44, output_7_5, output_6_44;
mixer gate_output_6_44(.a(output_7_44), .b(output_7_5), .y(output_6_44));
wire output_8_44, output_8_5, output_7_44;
mixer gate_output_7_44(.a(output_8_44), .b(output_8_5), .y(output_7_44));
wire output_1_45, output_1_6, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_6), .y(output_0_45));
wire output_2_45, output_2_6, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_6), .y(output_1_45));
wire output_3_45, output_3_6, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_6), .y(output_2_45));
wire output_4_45, output_4_6, output_3_45;
mixer gate_output_3_45(.a(output_4_45), .b(output_4_6), .y(output_3_45));
wire output_5_45, output_5_6, output_4_45;
mixer gate_output_4_45(.a(output_5_45), .b(output_5_6), .y(output_4_45));
wire output_6_45, output_6_6, output_5_45;
mixer gate_output_5_45(.a(output_6_45), .b(output_6_6), .y(output_5_45));
wire output_7_45, output_7_6, output_6_45;
mixer gate_output_6_45(.a(output_7_45), .b(output_7_6), .y(output_6_45));
wire output_8_45, output_8_6, output_7_45;
mixer gate_output_7_45(.a(output_8_45), .b(output_8_6), .y(output_7_45));
wire output_1_46, output_1_7, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_7), .y(output_0_46));
wire output_2_46, output_2_7, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_7), .y(output_1_46));
wire output_3_46, output_3_7, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_7), .y(output_2_46));
wire output_4_46, output_4_7, output_3_46;
mixer gate_output_3_46(.a(output_4_46), .b(output_4_7), .y(output_3_46));
wire output_5_46, output_5_7, output_4_46;
mixer gate_output_4_46(.a(output_5_46), .b(output_5_7), .y(output_4_46));
wire output_6_46, output_6_7, output_5_46;
mixer gate_output_5_46(.a(output_6_46), .b(output_6_7), .y(output_5_46));
wire output_7_46, output_7_7, output_6_46;
mixer gate_output_6_46(.a(output_7_46), .b(output_7_7), .y(output_6_46));
wire output_8_46, output_8_7, output_7_46;
mixer gate_output_7_46(.a(output_8_46), .b(output_8_7), .y(output_7_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_4_47, output_4_0, output_3_47;
mixer gate_output_3_47(.a(output_4_47), .b(output_4_0), .y(output_3_47));
wire output_5_47, output_5_0, output_4_47;
mixer gate_output_4_47(.a(output_5_47), .b(output_5_0), .y(output_4_47));
wire output_6_47, output_6_0, output_5_47;
mixer gate_output_5_47(.a(output_6_47), .b(output_6_0), .y(output_5_47));
wire output_7_47, output_7_0, output_6_47;
mixer gate_output_6_47(.a(output_7_47), .b(output_7_0), .y(output_6_47));
wire output_8_47, output_8_0, output_7_47;
mixer gate_output_7_47(.a(output_8_47), .b(output_8_0), .y(output_7_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_4_48, output_4_1, output_3_48;
mixer gate_output_3_48(.a(output_4_48), .b(output_4_1), .y(output_3_48));
wire output_5_48, output_5_1, output_4_48;
mixer gate_output_4_48(.a(output_5_48), .b(output_5_1), .y(output_4_48));
wire output_6_48, output_6_1, output_5_48;
mixer gate_output_5_48(.a(output_6_48), .b(output_6_1), .y(output_5_48));
wire output_7_48, output_7_1, output_6_48;
mixer gate_output_6_48(.a(output_7_48), .b(output_7_1), .y(output_6_48));
wire output_8_48, output_8_1, output_7_48;
mixer gate_output_7_48(.a(output_8_48), .b(output_8_1), .y(output_7_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_4_49, output_4_2, output_3_49;
mixer gate_output_3_49(.a(output_4_49), .b(output_4_2), .y(output_3_49));
wire output_5_49, output_5_2, output_4_49;
mixer gate_output_4_49(.a(output_5_49), .b(output_5_2), .y(output_4_49));
wire output_6_49, output_6_2, output_5_49;
mixer gate_output_5_49(.a(output_6_49), .b(output_6_2), .y(output_5_49));
wire output_7_49, output_7_2, output_6_49;
mixer gate_output_6_49(.a(output_7_49), .b(output_7_2), .y(output_6_49));
wire output_8_49, output_8_2, output_7_49;
mixer gate_output_7_49(.a(output_8_49), .b(output_8_2), .y(output_7_49));
wire output_1_50, output_1_3, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_3), .y(output_0_50));
wire output_2_50, output_2_3, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_3), .y(output_1_50));
wire output_3_50, output_3_3, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_3), .y(output_2_50));
wire output_4_50, output_4_3, output_3_50;
mixer gate_output_3_50(.a(output_4_50), .b(output_4_3), .y(output_3_50));
wire output_5_50, output_5_3, output_4_50;
mixer gate_output_4_50(.a(output_5_50), .b(output_5_3), .y(output_4_50));
wire output_6_50, output_6_3, output_5_50;
mixer gate_output_5_50(.a(output_6_50), .b(output_6_3), .y(output_5_50));
wire output_7_50, output_7_3, output_6_50;
mixer gate_output_6_50(.a(output_7_50), .b(output_7_3), .y(output_6_50));
wire output_8_50, output_8_3, output_7_50;
mixer gate_output_7_50(.a(output_8_50), .b(output_8_3), .y(output_7_50));
wire output_1_51, output_1_4, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_4), .y(output_0_51));
wire output_2_51, output_2_4, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_4), .y(output_1_51));
wire output_3_51, output_3_4, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_4), .y(output_2_51));
wire output_4_51, output_4_4, output_3_51;
mixer gate_output_3_51(.a(output_4_51), .b(output_4_4), .y(output_3_51));
wire output_5_51, output_5_4, output_4_51;
mixer gate_output_4_51(.a(output_5_51), .b(output_5_4), .y(output_4_51));
wire output_6_51, output_6_4, output_5_51;
mixer gate_output_5_51(.a(output_6_51), .b(output_6_4), .y(output_5_51));
wire output_7_51, output_7_4, output_6_51;
mixer gate_output_6_51(.a(output_7_51), .b(output_7_4), .y(output_6_51));
wire output_8_51, output_8_4, output_7_51;
mixer gate_output_7_51(.a(output_8_51), .b(output_8_4), .y(output_7_51));
wire output_1_52, output_1_5, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_5), .y(output_0_52));
wire output_2_52, output_2_5, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_5), .y(output_1_52));
wire output_3_52, output_3_5, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_5), .y(output_2_52));
wire output_4_52, output_4_5, output_3_52;
mixer gate_output_3_52(.a(output_4_52), .b(output_4_5), .y(output_3_52));
wire output_5_52, output_5_5, output_4_52;
mixer gate_output_4_52(.a(output_5_52), .b(output_5_5), .y(output_4_52));
wire output_6_52, output_6_5, output_5_52;
mixer gate_output_5_52(.a(output_6_52), .b(output_6_5), .y(output_5_52));
wire output_7_52, output_7_5, output_6_52;
mixer gate_output_6_52(.a(output_7_52), .b(output_7_5), .y(output_6_52));
wire output_8_52, output_8_5, output_7_52;
mixer gate_output_7_52(.a(output_8_52), .b(output_8_5), .y(output_7_52));
wire output_1_53, output_1_6, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_6), .y(output_0_53));
wire output_2_53, output_2_6, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_6), .y(output_1_53));
wire output_3_53, output_3_6, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_6), .y(output_2_53));
wire output_4_53, output_4_6, output_3_53;
mixer gate_output_3_53(.a(output_4_53), .b(output_4_6), .y(output_3_53));
wire output_5_53, output_5_6, output_4_53;
mixer gate_output_4_53(.a(output_5_53), .b(output_5_6), .y(output_4_53));
wire output_6_53, output_6_6, output_5_53;
mixer gate_output_5_53(.a(output_6_53), .b(output_6_6), .y(output_5_53));
wire output_7_53, output_7_6, output_6_53;
mixer gate_output_6_53(.a(output_7_53), .b(output_7_6), .y(output_6_53));
wire output_8_53, output_8_6, output_7_53;
mixer gate_output_7_53(.a(output_8_53), .b(output_8_6), .y(output_7_53));
wire output_1_54, output_1_7, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_7), .y(output_0_54));
wire output_2_54, output_2_7, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_7), .y(output_1_54));
wire output_3_54, output_3_7, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_7), .y(output_2_54));
wire output_4_54, output_4_7, output_3_54;
mixer gate_output_3_54(.a(output_4_54), .b(output_4_7), .y(output_3_54));
wire output_5_54, output_5_7, output_4_54;
mixer gate_output_4_54(.a(output_5_54), .b(output_5_7), .y(output_4_54));
wire output_6_54, output_6_7, output_5_54;
mixer gate_output_5_54(.a(output_6_54), .b(output_6_7), .y(output_5_54));
wire output_7_54, output_7_7, output_6_54;
mixer gate_output_6_54(.a(output_7_54), .b(output_7_7), .y(output_6_54));
wire output_8_54, output_8_7, output_7_54;
mixer gate_output_7_54(.a(output_8_54), .b(output_8_7), .y(output_7_54));
wire output_1_55, output_1_0, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_0), .y(output_0_55));
wire output_2_55, output_2_0, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_0), .y(output_1_55));
wire output_3_55, output_3_0, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_0), .y(output_2_55));
wire output_4_55, output_4_0, output_3_55;
mixer gate_output_3_55(.a(output_4_55), .b(output_4_0), .y(output_3_55));
wire output_5_55, output_5_0, output_4_55;
mixer gate_output_4_55(.a(output_5_55), .b(output_5_0), .y(output_4_55));
wire output_6_55, output_6_0, output_5_55;
mixer gate_output_5_55(.a(output_6_55), .b(output_6_0), .y(output_5_55));
wire output_7_55, output_7_0, output_6_55;
mixer gate_output_6_55(.a(output_7_55), .b(output_7_0), .y(output_6_55));
wire output_8_55, output_8_0, output_7_55;
mixer gate_output_7_55(.a(output_8_55), .b(output_8_0), .y(output_7_55));
wire output_1_56, output_1_1, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_1), .y(output_0_56));
wire output_2_56, output_2_1, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_1), .y(output_1_56));
wire output_3_56, output_3_1, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_1), .y(output_2_56));
wire output_4_56, output_4_1, output_3_56;
mixer gate_output_3_56(.a(output_4_56), .b(output_4_1), .y(output_3_56));
wire output_5_56, output_5_1, output_4_56;
mixer gate_output_4_56(.a(output_5_56), .b(output_5_1), .y(output_4_56));
wire output_6_56, output_6_1, output_5_56;
mixer gate_output_5_56(.a(output_6_56), .b(output_6_1), .y(output_5_56));
wire output_7_56, output_7_1, output_6_56;
mixer gate_output_6_56(.a(output_7_56), .b(output_7_1), .y(output_6_56));
wire output_8_56, output_8_1, output_7_56;
mixer gate_output_7_56(.a(output_8_56), .b(output_8_1), .y(output_7_56));
wire output_1_57, output_1_2, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_2), .y(output_0_57));
wire output_2_57, output_2_2, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_2), .y(output_1_57));
wire output_3_57, output_3_2, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_2), .y(output_2_57));
wire output_4_57, output_4_2, output_3_57;
mixer gate_output_3_57(.a(output_4_57), .b(output_4_2), .y(output_3_57));
wire output_5_57, output_5_2, output_4_57;
mixer gate_output_4_57(.a(output_5_57), .b(output_5_2), .y(output_4_57));
wire output_6_57, output_6_2, output_5_57;
mixer gate_output_5_57(.a(output_6_57), .b(output_6_2), .y(output_5_57));
wire output_7_57, output_7_2, output_6_57;
mixer gate_output_6_57(.a(output_7_57), .b(output_7_2), .y(output_6_57));
wire output_8_57, output_8_2, output_7_57;
mixer gate_output_7_57(.a(output_8_57), .b(output_8_2), .y(output_7_57));
wire output_1_58, output_1_3, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_3), .y(output_0_58));
wire output_2_58, output_2_3, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_3), .y(output_1_58));
wire output_3_58, output_3_3, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_3), .y(output_2_58));
wire output_4_58, output_4_3, output_3_58;
mixer gate_output_3_58(.a(output_4_58), .b(output_4_3), .y(output_3_58));
wire output_5_58, output_5_3, output_4_58;
mixer gate_output_4_58(.a(output_5_58), .b(output_5_3), .y(output_4_58));
wire output_6_58, output_6_3, output_5_58;
mixer gate_output_5_58(.a(output_6_58), .b(output_6_3), .y(output_5_58));
wire output_7_58, output_7_3, output_6_58;
mixer gate_output_6_58(.a(output_7_58), .b(output_7_3), .y(output_6_58));
wire output_8_58, output_8_3, output_7_58;
mixer gate_output_7_58(.a(output_8_58), .b(output_8_3), .y(output_7_58));
wire output_1_59, output_1_4, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_4), .y(output_0_59));
wire output_2_59, output_2_4, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_4), .y(output_1_59));
wire output_3_59, output_3_4, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_4), .y(output_2_59));
wire output_4_59, output_4_4, output_3_59;
mixer gate_output_3_59(.a(output_4_59), .b(output_4_4), .y(output_3_59));
wire output_5_59, output_5_4, output_4_59;
mixer gate_output_4_59(.a(output_5_59), .b(output_5_4), .y(output_4_59));
wire output_6_59, output_6_4, output_5_59;
mixer gate_output_5_59(.a(output_6_59), .b(output_6_4), .y(output_5_59));
wire output_7_59, output_7_4, output_6_59;
mixer gate_output_6_59(.a(output_7_59), .b(output_7_4), .y(output_6_59));
wire output_8_59, output_8_4, output_7_59;
mixer gate_output_7_59(.a(output_8_59), .b(output_8_4), .y(output_7_59));
wire output_1_60, output_1_5, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_5), .y(output_0_60));
wire output_2_60, output_2_5, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_5), .y(output_1_60));
wire output_3_60, output_3_5, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_5), .y(output_2_60));
wire output_4_60, output_4_5, output_3_60;
mixer gate_output_3_60(.a(output_4_60), .b(output_4_5), .y(output_3_60));
wire output_5_60, output_5_5, output_4_60;
mixer gate_output_4_60(.a(output_5_60), .b(output_5_5), .y(output_4_60));
wire output_6_60, output_6_5, output_5_60;
mixer gate_output_5_60(.a(output_6_60), .b(output_6_5), .y(output_5_60));
wire output_7_60, output_7_5, output_6_60;
mixer gate_output_6_60(.a(output_7_60), .b(output_7_5), .y(output_6_60));
wire output_8_60, output_8_5, output_7_60;
mixer gate_output_7_60(.a(output_8_60), .b(output_8_5), .y(output_7_60));
wire output_1_61, output_1_6, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_6), .y(output_0_61));
wire output_2_61, output_2_6, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_6), .y(output_1_61));
wire output_3_61, output_3_6, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_6), .y(output_2_61));
wire output_4_61, output_4_6, output_3_61;
mixer gate_output_3_61(.a(output_4_61), .b(output_4_6), .y(output_3_61));
wire output_5_61, output_5_6, output_4_61;
mixer gate_output_4_61(.a(output_5_61), .b(output_5_6), .y(output_4_61));
wire output_6_61, output_6_6, output_5_61;
mixer gate_output_5_61(.a(output_6_61), .b(output_6_6), .y(output_5_61));
wire output_7_61, output_7_6, output_6_61;
mixer gate_output_6_61(.a(output_7_61), .b(output_7_6), .y(output_6_61));
wire output_8_61, output_8_6, output_7_61;
mixer gate_output_7_61(.a(output_8_61), .b(output_8_6), .y(output_7_61));
wire output_1_62, output_1_7, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_7), .y(output_0_62));
wire output_2_62, output_2_7, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_7), .y(output_1_62));
wire output_3_62, output_3_7, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_7), .y(output_2_62));
wire output_4_62, output_4_7, output_3_62;
mixer gate_output_3_62(.a(output_4_62), .b(output_4_7), .y(output_3_62));
wire output_5_62, output_5_7, output_4_62;
mixer gate_output_4_62(.a(output_5_62), .b(output_5_7), .y(output_4_62));
wire output_6_62, output_6_7, output_5_62;
mixer gate_output_5_62(.a(output_6_62), .b(output_6_7), .y(output_5_62));
wire output_7_62, output_7_7, output_6_62;
mixer gate_output_6_62(.a(output_7_62), .b(output_7_7), .y(output_6_62));
wire output_8_62, output_8_7, output_7_62;
mixer gate_output_7_62(.a(output_8_62), .b(output_8_7), .y(output_7_62));
wire output_1_63, output_1_0, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_0), .y(output_0_63));
wire output_2_63, output_2_0, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_0), .y(output_1_63));
wire output_3_63, output_3_0, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_0), .y(output_2_63));
wire output_4_63, output_4_0, output_3_63;
mixer gate_output_3_63(.a(output_4_63), .b(output_4_0), .y(output_3_63));
wire output_5_63, output_5_0, output_4_63;
mixer gate_output_4_63(.a(output_5_63), .b(output_5_0), .y(output_4_63));
wire output_6_63, output_6_0, output_5_63;
mixer gate_output_5_63(.a(output_6_63), .b(output_6_0), .y(output_5_63));
wire output_7_63, output_7_0, output_6_63;
mixer gate_output_6_63(.a(output_7_63), .b(output_7_0), .y(output_6_63));
wire output_8_63, output_8_0, output_7_63;
mixer gate_output_7_63(.a(output_8_63), .b(output_8_0), .y(output_7_63));
wire output_1_64, output_1_1, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_1), .y(output_0_64));
wire output_2_64, output_2_1, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_1), .y(output_1_64));
wire output_3_64, output_3_1, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_1), .y(output_2_64));
wire output_4_64, output_4_1, output_3_64;
mixer gate_output_3_64(.a(output_4_64), .b(output_4_1), .y(output_3_64));
wire output_5_64, output_5_1, output_4_64;
mixer gate_output_4_64(.a(output_5_64), .b(output_5_1), .y(output_4_64));
wire output_6_64, output_6_1, output_5_64;
mixer gate_output_5_64(.a(output_6_64), .b(output_6_1), .y(output_5_64));
wire output_7_64, output_7_1, output_6_64;
mixer gate_output_6_64(.a(output_7_64), .b(output_7_1), .y(output_6_64));
wire output_8_64, output_8_1, output_7_64;
mixer gate_output_7_64(.a(output_8_64), .b(output_8_1), .y(output_7_64));
wire output_1_65, output_1_2, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_2), .y(output_0_65));
wire output_2_65, output_2_2, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_2), .y(output_1_65));
wire output_3_65, output_3_2, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_2), .y(output_2_65));
wire output_4_65, output_4_2, output_3_65;
mixer gate_output_3_65(.a(output_4_65), .b(output_4_2), .y(output_3_65));
wire output_5_65, output_5_2, output_4_65;
mixer gate_output_4_65(.a(output_5_65), .b(output_5_2), .y(output_4_65));
wire output_6_65, output_6_2, output_5_65;
mixer gate_output_5_65(.a(output_6_65), .b(output_6_2), .y(output_5_65));
wire output_7_65, output_7_2, output_6_65;
mixer gate_output_6_65(.a(output_7_65), .b(output_7_2), .y(output_6_65));
wire output_8_65, output_8_2, output_7_65;
mixer gate_output_7_65(.a(output_8_65), .b(output_8_2), .y(output_7_65));
wire output_1_66, output_1_3, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_3), .y(output_0_66));
wire output_2_66, output_2_3, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_3), .y(output_1_66));
wire output_3_66, output_3_3, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_3), .y(output_2_66));
wire output_4_66, output_4_3, output_3_66;
mixer gate_output_3_66(.a(output_4_66), .b(output_4_3), .y(output_3_66));
wire output_5_66, output_5_3, output_4_66;
mixer gate_output_4_66(.a(output_5_66), .b(output_5_3), .y(output_4_66));
wire output_6_66, output_6_3, output_5_66;
mixer gate_output_5_66(.a(output_6_66), .b(output_6_3), .y(output_5_66));
wire output_7_66, output_7_3, output_6_66;
mixer gate_output_6_66(.a(output_7_66), .b(output_7_3), .y(output_6_66));
wire output_8_66, output_8_3, output_7_66;
mixer gate_output_7_66(.a(output_8_66), .b(output_8_3), .y(output_7_66));
wire output_1_67, output_1_4, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_4), .y(output_0_67));
wire output_2_67, output_2_4, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_4), .y(output_1_67));
wire output_3_67, output_3_4, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_4), .y(output_2_67));
wire output_4_67, output_4_4, output_3_67;
mixer gate_output_3_67(.a(output_4_67), .b(output_4_4), .y(output_3_67));
wire output_5_67, output_5_4, output_4_67;
mixer gate_output_4_67(.a(output_5_67), .b(output_5_4), .y(output_4_67));
wire output_6_67, output_6_4, output_5_67;
mixer gate_output_5_67(.a(output_6_67), .b(output_6_4), .y(output_5_67));
wire output_7_67, output_7_4, output_6_67;
mixer gate_output_6_67(.a(output_7_67), .b(output_7_4), .y(output_6_67));
wire output_8_67, output_8_4, output_7_67;
mixer gate_output_7_67(.a(output_8_67), .b(output_8_4), .y(output_7_67));
wire output_1_68, output_1_5, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_5), .y(output_0_68));
wire output_2_68, output_2_5, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_5), .y(output_1_68));
wire output_3_68, output_3_5, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_5), .y(output_2_68));
wire output_4_68, output_4_5, output_3_68;
mixer gate_output_3_68(.a(output_4_68), .b(output_4_5), .y(output_3_68));
wire output_5_68, output_5_5, output_4_68;
mixer gate_output_4_68(.a(output_5_68), .b(output_5_5), .y(output_4_68));
wire output_6_68, output_6_5, output_5_68;
mixer gate_output_5_68(.a(output_6_68), .b(output_6_5), .y(output_5_68));
wire output_7_68, output_7_5, output_6_68;
mixer gate_output_6_68(.a(output_7_68), .b(output_7_5), .y(output_6_68));
wire output_8_68, output_8_5, output_7_68;
mixer gate_output_7_68(.a(output_8_68), .b(output_8_5), .y(output_7_68));
wire output_1_69, output_1_6, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_6), .y(output_0_69));
wire output_2_69, output_2_6, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_6), .y(output_1_69));
wire output_3_69, output_3_6, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_6), .y(output_2_69));
wire output_4_69, output_4_6, output_3_69;
mixer gate_output_3_69(.a(output_4_69), .b(output_4_6), .y(output_3_69));
wire output_5_69, output_5_6, output_4_69;
mixer gate_output_4_69(.a(output_5_69), .b(output_5_6), .y(output_4_69));
wire output_6_69, output_6_6, output_5_69;
mixer gate_output_5_69(.a(output_6_69), .b(output_6_6), .y(output_5_69));
wire output_7_69, output_7_6, output_6_69;
mixer gate_output_6_69(.a(output_7_69), .b(output_7_6), .y(output_6_69));
wire output_8_69, output_8_6, output_7_69;
mixer gate_output_7_69(.a(output_8_69), .b(output_8_6), .y(output_7_69));
wire output_1_70, output_1_7, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_7), .y(output_0_70));
wire output_2_70, output_2_7, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_7), .y(output_1_70));
wire output_3_70, output_3_7, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_7), .y(output_2_70));
wire output_4_70, output_4_7, output_3_70;
mixer gate_output_3_70(.a(output_4_70), .b(output_4_7), .y(output_3_70));
wire output_5_70, output_5_7, output_4_70;
mixer gate_output_4_70(.a(output_5_70), .b(output_5_7), .y(output_4_70));
wire output_6_70, output_6_7, output_5_70;
mixer gate_output_5_70(.a(output_6_70), .b(output_6_7), .y(output_5_70));
wire output_7_70, output_7_7, output_6_70;
mixer gate_output_6_70(.a(output_7_70), .b(output_7_7), .y(output_6_70));
wire output_8_70, output_8_7, output_7_70;
mixer gate_output_7_70(.a(output_8_70), .b(output_8_7), .y(output_7_70));
wire output_1_71, output_1_0, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_0), .y(output_0_71));
wire output_2_71, output_2_0, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_0), .y(output_1_71));
wire output_3_71, output_3_0, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_0), .y(output_2_71));
wire output_4_71, output_4_0, output_3_71;
mixer gate_output_3_71(.a(output_4_71), .b(output_4_0), .y(output_3_71));
wire output_5_71, output_5_0, output_4_71;
mixer gate_output_4_71(.a(output_5_71), .b(output_5_0), .y(output_4_71));
wire output_6_71, output_6_0, output_5_71;
mixer gate_output_5_71(.a(output_6_71), .b(output_6_0), .y(output_5_71));
wire output_7_71, output_7_0, output_6_71;
mixer gate_output_6_71(.a(output_7_71), .b(output_7_0), .y(output_6_71));
wire output_8_71, output_8_0, output_7_71;
mixer gate_output_7_71(.a(output_8_71), .b(output_8_0), .y(output_7_71));
wire output_1_72, output_1_1, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_1), .y(output_0_72));
wire output_2_72, output_2_1, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_1), .y(output_1_72));
wire output_3_72, output_3_1, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_1), .y(output_2_72));
wire output_4_72, output_4_1, output_3_72;
mixer gate_output_3_72(.a(output_4_72), .b(output_4_1), .y(output_3_72));
wire output_5_72, output_5_1, output_4_72;
mixer gate_output_4_72(.a(output_5_72), .b(output_5_1), .y(output_4_72));
wire output_6_72, output_6_1, output_5_72;
mixer gate_output_5_72(.a(output_6_72), .b(output_6_1), .y(output_5_72));
wire output_7_72, output_7_1, output_6_72;
mixer gate_output_6_72(.a(output_7_72), .b(output_7_1), .y(output_6_72));
wire output_8_72, output_8_1, output_7_72;
mixer gate_output_7_72(.a(output_8_72), .b(output_8_1), .y(output_7_72));
wire output_1_73, output_1_2, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_2), .y(output_0_73));
wire output_2_73, output_2_2, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_2), .y(output_1_73));
wire output_3_73, output_3_2, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_2), .y(output_2_73));
wire output_4_73, output_4_2, output_3_73;
mixer gate_output_3_73(.a(output_4_73), .b(output_4_2), .y(output_3_73));
wire output_5_73, output_5_2, output_4_73;
mixer gate_output_4_73(.a(output_5_73), .b(output_5_2), .y(output_4_73));
wire output_6_73, output_6_2, output_5_73;
mixer gate_output_5_73(.a(output_6_73), .b(output_6_2), .y(output_5_73));
wire output_7_73, output_7_2, output_6_73;
mixer gate_output_6_73(.a(output_7_73), .b(output_7_2), .y(output_6_73));
wire output_8_73, output_8_2, output_7_73;
mixer gate_output_7_73(.a(output_8_73), .b(output_8_2), .y(output_7_73));
wire output_1_74, output_1_3, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_3), .y(output_0_74));
wire output_2_74, output_2_3, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_3), .y(output_1_74));
wire output_3_74, output_3_3, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_3), .y(output_2_74));
wire output_4_74, output_4_3, output_3_74;
mixer gate_output_3_74(.a(output_4_74), .b(output_4_3), .y(output_3_74));
wire output_5_74, output_5_3, output_4_74;
mixer gate_output_4_74(.a(output_5_74), .b(output_5_3), .y(output_4_74));
wire output_6_74, output_6_3, output_5_74;
mixer gate_output_5_74(.a(output_6_74), .b(output_6_3), .y(output_5_74));
wire output_7_74, output_7_3, output_6_74;
mixer gate_output_6_74(.a(output_7_74), .b(output_7_3), .y(output_6_74));
wire output_8_74, output_8_3, output_7_74;
mixer gate_output_7_74(.a(output_8_74), .b(output_8_3), .y(output_7_74));
wire output_1_75, output_1_4, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_4), .y(output_0_75));
wire output_2_75, output_2_4, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_4), .y(output_1_75));
wire output_3_75, output_3_4, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_4), .y(output_2_75));
wire output_4_75, output_4_4, output_3_75;
mixer gate_output_3_75(.a(output_4_75), .b(output_4_4), .y(output_3_75));
wire output_5_75, output_5_4, output_4_75;
mixer gate_output_4_75(.a(output_5_75), .b(output_5_4), .y(output_4_75));
wire output_6_75, output_6_4, output_5_75;
mixer gate_output_5_75(.a(output_6_75), .b(output_6_4), .y(output_5_75));
wire output_7_75, output_7_4, output_6_75;
mixer gate_output_6_75(.a(output_7_75), .b(output_7_4), .y(output_6_75));
wire output_8_75, output_8_4, output_7_75;
mixer gate_output_7_75(.a(output_8_75), .b(output_8_4), .y(output_7_75));
wire output_1_76, output_1_5, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_5), .y(output_0_76));
wire output_2_76, output_2_5, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_5), .y(output_1_76));
wire output_3_76, output_3_5, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_5), .y(output_2_76));
wire output_4_76, output_4_5, output_3_76;
mixer gate_output_3_76(.a(output_4_76), .b(output_4_5), .y(output_3_76));
wire output_5_76, output_5_5, output_4_76;
mixer gate_output_4_76(.a(output_5_76), .b(output_5_5), .y(output_4_76));
wire output_6_76, output_6_5, output_5_76;
mixer gate_output_5_76(.a(output_6_76), .b(output_6_5), .y(output_5_76));
wire output_7_76, output_7_5, output_6_76;
mixer gate_output_6_76(.a(output_7_76), .b(output_7_5), .y(output_6_76));
wire output_8_76, output_8_5, output_7_76;
mixer gate_output_7_76(.a(output_8_76), .b(output_8_5), .y(output_7_76));
wire output_1_77, output_1_6, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_6), .y(output_0_77));
wire output_2_77, output_2_6, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_6), .y(output_1_77));
wire output_3_77, output_3_6, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_6), .y(output_2_77));
wire output_4_77, output_4_6, output_3_77;
mixer gate_output_3_77(.a(output_4_77), .b(output_4_6), .y(output_3_77));
wire output_5_77, output_5_6, output_4_77;
mixer gate_output_4_77(.a(output_5_77), .b(output_5_6), .y(output_4_77));
wire output_6_77, output_6_6, output_5_77;
mixer gate_output_5_77(.a(output_6_77), .b(output_6_6), .y(output_5_77));
wire output_7_77, output_7_6, output_6_77;
mixer gate_output_6_77(.a(output_7_77), .b(output_7_6), .y(output_6_77));
wire output_8_77, output_8_6, output_7_77;
mixer gate_output_7_77(.a(output_8_77), .b(output_8_6), .y(output_7_77));
wire output_1_78, output_1_7, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_7), .y(output_0_78));
wire output_2_78, output_2_7, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_7), .y(output_1_78));
wire output_3_78, output_3_7, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_7), .y(output_2_78));
wire output_4_78, output_4_7, output_3_78;
mixer gate_output_3_78(.a(output_4_78), .b(output_4_7), .y(output_3_78));
wire output_5_78, output_5_7, output_4_78;
mixer gate_output_4_78(.a(output_5_78), .b(output_5_7), .y(output_4_78));
wire output_6_78, output_6_7, output_5_78;
mixer gate_output_5_78(.a(output_6_78), .b(output_6_7), .y(output_5_78));
wire output_7_78, output_7_7, output_6_78;
mixer gate_output_6_78(.a(output_7_78), .b(output_7_7), .y(output_6_78));
wire output_8_78, output_8_7, output_7_78;
mixer gate_output_7_78(.a(output_8_78), .b(output_8_7), .y(output_7_78));
wire output_1_79, output_1_0, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_0), .y(output_0_79));
wire output_2_79, output_2_0, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_0), .y(output_1_79));
wire output_3_79, output_3_0, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_0), .y(output_2_79));
wire output_4_79, output_4_0, output_3_79;
mixer gate_output_3_79(.a(output_4_79), .b(output_4_0), .y(output_3_79));
wire output_5_79, output_5_0, output_4_79;
mixer gate_output_4_79(.a(output_5_79), .b(output_5_0), .y(output_4_79));
wire output_6_79, output_6_0, output_5_79;
mixer gate_output_5_79(.a(output_6_79), .b(output_6_0), .y(output_5_79));
wire output_7_79, output_7_0, output_6_79;
mixer gate_output_6_79(.a(output_7_79), .b(output_7_0), .y(output_6_79));
wire output_8_79, output_8_0, output_7_79;
mixer gate_output_7_79(.a(output_8_79), .b(output_8_0), .y(output_7_79));
wire output_1_80, output_1_1, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_1), .y(output_0_80));
wire output_2_80, output_2_1, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_1), .y(output_1_80));
wire output_3_80, output_3_1, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_1), .y(output_2_80));
wire output_4_80, output_4_1, output_3_80;
mixer gate_output_3_80(.a(output_4_80), .b(output_4_1), .y(output_3_80));
wire output_5_80, output_5_1, output_4_80;
mixer gate_output_4_80(.a(output_5_80), .b(output_5_1), .y(output_4_80));
wire output_6_80, output_6_1, output_5_80;
mixer gate_output_5_80(.a(output_6_80), .b(output_6_1), .y(output_5_80));
wire output_7_80, output_7_1, output_6_80;
mixer gate_output_6_80(.a(output_7_80), .b(output_7_1), .y(output_6_80));
wire output_8_80, output_8_1, output_7_80;
mixer gate_output_7_80(.a(output_8_80), .b(output_8_1), .y(output_7_80));
wire output_1_81, output_1_2, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_2), .y(output_0_81));
wire output_2_81, output_2_2, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_2), .y(output_1_81));
wire output_3_81, output_3_2, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_2), .y(output_2_81));
wire output_4_81, output_4_2, output_3_81;
mixer gate_output_3_81(.a(output_4_81), .b(output_4_2), .y(output_3_81));
wire output_5_81, output_5_2, output_4_81;
mixer gate_output_4_81(.a(output_5_81), .b(output_5_2), .y(output_4_81));
wire output_6_81, output_6_2, output_5_81;
mixer gate_output_5_81(.a(output_6_81), .b(output_6_2), .y(output_5_81));
wire output_7_81, output_7_2, output_6_81;
mixer gate_output_6_81(.a(output_7_81), .b(output_7_2), .y(output_6_81));
wire output_8_81, output_8_2, output_7_81;
mixer gate_output_7_81(.a(output_8_81), .b(output_8_2), .y(output_7_81));
wire output_1_82, output_1_3, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_3), .y(output_0_82));
wire output_2_82, output_2_3, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_3), .y(output_1_82));
wire output_3_82, output_3_3, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_3), .y(output_2_82));
wire output_4_82, output_4_3, output_3_82;
mixer gate_output_3_82(.a(output_4_82), .b(output_4_3), .y(output_3_82));
wire output_5_82, output_5_3, output_4_82;
mixer gate_output_4_82(.a(output_5_82), .b(output_5_3), .y(output_4_82));
wire output_6_82, output_6_3, output_5_82;
mixer gate_output_5_82(.a(output_6_82), .b(output_6_3), .y(output_5_82));
wire output_7_82, output_7_3, output_6_82;
mixer gate_output_6_82(.a(output_7_82), .b(output_7_3), .y(output_6_82));
wire output_8_82, output_8_3, output_7_82;
mixer gate_output_7_82(.a(output_8_82), .b(output_8_3), .y(output_7_82));
wire output_1_83, output_1_4, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_4), .y(output_0_83));
wire output_2_83, output_2_4, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_4), .y(output_1_83));
wire output_3_83, output_3_4, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_4), .y(output_2_83));
wire output_4_83, output_4_4, output_3_83;
mixer gate_output_3_83(.a(output_4_83), .b(output_4_4), .y(output_3_83));
wire output_5_83, output_5_4, output_4_83;
mixer gate_output_4_83(.a(output_5_83), .b(output_5_4), .y(output_4_83));
wire output_6_83, output_6_4, output_5_83;
mixer gate_output_5_83(.a(output_6_83), .b(output_6_4), .y(output_5_83));
wire output_7_83, output_7_4, output_6_83;
mixer gate_output_6_83(.a(output_7_83), .b(output_7_4), .y(output_6_83));
wire output_8_83, output_8_4, output_7_83;
mixer gate_output_7_83(.a(output_8_83), .b(output_8_4), .y(output_7_83));
wire output_1_84, output_1_5, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_5), .y(output_0_84));
wire output_2_84, output_2_5, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_5), .y(output_1_84));
wire output_3_84, output_3_5, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_5), .y(output_2_84));
wire output_4_84, output_4_5, output_3_84;
mixer gate_output_3_84(.a(output_4_84), .b(output_4_5), .y(output_3_84));
wire output_5_84, output_5_5, output_4_84;
mixer gate_output_4_84(.a(output_5_84), .b(output_5_5), .y(output_4_84));
wire output_6_84, output_6_5, output_5_84;
mixer gate_output_5_84(.a(output_6_84), .b(output_6_5), .y(output_5_84));
wire output_7_84, output_7_5, output_6_84;
mixer gate_output_6_84(.a(output_7_84), .b(output_7_5), .y(output_6_84));
wire output_8_84, output_8_5, output_7_84;
mixer gate_output_7_84(.a(output_8_84), .b(output_8_5), .y(output_7_84));
wire output_1_85, output_1_6, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_6), .y(output_0_85));
wire output_2_85, output_2_6, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_6), .y(output_1_85));
wire output_3_85, output_3_6, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_6), .y(output_2_85));
wire output_4_85, output_4_6, output_3_85;
mixer gate_output_3_85(.a(output_4_85), .b(output_4_6), .y(output_3_85));
wire output_5_85, output_5_6, output_4_85;
mixer gate_output_4_85(.a(output_5_85), .b(output_5_6), .y(output_4_85));
wire output_6_85, output_6_6, output_5_85;
mixer gate_output_5_85(.a(output_6_85), .b(output_6_6), .y(output_5_85));
wire output_7_85, output_7_6, output_6_85;
mixer gate_output_6_85(.a(output_7_85), .b(output_7_6), .y(output_6_85));
wire output_8_85, output_8_6, output_7_85;
mixer gate_output_7_85(.a(output_8_85), .b(output_8_6), .y(output_7_85));
wire output_1_86, output_1_7, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_7), .y(output_0_86));
wire output_2_86, output_2_7, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_7), .y(output_1_86));
wire output_3_86, output_3_7, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_7), .y(output_2_86));
wire output_4_86, output_4_7, output_3_86;
mixer gate_output_3_86(.a(output_4_86), .b(output_4_7), .y(output_3_86));
wire output_5_86, output_5_7, output_4_86;
mixer gate_output_4_86(.a(output_5_86), .b(output_5_7), .y(output_4_86));
wire output_6_86, output_6_7, output_5_86;
mixer gate_output_5_86(.a(output_6_86), .b(output_6_7), .y(output_5_86));
wire output_7_86, output_7_7, output_6_86;
mixer gate_output_6_86(.a(output_7_86), .b(output_7_7), .y(output_6_86));
wire output_8_86, output_8_7, output_7_86;
mixer gate_output_7_86(.a(output_8_86), .b(output_8_7), .y(output_7_86));
wire output_1_87, output_1_0, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_0), .y(output_0_87));
wire output_2_87, output_2_0, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_0), .y(output_1_87));
wire output_3_87, output_3_0, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_0), .y(output_2_87));
wire output_4_87, output_4_0, output_3_87;
mixer gate_output_3_87(.a(output_4_87), .b(output_4_0), .y(output_3_87));
wire output_5_87, output_5_0, output_4_87;
mixer gate_output_4_87(.a(output_5_87), .b(output_5_0), .y(output_4_87));
wire output_6_87, output_6_0, output_5_87;
mixer gate_output_5_87(.a(output_6_87), .b(output_6_0), .y(output_5_87));
wire output_7_87, output_7_0, output_6_87;
mixer gate_output_6_87(.a(output_7_87), .b(output_7_0), .y(output_6_87));
wire output_8_87, output_8_0, output_7_87;
mixer gate_output_7_87(.a(output_8_87), .b(output_8_0), .y(output_7_87));
wire output_1_88, output_1_1, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_1), .y(output_0_88));
wire output_2_88, output_2_1, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_1), .y(output_1_88));
wire output_3_88, output_3_1, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_1), .y(output_2_88));
wire output_4_88, output_4_1, output_3_88;
mixer gate_output_3_88(.a(output_4_88), .b(output_4_1), .y(output_3_88));
wire output_5_88, output_5_1, output_4_88;
mixer gate_output_4_88(.a(output_5_88), .b(output_5_1), .y(output_4_88));
wire output_6_88, output_6_1, output_5_88;
mixer gate_output_5_88(.a(output_6_88), .b(output_6_1), .y(output_5_88));
wire output_7_88, output_7_1, output_6_88;
mixer gate_output_6_88(.a(output_7_88), .b(output_7_1), .y(output_6_88));
wire output_8_88, output_8_1, output_7_88;
mixer gate_output_7_88(.a(output_8_88), .b(output_8_1), .y(output_7_88));
wire output_1_89, output_1_2, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_2), .y(output_0_89));
wire output_2_89, output_2_2, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_2), .y(output_1_89));
wire output_3_89, output_3_2, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_2), .y(output_2_89));
wire output_4_89, output_4_2, output_3_89;
mixer gate_output_3_89(.a(output_4_89), .b(output_4_2), .y(output_3_89));
wire output_5_89, output_5_2, output_4_89;
mixer gate_output_4_89(.a(output_5_89), .b(output_5_2), .y(output_4_89));
wire output_6_89, output_6_2, output_5_89;
mixer gate_output_5_89(.a(output_6_89), .b(output_6_2), .y(output_5_89));
wire output_7_89, output_7_2, output_6_89;
mixer gate_output_6_89(.a(output_7_89), .b(output_7_2), .y(output_6_89));
wire output_8_89, output_8_2, output_7_89;
mixer gate_output_7_89(.a(output_8_89), .b(output_8_2), .y(output_7_89));
wire output_1_90, output_1_3, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_3), .y(output_0_90));
wire output_2_90, output_2_3, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_3), .y(output_1_90));
wire output_3_90, output_3_3, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_3), .y(output_2_90));
wire output_4_90, output_4_3, output_3_90;
mixer gate_output_3_90(.a(output_4_90), .b(output_4_3), .y(output_3_90));
wire output_5_90, output_5_3, output_4_90;
mixer gate_output_4_90(.a(output_5_90), .b(output_5_3), .y(output_4_90));
wire output_6_90, output_6_3, output_5_90;
mixer gate_output_5_90(.a(output_6_90), .b(output_6_3), .y(output_5_90));
wire output_7_90, output_7_3, output_6_90;
mixer gate_output_6_90(.a(output_7_90), .b(output_7_3), .y(output_6_90));
wire output_8_90, output_8_3, output_7_90;
mixer gate_output_7_90(.a(output_8_90), .b(output_8_3), .y(output_7_90));
wire output_1_91, output_1_4, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_4), .y(output_0_91));
wire output_2_91, output_2_4, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_4), .y(output_1_91));
wire output_3_91, output_3_4, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_4), .y(output_2_91));
wire output_4_91, output_4_4, output_3_91;
mixer gate_output_3_91(.a(output_4_91), .b(output_4_4), .y(output_3_91));
wire output_5_91, output_5_4, output_4_91;
mixer gate_output_4_91(.a(output_5_91), .b(output_5_4), .y(output_4_91));
wire output_6_91, output_6_4, output_5_91;
mixer gate_output_5_91(.a(output_6_91), .b(output_6_4), .y(output_5_91));
wire output_7_91, output_7_4, output_6_91;
mixer gate_output_6_91(.a(output_7_91), .b(output_7_4), .y(output_6_91));
wire output_8_91, output_8_4, output_7_91;
mixer gate_output_7_91(.a(output_8_91), .b(output_8_4), .y(output_7_91));
wire output_1_92, output_1_5, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_5), .y(output_0_92));
wire output_2_92, output_2_5, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_5), .y(output_1_92));
wire output_3_92, output_3_5, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_5), .y(output_2_92));
wire output_4_92, output_4_5, output_3_92;
mixer gate_output_3_92(.a(output_4_92), .b(output_4_5), .y(output_3_92));
wire output_5_92, output_5_5, output_4_92;
mixer gate_output_4_92(.a(output_5_92), .b(output_5_5), .y(output_4_92));
wire output_6_92, output_6_5, output_5_92;
mixer gate_output_5_92(.a(output_6_92), .b(output_6_5), .y(output_5_92));
wire output_7_92, output_7_5, output_6_92;
mixer gate_output_6_92(.a(output_7_92), .b(output_7_5), .y(output_6_92));
wire output_8_92, output_8_5, output_7_92;
mixer gate_output_7_92(.a(output_8_92), .b(output_8_5), .y(output_7_92));
wire output_1_93, output_1_6, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_6), .y(output_0_93));
wire output_2_93, output_2_6, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_6), .y(output_1_93));
wire output_3_93, output_3_6, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_6), .y(output_2_93));
wire output_4_93, output_4_6, output_3_93;
mixer gate_output_3_93(.a(output_4_93), .b(output_4_6), .y(output_3_93));
wire output_5_93, output_5_6, output_4_93;
mixer gate_output_4_93(.a(output_5_93), .b(output_5_6), .y(output_4_93));
wire output_6_93, output_6_6, output_5_93;
mixer gate_output_5_93(.a(output_6_93), .b(output_6_6), .y(output_5_93));
wire output_7_93, output_7_6, output_6_93;
mixer gate_output_6_93(.a(output_7_93), .b(output_7_6), .y(output_6_93));
wire output_8_93, output_8_6, output_7_93;
mixer gate_output_7_93(.a(output_8_93), .b(output_8_6), .y(output_7_93));
wire output_1_94, output_1_7, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_7), .y(output_0_94));
wire output_2_94, output_2_7, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_7), .y(output_1_94));
wire output_3_94, output_3_7, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_7), .y(output_2_94));
wire output_4_94, output_4_7, output_3_94;
mixer gate_output_3_94(.a(output_4_94), .b(output_4_7), .y(output_3_94));
wire output_5_94, output_5_7, output_4_94;
mixer gate_output_4_94(.a(output_5_94), .b(output_5_7), .y(output_4_94));
wire output_6_94, output_6_7, output_5_94;
mixer gate_output_5_94(.a(output_6_94), .b(output_6_7), .y(output_5_94));
wire output_7_94, output_7_7, output_6_94;
mixer gate_output_6_94(.a(output_7_94), .b(output_7_7), .y(output_6_94));
wire output_8_94, output_8_7, output_7_94;
mixer gate_output_7_94(.a(output_8_94), .b(output_8_7), .y(output_7_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_4_95, output_4_0, output_3_95;
mixer gate_output_3_95(.a(output_4_95), .b(output_4_0), .y(output_3_95));
wire output_5_95, output_5_0, output_4_95;
mixer gate_output_4_95(.a(output_5_95), .b(output_5_0), .y(output_4_95));
wire output_6_95, output_6_0, output_5_95;
mixer gate_output_5_95(.a(output_6_95), .b(output_6_0), .y(output_5_95));
wire output_7_95, output_7_0, output_6_95;
mixer gate_output_6_95(.a(output_7_95), .b(output_7_0), .y(output_6_95));
wire output_8_95, output_8_0, output_7_95;
mixer gate_output_7_95(.a(output_8_95), .b(output_8_0), .y(output_7_95));
wire output_1_96, output_1_1, output_0_96;
mixer gate_output_0_96(.a(output_1_96), .b(output_1_1), .y(output_0_96));
wire output_2_96, output_2_1, output_1_96;
mixer gate_output_1_96(.a(output_2_96), .b(output_2_1), .y(output_1_96));
wire output_3_96, output_3_1, output_2_96;
mixer gate_output_2_96(.a(output_3_96), .b(output_3_1), .y(output_2_96));
wire output_4_96, output_4_1, output_3_96;
mixer gate_output_3_96(.a(output_4_96), .b(output_4_1), .y(output_3_96));
wire output_5_96, output_5_1, output_4_96;
mixer gate_output_4_96(.a(output_5_96), .b(output_5_1), .y(output_4_96));
wire output_6_96, output_6_1, output_5_96;
mixer gate_output_5_96(.a(output_6_96), .b(output_6_1), .y(output_5_96));
wire output_7_96, output_7_1, output_6_96;
mixer gate_output_6_96(.a(output_7_96), .b(output_7_1), .y(output_6_96));
wire output_8_96, output_8_1, output_7_96;
mixer gate_output_7_96(.a(output_8_96), .b(output_8_1), .y(output_7_96));
wire output_1_97, output_1_2, output_0_97;
mixer gate_output_0_97(.a(output_1_97), .b(output_1_2), .y(output_0_97));
wire output_2_97, output_2_2, output_1_97;
mixer gate_output_1_97(.a(output_2_97), .b(output_2_2), .y(output_1_97));
wire output_3_97, output_3_2, output_2_97;
mixer gate_output_2_97(.a(output_3_97), .b(output_3_2), .y(output_2_97));
wire output_4_97, output_4_2, output_3_97;
mixer gate_output_3_97(.a(output_4_97), .b(output_4_2), .y(output_3_97));
wire output_5_97, output_5_2, output_4_97;
mixer gate_output_4_97(.a(output_5_97), .b(output_5_2), .y(output_4_97));
wire output_6_97, output_6_2, output_5_97;
mixer gate_output_5_97(.a(output_6_97), .b(output_6_2), .y(output_5_97));
wire output_7_97, output_7_2, output_6_97;
mixer gate_output_6_97(.a(output_7_97), .b(output_7_2), .y(output_6_97));
wire output_8_97, output_8_2, output_7_97;
mixer gate_output_7_97(.a(output_8_97), .b(output_8_2), .y(output_7_97));
wire output_1_98, output_1_3, output_0_98;
mixer gate_output_0_98(.a(output_1_98), .b(output_1_3), .y(output_0_98));
wire output_2_98, output_2_3, output_1_98;
mixer gate_output_1_98(.a(output_2_98), .b(output_2_3), .y(output_1_98));
wire output_3_98, output_3_3, output_2_98;
mixer gate_output_2_98(.a(output_3_98), .b(output_3_3), .y(output_2_98));
wire output_4_98, output_4_3, output_3_98;
mixer gate_output_3_98(.a(output_4_98), .b(output_4_3), .y(output_3_98));
wire output_5_98, output_5_3, output_4_98;
mixer gate_output_4_98(.a(output_5_98), .b(output_5_3), .y(output_4_98));
wire output_6_98, output_6_3, output_5_98;
mixer gate_output_5_98(.a(output_6_98), .b(output_6_3), .y(output_5_98));
wire output_7_98, output_7_3, output_6_98;
mixer gate_output_6_98(.a(output_7_98), .b(output_7_3), .y(output_6_98));
wire output_8_98, output_8_3, output_7_98;
mixer gate_output_7_98(.a(output_8_98), .b(output_8_3), .y(output_7_98));
wire output_1_99, output_1_4, output_0_99;
mixer gate_output_0_99(.a(output_1_99), .b(output_1_4), .y(output_0_99));
wire output_2_99, output_2_4, output_1_99;
mixer gate_output_1_99(.a(output_2_99), .b(output_2_4), .y(output_1_99));
wire output_3_99, output_3_4, output_2_99;
mixer gate_output_2_99(.a(output_3_99), .b(output_3_4), .y(output_2_99));
wire output_4_99, output_4_4, output_3_99;
mixer gate_output_3_99(.a(output_4_99), .b(output_4_4), .y(output_3_99));
wire output_5_99, output_5_4, output_4_99;
mixer gate_output_4_99(.a(output_5_99), .b(output_5_4), .y(output_4_99));
wire output_6_99, output_6_4, output_5_99;
mixer gate_output_5_99(.a(output_6_99), .b(output_6_4), .y(output_5_99));
wire output_7_99, output_7_4, output_6_99;
mixer gate_output_6_99(.a(output_7_99), .b(output_7_4), .y(output_6_99));
wire output_8_99, output_8_4, output_7_99;
mixer gate_output_7_99(.a(output_8_99), .b(output_8_4), .y(output_7_99));
wire output_1_100, output_1_5, output_0_100;
mixer gate_output_0_100(.a(output_1_100), .b(output_1_5), .y(output_0_100));
wire output_2_100, output_2_5, output_1_100;
mixer gate_output_1_100(.a(output_2_100), .b(output_2_5), .y(output_1_100));
wire output_3_100, output_3_5, output_2_100;
mixer gate_output_2_100(.a(output_3_100), .b(output_3_5), .y(output_2_100));
wire output_4_100, output_4_5, output_3_100;
mixer gate_output_3_100(.a(output_4_100), .b(output_4_5), .y(output_3_100));
wire output_5_100, output_5_5, output_4_100;
mixer gate_output_4_100(.a(output_5_100), .b(output_5_5), .y(output_4_100));
wire output_6_100, output_6_5, output_5_100;
mixer gate_output_5_100(.a(output_6_100), .b(output_6_5), .y(output_5_100));
wire output_7_100, output_7_5, output_6_100;
mixer gate_output_6_100(.a(output_7_100), .b(output_7_5), .y(output_6_100));
wire output_8_100, output_8_5, output_7_100;
mixer gate_output_7_100(.a(output_8_100), .b(output_8_5), .y(output_7_100));
wire output_1_101, output_1_6, output_0_101;
mixer gate_output_0_101(.a(output_1_101), .b(output_1_6), .y(output_0_101));
wire output_2_101, output_2_6, output_1_101;
mixer gate_output_1_101(.a(output_2_101), .b(output_2_6), .y(output_1_101));
wire output_3_101, output_3_6, output_2_101;
mixer gate_output_2_101(.a(output_3_101), .b(output_3_6), .y(output_2_101));
wire output_4_101, output_4_6, output_3_101;
mixer gate_output_3_101(.a(output_4_101), .b(output_4_6), .y(output_3_101));
wire output_5_101, output_5_6, output_4_101;
mixer gate_output_4_101(.a(output_5_101), .b(output_5_6), .y(output_4_101));
wire output_6_101, output_6_6, output_5_101;
mixer gate_output_5_101(.a(output_6_101), .b(output_6_6), .y(output_5_101));
wire output_7_101, output_7_6, output_6_101;
mixer gate_output_6_101(.a(output_7_101), .b(output_7_6), .y(output_6_101));
wire output_8_101, output_8_6, output_7_101;
mixer gate_output_7_101(.a(output_8_101), .b(output_8_6), .y(output_7_101));
wire output_1_102, output_1_7, output_0_102;
mixer gate_output_0_102(.a(output_1_102), .b(output_1_7), .y(output_0_102));
wire output_2_102, output_2_7, output_1_102;
mixer gate_output_1_102(.a(output_2_102), .b(output_2_7), .y(output_1_102));
wire output_3_102, output_3_7, output_2_102;
mixer gate_output_2_102(.a(output_3_102), .b(output_3_7), .y(output_2_102));
wire output_4_102, output_4_7, output_3_102;
mixer gate_output_3_102(.a(output_4_102), .b(output_4_7), .y(output_3_102));
wire output_5_102, output_5_7, output_4_102;
mixer gate_output_4_102(.a(output_5_102), .b(output_5_7), .y(output_4_102));
wire output_6_102, output_6_7, output_5_102;
mixer gate_output_5_102(.a(output_6_102), .b(output_6_7), .y(output_5_102));
wire output_7_102, output_7_7, output_6_102;
mixer gate_output_6_102(.a(output_7_102), .b(output_7_7), .y(output_6_102));
wire output_8_102, output_8_7, output_7_102;
mixer gate_output_7_102(.a(output_8_102), .b(output_8_7), .y(output_7_102));
wire output_1_103, output_1_0, output_0_103;
mixer gate_output_0_103(.a(output_1_103), .b(output_1_0), .y(output_0_103));
wire output_2_103, output_2_0, output_1_103;
mixer gate_output_1_103(.a(output_2_103), .b(output_2_0), .y(output_1_103));
wire output_3_103, output_3_0, output_2_103;
mixer gate_output_2_103(.a(output_3_103), .b(output_3_0), .y(output_2_103));
wire output_4_103, output_4_0, output_3_103;
mixer gate_output_3_103(.a(output_4_103), .b(output_4_0), .y(output_3_103));
wire output_5_103, output_5_0, output_4_103;
mixer gate_output_4_103(.a(output_5_103), .b(output_5_0), .y(output_4_103));
wire output_6_103, output_6_0, output_5_103;
mixer gate_output_5_103(.a(output_6_103), .b(output_6_0), .y(output_5_103));
wire output_7_103, output_7_0, output_6_103;
mixer gate_output_6_103(.a(output_7_103), .b(output_7_0), .y(output_6_103));
wire output_8_103, output_8_0, output_7_103;
mixer gate_output_7_103(.a(output_8_103), .b(output_8_0), .y(output_7_103));
wire output_1_104, output_1_1, output_0_104;
mixer gate_output_0_104(.a(output_1_104), .b(output_1_1), .y(output_0_104));
wire output_2_104, output_2_1, output_1_104;
mixer gate_output_1_104(.a(output_2_104), .b(output_2_1), .y(output_1_104));
wire output_3_104, output_3_1, output_2_104;
mixer gate_output_2_104(.a(output_3_104), .b(output_3_1), .y(output_2_104));
wire output_4_104, output_4_1, output_3_104;
mixer gate_output_3_104(.a(output_4_104), .b(output_4_1), .y(output_3_104));
wire output_5_104, output_5_1, output_4_104;
mixer gate_output_4_104(.a(output_5_104), .b(output_5_1), .y(output_4_104));
wire output_6_104, output_6_1, output_5_104;
mixer gate_output_5_104(.a(output_6_104), .b(output_6_1), .y(output_5_104));
wire output_7_104, output_7_1, output_6_104;
mixer gate_output_6_104(.a(output_7_104), .b(output_7_1), .y(output_6_104));
wire output_8_104, output_8_1, output_7_104;
mixer gate_output_7_104(.a(output_8_104), .b(output_8_1), .y(output_7_104));
wire output_1_105, output_1_2, output_0_105;
mixer gate_output_0_105(.a(output_1_105), .b(output_1_2), .y(output_0_105));
wire output_2_105, output_2_2, output_1_105;
mixer gate_output_1_105(.a(output_2_105), .b(output_2_2), .y(output_1_105));
wire output_3_105, output_3_2, output_2_105;
mixer gate_output_2_105(.a(output_3_105), .b(output_3_2), .y(output_2_105));
wire output_4_105, output_4_2, output_3_105;
mixer gate_output_3_105(.a(output_4_105), .b(output_4_2), .y(output_3_105));
wire output_5_105, output_5_2, output_4_105;
mixer gate_output_4_105(.a(output_5_105), .b(output_5_2), .y(output_4_105));
wire output_6_105, output_6_2, output_5_105;
mixer gate_output_5_105(.a(output_6_105), .b(output_6_2), .y(output_5_105));
wire output_7_105, output_7_2, output_6_105;
mixer gate_output_6_105(.a(output_7_105), .b(output_7_2), .y(output_6_105));
wire output_8_105, output_8_2, output_7_105;
mixer gate_output_7_105(.a(output_8_105), .b(output_8_2), .y(output_7_105));
wire output_1_106, output_1_3, output_0_106;
mixer gate_output_0_106(.a(output_1_106), .b(output_1_3), .y(output_0_106));
wire output_2_106, output_2_3, output_1_106;
mixer gate_output_1_106(.a(output_2_106), .b(output_2_3), .y(output_1_106));
wire output_3_106, output_3_3, output_2_106;
mixer gate_output_2_106(.a(output_3_106), .b(output_3_3), .y(output_2_106));
wire output_4_106, output_4_3, output_3_106;
mixer gate_output_3_106(.a(output_4_106), .b(output_4_3), .y(output_3_106));
wire output_5_106, output_5_3, output_4_106;
mixer gate_output_4_106(.a(output_5_106), .b(output_5_3), .y(output_4_106));
wire output_6_106, output_6_3, output_5_106;
mixer gate_output_5_106(.a(output_6_106), .b(output_6_3), .y(output_5_106));
wire output_7_106, output_7_3, output_6_106;
mixer gate_output_6_106(.a(output_7_106), .b(output_7_3), .y(output_6_106));
wire output_8_106, output_8_3, output_7_106;
mixer gate_output_7_106(.a(output_8_106), .b(output_8_3), .y(output_7_106));
wire output_1_107, output_1_4, output_0_107;
mixer gate_output_0_107(.a(output_1_107), .b(output_1_4), .y(output_0_107));
wire output_2_107, output_2_4, output_1_107;
mixer gate_output_1_107(.a(output_2_107), .b(output_2_4), .y(output_1_107));
wire output_3_107, output_3_4, output_2_107;
mixer gate_output_2_107(.a(output_3_107), .b(output_3_4), .y(output_2_107));
wire output_4_107, output_4_4, output_3_107;
mixer gate_output_3_107(.a(output_4_107), .b(output_4_4), .y(output_3_107));
wire output_5_107, output_5_4, output_4_107;
mixer gate_output_4_107(.a(output_5_107), .b(output_5_4), .y(output_4_107));
wire output_6_107, output_6_4, output_5_107;
mixer gate_output_5_107(.a(output_6_107), .b(output_6_4), .y(output_5_107));
wire output_7_107, output_7_4, output_6_107;
mixer gate_output_6_107(.a(output_7_107), .b(output_7_4), .y(output_6_107));
wire output_8_107, output_8_4, output_7_107;
mixer gate_output_7_107(.a(output_8_107), .b(output_8_4), .y(output_7_107));
wire output_1_108, output_1_5, output_0_108;
mixer gate_output_0_108(.a(output_1_108), .b(output_1_5), .y(output_0_108));
wire output_2_108, output_2_5, output_1_108;
mixer gate_output_1_108(.a(output_2_108), .b(output_2_5), .y(output_1_108));
wire output_3_108, output_3_5, output_2_108;
mixer gate_output_2_108(.a(output_3_108), .b(output_3_5), .y(output_2_108));
wire output_4_108, output_4_5, output_3_108;
mixer gate_output_3_108(.a(output_4_108), .b(output_4_5), .y(output_3_108));
wire output_5_108, output_5_5, output_4_108;
mixer gate_output_4_108(.a(output_5_108), .b(output_5_5), .y(output_4_108));
wire output_6_108, output_6_5, output_5_108;
mixer gate_output_5_108(.a(output_6_108), .b(output_6_5), .y(output_5_108));
wire output_7_108, output_7_5, output_6_108;
mixer gate_output_6_108(.a(output_7_108), .b(output_7_5), .y(output_6_108));
wire output_8_108, output_8_5, output_7_108;
mixer gate_output_7_108(.a(output_8_108), .b(output_8_5), .y(output_7_108));
wire output_1_109, output_1_6, output_0_109;
mixer gate_output_0_109(.a(output_1_109), .b(output_1_6), .y(output_0_109));
wire output_2_109, output_2_6, output_1_109;
mixer gate_output_1_109(.a(output_2_109), .b(output_2_6), .y(output_1_109));
wire output_3_109, output_3_6, output_2_109;
mixer gate_output_2_109(.a(output_3_109), .b(output_3_6), .y(output_2_109));
wire output_4_109, output_4_6, output_3_109;
mixer gate_output_3_109(.a(output_4_109), .b(output_4_6), .y(output_3_109));
wire output_5_109, output_5_6, output_4_109;
mixer gate_output_4_109(.a(output_5_109), .b(output_5_6), .y(output_4_109));
wire output_6_109, output_6_6, output_5_109;
mixer gate_output_5_109(.a(output_6_109), .b(output_6_6), .y(output_5_109));
wire output_7_109, output_7_6, output_6_109;
mixer gate_output_6_109(.a(output_7_109), .b(output_7_6), .y(output_6_109));
wire output_8_109, output_8_6, output_7_109;
mixer gate_output_7_109(.a(output_8_109), .b(output_8_6), .y(output_7_109));
wire output_1_110, output_1_7, output_0_110;
mixer gate_output_0_110(.a(output_1_110), .b(output_1_7), .y(output_0_110));
wire output_2_110, output_2_7, output_1_110;
mixer gate_output_1_110(.a(output_2_110), .b(output_2_7), .y(output_1_110));
wire output_3_110, output_3_7, output_2_110;
mixer gate_output_2_110(.a(output_3_110), .b(output_3_7), .y(output_2_110));
wire output_4_110, output_4_7, output_3_110;
mixer gate_output_3_110(.a(output_4_110), .b(output_4_7), .y(output_3_110));
wire output_5_110, output_5_7, output_4_110;
mixer gate_output_4_110(.a(output_5_110), .b(output_5_7), .y(output_4_110));
wire output_6_110, output_6_7, output_5_110;
mixer gate_output_5_110(.a(output_6_110), .b(output_6_7), .y(output_5_110));
wire output_7_110, output_7_7, output_6_110;
mixer gate_output_6_110(.a(output_7_110), .b(output_7_7), .y(output_6_110));
wire output_8_110, output_8_7, output_7_110;
mixer gate_output_7_110(.a(output_8_110), .b(output_8_7), .y(output_7_110));
wire output_1_111, output_1_0, output_0_111;
mixer gate_output_0_111(.a(output_1_111), .b(output_1_0), .y(output_0_111));
wire output_2_111, output_2_0, output_1_111;
mixer gate_output_1_111(.a(output_2_111), .b(output_2_0), .y(output_1_111));
wire output_3_111, output_3_0, output_2_111;
mixer gate_output_2_111(.a(output_3_111), .b(output_3_0), .y(output_2_111));
wire output_4_111, output_4_0, output_3_111;
mixer gate_output_3_111(.a(output_4_111), .b(output_4_0), .y(output_3_111));
wire output_5_111, output_5_0, output_4_111;
mixer gate_output_4_111(.a(output_5_111), .b(output_5_0), .y(output_4_111));
wire output_6_111, output_6_0, output_5_111;
mixer gate_output_5_111(.a(output_6_111), .b(output_6_0), .y(output_5_111));
wire output_7_111, output_7_0, output_6_111;
mixer gate_output_6_111(.a(output_7_111), .b(output_7_0), .y(output_6_111));
wire output_8_111, output_8_0, output_7_111;
mixer gate_output_7_111(.a(output_8_111), .b(output_8_0), .y(output_7_111));
wire output_1_112, output_1_1, output_0_112;
mixer gate_output_0_112(.a(output_1_112), .b(output_1_1), .y(output_0_112));
wire output_2_112, output_2_1, output_1_112;
mixer gate_output_1_112(.a(output_2_112), .b(output_2_1), .y(output_1_112));
wire output_3_112, output_3_1, output_2_112;
mixer gate_output_2_112(.a(output_3_112), .b(output_3_1), .y(output_2_112));
wire output_4_112, output_4_1, output_3_112;
mixer gate_output_3_112(.a(output_4_112), .b(output_4_1), .y(output_3_112));
wire output_5_112, output_5_1, output_4_112;
mixer gate_output_4_112(.a(output_5_112), .b(output_5_1), .y(output_4_112));
wire output_6_112, output_6_1, output_5_112;
mixer gate_output_5_112(.a(output_6_112), .b(output_6_1), .y(output_5_112));
wire output_7_112, output_7_1, output_6_112;
mixer gate_output_6_112(.a(output_7_112), .b(output_7_1), .y(output_6_112));
wire output_8_112, output_8_1, output_7_112;
mixer gate_output_7_112(.a(output_8_112), .b(output_8_1), .y(output_7_112));
wire output_1_113, output_1_2, output_0_113;
mixer gate_output_0_113(.a(output_1_113), .b(output_1_2), .y(output_0_113));
wire output_2_113, output_2_2, output_1_113;
mixer gate_output_1_113(.a(output_2_113), .b(output_2_2), .y(output_1_113));
wire output_3_113, output_3_2, output_2_113;
mixer gate_output_2_113(.a(output_3_113), .b(output_3_2), .y(output_2_113));
wire output_4_113, output_4_2, output_3_113;
mixer gate_output_3_113(.a(output_4_113), .b(output_4_2), .y(output_3_113));
wire output_5_113, output_5_2, output_4_113;
mixer gate_output_4_113(.a(output_5_113), .b(output_5_2), .y(output_4_113));
wire output_6_113, output_6_2, output_5_113;
mixer gate_output_5_113(.a(output_6_113), .b(output_6_2), .y(output_5_113));
wire output_7_113, output_7_2, output_6_113;
mixer gate_output_6_113(.a(output_7_113), .b(output_7_2), .y(output_6_113));
wire output_8_113, output_8_2, output_7_113;
mixer gate_output_7_113(.a(output_8_113), .b(output_8_2), .y(output_7_113));
wire output_1_114, output_1_3, output_0_114;
mixer gate_output_0_114(.a(output_1_114), .b(output_1_3), .y(output_0_114));
wire output_2_114, output_2_3, output_1_114;
mixer gate_output_1_114(.a(output_2_114), .b(output_2_3), .y(output_1_114));
wire output_3_114, output_3_3, output_2_114;
mixer gate_output_2_114(.a(output_3_114), .b(output_3_3), .y(output_2_114));
wire output_4_114, output_4_3, output_3_114;
mixer gate_output_3_114(.a(output_4_114), .b(output_4_3), .y(output_3_114));
wire output_5_114, output_5_3, output_4_114;
mixer gate_output_4_114(.a(output_5_114), .b(output_5_3), .y(output_4_114));
wire output_6_114, output_6_3, output_5_114;
mixer gate_output_5_114(.a(output_6_114), .b(output_6_3), .y(output_5_114));
wire output_7_114, output_7_3, output_6_114;
mixer gate_output_6_114(.a(output_7_114), .b(output_7_3), .y(output_6_114));
wire output_8_114, output_8_3, output_7_114;
mixer gate_output_7_114(.a(output_8_114), .b(output_8_3), .y(output_7_114));
wire output_1_115, output_1_4, output_0_115;
mixer gate_output_0_115(.a(output_1_115), .b(output_1_4), .y(output_0_115));
wire output_2_115, output_2_4, output_1_115;
mixer gate_output_1_115(.a(output_2_115), .b(output_2_4), .y(output_1_115));
wire output_3_115, output_3_4, output_2_115;
mixer gate_output_2_115(.a(output_3_115), .b(output_3_4), .y(output_2_115));
wire output_4_115, output_4_4, output_3_115;
mixer gate_output_3_115(.a(output_4_115), .b(output_4_4), .y(output_3_115));
wire output_5_115, output_5_4, output_4_115;
mixer gate_output_4_115(.a(output_5_115), .b(output_5_4), .y(output_4_115));
wire output_6_115, output_6_4, output_5_115;
mixer gate_output_5_115(.a(output_6_115), .b(output_6_4), .y(output_5_115));
wire output_7_115, output_7_4, output_6_115;
mixer gate_output_6_115(.a(output_7_115), .b(output_7_4), .y(output_6_115));
wire output_8_115, output_8_4, output_7_115;
mixer gate_output_7_115(.a(output_8_115), .b(output_8_4), .y(output_7_115));
wire output_1_116, output_1_5, output_0_116;
mixer gate_output_0_116(.a(output_1_116), .b(output_1_5), .y(output_0_116));
wire output_2_116, output_2_5, output_1_116;
mixer gate_output_1_116(.a(output_2_116), .b(output_2_5), .y(output_1_116));
wire output_3_116, output_3_5, output_2_116;
mixer gate_output_2_116(.a(output_3_116), .b(output_3_5), .y(output_2_116));
wire output_4_116, output_4_5, output_3_116;
mixer gate_output_3_116(.a(output_4_116), .b(output_4_5), .y(output_3_116));
wire output_5_116, output_5_5, output_4_116;
mixer gate_output_4_116(.a(output_5_116), .b(output_5_5), .y(output_4_116));
wire output_6_116, output_6_5, output_5_116;
mixer gate_output_5_116(.a(output_6_116), .b(output_6_5), .y(output_5_116));
wire output_7_116, output_7_5, output_6_116;
mixer gate_output_6_116(.a(output_7_116), .b(output_7_5), .y(output_6_116));
wire output_8_116, output_8_5, output_7_116;
mixer gate_output_7_116(.a(output_8_116), .b(output_8_5), .y(output_7_116));
wire output_1_117, output_1_6, output_0_117;
mixer gate_output_0_117(.a(output_1_117), .b(output_1_6), .y(output_0_117));
wire output_2_117, output_2_6, output_1_117;
mixer gate_output_1_117(.a(output_2_117), .b(output_2_6), .y(output_1_117));
wire output_3_117, output_3_6, output_2_117;
mixer gate_output_2_117(.a(output_3_117), .b(output_3_6), .y(output_2_117));
wire output_4_117, output_4_6, output_3_117;
mixer gate_output_3_117(.a(output_4_117), .b(output_4_6), .y(output_3_117));
wire output_5_117, output_5_6, output_4_117;
mixer gate_output_4_117(.a(output_5_117), .b(output_5_6), .y(output_4_117));
wire output_6_117, output_6_6, output_5_117;
mixer gate_output_5_117(.a(output_6_117), .b(output_6_6), .y(output_5_117));
wire output_7_117, output_7_6, output_6_117;
mixer gate_output_6_117(.a(output_7_117), .b(output_7_6), .y(output_6_117));
wire output_8_117, output_8_6, output_7_117;
mixer gate_output_7_117(.a(output_8_117), .b(output_8_6), .y(output_7_117));
wire output_1_118, output_1_7, output_0_118;
mixer gate_output_0_118(.a(output_1_118), .b(output_1_7), .y(output_0_118));
wire output_2_118, output_2_7, output_1_118;
mixer gate_output_1_118(.a(output_2_118), .b(output_2_7), .y(output_1_118));
wire output_3_118, output_3_7, output_2_118;
mixer gate_output_2_118(.a(output_3_118), .b(output_3_7), .y(output_2_118));
wire output_4_118, output_4_7, output_3_118;
mixer gate_output_3_118(.a(output_4_118), .b(output_4_7), .y(output_3_118));
wire output_5_118, output_5_7, output_4_118;
mixer gate_output_4_118(.a(output_5_118), .b(output_5_7), .y(output_4_118));
wire output_6_118, output_6_7, output_5_118;
mixer gate_output_5_118(.a(output_6_118), .b(output_6_7), .y(output_5_118));
wire output_7_118, output_7_7, output_6_118;
mixer gate_output_6_118(.a(output_7_118), .b(output_7_7), .y(output_6_118));
wire output_8_118, output_8_7, output_7_118;
mixer gate_output_7_118(.a(output_8_118), .b(output_8_7), .y(output_7_118));
wire output_1_119, output_1_0, output_0_119;
mixer gate_output_0_119(.a(output_1_119), .b(output_1_0), .y(output_0_119));
wire output_2_119, output_2_0, output_1_119;
mixer gate_output_1_119(.a(output_2_119), .b(output_2_0), .y(output_1_119));
wire output_3_119, output_3_0, output_2_119;
mixer gate_output_2_119(.a(output_3_119), .b(output_3_0), .y(output_2_119));
wire output_4_119, output_4_0, output_3_119;
mixer gate_output_3_119(.a(output_4_119), .b(output_4_0), .y(output_3_119));
wire output_5_119, output_5_0, output_4_119;
mixer gate_output_4_119(.a(output_5_119), .b(output_5_0), .y(output_4_119));
wire output_6_119, output_6_0, output_5_119;
mixer gate_output_5_119(.a(output_6_119), .b(output_6_0), .y(output_5_119));
wire output_7_119, output_7_0, output_6_119;
mixer gate_output_6_119(.a(output_7_119), .b(output_7_0), .y(output_6_119));
wire output_8_119, output_8_0, output_7_119;
mixer gate_output_7_119(.a(output_8_119), .b(output_8_0), .y(output_7_119));
wire output_1_120, output_1_1, output_0_120;
mixer gate_output_0_120(.a(output_1_120), .b(output_1_1), .y(output_0_120));
wire output_2_120, output_2_1, output_1_120;
mixer gate_output_1_120(.a(output_2_120), .b(output_2_1), .y(output_1_120));
wire output_3_120, output_3_1, output_2_120;
mixer gate_output_2_120(.a(output_3_120), .b(output_3_1), .y(output_2_120));
wire output_4_120, output_4_1, output_3_120;
mixer gate_output_3_120(.a(output_4_120), .b(output_4_1), .y(output_3_120));
wire output_5_120, output_5_1, output_4_120;
mixer gate_output_4_120(.a(output_5_120), .b(output_5_1), .y(output_4_120));
wire output_6_120, output_6_1, output_5_120;
mixer gate_output_5_120(.a(output_6_120), .b(output_6_1), .y(output_5_120));
wire output_7_120, output_7_1, output_6_120;
mixer gate_output_6_120(.a(output_7_120), .b(output_7_1), .y(output_6_120));
wire output_8_120, output_8_1, output_7_120;
mixer gate_output_7_120(.a(output_8_120), .b(output_8_1), .y(output_7_120));
wire output_1_121, output_1_2, output_0_121;
mixer gate_output_0_121(.a(output_1_121), .b(output_1_2), .y(output_0_121));
wire output_2_121, output_2_2, output_1_121;
mixer gate_output_1_121(.a(output_2_121), .b(output_2_2), .y(output_1_121));
wire output_3_121, output_3_2, output_2_121;
mixer gate_output_2_121(.a(output_3_121), .b(output_3_2), .y(output_2_121));
wire output_4_121, output_4_2, output_3_121;
mixer gate_output_3_121(.a(output_4_121), .b(output_4_2), .y(output_3_121));
wire output_5_121, output_5_2, output_4_121;
mixer gate_output_4_121(.a(output_5_121), .b(output_5_2), .y(output_4_121));
wire output_6_121, output_6_2, output_5_121;
mixer gate_output_5_121(.a(output_6_121), .b(output_6_2), .y(output_5_121));
wire output_7_121, output_7_2, output_6_121;
mixer gate_output_6_121(.a(output_7_121), .b(output_7_2), .y(output_6_121));
wire output_8_121, output_8_2, output_7_121;
mixer gate_output_7_121(.a(output_8_121), .b(output_8_2), .y(output_7_121));
wire output_1_122, output_1_3, output_0_122;
mixer gate_output_0_122(.a(output_1_122), .b(output_1_3), .y(output_0_122));
wire output_2_122, output_2_3, output_1_122;
mixer gate_output_1_122(.a(output_2_122), .b(output_2_3), .y(output_1_122));
wire output_3_122, output_3_3, output_2_122;
mixer gate_output_2_122(.a(output_3_122), .b(output_3_3), .y(output_2_122));
wire output_4_122, output_4_3, output_3_122;
mixer gate_output_3_122(.a(output_4_122), .b(output_4_3), .y(output_3_122));
wire output_5_122, output_5_3, output_4_122;
mixer gate_output_4_122(.a(output_5_122), .b(output_5_3), .y(output_4_122));
wire output_6_122, output_6_3, output_5_122;
mixer gate_output_5_122(.a(output_6_122), .b(output_6_3), .y(output_5_122));
wire output_7_122, output_7_3, output_6_122;
mixer gate_output_6_122(.a(output_7_122), .b(output_7_3), .y(output_6_122));
wire output_8_122, output_8_3, output_7_122;
mixer gate_output_7_122(.a(output_8_122), .b(output_8_3), .y(output_7_122));
wire output_1_123, output_1_4, output_0_123;
mixer gate_output_0_123(.a(output_1_123), .b(output_1_4), .y(output_0_123));
wire output_2_123, output_2_4, output_1_123;
mixer gate_output_1_123(.a(output_2_123), .b(output_2_4), .y(output_1_123));
wire output_3_123, output_3_4, output_2_123;
mixer gate_output_2_123(.a(output_3_123), .b(output_3_4), .y(output_2_123));
wire output_4_123, output_4_4, output_3_123;
mixer gate_output_3_123(.a(output_4_123), .b(output_4_4), .y(output_3_123));
wire output_5_123, output_5_4, output_4_123;
mixer gate_output_4_123(.a(output_5_123), .b(output_5_4), .y(output_4_123));
wire output_6_123, output_6_4, output_5_123;
mixer gate_output_5_123(.a(output_6_123), .b(output_6_4), .y(output_5_123));
wire output_7_123, output_7_4, output_6_123;
mixer gate_output_6_123(.a(output_7_123), .b(output_7_4), .y(output_6_123));
wire output_8_123, output_8_4, output_7_123;
mixer gate_output_7_123(.a(output_8_123), .b(output_8_4), .y(output_7_123));
wire output_1_124, output_1_5, output_0_124;
mixer gate_output_0_124(.a(output_1_124), .b(output_1_5), .y(output_0_124));
wire output_2_124, output_2_5, output_1_124;
mixer gate_output_1_124(.a(output_2_124), .b(output_2_5), .y(output_1_124));
wire output_3_124, output_3_5, output_2_124;
mixer gate_output_2_124(.a(output_3_124), .b(output_3_5), .y(output_2_124));
wire output_4_124, output_4_5, output_3_124;
mixer gate_output_3_124(.a(output_4_124), .b(output_4_5), .y(output_3_124));
wire output_5_124, output_5_5, output_4_124;
mixer gate_output_4_124(.a(output_5_124), .b(output_5_5), .y(output_4_124));
wire output_6_124, output_6_5, output_5_124;
mixer gate_output_5_124(.a(output_6_124), .b(output_6_5), .y(output_5_124));
wire output_7_124, output_7_5, output_6_124;
mixer gate_output_6_124(.a(output_7_124), .b(output_7_5), .y(output_6_124));
wire output_8_124, output_8_5, output_7_124;
mixer gate_output_7_124(.a(output_8_124), .b(output_8_5), .y(output_7_124));
wire output_1_125, output_1_6, output_0_125;
mixer gate_output_0_125(.a(output_1_125), .b(output_1_6), .y(output_0_125));
wire output_2_125, output_2_6, output_1_125;
mixer gate_output_1_125(.a(output_2_125), .b(output_2_6), .y(output_1_125));
wire output_3_125, output_3_6, output_2_125;
mixer gate_output_2_125(.a(output_3_125), .b(output_3_6), .y(output_2_125));
wire output_4_125, output_4_6, output_3_125;
mixer gate_output_3_125(.a(output_4_125), .b(output_4_6), .y(output_3_125));
wire output_5_125, output_5_6, output_4_125;
mixer gate_output_4_125(.a(output_5_125), .b(output_5_6), .y(output_4_125));
wire output_6_125, output_6_6, output_5_125;
mixer gate_output_5_125(.a(output_6_125), .b(output_6_6), .y(output_5_125));
wire output_7_125, output_7_6, output_6_125;
mixer gate_output_6_125(.a(output_7_125), .b(output_7_6), .y(output_6_125));
wire output_8_125, output_8_6, output_7_125;
mixer gate_output_7_125(.a(output_8_125), .b(output_8_6), .y(output_7_125));
wire output_1_126, output_1_7, output_0_126;
mixer gate_output_0_126(.a(output_1_126), .b(output_1_7), .y(output_0_126));
wire output_2_126, output_2_7, output_1_126;
mixer gate_output_1_126(.a(output_2_126), .b(output_2_7), .y(output_1_126));
wire output_3_126, output_3_7, output_2_126;
mixer gate_output_2_126(.a(output_3_126), .b(output_3_7), .y(output_2_126));
wire output_4_126, output_4_7, output_3_126;
mixer gate_output_3_126(.a(output_4_126), .b(output_4_7), .y(output_3_126));
wire output_5_126, output_5_7, output_4_126;
mixer gate_output_4_126(.a(output_5_126), .b(output_5_7), .y(output_4_126));
wire output_6_126, output_6_7, output_5_126;
mixer gate_output_5_126(.a(output_6_126), .b(output_6_7), .y(output_5_126));
wire output_7_126, output_7_7, output_6_126;
mixer gate_output_6_126(.a(output_7_126), .b(output_7_7), .y(output_6_126));
wire output_8_126, output_8_7, output_7_126;
mixer gate_output_7_126(.a(output_8_126), .b(output_8_7), .y(output_7_126));
wire output_1_127, output_1_0, output_0_127;
mixer gate_output_0_127(.a(output_1_127), .b(output_1_0), .y(output_0_127));
wire output_2_127, output_2_0, output_1_127;
mixer gate_output_1_127(.a(output_2_127), .b(output_2_0), .y(output_1_127));
wire output_3_127, output_3_0, output_2_127;
mixer gate_output_2_127(.a(output_3_127), .b(output_3_0), .y(output_2_127));
wire output_4_127, output_4_0, output_3_127;
mixer gate_output_3_127(.a(output_4_127), .b(output_4_0), .y(output_3_127));
wire output_5_127, output_5_0, output_4_127;
mixer gate_output_4_127(.a(output_5_127), .b(output_5_0), .y(output_4_127));
wire output_6_127, output_6_0, output_5_127;
mixer gate_output_5_127(.a(output_6_127), .b(output_6_0), .y(output_5_127));
wire output_7_127, output_7_0, output_6_127;
mixer gate_output_6_127(.a(output_7_127), .b(output_7_0), .y(output_6_127));
wire output_8_127, output_8_0, output_7_127;
mixer gate_output_7_127(.a(output_8_127), .b(output_8_0), .y(output_7_127));
wire output_1_128, output_1_1, output_0_128;
mixer gate_output_0_128(.a(output_1_128), .b(output_1_1), .y(output_0_128));
wire output_2_128, output_2_1, output_1_128;
mixer gate_output_1_128(.a(output_2_128), .b(output_2_1), .y(output_1_128));
wire output_3_128, output_3_1, output_2_128;
mixer gate_output_2_128(.a(output_3_128), .b(output_3_1), .y(output_2_128));
wire output_4_128, output_4_1, output_3_128;
mixer gate_output_3_128(.a(output_4_128), .b(output_4_1), .y(output_3_128));
wire output_5_128, output_5_1, output_4_128;
mixer gate_output_4_128(.a(output_5_128), .b(output_5_1), .y(output_4_128));
wire output_6_128, output_6_1, output_5_128;
mixer gate_output_5_128(.a(output_6_128), .b(output_6_1), .y(output_5_128));
wire output_7_128, output_7_1, output_6_128;
mixer gate_output_6_128(.a(output_7_128), .b(output_7_1), .y(output_6_128));
wire output_8_128, output_8_1, output_7_128;
mixer gate_output_7_128(.a(output_8_128), .b(output_8_1), .y(output_7_128));
wire output_1_129, output_1_2, output_0_129;
mixer gate_output_0_129(.a(output_1_129), .b(output_1_2), .y(output_0_129));
wire output_2_129, output_2_2, output_1_129;
mixer gate_output_1_129(.a(output_2_129), .b(output_2_2), .y(output_1_129));
wire output_3_129, output_3_2, output_2_129;
mixer gate_output_2_129(.a(output_3_129), .b(output_3_2), .y(output_2_129));
wire output_4_129, output_4_2, output_3_129;
mixer gate_output_3_129(.a(output_4_129), .b(output_4_2), .y(output_3_129));
wire output_5_129, output_5_2, output_4_129;
mixer gate_output_4_129(.a(output_5_129), .b(output_5_2), .y(output_4_129));
wire output_6_129, output_6_2, output_5_129;
mixer gate_output_5_129(.a(output_6_129), .b(output_6_2), .y(output_5_129));
wire output_7_129, output_7_2, output_6_129;
mixer gate_output_6_129(.a(output_7_129), .b(output_7_2), .y(output_6_129));
wire output_8_129, output_8_2, output_7_129;
mixer gate_output_7_129(.a(output_8_129), .b(output_8_2), .y(output_7_129));
wire output_1_130, output_1_3, output_0_130;
mixer gate_output_0_130(.a(output_1_130), .b(output_1_3), .y(output_0_130));
wire output_2_130, output_2_3, output_1_130;
mixer gate_output_1_130(.a(output_2_130), .b(output_2_3), .y(output_1_130));
wire output_3_130, output_3_3, output_2_130;
mixer gate_output_2_130(.a(output_3_130), .b(output_3_3), .y(output_2_130));
wire output_4_130, output_4_3, output_3_130;
mixer gate_output_3_130(.a(output_4_130), .b(output_4_3), .y(output_3_130));
wire output_5_130, output_5_3, output_4_130;
mixer gate_output_4_130(.a(output_5_130), .b(output_5_3), .y(output_4_130));
wire output_6_130, output_6_3, output_5_130;
mixer gate_output_5_130(.a(output_6_130), .b(output_6_3), .y(output_5_130));
wire output_7_130, output_7_3, output_6_130;
mixer gate_output_6_130(.a(output_7_130), .b(output_7_3), .y(output_6_130));
wire output_8_130, output_8_3, output_7_130;
mixer gate_output_7_130(.a(output_8_130), .b(output_8_3), .y(output_7_130));
wire output_1_131, output_1_4, output_0_131;
mixer gate_output_0_131(.a(output_1_131), .b(output_1_4), .y(output_0_131));
wire output_2_131, output_2_4, output_1_131;
mixer gate_output_1_131(.a(output_2_131), .b(output_2_4), .y(output_1_131));
wire output_3_131, output_3_4, output_2_131;
mixer gate_output_2_131(.a(output_3_131), .b(output_3_4), .y(output_2_131));
wire output_4_131, output_4_4, output_3_131;
mixer gate_output_3_131(.a(output_4_131), .b(output_4_4), .y(output_3_131));
wire output_5_131, output_5_4, output_4_131;
mixer gate_output_4_131(.a(output_5_131), .b(output_5_4), .y(output_4_131));
wire output_6_131, output_6_4, output_5_131;
mixer gate_output_5_131(.a(output_6_131), .b(output_6_4), .y(output_5_131));
wire output_7_131, output_7_4, output_6_131;
mixer gate_output_6_131(.a(output_7_131), .b(output_7_4), .y(output_6_131));
wire output_8_131, output_8_4, output_7_131;
mixer gate_output_7_131(.a(output_8_131), .b(output_8_4), .y(output_7_131));
wire output_1_132, output_1_5, output_0_132;
mixer gate_output_0_132(.a(output_1_132), .b(output_1_5), .y(output_0_132));
wire output_2_132, output_2_5, output_1_132;
mixer gate_output_1_132(.a(output_2_132), .b(output_2_5), .y(output_1_132));
wire output_3_132, output_3_5, output_2_132;
mixer gate_output_2_132(.a(output_3_132), .b(output_3_5), .y(output_2_132));
wire output_4_132, output_4_5, output_3_132;
mixer gate_output_3_132(.a(output_4_132), .b(output_4_5), .y(output_3_132));
wire output_5_132, output_5_5, output_4_132;
mixer gate_output_4_132(.a(output_5_132), .b(output_5_5), .y(output_4_132));
wire output_6_132, output_6_5, output_5_132;
mixer gate_output_5_132(.a(output_6_132), .b(output_6_5), .y(output_5_132));
wire output_7_132, output_7_5, output_6_132;
mixer gate_output_6_132(.a(output_7_132), .b(output_7_5), .y(output_6_132));
wire output_8_132, output_8_5, output_7_132;
mixer gate_output_7_132(.a(output_8_132), .b(output_8_5), .y(output_7_132));
wire output_1_133, output_1_6, output_0_133;
mixer gate_output_0_133(.a(output_1_133), .b(output_1_6), .y(output_0_133));
wire output_2_133, output_2_6, output_1_133;
mixer gate_output_1_133(.a(output_2_133), .b(output_2_6), .y(output_1_133));
wire output_3_133, output_3_6, output_2_133;
mixer gate_output_2_133(.a(output_3_133), .b(output_3_6), .y(output_2_133));
wire output_4_133, output_4_6, output_3_133;
mixer gate_output_3_133(.a(output_4_133), .b(output_4_6), .y(output_3_133));
wire output_5_133, output_5_6, output_4_133;
mixer gate_output_4_133(.a(output_5_133), .b(output_5_6), .y(output_4_133));
wire output_6_133, output_6_6, output_5_133;
mixer gate_output_5_133(.a(output_6_133), .b(output_6_6), .y(output_5_133));
wire output_7_133, output_7_6, output_6_133;
mixer gate_output_6_133(.a(output_7_133), .b(output_7_6), .y(output_6_133));
wire output_8_133, output_8_6, output_7_133;
mixer gate_output_7_133(.a(output_8_133), .b(output_8_6), .y(output_7_133));
wire output_1_134, output_1_7, output_0_134;
mixer gate_output_0_134(.a(output_1_134), .b(output_1_7), .y(output_0_134));
wire output_2_134, output_2_7, output_1_134;
mixer gate_output_1_134(.a(output_2_134), .b(output_2_7), .y(output_1_134));
wire output_3_134, output_3_7, output_2_134;
mixer gate_output_2_134(.a(output_3_134), .b(output_3_7), .y(output_2_134));
wire output_4_134, output_4_7, output_3_134;
mixer gate_output_3_134(.a(output_4_134), .b(output_4_7), .y(output_3_134));
wire output_5_134, output_5_7, output_4_134;
mixer gate_output_4_134(.a(output_5_134), .b(output_5_7), .y(output_4_134));
wire output_6_134, output_6_7, output_5_134;
mixer gate_output_5_134(.a(output_6_134), .b(output_6_7), .y(output_5_134));
wire output_7_134, output_7_7, output_6_134;
mixer gate_output_6_134(.a(output_7_134), .b(output_7_7), .y(output_6_134));
wire output_8_134, output_8_7, output_7_134;
mixer gate_output_7_134(.a(output_8_134), .b(output_8_7), .y(output_7_134));
wire output_1_135, output_1_0, output_0_135;
mixer gate_output_0_135(.a(output_1_135), .b(output_1_0), .y(output_0_135));
wire output_2_135, output_2_0, output_1_135;
mixer gate_output_1_135(.a(output_2_135), .b(output_2_0), .y(output_1_135));
wire output_3_135, output_3_0, output_2_135;
mixer gate_output_2_135(.a(output_3_135), .b(output_3_0), .y(output_2_135));
wire output_4_135, output_4_0, output_3_135;
mixer gate_output_3_135(.a(output_4_135), .b(output_4_0), .y(output_3_135));
wire output_5_135, output_5_0, output_4_135;
mixer gate_output_4_135(.a(output_5_135), .b(output_5_0), .y(output_4_135));
wire output_6_135, output_6_0, output_5_135;
mixer gate_output_5_135(.a(output_6_135), .b(output_6_0), .y(output_5_135));
wire output_7_135, output_7_0, output_6_135;
mixer gate_output_6_135(.a(output_7_135), .b(output_7_0), .y(output_6_135));
wire output_8_135, output_8_0, output_7_135;
mixer gate_output_7_135(.a(output_8_135), .b(output_8_0), .y(output_7_135));
wire output_1_136, output_1_1, output_0_136;
mixer gate_output_0_136(.a(output_1_136), .b(output_1_1), .y(output_0_136));
wire output_2_136, output_2_1, output_1_136;
mixer gate_output_1_136(.a(output_2_136), .b(output_2_1), .y(output_1_136));
wire output_3_136, output_3_1, output_2_136;
mixer gate_output_2_136(.a(output_3_136), .b(output_3_1), .y(output_2_136));
wire output_4_136, output_4_1, output_3_136;
mixer gate_output_3_136(.a(output_4_136), .b(output_4_1), .y(output_3_136));
wire output_5_136, output_5_1, output_4_136;
mixer gate_output_4_136(.a(output_5_136), .b(output_5_1), .y(output_4_136));
wire output_6_136, output_6_1, output_5_136;
mixer gate_output_5_136(.a(output_6_136), .b(output_6_1), .y(output_5_136));
wire output_7_136, output_7_1, output_6_136;
mixer gate_output_6_136(.a(output_7_136), .b(output_7_1), .y(output_6_136));
wire output_8_136, output_8_1, output_7_136;
mixer gate_output_7_136(.a(output_8_136), .b(output_8_1), .y(output_7_136));
wire output_1_137, output_1_2, output_0_137;
mixer gate_output_0_137(.a(output_1_137), .b(output_1_2), .y(output_0_137));
wire output_2_137, output_2_2, output_1_137;
mixer gate_output_1_137(.a(output_2_137), .b(output_2_2), .y(output_1_137));
wire output_3_137, output_3_2, output_2_137;
mixer gate_output_2_137(.a(output_3_137), .b(output_3_2), .y(output_2_137));
wire output_4_137, output_4_2, output_3_137;
mixer gate_output_3_137(.a(output_4_137), .b(output_4_2), .y(output_3_137));
wire output_5_137, output_5_2, output_4_137;
mixer gate_output_4_137(.a(output_5_137), .b(output_5_2), .y(output_4_137));
wire output_6_137, output_6_2, output_5_137;
mixer gate_output_5_137(.a(output_6_137), .b(output_6_2), .y(output_5_137));
wire output_7_137, output_7_2, output_6_137;
mixer gate_output_6_137(.a(output_7_137), .b(output_7_2), .y(output_6_137));
wire output_8_137, output_8_2, output_7_137;
mixer gate_output_7_137(.a(output_8_137), .b(output_8_2), .y(output_7_137));
wire output_1_138, output_1_3, output_0_138;
mixer gate_output_0_138(.a(output_1_138), .b(output_1_3), .y(output_0_138));
wire output_2_138, output_2_3, output_1_138;
mixer gate_output_1_138(.a(output_2_138), .b(output_2_3), .y(output_1_138));
wire output_3_138, output_3_3, output_2_138;
mixer gate_output_2_138(.a(output_3_138), .b(output_3_3), .y(output_2_138));
wire output_4_138, output_4_3, output_3_138;
mixer gate_output_3_138(.a(output_4_138), .b(output_4_3), .y(output_3_138));
wire output_5_138, output_5_3, output_4_138;
mixer gate_output_4_138(.a(output_5_138), .b(output_5_3), .y(output_4_138));
wire output_6_138, output_6_3, output_5_138;
mixer gate_output_5_138(.a(output_6_138), .b(output_6_3), .y(output_5_138));
wire output_7_138, output_7_3, output_6_138;
mixer gate_output_6_138(.a(output_7_138), .b(output_7_3), .y(output_6_138));
wire output_8_138, output_8_3, output_7_138;
mixer gate_output_7_138(.a(output_8_138), .b(output_8_3), .y(output_7_138));
wire output_1_139, output_1_4, output_0_139;
mixer gate_output_0_139(.a(output_1_139), .b(output_1_4), .y(output_0_139));
wire output_2_139, output_2_4, output_1_139;
mixer gate_output_1_139(.a(output_2_139), .b(output_2_4), .y(output_1_139));
wire output_3_139, output_3_4, output_2_139;
mixer gate_output_2_139(.a(output_3_139), .b(output_3_4), .y(output_2_139));
wire output_4_139, output_4_4, output_3_139;
mixer gate_output_3_139(.a(output_4_139), .b(output_4_4), .y(output_3_139));
wire output_5_139, output_5_4, output_4_139;
mixer gate_output_4_139(.a(output_5_139), .b(output_5_4), .y(output_4_139));
wire output_6_139, output_6_4, output_5_139;
mixer gate_output_5_139(.a(output_6_139), .b(output_6_4), .y(output_5_139));
wire output_7_139, output_7_4, output_6_139;
mixer gate_output_6_139(.a(output_7_139), .b(output_7_4), .y(output_6_139));
wire output_8_139, output_8_4, output_7_139;
mixer gate_output_7_139(.a(output_8_139), .b(output_8_4), .y(output_7_139));
wire output_1_140, output_1_5, output_0_140;
mixer gate_output_0_140(.a(output_1_140), .b(output_1_5), .y(output_0_140));
wire output_2_140, output_2_5, output_1_140;
mixer gate_output_1_140(.a(output_2_140), .b(output_2_5), .y(output_1_140));
wire output_3_140, output_3_5, output_2_140;
mixer gate_output_2_140(.a(output_3_140), .b(output_3_5), .y(output_2_140));
wire output_4_140, output_4_5, output_3_140;
mixer gate_output_3_140(.a(output_4_140), .b(output_4_5), .y(output_3_140));
wire output_5_140, output_5_5, output_4_140;
mixer gate_output_4_140(.a(output_5_140), .b(output_5_5), .y(output_4_140));
wire output_6_140, output_6_5, output_5_140;
mixer gate_output_5_140(.a(output_6_140), .b(output_6_5), .y(output_5_140));
wire output_7_140, output_7_5, output_6_140;
mixer gate_output_6_140(.a(output_7_140), .b(output_7_5), .y(output_6_140));
wire output_8_140, output_8_5, output_7_140;
mixer gate_output_7_140(.a(output_8_140), .b(output_8_5), .y(output_7_140));
wire output_1_141, output_1_6, output_0_141;
mixer gate_output_0_141(.a(output_1_141), .b(output_1_6), .y(output_0_141));
wire output_2_141, output_2_6, output_1_141;
mixer gate_output_1_141(.a(output_2_141), .b(output_2_6), .y(output_1_141));
wire output_3_141, output_3_6, output_2_141;
mixer gate_output_2_141(.a(output_3_141), .b(output_3_6), .y(output_2_141));
wire output_4_141, output_4_6, output_3_141;
mixer gate_output_3_141(.a(output_4_141), .b(output_4_6), .y(output_3_141));
wire output_5_141, output_5_6, output_4_141;
mixer gate_output_4_141(.a(output_5_141), .b(output_5_6), .y(output_4_141));
wire output_6_141, output_6_6, output_5_141;
mixer gate_output_5_141(.a(output_6_141), .b(output_6_6), .y(output_5_141));
wire output_7_141, output_7_6, output_6_141;
mixer gate_output_6_141(.a(output_7_141), .b(output_7_6), .y(output_6_141));
wire output_8_141, output_8_6, output_7_141;
mixer gate_output_7_141(.a(output_8_141), .b(output_8_6), .y(output_7_141));
wire output_1_142, output_1_7, output_0_142;
mixer gate_output_0_142(.a(output_1_142), .b(output_1_7), .y(output_0_142));
wire output_2_142, output_2_7, output_1_142;
mixer gate_output_1_142(.a(output_2_142), .b(output_2_7), .y(output_1_142));
wire output_3_142, output_3_7, output_2_142;
mixer gate_output_2_142(.a(output_3_142), .b(output_3_7), .y(output_2_142));
wire output_4_142, output_4_7, output_3_142;
mixer gate_output_3_142(.a(output_4_142), .b(output_4_7), .y(output_3_142));
wire output_5_142, output_5_7, output_4_142;
mixer gate_output_4_142(.a(output_5_142), .b(output_5_7), .y(output_4_142));
wire output_6_142, output_6_7, output_5_142;
mixer gate_output_5_142(.a(output_6_142), .b(output_6_7), .y(output_5_142));
wire output_7_142, output_7_7, output_6_142;
mixer gate_output_6_142(.a(output_7_142), .b(output_7_7), .y(output_6_142));
wire output_8_142, output_8_7, output_7_142;
mixer gate_output_7_142(.a(output_8_142), .b(output_8_7), .y(output_7_142));
wire output_1_143, output_1_0, output_0_143;
mixer gate_output_0_143(.a(output_1_143), .b(output_1_0), .y(output_0_143));
wire output_2_143, output_2_0, output_1_143;
mixer gate_output_1_143(.a(output_2_143), .b(output_2_0), .y(output_1_143));
wire output_3_143, output_3_0, output_2_143;
mixer gate_output_2_143(.a(output_3_143), .b(output_3_0), .y(output_2_143));
wire output_4_143, output_4_0, output_3_143;
mixer gate_output_3_143(.a(output_4_143), .b(output_4_0), .y(output_3_143));
wire output_5_143, output_5_0, output_4_143;
mixer gate_output_4_143(.a(output_5_143), .b(output_5_0), .y(output_4_143));
wire output_6_143, output_6_0, output_5_143;
mixer gate_output_5_143(.a(output_6_143), .b(output_6_0), .y(output_5_143));
wire output_7_143, output_7_0, output_6_143;
mixer gate_output_6_143(.a(output_7_143), .b(output_7_0), .y(output_6_143));
wire output_8_143, output_8_0, output_7_143;
mixer gate_output_7_143(.a(output_8_143), .b(output_8_0), .y(output_7_143));
wire output_1_144, output_1_1, output_0_144;
mixer gate_output_0_144(.a(output_1_144), .b(output_1_1), .y(output_0_144));
wire output_2_144, output_2_1, output_1_144;
mixer gate_output_1_144(.a(output_2_144), .b(output_2_1), .y(output_1_144));
wire output_3_144, output_3_1, output_2_144;
mixer gate_output_2_144(.a(output_3_144), .b(output_3_1), .y(output_2_144));
wire output_4_144, output_4_1, output_3_144;
mixer gate_output_3_144(.a(output_4_144), .b(output_4_1), .y(output_3_144));
wire output_5_144, output_5_1, output_4_144;
mixer gate_output_4_144(.a(output_5_144), .b(output_5_1), .y(output_4_144));
wire output_6_144, output_6_1, output_5_144;
mixer gate_output_5_144(.a(output_6_144), .b(output_6_1), .y(output_5_144));
wire output_7_144, output_7_1, output_6_144;
mixer gate_output_6_144(.a(output_7_144), .b(output_7_1), .y(output_6_144));
wire output_8_144, output_8_1, output_7_144;
mixer gate_output_7_144(.a(output_8_144), .b(output_8_1), .y(output_7_144));
wire output_1_145, output_1_2, output_0_145;
mixer gate_output_0_145(.a(output_1_145), .b(output_1_2), .y(output_0_145));
wire output_2_145, output_2_2, output_1_145;
mixer gate_output_1_145(.a(output_2_145), .b(output_2_2), .y(output_1_145));
wire output_3_145, output_3_2, output_2_145;
mixer gate_output_2_145(.a(output_3_145), .b(output_3_2), .y(output_2_145));
wire output_4_145, output_4_2, output_3_145;
mixer gate_output_3_145(.a(output_4_145), .b(output_4_2), .y(output_3_145));
wire output_5_145, output_5_2, output_4_145;
mixer gate_output_4_145(.a(output_5_145), .b(output_5_2), .y(output_4_145));
wire output_6_145, output_6_2, output_5_145;
mixer gate_output_5_145(.a(output_6_145), .b(output_6_2), .y(output_5_145));
wire output_7_145, output_7_2, output_6_145;
mixer gate_output_6_145(.a(output_7_145), .b(output_7_2), .y(output_6_145));
wire output_8_145, output_8_2, output_7_145;
mixer gate_output_7_145(.a(output_8_145), .b(output_8_2), .y(output_7_145));
wire output_1_146, output_1_3, output_0_146;
mixer gate_output_0_146(.a(output_1_146), .b(output_1_3), .y(output_0_146));
wire output_2_146, output_2_3, output_1_146;
mixer gate_output_1_146(.a(output_2_146), .b(output_2_3), .y(output_1_146));
wire output_3_146, output_3_3, output_2_146;
mixer gate_output_2_146(.a(output_3_146), .b(output_3_3), .y(output_2_146));
wire output_4_146, output_4_3, output_3_146;
mixer gate_output_3_146(.a(output_4_146), .b(output_4_3), .y(output_3_146));
wire output_5_146, output_5_3, output_4_146;
mixer gate_output_4_146(.a(output_5_146), .b(output_5_3), .y(output_4_146));
wire output_6_146, output_6_3, output_5_146;
mixer gate_output_5_146(.a(output_6_146), .b(output_6_3), .y(output_5_146));
wire output_7_146, output_7_3, output_6_146;
mixer gate_output_6_146(.a(output_7_146), .b(output_7_3), .y(output_6_146));
wire output_8_146, output_8_3, output_7_146;
mixer gate_output_7_146(.a(output_8_146), .b(output_8_3), .y(output_7_146));
wire output_1_147, output_1_4, output_0_147;
mixer gate_output_0_147(.a(output_1_147), .b(output_1_4), .y(output_0_147));
wire output_2_147, output_2_4, output_1_147;
mixer gate_output_1_147(.a(output_2_147), .b(output_2_4), .y(output_1_147));
wire output_3_147, output_3_4, output_2_147;
mixer gate_output_2_147(.a(output_3_147), .b(output_3_4), .y(output_2_147));
wire output_4_147, output_4_4, output_3_147;
mixer gate_output_3_147(.a(output_4_147), .b(output_4_4), .y(output_3_147));
wire output_5_147, output_5_4, output_4_147;
mixer gate_output_4_147(.a(output_5_147), .b(output_5_4), .y(output_4_147));
wire output_6_147, output_6_4, output_5_147;
mixer gate_output_5_147(.a(output_6_147), .b(output_6_4), .y(output_5_147));
wire output_7_147, output_7_4, output_6_147;
mixer gate_output_6_147(.a(output_7_147), .b(output_7_4), .y(output_6_147));
wire output_8_147, output_8_4, output_7_147;
mixer gate_output_7_147(.a(output_8_147), .b(output_8_4), .y(output_7_147));
wire output_1_148, output_1_5, output_0_148;
mixer gate_output_0_148(.a(output_1_148), .b(output_1_5), .y(output_0_148));
wire output_2_148, output_2_5, output_1_148;
mixer gate_output_1_148(.a(output_2_148), .b(output_2_5), .y(output_1_148));
wire output_3_148, output_3_5, output_2_148;
mixer gate_output_2_148(.a(output_3_148), .b(output_3_5), .y(output_2_148));
wire output_4_148, output_4_5, output_3_148;
mixer gate_output_3_148(.a(output_4_148), .b(output_4_5), .y(output_3_148));
wire output_5_148, output_5_5, output_4_148;
mixer gate_output_4_148(.a(output_5_148), .b(output_5_5), .y(output_4_148));
wire output_6_148, output_6_5, output_5_148;
mixer gate_output_5_148(.a(output_6_148), .b(output_6_5), .y(output_5_148));
wire output_7_148, output_7_5, output_6_148;
mixer gate_output_6_148(.a(output_7_148), .b(output_7_5), .y(output_6_148));
wire output_8_148, output_8_5, output_7_148;
mixer gate_output_7_148(.a(output_8_148), .b(output_8_5), .y(output_7_148));
wire output_1_149, output_1_6, output_0_149;
mixer gate_output_0_149(.a(output_1_149), .b(output_1_6), .y(output_0_149));
wire output_2_149, output_2_6, output_1_149;
mixer gate_output_1_149(.a(output_2_149), .b(output_2_6), .y(output_1_149));
wire output_3_149, output_3_6, output_2_149;
mixer gate_output_2_149(.a(output_3_149), .b(output_3_6), .y(output_2_149));
wire output_4_149, output_4_6, output_3_149;
mixer gate_output_3_149(.a(output_4_149), .b(output_4_6), .y(output_3_149));
wire output_5_149, output_5_6, output_4_149;
mixer gate_output_4_149(.a(output_5_149), .b(output_5_6), .y(output_4_149));
wire output_6_149, output_6_6, output_5_149;
mixer gate_output_5_149(.a(output_6_149), .b(output_6_6), .y(output_5_149));
wire output_7_149, output_7_6, output_6_149;
mixer gate_output_6_149(.a(output_7_149), .b(output_7_6), .y(output_6_149));
wire output_8_149, output_8_6, output_7_149;
mixer gate_output_7_149(.a(output_8_149), .b(output_8_6), .y(output_7_149));
wire output_1_150, output_1_7, output_0_150;
mixer gate_output_0_150(.a(output_1_150), .b(output_1_7), .y(output_0_150));
wire output_2_150, output_2_7, output_1_150;
mixer gate_output_1_150(.a(output_2_150), .b(output_2_7), .y(output_1_150));
wire output_3_150, output_3_7, output_2_150;
mixer gate_output_2_150(.a(output_3_150), .b(output_3_7), .y(output_2_150));
wire output_4_150, output_4_7, output_3_150;
mixer gate_output_3_150(.a(output_4_150), .b(output_4_7), .y(output_3_150));
wire output_5_150, output_5_7, output_4_150;
mixer gate_output_4_150(.a(output_5_150), .b(output_5_7), .y(output_4_150));
wire output_6_150, output_6_7, output_5_150;
mixer gate_output_5_150(.a(output_6_150), .b(output_6_7), .y(output_5_150));
wire output_7_150, output_7_7, output_6_150;
mixer gate_output_6_150(.a(output_7_150), .b(output_7_7), .y(output_6_150));
wire output_8_150, output_8_7, output_7_150;
mixer gate_output_7_150(.a(output_8_150), .b(output_8_7), .y(output_7_150));
wire output_1_151, output_1_0, output_0_151;
mixer gate_output_0_151(.a(output_1_151), .b(output_1_0), .y(output_0_151));
wire output_2_151, output_2_0, output_1_151;
mixer gate_output_1_151(.a(output_2_151), .b(output_2_0), .y(output_1_151));
wire output_3_151, output_3_0, output_2_151;
mixer gate_output_2_151(.a(output_3_151), .b(output_3_0), .y(output_2_151));
wire output_4_151, output_4_0, output_3_151;
mixer gate_output_3_151(.a(output_4_151), .b(output_4_0), .y(output_3_151));
wire output_5_151, output_5_0, output_4_151;
mixer gate_output_4_151(.a(output_5_151), .b(output_5_0), .y(output_4_151));
wire output_6_151, output_6_0, output_5_151;
mixer gate_output_5_151(.a(output_6_151), .b(output_6_0), .y(output_5_151));
wire output_7_151, output_7_0, output_6_151;
mixer gate_output_6_151(.a(output_7_151), .b(output_7_0), .y(output_6_151));
wire output_8_151, output_8_0, output_7_151;
mixer gate_output_7_151(.a(output_8_151), .b(output_8_0), .y(output_7_151));
wire output_1_152, output_1_1, output_0_152;
mixer gate_output_0_152(.a(output_1_152), .b(output_1_1), .y(output_0_152));
wire output_2_152, output_2_1, output_1_152;
mixer gate_output_1_152(.a(output_2_152), .b(output_2_1), .y(output_1_152));
wire output_3_152, output_3_1, output_2_152;
mixer gate_output_2_152(.a(output_3_152), .b(output_3_1), .y(output_2_152));
wire output_4_152, output_4_1, output_3_152;
mixer gate_output_3_152(.a(output_4_152), .b(output_4_1), .y(output_3_152));
wire output_5_152, output_5_1, output_4_152;
mixer gate_output_4_152(.a(output_5_152), .b(output_5_1), .y(output_4_152));
wire output_6_152, output_6_1, output_5_152;
mixer gate_output_5_152(.a(output_6_152), .b(output_6_1), .y(output_5_152));
wire output_7_152, output_7_1, output_6_152;
mixer gate_output_6_152(.a(output_7_152), .b(output_7_1), .y(output_6_152));
wire output_8_152, output_8_1, output_7_152;
mixer gate_output_7_152(.a(output_8_152), .b(output_8_1), .y(output_7_152));
wire output_1_153, output_1_2, output_0_153;
mixer gate_output_0_153(.a(output_1_153), .b(output_1_2), .y(output_0_153));
wire output_2_153, output_2_2, output_1_153;
mixer gate_output_1_153(.a(output_2_153), .b(output_2_2), .y(output_1_153));
wire output_3_153, output_3_2, output_2_153;
mixer gate_output_2_153(.a(output_3_153), .b(output_3_2), .y(output_2_153));
wire output_4_153, output_4_2, output_3_153;
mixer gate_output_3_153(.a(output_4_153), .b(output_4_2), .y(output_3_153));
wire output_5_153, output_5_2, output_4_153;
mixer gate_output_4_153(.a(output_5_153), .b(output_5_2), .y(output_4_153));
wire output_6_153, output_6_2, output_5_153;
mixer gate_output_5_153(.a(output_6_153), .b(output_6_2), .y(output_5_153));
wire output_7_153, output_7_2, output_6_153;
mixer gate_output_6_153(.a(output_7_153), .b(output_7_2), .y(output_6_153));
wire output_8_153, output_8_2, output_7_153;
mixer gate_output_7_153(.a(output_8_153), .b(output_8_2), .y(output_7_153));
wire output_1_154, output_1_3, output_0_154;
mixer gate_output_0_154(.a(output_1_154), .b(output_1_3), .y(output_0_154));
wire output_2_154, output_2_3, output_1_154;
mixer gate_output_1_154(.a(output_2_154), .b(output_2_3), .y(output_1_154));
wire output_3_154, output_3_3, output_2_154;
mixer gate_output_2_154(.a(output_3_154), .b(output_3_3), .y(output_2_154));
wire output_4_154, output_4_3, output_3_154;
mixer gate_output_3_154(.a(output_4_154), .b(output_4_3), .y(output_3_154));
wire output_5_154, output_5_3, output_4_154;
mixer gate_output_4_154(.a(output_5_154), .b(output_5_3), .y(output_4_154));
wire output_6_154, output_6_3, output_5_154;
mixer gate_output_5_154(.a(output_6_154), .b(output_6_3), .y(output_5_154));
wire output_7_154, output_7_3, output_6_154;
mixer gate_output_6_154(.a(output_7_154), .b(output_7_3), .y(output_6_154));
wire output_8_154, output_8_3, output_7_154;
mixer gate_output_7_154(.a(output_8_154), .b(output_8_3), .y(output_7_154));
wire output_1_155, output_1_4, output_0_155;
mixer gate_output_0_155(.a(output_1_155), .b(output_1_4), .y(output_0_155));
wire output_2_155, output_2_4, output_1_155;
mixer gate_output_1_155(.a(output_2_155), .b(output_2_4), .y(output_1_155));
wire output_3_155, output_3_4, output_2_155;
mixer gate_output_2_155(.a(output_3_155), .b(output_3_4), .y(output_2_155));
wire output_4_155, output_4_4, output_3_155;
mixer gate_output_3_155(.a(output_4_155), .b(output_4_4), .y(output_3_155));
wire output_5_155, output_5_4, output_4_155;
mixer gate_output_4_155(.a(output_5_155), .b(output_5_4), .y(output_4_155));
wire output_6_155, output_6_4, output_5_155;
mixer gate_output_5_155(.a(output_6_155), .b(output_6_4), .y(output_5_155));
wire output_7_155, output_7_4, output_6_155;
mixer gate_output_6_155(.a(output_7_155), .b(output_7_4), .y(output_6_155));
wire output_8_155, output_8_4, output_7_155;
mixer gate_output_7_155(.a(output_8_155), .b(output_8_4), .y(output_7_155));
wire output_1_156, output_1_5, output_0_156;
mixer gate_output_0_156(.a(output_1_156), .b(output_1_5), .y(output_0_156));
wire output_2_156, output_2_5, output_1_156;
mixer gate_output_1_156(.a(output_2_156), .b(output_2_5), .y(output_1_156));
wire output_3_156, output_3_5, output_2_156;
mixer gate_output_2_156(.a(output_3_156), .b(output_3_5), .y(output_2_156));
wire output_4_156, output_4_5, output_3_156;
mixer gate_output_3_156(.a(output_4_156), .b(output_4_5), .y(output_3_156));
wire output_5_156, output_5_5, output_4_156;
mixer gate_output_4_156(.a(output_5_156), .b(output_5_5), .y(output_4_156));
wire output_6_156, output_6_5, output_5_156;
mixer gate_output_5_156(.a(output_6_156), .b(output_6_5), .y(output_5_156));
wire output_7_156, output_7_5, output_6_156;
mixer gate_output_6_156(.a(output_7_156), .b(output_7_5), .y(output_6_156));
wire output_8_156, output_8_5, output_7_156;
mixer gate_output_7_156(.a(output_8_156), .b(output_8_5), .y(output_7_156));
wire output_1_157, output_1_6, output_0_157;
mixer gate_output_0_157(.a(output_1_157), .b(output_1_6), .y(output_0_157));
wire output_2_157, output_2_6, output_1_157;
mixer gate_output_1_157(.a(output_2_157), .b(output_2_6), .y(output_1_157));
wire output_3_157, output_3_6, output_2_157;
mixer gate_output_2_157(.a(output_3_157), .b(output_3_6), .y(output_2_157));
wire output_4_157, output_4_6, output_3_157;
mixer gate_output_3_157(.a(output_4_157), .b(output_4_6), .y(output_3_157));
wire output_5_157, output_5_6, output_4_157;
mixer gate_output_4_157(.a(output_5_157), .b(output_5_6), .y(output_4_157));
wire output_6_157, output_6_6, output_5_157;
mixer gate_output_5_157(.a(output_6_157), .b(output_6_6), .y(output_5_157));
wire output_7_157, output_7_6, output_6_157;
mixer gate_output_6_157(.a(output_7_157), .b(output_7_6), .y(output_6_157));
wire output_8_157, output_8_6, output_7_157;
mixer gate_output_7_157(.a(output_8_157), .b(output_8_6), .y(output_7_157));
wire output_1_158, output_1_7, output_0_158;
mixer gate_output_0_158(.a(output_1_158), .b(output_1_7), .y(output_0_158));
wire output_2_158, output_2_7, output_1_158;
mixer gate_output_1_158(.a(output_2_158), .b(output_2_7), .y(output_1_158));
wire output_3_158, output_3_7, output_2_158;
mixer gate_output_2_158(.a(output_3_158), .b(output_3_7), .y(output_2_158));
wire output_4_158, output_4_7, output_3_158;
mixer gate_output_3_158(.a(output_4_158), .b(output_4_7), .y(output_3_158));
wire output_5_158, output_5_7, output_4_158;
mixer gate_output_4_158(.a(output_5_158), .b(output_5_7), .y(output_4_158));
wire output_6_158, output_6_7, output_5_158;
mixer gate_output_5_158(.a(output_6_158), .b(output_6_7), .y(output_5_158));
wire output_7_158, output_7_7, output_6_158;
mixer gate_output_6_158(.a(output_7_158), .b(output_7_7), .y(output_6_158));
wire output_8_158, output_8_7, output_7_158;
mixer gate_output_7_158(.a(output_8_158), .b(output_8_7), .y(output_7_158));
wire output_1_159, output_1_0, output_0_159;
mixer gate_output_0_159(.a(output_1_159), .b(output_1_0), .y(output_0_159));
wire output_2_159, output_2_0, output_1_159;
mixer gate_output_1_159(.a(output_2_159), .b(output_2_0), .y(output_1_159));
wire output_3_159, output_3_0, output_2_159;
mixer gate_output_2_159(.a(output_3_159), .b(output_3_0), .y(output_2_159));
wire output_4_159, output_4_0, output_3_159;
mixer gate_output_3_159(.a(output_4_159), .b(output_4_0), .y(output_3_159));
wire output_5_159, output_5_0, output_4_159;
mixer gate_output_4_159(.a(output_5_159), .b(output_5_0), .y(output_4_159));
wire output_6_159, output_6_0, output_5_159;
mixer gate_output_5_159(.a(output_6_159), .b(output_6_0), .y(output_5_159));
wire output_7_159, output_7_0, output_6_159;
mixer gate_output_6_159(.a(output_7_159), .b(output_7_0), .y(output_6_159));
wire output_8_159, output_8_0, output_7_159;
mixer gate_output_7_159(.a(output_8_159), .b(output_8_0), .y(output_7_159));
wire output_1_160, output_1_1, output_0_160;
mixer gate_output_0_160(.a(output_1_160), .b(output_1_1), .y(output_0_160));
wire output_2_160, output_2_1, output_1_160;
mixer gate_output_1_160(.a(output_2_160), .b(output_2_1), .y(output_1_160));
wire output_3_160, output_3_1, output_2_160;
mixer gate_output_2_160(.a(output_3_160), .b(output_3_1), .y(output_2_160));
wire output_4_160, output_4_1, output_3_160;
mixer gate_output_3_160(.a(output_4_160), .b(output_4_1), .y(output_3_160));
wire output_5_160, output_5_1, output_4_160;
mixer gate_output_4_160(.a(output_5_160), .b(output_5_1), .y(output_4_160));
wire output_6_160, output_6_1, output_5_160;
mixer gate_output_5_160(.a(output_6_160), .b(output_6_1), .y(output_5_160));
wire output_7_160, output_7_1, output_6_160;
mixer gate_output_6_160(.a(output_7_160), .b(output_7_1), .y(output_6_160));
wire output_8_160, output_8_1, output_7_160;
mixer gate_output_7_160(.a(output_8_160), .b(output_8_1), .y(output_7_160));
wire output_1_161, output_1_2, output_0_161;
mixer gate_output_0_161(.a(output_1_161), .b(output_1_2), .y(output_0_161));
wire output_2_161, output_2_2, output_1_161;
mixer gate_output_1_161(.a(output_2_161), .b(output_2_2), .y(output_1_161));
wire output_3_161, output_3_2, output_2_161;
mixer gate_output_2_161(.a(output_3_161), .b(output_3_2), .y(output_2_161));
wire output_4_161, output_4_2, output_3_161;
mixer gate_output_3_161(.a(output_4_161), .b(output_4_2), .y(output_3_161));
wire output_5_161, output_5_2, output_4_161;
mixer gate_output_4_161(.a(output_5_161), .b(output_5_2), .y(output_4_161));
wire output_6_161, output_6_2, output_5_161;
mixer gate_output_5_161(.a(output_6_161), .b(output_6_2), .y(output_5_161));
wire output_7_161, output_7_2, output_6_161;
mixer gate_output_6_161(.a(output_7_161), .b(output_7_2), .y(output_6_161));
wire output_8_161, output_8_2, output_7_161;
mixer gate_output_7_161(.a(output_8_161), .b(output_8_2), .y(output_7_161));
wire output_1_162, output_1_3, output_0_162;
mixer gate_output_0_162(.a(output_1_162), .b(output_1_3), .y(output_0_162));
wire output_2_162, output_2_3, output_1_162;
mixer gate_output_1_162(.a(output_2_162), .b(output_2_3), .y(output_1_162));
wire output_3_162, output_3_3, output_2_162;
mixer gate_output_2_162(.a(output_3_162), .b(output_3_3), .y(output_2_162));
wire output_4_162, output_4_3, output_3_162;
mixer gate_output_3_162(.a(output_4_162), .b(output_4_3), .y(output_3_162));
wire output_5_162, output_5_3, output_4_162;
mixer gate_output_4_162(.a(output_5_162), .b(output_5_3), .y(output_4_162));
wire output_6_162, output_6_3, output_5_162;
mixer gate_output_5_162(.a(output_6_162), .b(output_6_3), .y(output_5_162));
wire output_7_162, output_7_3, output_6_162;
mixer gate_output_6_162(.a(output_7_162), .b(output_7_3), .y(output_6_162));
wire output_8_162, output_8_3, output_7_162;
mixer gate_output_7_162(.a(output_8_162), .b(output_8_3), .y(output_7_162));
wire output_1_163, output_1_4, output_0_163;
mixer gate_output_0_163(.a(output_1_163), .b(output_1_4), .y(output_0_163));
wire output_2_163, output_2_4, output_1_163;
mixer gate_output_1_163(.a(output_2_163), .b(output_2_4), .y(output_1_163));
wire output_3_163, output_3_4, output_2_163;
mixer gate_output_2_163(.a(output_3_163), .b(output_3_4), .y(output_2_163));
wire output_4_163, output_4_4, output_3_163;
mixer gate_output_3_163(.a(output_4_163), .b(output_4_4), .y(output_3_163));
wire output_5_163, output_5_4, output_4_163;
mixer gate_output_4_163(.a(output_5_163), .b(output_5_4), .y(output_4_163));
wire output_6_163, output_6_4, output_5_163;
mixer gate_output_5_163(.a(output_6_163), .b(output_6_4), .y(output_5_163));
wire output_7_163, output_7_4, output_6_163;
mixer gate_output_6_163(.a(output_7_163), .b(output_7_4), .y(output_6_163));
wire output_8_163, output_8_4, output_7_163;
mixer gate_output_7_163(.a(output_8_163), .b(output_8_4), .y(output_7_163));
wire output_1_164, output_1_5, output_0_164;
mixer gate_output_0_164(.a(output_1_164), .b(output_1_5), .y(output_0_164));
wire output_2_164, output_2_5, output_1_164;
mixer gate_output_1_164(.a(output_2_164), .b(output_2_5), .y(output_1_164));
wire output_3_164, output_3_5, output_2_164;
mixer gate_output_2_164(.a(output_3_164), .b(output_3_5), .y(output_2_164));
wire output_4_164, output_4_5, output_3_164;
mixer gate_output_3_164(.a(output_4_164), .b(output_4_5), .y(output_3_164));
wire output_5_164, output_5_5, output_4_164;
mixer gate_output_4_164(.a(output_5_164), .b(output_5_5), .y(output_4_164));
wire output_6_164, output_6_5, output_5_164;
mixer gate_output_5_164(.a(output_6_164), .b(output_6_5), .y(output_5_164));
wire output_7_164, output_7_5, output_6_164;
mixer gate_output_6_164(.a(output_7_164), .b(output_7_5), .y(output_6_164));
wire output_8_164, output_8_5, output_7_164;
mixer gate_output_7_164(.a(output_8_164), .b(output_8_5), .y(output_7_164));
wire output_1_165, output_1_6, output_0_165;
mixer gate_output_0_165(.a(output_1_165), .b(output_1_6), .y(output_0_165));
wire output_2_165, output_2_6, output_1_165;
mixer gate_output_1_165(.a(output_2_165), .b(output_2_6), .y(output_1_165));
wire output_3_165, output_3_6, output_2_165;
mixer gate_output_2_165(.a(output_3_165), .b(output_3_6), .y(output_2_165));
wire output_4_165, output_4_6, output_3_165;
mixer gate_output_3_165(.a(output_4_165), .b(output_4_6), .y(output_3_165));
wire output_5_165, output_5_6, output_4_165;
mixer gate_output_4_165(.a(output_5_165), .b(output_5_6), .y(output_4_165));
wire output_6_165, output_6_6, output_5_165;
mixer gate_output_5_165(.a(output_6_165), .b(output_6_6), .y(output_5_165));
wire output_7_165, output_7_6, output_6_165;
mixer gate_output_6_165(.a(output_7_165), .b(output_7_6), .y(output_6_165));
wire output_8_165, output_8_6, output_7_165;
mixer gate_output_7_165(.a(output_8_165), .b(output_8_6), .y(output_7_165));
wire output_1_166, output_1_7, output_0_166;
mixer gate_output_0_166(.a(output_1_166), .b(output_1_7), .y(output_0_166));
wire output_2_166, output_2_7, output_1_166;
mixer gate_output_1_166(.a(output_2_166), .b(output_2_7), .y(output_1_166));
wire output_3_166, output_3_7, output_2_166;
mixer gate_output_2_166(.a(output_3_166), .b(output_3_7), .y(output_2_166));
wire output_4_166, output_4_7, output_3_166;
mixer gate_output_3_166(.a(output_4_166), .b(output_4_7), .y(output_3_166));
wire output_5_166, output_5_7, output_4_166;
mixer gate_output_4_166(.a(output_5_166), .b(output_5_7), .y(output_4_166));
wire output_6_166, output_6_7, output_5_166;
mixer gate_output_5_166(.a(output_6_166), .b(output_6_7), .y(output_5_166));
wire output_7_166, output_7_7, output_6_166;
mixer gate_output_6_166(.a(output_7_166), .b(output_7_7), .y(output_6_166));
wire output_8_166, output_8_7, output_7_166;
mixer gate_output_7_166(.a(output_8_166), .b(output_8_7), .y(output_7_166));
wire output_1_167, output_1_0, output_0_167;
mixer gate_output_0_167(.a(output_1_167), .b(output_1_0), .y(output_0_167));
wire output_2_167, output_2_0, output_1_167;
mixer gate_output_1_167(.a(output_2_167), .b(output_2_0), .y(output_1_167));
wire output_3_167, output_3_0, output_2_167;
mixer gate_output_2_167(.a(output_3_167), .b(output_3_0), .y(output_2_167));
wire output_4_167, output_4_0, output_3_167;
mixer gate_output_3_167(.a(output_4_167), .b(output_4_0), .y(output_3_167));
wire output_5_167, output_5_0, output_4_167;
mixer gate_output_4_167(.a(output_5_167), .b(output_5_0), .y(output_4_167));
wire output_6_167, output_6_0, output_5_167;
mixer gate_output_5_167(.a(output_6_167), .b(output_6_0), .y(output_5_167));
wire output_7_167, output_7_0, output_6_167;
mixer gate_output_6_167(.a(output_7_167), .b(output_7_0), .y(output_6_167));
wire output_8_167, output_8_0, output_7_167;
mixer gate_output_7_167(.a(output_8_167), .b(output_8_0), .y(output_7_167));
wire output_1_168, output_1_1, output_0_168;
mixer gate_output_0_168(.a(output_1_168), .b(output_1_1), .y(output_0_168));
wire output_2_168, output_2_1, output_1_168;
mixer gate_output_1_168(.a(output_2_168), .b(output_2_1), .y(output_1_168));
wire output_3_168, output_3_1, output_2_168;
mixer gate_output_2_168(.a(output_3_168), .b(output_3_1), .y(output_2_168));
wire output_4_168, output_4_1, output_3_168;
mixer gate_output_3_168(.a(output_4_168), .b(output_4_1), .y(output_3_168));
wire output_5_168, output_5_1, output_4_168;
mixer gate_output_4_168(.a(output_5_168), .b(output_5_1), .y(output_4_168));
wire output_6_168, output_6_1, output_5_168;
mixer gate_output_5_168(.a(output_6_168), .b(output_6_1), .y(output_5_168));
wire output_7_168, output_7_1, output_6_168;
mixer gate_output_6_168(.a(output_7_168), .b(output_7_1), .y(output_6_168));
wire output_8_168, output_8_1, output_7_168;
mixer gate_output_7_168(.a(output_8_168), .b(output_8_1), .y(output_7_168));
wire output_1_169, output_1_2, output_0_169;
mixer gate_output_0_169(.a(output_1_169), .b(output_1_2), .y(output_0_169));
wire output_2_169, output_2_2, output_1_169;
mixer gate_output_1_169(.a(output_2_169), .b(output_2_2), .y(output_1_169));
wire output_3_169, output_3_2, output_2_169;
mixer gate_output_2_169(.a(output_3_169), .b(output_3_2), .y(output_2_169));
wire output_4_169, output_4_2, output_3_169;
mixer gate_output_3_169(.a(output_4_169), .b(output_4_2), .y(output_3_169));
wire output_5_169, output_5_2, output_4_169;
mixer gate_output_4_169(.a(output_5_169), .b(output_5_2), .y(output_4_169));
wire output_6_169, output_6_2, output_5_169;
mixer gate_output_5_169(.a(output_6_169), .b(output_6_2), .y(output_5_169));
wire output_7_169, output_7_2, output_6_169;
mixer gate_output_6_169(.a(output_7_169), .b(output_7_2), .y(output_6_169));
wire output_8_169, output_8_2, output_7_169;
mixer gate_output_7_169(.a(output_8_169), .b(output_8_2), .y(output_7_169));
wire output_1_170, output_1_3, output_0_170;
mixer gate_output_0_170(.a(output_1_170), .b(output_1_3), .y(output_0_170));
wire output_2_170, output_2_3, output_1_170;
mixer gate_output_1_170(.a(output_2_170), .b(output_2_3), .y(output_1_170));
wire output_3_170, output_3_3, output_2_170;
mixer gate_output_2_170(.a(output_3_170), .b(output_3_3), .y(output_2_170));
wire output_4_170, output_4_3, output_3_170;
mixer gate_output_3_170(.a(output_4_170), .b(output_4_3), .y(output_3_170));
wire output_5_170, output_5_3, output_4_170;
mixer gate_output_4_170(.a(output_5_170), .b(output_5_3), .y(output_4_170));
wire output_6_170, output_6_3, output_5_170;
mixer gate_output_5_170(.a(output_6_170), .b(output_6_3), .y(output_5_170));
wire output_7_170, output_7_3, output_6_170;
mixer gate_output_6_170(.a(output_7_170), .b(output_7_3), .y(output_6_170));
wire output_8_170, output_8_3, output_7_170;
mixer gate_output_7_170(.a(output_8_170), .b(output_8_3), .y(output_7_170));
wire output_1_171, output_1_4, output_0_171;
mixer gate_output_0_171(.a(output_1_171), .b(output_1_4), .y(output_0_171));
wire output_2_171, output_2_4, output_1_171;
mixer gate_output_1_171(.a(output_2_171), .b(output_2_4), .y(output_1_171));
wire output_3_171, output_3_4, output_2_171;
mixer gate_output_2_171(.a(output_3_171), .b(output_3_4), .y(output_2_171));
wire output_4_171, output_4_4, output_3_171;
mixer gate_output_3_171(.a(output_4_171), .b(output_4_4), .y(output_3_171));
wire output_5_171, output_5_4, output_4_171;
mixer gate_output_4_171(.a(output_5_171), .b(output_5_4), .y(output_4_171));
wire output_6_171, output_6_4, output_5_171;
mixer gate_output_5_171(.a(output_6_171), .b(output_6_4), .y(output_5_171));
wire output_7_171, output_7_4, output_6_171;
mixer gate_output_6_171(.a(output_7_171), .b(output_7_4), .y(output_6_171));
wire output_8_171, output_8_4, output_7_171;
mixer gate_output_7_171(.a(output_8_171), .b(output_8_4), .y(output_7_171));
wire output_1_172, output_1_5, output_0_172;
mixer gate_output_0_172(.a(output_1_172), .b(output_1_5), .y(output_0_172));
wire output_2_172, output_2_5, output_1_172;
mixer gate_output_1_172(.a(output_2_172), .b(output_2_5), .y(output_1_172));
wire output_3_172, output_3_5, output_2_172;
mixer gate_output_2_172(.a(output_3_172), .b(output_3_5), .y(output_2_172));
wire output_4_172, output_4_5, output_3_172;
mixer gate_output_3_172(.a(output_4_172), .b(output_4_5), .y(output_3_172));
wire output_5_172, output_5_5, output_4_172;
mixer gate_output_4_172(.a(output_5_172), .b(output_5_5), .y(output_4_172));
wire output_6_172, output_6_5, output_5_172;
mixer gate_output_5_172(.a(output_6_172), .b(output_6_5), .y(output_5_172));
wire output_7_172, output_7_5, output_6_172;
mixer gate_output_6_172(.a(output_7_172), .b(output_7_5), .y(output_6_172));
wire output_8_172, output_8_5, output_7_172;
mixer gate_output_7_172(.a(output_8_172), .b(output_8_5), .y(output_7_172));
wire output_1_173, output_1_6, output_0_173;
mixer gate_output_0_173(.a(output_1_173), .b(output_1_6), .y(output_0_173));
wire output_2_173, output_2_6, output_1_173;
mixer gate_output_1_173(.a(output_2_173), .b(output_2_6), .y(output_1_173));
wire output_3_173, output_3_6, output_2_173;
mixer gate_output_2_173(.a(output_3_173), .b(output_3_6), .y(output_2_173));
wire output_4_173, output_4_6, output_3_173;
mixer gate_output_3_173(.a(output_4_173), .b(output_4_6), .y(output_3_173));
wire output_5_173, output_5_6, output_4_173;
mixer gate_output_4_173(.a(output_5_173), .b(output_5_6), .y(output_4_173));
wire output_6_173, output_6_6, output_5_173;
mixer gate_output_5_173(.a(output_6_173), .b(output_6_6), .y(output_5_173));
wire output_7_173, output_7_6, output_6_173;
mixer gate_output_6_173(.a(output_7_173), .b(output_7_6), .y(output_6_173));
wire output_8_173, output_8_6, output_7_173;
mixer gate_output_7_173(.a(output_8_173), .b(output_8_6), .y(output_7_173));
wire output_1_174, output_1_7, output_0_174;
mixer gate_output_0_174(.a(output_1_174), .b(output_1_7), .y(output_0_174));
wire output_2_174, output_2_7, output_1_174;
mixer gate_output_1_174(.a(output_2_174), .b(output_2_7), .y(output_1_174));
wire output_3_174, output_3_7, output_2_174;
mixer gate_output_2_174(.a(output_3_174), .b(output_3_7), .y(output_2_174));
wire output_4_174, output_4_7, output_3_174;
mixer gate_output_3_174(.a(output_4_174), .b(output_4_7), .y(output_3_174));
wire output_5_174, output_5_7, output_4_174;
mixer gate_output_4_174(.a(output_5_174), .b(output_5_7), .y(output_4_174));
wire output_6_174, output_6_7, output_5_174;
mixer gate_output_5_174(.a(output_6_174), .b(output_6_7), .y(output_5_174));
wire output_7_174, output_7_7, output_6_174;
mixer gate_output_6_174(.a(output_7_174), .b(output_7_7), .y(output_6_174));
wire output_8_174, output_8_7, output_7_174;
mixer gate_output_7_174(.a(output_8_174), .b(output_8_7), .y(output_7_174));
wire output_1_175, output_1_0, output_0_175;
mixer gate_output_0_175(.a(output_1_175), .b(output_1_0), .y(output_0_175));
wire output_2_175, output_2_0, output_1_175;
mixer gate_output_1_175(.a(output_2_175), .b(output_2_0), .y(output_1_175));
wire output_3_175, output_3_0, output_2_175;
mixer gate_output_2_175(.a(output_3_175), .b(output_3_0), .y(output_2_175));
wire output_4_175, output_4_0, output_3_175;
mixer gate_output_3_175(.a(output_4_175), .b(output_4_0), .y(output_3_175));
wire output_5_175, output_5_0, output_4_175;
mixer gate_output_4_175(.a(output_5_175), .b(output_5_0), .y(output_4_175));
wire output_6_175, output_6_0, output_5_175;
mixer gate_output_5_175(.a(output_6_175), .b(output_6_0), .y(output_5_175));
wire output_7_175, output_7_0, output_6_175;
mixer gate_output_6_175(.a(output_7_175), .b(output_7_0), .y(output_6_175));
wire output_8_175, output_8_0, output_7_175;
mixer gate_output_7_175(.a(output_8_175), .b(output_8_0), .y(output_7_175));
wire output_1_176, output_1_1, output_0_176;
mixer gate_output_0_176(.a(output_1_176), .b(output_1_1), .y(output_0_176));
wire output_2_176, output_2_1, output_1_176;
mixer gate_output_1_176(.a(output_2_176), .b(output_2_1), .y(output_1_176));
wire output_3_176, output_3_1, output_2_176;
mixer gate_output_2_176(.a(output_3_176), .b(output_3_1), .y(output_2_176));
wire output_4_176, output_4_1, output_3_176;
mixer gate_output_3_176(.a(output_4_176), .b(output_4_1), .y(output_3_176));
wire output_5_176, output_5_1, output_4_176;
mixer gate_output_4_176(.a(output_5_176), .b(output_5_1), .y(output_4_176));
wire output_6_176, output_6_1, output_5_176;
mixer gate_output_5_176(.a(output_6_176), .b(output_6_1), .y(output_5_176));
wire output_7_176, output_7_1, output_6_176;
mixer gate_output_6_176(.a(output_7_176), .b(output_7_1), .y(output_6_176));
wire output_8_176, output_8_1, output_7_176;
mixer gate_output_7_176(.a(output_8_176), .b(output_8_1), .y(output_7_176));
wire output_1_177, output_1_2, output_0_177;
mixer gate_output_0_177(.a(output_1_177), .b(output_1_2), .y(output_0_177));
wire output_2_177, output_2_2, output_1_177;
mixer gate_output_1_177(.a(output_2_177), .b(output_2_2), .y(output_1_177));
wire output_3_177, output_3_2, output_2_177;
mixer gate_output_2_177(.a(output_3_177), .b(output_3_2), .y(output_2_177));
wire output_4_177, output_4_2, output_3_177;
mixer gate_output_3_177(.a(output_4_177), .b(output_4_2), .y(output_3_177));
wire output_5_177, output_5_2, output_4_177;
mixer gate_output_4_177(.a(output_5_177), .b(output_5_2), .y(output_4_177));
wire output_6_177, output_6_2, output_5_177;
mixer gate_output_5_177(.a(output_6_177), .b(output_6_2), .y(output_5_177));
wire output_7_177, output_7_2, output_6_177;
mixer gate_output_6_177(.a(output_7_177), .b(output_7_2), .y(output_6_177));
wire output_8_177, output_8_2, output_7_177;
mixer gate_output_7_177(.a(output_8_177), .b(output_8_2), .y(output_7_177));
wire output_1_178, output_1_3, output_0_178;
mixer gate_output_0_178(.a(output_1_178), .b(output_1_3), .y(output_0_178));
wire output_2_178, output_2_3, output_1_178;
mixer gate_output_1_178(.a(output_2_178), .b(output_2_3), .y(output_1_178));
wire output_3_178, output_3_3, output_2_178;
mixer gate_output_2_178(.a(output_3_178), .b(output_3_3), .y(output_2_178));
wire output_4_178, output_4_3, output_3_178;
mixer gate_output_3_178(.a(output_4_178), .b(output_4_3), .y(output_3_178));
wire output_5_178, output_5_3, output_4_178;
mixer gate_output_4_178(.a(output_5_178), .b(output_5_3), .y(output_4_178));
wire output_6_178, output_6_3, output_5_178;
mixer gate_output_5_178(.a(output_6_178), .b(output_6_3), .y(output_5_178));
wire output_7_178, output_7_3, output_6_178;
mixer gate_output_6_178(.a(output_7_178), .b(output_7_3), .y(output_6_178));
wire output_8_178, output_8_3, output_7_178;
mixer gate_output_7_178(.a(output_8_178), .b(output_8_3), .y(output_7_178));
wire output_1_179, output_1_4, output_0_179;
mixer gate_output_0_179(.a(output_1_179), .b(output_1_4), .y(output_0_179));
wire output_2_179, output_2_4, output_1_179;
mixer gate_output_1_179(.a(output_2_179), .b(output_2_4), .y(output_1_179));
wire output_3_179, output_3_4, output_2_179;
mixer gate_output_2_179(.a(output_3_179), .b(output_3_4), .y(output_2_179));
wire output_4_179, output_4_4, output_3_179;
mixer gate_output_3_179(.a(output_4_179), .b(output_4_4), .y(output_3_179));
wire output_5_179, output_5_4, output_4_179;
mixer gate_output_4_179(.a(output_5_179), .b(output_5_4), .y(output_4_179));
wire output_6_179, output_6_4, output_5_179;
mixer gate_output_5_179(.a(output_6_179), .b(output_6_4), .y(output_5_179));
wire output_7_179, output_7_4, output_6_179;
mixer gate_output_6_179(.a(output_7_179), .b(output_7_4), .y(output_6_179));
wire output_8_179, output_8_4, output_7_179;
mixer gate_output_7_179(.a(output_8_179), .b(output_8_4), .y(output_7_179));
wire output_1_180, output_1_5, output_0_180;
mixer gate_output_0_180(.a(output_1_180), .b(output_1_5), .y(output_0_180));
wire output_2_180, output_2_5, output_1_180;
mixer gate_output_1_180(.a(output_2_180), .b(output_2_5), .y(output_1_180));
wire output_3_180, output_3_5, output_2_180;
mixer gate_output_2_180(.a(output_3_180), .b(output_3_5), .y(output_2_180));
wire output_4_180, output_4_5, output_3_180;
mixer gate_output_3_180(.a(output_4_180), .b(output_4_5), .y(output_3_180));
wire output_5_180, output_5_5, output_4_180;
mixer gate_output_4_180(.a(output_5_180), .b(output_5_5), .y(output_4_180));
wire output_6_180, output_6_5, output_5_180;
mixer gate_output_5_180(.a(output_6_180), .b(output_6_5), .y(output_5_180));
wire output_7_180, output_7_5, output_6_180;
mixer gate_output_6_180(.a(output_7_180), .b(output_7_5), .y(output_6_180));
wire output_8_180, output_8_5, output_7_180;
mixer gate_output_7_180(.a(output_8_180), .b(output_8_5), .y(output_7_180));
wire output_1_181, output_1_6, output_0_181;
mixer gate_output_0_181(.a(output_1_181), .b(output_1_6), .y(output_0_181));
wire output_2_181, output_2_6, output_1_181;
mixer gate_output_1_181(.a(output_2_181), .b(output_2_6), .y(output_1_181));
wire output_3_181, output_3_6, output_2_181;
mixer gate_output_2_181(.a(output_3_181), .b(output_3_6), .y(output_2_181));
wire output_4_181, output_4_6, output_3_181;
mixer gate_output_3_181(.a(output_4_181), .b(output_4_6), .y(output_3_181));
wire output_5_181, output_5_6, output_4_181;
mixer gate_output_4_181(.a(output_5_181), .b(output_5_6), .y(output_4_181));
wire output_6_181, output_6_6, output_5_181;
mixer gate_output_5_181(.a(output_6_181), .b(output_6_6), .y(output_5_181));
wire output_7_181, output_7_6, output_6_181;
mixer gate_output_6_181(.a(output_7_181), .b(output_7_6), .y(output_6_181));
wire output_8_181, output_8_6, output_7_181;
mixer gate_output_7_181(.a(output_8_181), .b(output_8_6), .y(output_7_181));
wire output_1_182, output_1_7, output_0_182;
mixer gate_output_0_182(.a(output_1_182), .b(output_1_7), .y(output_0_182));
wire output_2_182, output_2_7, output_1_182;
mixer gate_output_1_182(.a(output_2_182), .b(output_2_7), .y(output_1_182));
wire output_3_182, output_3_7, output_2_182;
mixer gate_output_2_182(.a(output_3_182), .b(output_3_7), .y(output_2_182));
wire output_4_182, output_4_7, output_3_182;
mixer gate_output_3_182(.a(output_4_182), .b(output_4_7), .y(output_3_182));
wire output_5_182, output_5_7, output_4_182;
mixer gate_output_4_182(.a(output_5_182), .b(output_5_7), .y(output_4_182));
wire output_6_182, output_6_7, output_5_182;
mixer gate_output_5_182(.a(output_6_182), .b(output_6_7), .y(output_5_182));
wire output_7_182, output_7_7, output_6_182;
mixer gate_output_6_182(.a(output_7_182), .b(output_7_7), .y(output_6_182));
wire output_8_182, output_8_7, output_7_182;
mixer gate_output_7_182(.a(output_8_182), .b(output_8_7), .y(output_7_182));
wire output_1_183, output_1_0, output_0_183;
mixer gate_output_0_183(.a(output_1_183), .b(output_1_0), .y(output_0_183));
wire output_2_183, output_2_0, output_1_183;
mixer gate_output_1_183(.a(output_2_183), .b(output_2_0), .y(output_1_183));
wire output_3_183, output_3_0, output_2_183;
mixer gate_output_2_183(.a(output_3_183), .b(output_3_0), .y(output_2_183));
wire output_4_183, output_4_0, output_3_183;
mixer gate_output_3_183(.a(output_4_183), .b(output_4_0), .y(output_3_183));
wire output_5_183, output_5_0, output_4_183;
mixer gate_output_4_183(.a(output_5_183), .b(output_5_0), .y(output_4_183));
wire output_6_183, output_6_0, output_5_183;
mixer gate_output_5_183(.a(output_6_183), .b(output_6_0), .y(output_5_183));
wire output_7_183, output_7_0, output_6_183;
mixer gate_output_6_183(.a(output_7_183), .b(output_7_0), .y(output_6_183));
wire output_8_183, output_8_0, output_7_183;
mixer gate_output_7_183(.a(output_8_183), .b(output_8_0), .y(output_7_183));
wire output_1_184, output_1_1, output_0_184;
mixer gate_output_0_184(.a(output_1_184), .b(output_1_1), .y(output_0_184));
wire output_2_184, output_2_1, output_1_184;
mixer gate_output_1_184(.a(output_2_184), .b(output_2_1), .y(output_1_184));
wire output_3_184, output_3_1, output_2_184;
mixer gate_output_2_184(.a(output_3_184), .b(output_3_1), .y(output_2_184));
wire output_4_184, output_4_1, output_3_184;
mixer gate_output_3_184(.a(output_4_184), .b(output_4_1), .y(output_3_184));
wire output_5_184, output_5_1, output_4_184;
mixer gate_output_4_184(.a(output_5_184), .b(output_5_1), .y(output_4_184));
wire output_6_184, output_6_1, output_5_184;
mixer gate_output_5_184(.a(output_6_184), .b(output_6_1), .y(output_5_184));
wire output_7_184, output_7_1, output_6_184;
mixer gate_output_6_184(.a(output_7_184), .b(output_7_1), .y(output_6_184));
wire output_8_184, output_8_1, output_7_184;
mixer gate_output_7_184(.a(output_8_184), .b(output_8_1), .y(output_7_184));
wire output_1_185, output_1_2, output_0_185;
mixer gate_output_0_185(.a(output_1_185), .b(output_1_2), .y(output_0_185));
wire output_2_185, output_2_2, output_1_185;
mixer gate_output_1_185(.a(output_2_185), .b(output_2_2), .y(output_1_185));
wire output_3_185, output_3_2, output_2_185;
mixer gate_output_2_185(.a(output_3_185), .b(output_3_2), .y(output_2_185));
wire output_4_185, output_4_2, output_3_185;
mixer gate_output_3_185(.a(output_4_185), .b(output_4_2), .y(output_3_185));
wire output_5_185, output_5_2, output_4_185;
mixer gate_output_4_185(.a(output_5_185), .b(output_5_2), .y(output_4_185));
wire output_6_185, output_6_2, output_5_185;
mixer gate_output_5_185(.a(output_6_185), .b(output_6_2), .y(output_5_185));
wire output_7_185, output_7_2, output_6_185;
mixer gate_output_6_185(.a(output_7_185), .b(output_7_2), .y(output_6_185));
wire output_8_185, output_8_2, output_7_185;
mixer gate_output_7_185(.a(output_8_185), .b(output_8_2), .y(output_7_185));
wire output_1_186, output_1_3, output_0_186;
mixer gate_output_0_186(.a(output_1_186), .b(output_1_3), .y(output_0_186));
wire output_2_186, output_2_3, output_1_186;
mixer gate_output_1_186(.a(output_2_186), .b(output_2_3), .y(output_1_186));
wire output_3_186, output_3_3, output_2_186;
mixer gate_output_2_186(.a(output_3_186), .b(output_3_3), .y(output_2_186));
wire output_4_186, output_4_3, output_3_186;
mixer gate_output_3_186(.a(output_4_186), .b(output_4_3), .y(output_3_186));
wire output_5_186, output_5_3, output_4_186;
mixer gate_output_4_186(.a(output_5_186), .b(output_5_3), .y(output_4_186));
wire output_6_186, output_6_3, output_5_186;
mixer gate_output_5_186(.a(output_6_186), .b(output_6_3), .y(output_5_186));
wire output_7_186, output_7_3, output_6_186;
mixer gate_output_6_186(.a(output_7_186), .b(output_7_3), .y(output_6_186));
wire output_8_186, output_8_3, output_7_186;
mixer gate_output_7_186(.a(output_8_186), .b(output_8_3), .y(output_7_186));
wire output_1_187, output_1_4, output_0_187;
mixer gate_output_0_187(.a(output_1_187), .b(output_1_4), .y(output_0_187));
wire output_2_187, output_2_4, output_1_187;
mixer gate_output_1_187(.a(output_2_187), .b(output_2_4), .y(output_1_187));
wire output_3_187, output_3_4, output_2_187;
mixer gate_output_2_187(.a(output_3_187), .b(output_3_4), .y(output_2_187));
wire output_4_187, output_4_4, output_3_187;
mixer gate_output_3_187(.a(output_4_187), .b(output_4_4), .y(output_3_187));
wire output_5_187, output_5_4, output_4_187;
mixer gate_output_4_187(.a(output_5_187), .b(output_5_4), .y(output_4_187));
wire output_6_187, output_6_4, output_5_187;
mixer gate_output_5_187(.a(output_6_187), .b(output_6_4), .y(output_5_187));
wire output_7_187, output_7_4, output_6_187;
mixer gate_output_6_187(.a(output_7_187), .b(output_7_4), .y(output_6_187));
wire output_8_187, output_8_4, output_7_187;
mixer gate_output_7_187(.a(output_8_187), .b(output_8_4), .y(output_7_187));
wire output_1_188, output_1_5, output_0_188;
mixer gate_output_0_188(.a(output_1_188), .b(output_1_5), .y(output_0_188));
wire output_2_188, output_2_5, output_1_188;
mixer gate_output_1_188(.a(output_2_188), .b(output_2_5), .y(output_1_188));
wire output_3_188, output_3_5, output_2_188;
mixer gate_output_2_188(.a(output_3_188), .b(output_3_5), .y(output_2_188));
wire output_4_188, output_4_5, output_3_188;
mixer gate_output_3_188(.a(output_4_188), .b(output_4_5), .y(output_3_188));
wire output_5_188, output_5_5, output_4_188;
mixer gate_output_4_188(.a(output_5_188), .b(output_5_5), .y(output_4_188));
wire output_6_188, output_6_5, output_5_188;
mixer gate_output_5_188(.a(output_6_188), .b(output_6_5), .y(output_5_188));
wire output_7_188, output_7_5, output_6_188;
mixer gate_output_6_188(.a(output_7_188), .b(output_7_5), .y(output_6_188));
wire output_8_188, output_8_5, output_7_188;
mixer gate_output_7_188(.a(output_8_188), .b(output_8_5), .y(output_7_188));
wire output_1_189, output_1_6, output_0_189;
mixer gate_output_0_189(.a(output_1_189), .b(output_1_6), .y(output_0_189));
wire output_2_189, output_2_6, output_1_189;
mixer gate_output_1_189(.a(output_2_189), .b(output_2_6), .y(output_1_189));
wire output_3_189, output_3_6, output_2_189;
mixer gate_output_2_189(.a(output_3_189), .b(output_3_6), .y(output_2_189));
wire output_4_189, output_4_6, output_3_189;
mixer gate_output_3_189(.a(output_4_189), .b(output_4_6), .y(output_3_189));
wire output_5_189, output_5_6, output_4_189;
mixer gate_output_4_189(.a(output_5_189), .b(output_5_6), .y(output_4_189));
wire output_6_189, output_6_6, output_5_189;
mixer gate_output_5_189(.a(output_6_189), .b(output_6_6), .y(output_5_189));
wire output_7_189, output_7_6, output_6_189;
mixer gate_output_6_189(.a(output_7_189), .b(output_7_6), .y(output_6_189));
wire output_8_189, output_8_6, output_7_189;
mixer gate_output_7_189(.a(output_8_189), .b(output_8_6), .y(output_7_189));
wire output_1_190, output_1_7, output_0_190;
mixer gate_output_0_190(.a(output_1_190), .b(output_1_7), .y(output_0_190));
wire output_2_190, output_2_7, output_1_190;
mixer gate_output_1_190(.a(output_2_190), .b(output_2_7), .y(output_1_190));
wire output_3_190, output_3_7, output_2_190;
mixer gate_output_2_190(.a(output_3_190), .b(output_3_7), .y(output_2_190));
wire output_4_190, output_4_7, output_3_190;
mixer gate_output_3_190(.a(output_4_190), .b(output_4_7), .y(output_3_190));
wire output_5_190, output_5_7, output_4_190;
mixer gate_output_4_190(.a(output_5_190), .b(output_5_7), .y(output_4_190));
wire output_6_190, output_6_7, output_5_190;
mixer gate_output_5_190(.a(output_6_190), .b(output_6_7), .y(output_5_190));
wire output_7_190, output_7_7, output_6_190;
mixer gate_output_6_190(.a(output_7_190), .b(output_7_7), .y(output_6_190));
wire output_8_190, output_8_7, output_7_190;
mixer gate_output_7_190(.a(output_8_190), .b(output_8_7), .y(output_7_190));
wire output_1_191, output_1_0, output_0_191;
mixer gate_output_0_191(.a(output_1_191), .b(output_1_0), .y(output_0_191));
wire output_2_191, output_2_0, output_1_191;
mixer gate_output_1_191(.a(output_2_191), .b(output_2_0), .y(output_1_191));
wire output_3_191, output_3_0, output_2_191;
mixer gate_output_2_191(.a(output_3_191), .b(output_3_0), .y(output_2_191));
wire output_4_191, output_4_0, output_3_191;
mixer gate_output_3_191(.a(output_4_191), .b(output_4_0), .y(output_3_191));
wire output_5_191, output_5_0, output_4_191;
mixer gate_output_4_191(.a(output_5_191), .b(output_5_0), .y(output_4_191));
wire output_6_191, output_6_0, output_5_191;
mixer gate_output_5_191(.a(output_6_191), .b(output_6_0), .y(output_5_191));
wire output_7_191, output_7_0, output_6_191;
mixer gate_output_6_191(.a(output_7_191), .b(output_7_0), .y(output_6_191));
wire output_8_191, output_8_0, output_7_191;
mixer gate_output_7_191(.a(output_8_191), .b(output_8_0), .y(output_7_191));
wire output_1_192, output_1_1, output_0_192;
mixer gate_output_0_192(.a(output_1_192), .b(output_1_1), .y(output_0_192));
wire output_2_192, output_2_1, output_1_192;
mixer gate_output_1_192(.a(output_2_192), .b(output_2_1), .y(output_1_192));
wire output_3_192, output_3_1, output_2_192;
mixer gate_output_2_192(.a(output_3_192), .b(output_3_1), .y(output_2_192));
wire output_4_192, output_4_1, output_3_192;
mixer gate_output_3_192(.a(output_4_192), .b(output_4_1), .y(output_3_192));
wire output_5_192, output_5_1, output_4_192;
mixer gate_output_4_192(.a(output_5_192), .b(output_5_1), .y(output_4_192));
wire output_6_192, output_6_1, output_5_192;
mixer gate_output_5_192(.a(output_6_192), .b(output_6_1), .y(output_5_192));
wire output_7_192, output_7_1, output_6_192;
mixer gate_output_6_192(.a(output_7_192), .b(output_7_1), .y(output_6_192));
wire output_8_192, output_8_1, output_7_192;
mixer gate_output_7_192(.a(output_8_192), .b(output_8_1), .y(output_7_192));
wire output_1_193, output_1_2, output_0_193;
mixer gate_output_0_193(.a(output_1_193), .b(output_1_2), .y(output_0_193));
wire output_2_193, output_2_2, output_1_193;
mixer gate_output_1_193(.a(output_2_193), .b(output_2_2), .y(output_1_193));
wire output_3_193, output_3_2, output_2_193;
mixer gate_output_2_193(.a(output_3_193), .b(output_3_2), .y(output_2_193));
wire output_4_193, output_4_2, output_3_193;
mixer gate_output_3_193(.a(output_4_193), .b(output_4_2), .y(output_3_193));
wire output_5_193, output_5_2, output_4_193;
mixer gate_output_4_193(.a(output_5_193), .b(output_5_2), .y(output_4_193));
wire output_6_193, output_6_2, output_5_193;
mixer gate_output_5_193(.a(output_6_193), .b(output_6_2), .y(output_5_193));
wire output_7_193, output_7_2, output_6_193;
mixer gate_output_6_193(.a(output_7_193), .b(output_7_2), .y(output_6_193));
wire output_8_193, output_8_2, output_7_193;
mixer gate_output_7_193(.a(output_8_193), .b(output_8_2), .y(output_7_193));
wire output_1_194, output_1_3, output_0_194;
mixer gate_output_0_194(.a(output_1_194), .b(output_1_3), .y(output_0_194));
wire output_2_194, output_2_3, output_1_194;
mixer gate_output_1_194(.a(output_2_194), .b(output_2_3), .y(output_1_194));
wire output_3_194, output_3_3, output_2_194;
mixer gate_output_2_194(.a(output_3_194), .b(output_3_3), .y(output_2_194));
wire output_4_194, output_4_3, output_3_194;
mixer gate_output_3_194(.a(output_4_194), .b(output_4_3), .y(output_3_194));
wire output_5_194, output_5_3, output_4_194;
mixer gate_output_4_194(.a(output_5_194), .b(output_5_3), .y(output_4_194));
wire output_6_194, output_6_3, output_5_194;
mixer gate_output_5_194(.a(output_6_194), .b(output_6_3), .y(output_5_194));
wire output_7_194, output_7_3, output_6_194;
mixer gate_output_6_194(.a(output_7_194), .b(output_7_3), .y(output_6_194));
wire output_8_194, output_8_3, output_7_194;
mixer gate_output_7_194(.a(output_8_194), .b(output_8_3), .y(output_7_194));
wire output_1_195, output_1_4, output_0_195;
mixer gate_output_0_195(.a(output_1_195), .b(output_1_4), .y(output_0_195));
wire output_2_195, output_2_4, output_1_195;
mixer gate_output_1_195(.a(output_2_195), .b(output_2_4), .y(output_1_195));
wire output_3_195, output_3_4, output_2_195;
mixer gate_output_2_195(.a(output_3_195), .b(output_3_4), .y(output_2_195));
wire output_4_195, output_4_4, output_3_195;
mixer gate_output_3_195(.a(output_4_195), .b(output_4_4), .y(output_3_195));
wire output_5_195, output_5_4, output_4_195;
mixer gate_output_4_195(.a(output_5_195), .b(output_5_4), .y(output_4_195));
wire output_6_195, output_6_4, output_5_195;
mixer gate_output_5_195(.a(output_6_195), .b(output_6_4), .y(output_5_195));
wire output_7_195, output_7_4, output_6_195;
mixer gate_output_6_195(.a(output_7_195), .b(output_7_4), .y(output_6_195));
wire output_8_195, output_8_4, output_7_195;
mixer gate_output_7_195(.a(output_8_195), .b(output_8_4), .y(output_7_195));
wire output_1_196, output_1_5, output_0_196;
mixer gate_output_0_196(.a(output_1_196), .b(output_1_5), .y(output_0_196));
wire output_2_196, output_2_5, output_1_196;
mixer gate_output_1_196(.a(output_2_196), .b(output_2_5), .y(output_1_196));
wire output_3_196, output_3_5, output_2_196;
mixer gate_output_2_196(.a(output_3_196), .b(output_3_5), .y(output_2_196));
wire output_4_196, output_4_5, output_3_196;
mixer gate_output_3_196(.a(output_4_196), .b(output_4_5), .y(output_3_196));
wire output_5_196, output_5_5, output_4_196;
mixer gate_output_4_196(.a(output_5_196), .b(output_5_5), .y(output_4_196));
wire output_6_196, output_6_5, output_5_196;
mixer gate_output_5_196(.a(output_6_196), .b(output_6_5), .y(output_5_196));
wire output_7_196, output_7_5, output_6_196;
mixer gate_output_6_196(.a(output_7_196), .b(output_7_5), .y(output_6_196));
wire output_8_196, output_8_5, output_7_196;
mixer gate_output_7_196(.a(output_8_196), .b(output_8_5), .y(output_7_196));
wire output_1_197, output_1_6, output_0_197;
mixer gate_output_0_197(.a(output_1_197), .b(output_1_6), .y(output_0_197));
wire output_2_197, output_2_6, output_1_197;
mixer gate_output_1_197(.a(output_2_197), .b(output_2_6), .y(output_1_197));
wire output_3_197, output_3_6, output_2_197;
mixer gate_output_2_197(.a(output_3_197), .b(output_3_6), .y(output_2_197));
wire output_4_197, output_4_6, output_3_197;
mixer gate_output_3_197(.a(output_4_197), .b(output_4_6), .y(output_3_197));
wire output_5_197, output_5_6, output_4_197;
mixer gate_output_4_197(.a(output_5_197), .b(output_5_6), .y(output_4_197));
wire output_6_197, output_6_6, output_5_197;
mixer gate_output_5_197(.a(output_6_197), .b(output_6_6), .y(output_5_197));
wire output_7_197, output_7_6, output_6_197;
mixer gate_output_6_197(.a(output_7_197), .b(output_7_6), .y(output_6_197));
wire output_8_197, output_8_6, output_7_197;
mixer gate_output_7_197(.a(output_8_197), .b(output_8_6), .y(output_7_197));
wire output_1_198, output_1_7, output_0_198;
mixer gate_output_0_198(.a(output_1_198), .b(output_1_7), .y(output_0_198));
wire output_2_198, output_2_7, output_1_198;
mixer gate_output_1_198(.a(output_2_198), .b(output_2_7), .y(output_1_198));
wire output_3_198, output_3_7, output_2_198;
mixer gate_output_2_198(.a(output_3_198), .b(output_3_7), .y(output_2_198));
wire output_4_198, output_4_7, output_3_198;
mixer gate_output_3_198(.a(output_4_198), .b(output_4_7), .y(output_3_198));
wire output_5_198, output_5_7, output_4_198;
mixer gate_output_4_198(.a(output_5_198), .b(output_5_7), .y(output_4_198));
wire output_6_198, output_6_7, output_5_198;
mixer gate_output_5_198(.a(output_6_198), .b(output_6_7), .y(output_5_198));
wire output_7_198, output_7_7, output_6_198;
mixer gate_output_6_198(.a(output_7_198), .b(output_7_7), .y(output_6_198));
wire output_8_198, output_8_7, output_7_198;
mixer gate_output_7_198(.a(output_8_198), .b(output_8_7), .y(output_7_198));
wire output_1_199, output_1_0, output_0_199;
mixer gate_output_0_199(.a(output_1_199), .b(output_1_0), .y(output_0_199));
wire output_2_199, output_2_0, output_1_199;
mixer gate_output_1_199(.a(output_2_199), .b(output_2_0), .y(output_1_199));
wire output_3_199, output_3_0, output_2_199;
mixer gate_output_2_199(.a(output_3_199), .b(output_3_0), .y(output_2_199));
wire output_4_199, output_4_0, output_3_199;
mixer gate_output_3_199(.a(output_4_199), .b(output_4_0), .y(output_3_199));
wire output_5_199, output_5_0, output_4_199;
mixer gate_output_4_199(.a(output_5_199), .b(output_5_0), .y(output_4_199));
wire output_6_199, output_6_0, output_5_199;
mixer gate_output_5_199(.a(output_6_199), .b(output_6_0), .y(output_5_199));
wire output_7_199, output_7_0, output_6_199;
mixer gate_output_6_199(.a(output_7_199), .b(output_7_0), .y(output_6_199));
wire output_8_199, output_8_0, output_7_199;
mixer gate_output_7_199(.a(output_8_199), .b(output_8_0), .y(output_7_199));
wire output_1_200, output_1_1, output_0_200;
mixer gate_output_0_200(.a(output_1_200), .b(output_1_1), .y(output_0_200));
wire output_2_200, output_2_1, output_1_200;
mixer gate_output_1_200(.a(output_2_200), .b(output_2_1), .y(output_1_200));
wire output_3_200, output_3_1, output_2_200;
mixer gate_output_2_200(.a(output_3_200), .b(output_3_1), .y(output_2_200));
wire output_4_200, output_4_1, output_3_200;
mixer gate_output_3_200(.a(output_4_200), .b(output_4_1), .y(output_3_200));
wire output_5_200, output_5_1, output_4_200;
mixer gate_output_4_200(.a(output_5_200), .b(output_5_1), .y(output_4_200));
wire output_6_200, output_6_1, output_5_200;
mixer gate_output_5_200(.a(output_6_200), .b(output_6_1), .y(output_5_200));
wire output_7_200, output_7_1, output_6_200;
mixer gate_output_6_200(.a(output_7_200), .b(output_7_1), .y(output_6_200));
wire output_8_200, output_8_1, output_7_200;
mixer gate_output_7_200(.a(output_8_200), .b(output_8_1), .y(output_7_200));
wire output_1_201, output_1_2, output_0_201;
mixer gate_output_0_201(.a(output_1_201), .b(output_1_2), .y(output_0_201));
wire output_2_201, output_2_2, output_1_201;
mixer gate_output_1_201(.a(output_2_201), .b(output_2_2), .y(output_1_201));
wire output_3_201, output_3_2, output_2_201;
mixer gate_output_2_201(.a(output_3_201), .b(output_3_2), .y(output_2_201));
wire output_4_201, output_4_2, output_3_201;
mixer gate_output_3_201(.a(output_4_201), .b(output_4_2), .y(output_3_201));
wire output_5_201, output_5_2, output_4_201;
mixer gate_output_4_201(.a(output_5_201), .b(output_5_2), .y(output_4_201));
wire output_6_201, output_6_2, output_5_201;
mixer gate_output_5_201(.a(output_6_201), .b(output_6_2), .y(output_5_201));
wire output_7_201, output_7_2, output_6_201;
mixer gate_output_6_201(.a(output_7_201), .b(output_7_2), .y(output_6_201));
wire output_8_201, output_8_2, output_7_201;
mixer gate_output_7_201(.a(output_8_201), .b(output_8_2), .y(output_7_201));
wire output_1_202, output_1_3, output_0_202;
mixer gate_output_0_202(.a(output_1_202), .b(output_1_3), .y(output_0_202));
wire output_2_202, output_2_3, output_1_202;
mixer gate_output_1_202(.a(output_2_202), .b(output_2_3), .y(output_1_202));
wire output_3_202, output_3_3, output_2_202;
mixer gate_output_2_202(.a(output_3_202), .b(output_3_3), .y(output_2_202));
wire output_4_202, output_4_3, output_3_202;
mixer gate_output_3_202(.a(output_4_202), .b(output_4_3), .y(output_3_202));
wire output_5_202, output_5_3, output_4_202;
mixer gate_output_4_202(.a(output_5_202), .b(output_5_3), .y(output_4_202));
wire output_6_202, output_6_3, output_5_202;
mixer gate_output_5_202(.a(output_6_202), .b(output_6_3), .y(output_5_202));
wire output_7_202, output_7_3, output_6_202;
mixer gate_output_6_202(.a(output_7_202), .b(output_7_3), .y(output_6_202));
wire output_8_202, output_8_3, output_7_202;
mixer gate_output_7_202(.a(output_8_202), .b(output_8_3), .y(output_7_202));
wire output_1_203, output_1_4, output_0_203;
mixer gate_output_0_203(.a(output_1_203), .b(output_1_4), .y(output_0_203));
wire output_2_203, output_2_4, output_1_203;
mixer gate_output_1_203(.a(output_2_203), .b(output_2_4), .y(output_1_203));
wire output_3_203, output_3_4, output_2_203;
mixer gate_output_2_203(.a(output_3_203), .b(output_3_4), .y(output_2_203));
wire output_4_203, output_4_4, output_3_203;
mixer gate_output_3_203(.a(output_4_203), .b(output_4_4), .y(output_3_203));
wire output_5_203, output_5_4, output_4_203;
mixer gate_output_4_203(.a(output_5_203), .b(output_5_4), .y(output_4_203));
wire output_6_203, output_6_4, output_5_203;
mixer gate_output_5_203(.a(output_6_203), .b(output_6_4), .y(output_5_203));
wire output_7_203, output_7_4, output_6_203;
mixer gate_output_6_203(.a(output_7_203), .b(output_7_4), .y(output_6_203));
wire output_8_203, output_8_4, output_7_203;
mixer gate_output_7_203(.a(output_8_203), .b(output_8_4), .y(output_7_203));
wire output_1_204, output_1_5, output_0_204;
mixer gate_output_0_204(.a(output_1_204), .b(output_1_5), .y(output_0_204));
wire output_2_204, output_2_5, output_1_204;
mixer gate_output_1_204(.a(output_2_204), .b(output_2_5), .y(output_1_204));
wire output_3_204, output_3_5, output_2_204;
mixer gate_output_2_204(.a(output_3_204), .b(output_3_5), .y(output_2_204));
wire output_4_204, output_4_5, output_3_204;
mixer gate_output_3_204(.a(output_4_204), .b(output_4_5), .y(output_3_204));
wire output_5_204, output_5_5, output_4_204;
mixer gate_output_4_204(.a(output_5_204), .b(output_5_5), .y(output_4_204));
wire output_6_204, output_6_5, output_5_204;
mixer gate_output_5_204(.a(output_6_204), .b(output_6_5), .y(output_5_204));
wire output_7_204, output_7_5, output_6_204;
mixer gate_output_6_204(.a(output_7_204), .b(output_7_5), .y(output_6_204));
wire output_8_204, output_8_5, output_7_204;
mixer gate_output_7_204(.a(output_8_204), .b(output_8_5), .y(output_7_204));
wire output_1_205, output_1_6, output_0_205;
mixer gate_output_0_205(.a(output_1_205), .b(output_1_6), .y(output_0_205));
wire output_2_205, output_2_6, output_1_205;
mixer gate_output_1_205(.a(output_2_205), .b(output_2_6), .y(output_1_205));
wire output_3_205, output_3_6, output_2_205;
mixer gate_output_2_205(.a(output_3_205), .b(output_3_6), .y(output_2_205));
wire output_4_205, output_4_6, output_3_205;
mixer gate_output_3_205(.a(output_4_205), .b(output_4_6), .y(output_3_205));
wire output_5_205, output_5_6, output_4_205;
mixer gate_output_4_205(.a(output_5_205), .b(output_5_6), .y(output_4_205));
wire output_6_205, output_6_6, output_5_205;
mixer gate_output_5_205(.a(output_6_205), .b(output_6_6), .y(output_5_205));
wire output_7_205, output_7_6, output_6_205;
mixer gate_output_6_205(.a(output_7_205), .b(output_7_6), .y(output_6_205));
wire output_8_205, output_8_6, output_7_205;
mixer gate_output_7_205(.a(output_8_205), .b(output_8_6), .y(output_7_205));
wire output_1_206, output_1_7, output_0_206;
mixer gate_output_0_206(.a(output_1_206), .b(output_1_7), .y(output_0_206));
wire output_2_206, output_2_7, output_1_206;
mixer gate_output_1_206(.a(output_2_206), .b(output_2_7), .y(output_1_206));
wire output_3_206, output_3_7, output_2_206;
mixer gate_output_2_206(.a(output_3_206), .b(output_3_7), .y(output_2_206));
wire output_4_206, output_4_7, output_3_206;
mixer gate_output_3_206(.a(output_4_206), .b(output_4_7), .y(output_3_206));
wire output_5_206, output_5_7, output_4_206;
mixer gate_output_4_206(.a(output_5_206), .b(output_5_7), .y(output_4_206));
wire output_6_206, output_6_7, output_5_206;
mixer gate_output_5_206(.a(output_6_206), .b(output_6_7), .y(output_5_206));
wire output_7_206, output_7_7, output_6_206;
mixer gate_output_6_206(.a(output_7_206), .b(output_7_7), .y(output_6_206));
wire output_8_206, output_8_7, output_7_206;
mixer gate_output_7_206(.a(output_8_206), .b(output_8_7), .y(output_7_206));
wire output_1_207, output_1_0, output_0_207;
mixer gate_output_0_207(.a(output_1_207), .b(output_1_0), .y(output_0_207));
wire output_2_207, output_2_0, output_1_207;
mixer gate_output_1_207(.a(output_2_207), .b(output_2_0), .y(output_1_207));
wire output_3_207, output_3_0, output_2_207;
mixer gate_output_2_207(.a(output_3_207), .b(output_3_0), .y(output_2_207));
wire output_4_207, output_4_0, output_3_207;
mixer gate_output_3_207(.a(output_4_207), .b(output_4_0), .y(output_3_207));
wire output_5_207, output_5_0, output_4_207;
mixer gate_output_4_207(.a(output_5_207), .b(output_5_0), .y(output_4_207));
wire output_6_207, output_6_0, output_5_207;
mixer gate_output_5_207(.a(output_6_207), .b(output_6_0), .y(output_5_207));
wire output_7_207, output_7_0, output_6_207;
mixer gate_output_6_207(.a(output_7_207), .b(output_7_0), .y(output_6_207));
wire output_8_207, output_8_0, output_7_207;
mixer gate_output_7_207(.a(output_8_207), .b(output_8_0), .y(output_7_207));
wire output_1_208, output_1_1, output_0_208;
mixer gate_output_0_208(.a(output_1_208), .b(output_1_1), .y(output_0_208));
wire output_2_208, output_2_1, output_1_208;
mixer gate_output_1_208(.a(output_2_208), .b(output_2_1), .y(output_1_208));
wire output_3_208, output_3_1, output_2_208;
mixer gate_output_2_208(.a(output_3_208), .b(output_3_1), .y(output_2_208));
wire output_4_208, output_4_1, output_3_208;
mixer gate_output_3_208(.a(output_4_208), .b(output_4_1), .y(output_3_208));
wire output_5_208, output_5_1, output_4_208;
mixer gate_output_4_208(.a(output_5_208), .b(output_5_1), .y(output_4_208));
wire output_6_208, output_6_1, output_5_208;
mixer gate_output_5_208(.a(output_6_208), .b(output_6_1), .y(output_5_208));
wire output_7_208, output_7_1, output_6_208;
mixer gate_output_6_208(.a(output_7_208), .b(output_7_1), .y(output_6_208));
wire output_8_208, output_8_1, output_7_208;
mixer gate_output_7_208(.a(output_8_208), .b(output_8_1), .y(output_7_208));
wire output_1_209, output_1_2, output_0_209;
mixer gate_output_0_209(.a(output_1_209), .b(output_1_2), .y(output_0_209));
wire output_2_209, output_2_2, output_1_209;
mixer gate_output_1_209(.a(output_2_209), .b(output_2_2), .y(output_1_209));
wire output_3_209, output_3_2, output_2_209;
mixer gate_output_2_209(.a(output_3_209), .b(output_3_2), .y(output_2_209));
wire output_4_209, output_4_2, output_3_209;
mixer gate_output_3_209(.a(output_4_209), .b(output_4_2), .y(output_3_209));
wire output_5_209, output_5_2, output_4_209;
mixer gate_output_4_209(.a(output_5_209), .b(output_5_2), .y(output_4_209));
wire output_6_209, output_6_2, output_5_209;
mixer gate_output_5_209(.a(output_6_209), .b(output_6_2), .y(output_5_209));
wire output_7_209, output_7_2, output_6_209;
mixer gate_output_6_209(.a(output_7_209), .b(output_7_2), .y(output_6_209));
wire output_8_209, output_8_2, output_7_209;
mixer gate_output_7_209(.a(output_8_209), .b(output_8_2), .y(output_7_209));
wire output_1_210, output_1_3, output_0_210;
mixer gate_output_0_210(.a(output_1_210), .b(output_1_3), .y(output_0_210));
wire output_2_210, output_2_3, output_1_210;
mixer gate_output_1_210(.a(output_2_210), .b(output_2_3), .y(output_1_210));
wire output_3_210, output_3_3, output_2_210;
mixer gate_output_2_210(.a(output_3_210), .b(output_3_3), .y(output_2_210));
wire output_4_210, output_4_3, output_3_210;
mixer gate_output_3_210(.a(output_4_210), .b(output_4_3), .y(output_3_210));
wire output_5_210, output_5_3, output_4_210;
mixer gate_output_4_210(.a(output_5_210), .b(output_5_3), .y(output_4_210));
wire output_6_210, output_6_3, output_5_210;
mixer gate_output_5_210(.a(output_6_210), .b(output_6_3), .y(output_5_210));
wire output_7_210, output_7_3, output_6_210;
mixer gate_output_6_210(.a(output_7_210), .b(output_7_3), .y(output_6_210));
wire output_8_210, output_8_3, output_7_210;
mixer gate_output_7_210(.a(output_8_210), .b(output_8_3), .y(output_7_210));
wire output_1_211, output_1_4, output_0_211;
mixer gate_output_0_211(.a(output_1_211), .b(output_1_4), .y(output_0_211));
wire output_2_211, output_2_4, output_1_211;
mixer gate_output_1_211(.a(output_2_211), .b(output_2_4), .y(output_1_211));
wire output_3_211, output_3_4, output_2_211;
mixer gate_output_2_211(.a(output_3_211), .b(output_3_4), .y(output_2_211));
wire output_4_211, output_4_4, output_3_211;
mixer gate_output_3_211(.a(output_4_211), .b(output_4_4), .y(output_3_211));
wire output_5_211, output_5_4, output_4_211;
mixer gate_output_4_211(.a(output_5_211), .b(output_5_4), .y(output_4_211));
wire output_6_211, output_6_4, output_5_211;
mixer gate_output_5_211(.a(output_6_211), .b(output_6_4), .y(output_5_211));
wire output_7_211, output_7_4, output_6_211;
mixer gate_output_6_211(.a(output_7_211), .b(output_7_4), .y(output_6_211));
wire output_8_211, output_8_4, output_7_211;
mixer gate_output_7_211(.a(output_8_211), .b(output_8_4), .y(output_7_211));
wire output_1_212, output_1_5, output_0_212;
mixer gate_output_0_212(.a(output_1_212), .b(output_1_5), .y(output_0_212));
wire output_2_212, output_2_5, output_1_212;
mixer gate_output_1_212(.a(output_2_212), .b(output_2_5), .y(output_1_212));
wire output_3_212, output_3_5, output_2_212;
mixer gate_output_2_212(.a(output_3_212), .b(output_3_5), .y(output_2_212));
wire output_4_212, output_4_5, output_3_212;
mixer gate_output_3_212(.a(output_4_212), .b(output_4_5), .y(output_3_212));
wire output_5_212, output_5_5, output_4_212;
mixer gate_output_4_212(.a(output_5_212), .b(output_5_5), .y(output_4_212));
wire output_6_212, output_6_5, output_5_212;
mixer gate_output_5_212(.a(output_6_212), .b(output_6_5), .y(output_5_212));
wire output_7_212, output_7_5, output_6_212;
mixer gate_output_6_212(.a(output_7_212), .b(output_7_5), .y(output_6_212));
wire output_8_212, output_8_5, output_7_212;
mixer gate_output_7_212(.a(output_8_212), .b(output_8_5), .y(output_7_212));
wire output_1_213, output_1_6, output_0_213;
mixer gate_output_0_213(.a(output_1_213), .b(output_1_6), .y(output_0_213));
wire output_2_213, output_2_6, output_1_213;
mixer gate_output_1_213(.a(output_2_213), .b(output_2_6), .y(output_1_213));
wire output_3_213, output_3_6, output_2_213;
mixer gate_output_2_213(.a(output_3_213), .b(output_3_6), .y(output_2_213));
wire output_4_213, output_4_6, output_3_213;
mixer gate_output_3_213(.a(output_4_213), .b(output_4_6), .y(output_3_213));
wire output_5_213, output_5_6, output_4_213;
mixer gate_output_4_213(.a(output_5_213), .b(output_5_6), .y(output_4_213));
wire output_6_213, output_6_6, output_5_213;
mixer gate_output_5_213(.a(output_6_213), .b(output_6_6), .y(output_5_213));
wire output_7_213, output_7_6, output_6_213;
mixer gate_output_6_213(.a(output_7_213), .b(output_7_6), .y(output_6_213));
wire output_8_213, output_8_6, output_7_213;
mixer gate_output_7_213(.a(output_8_213), .b(output_8_6), .y(output_7_213));
wire output_1_214, output_1_7, output_0_214;
mixer gate_output_0_214(.a(output_1_214), .b(output_1_7), .y(output_0_214));
wire output_2_214, output_2_7, output_1_214;
mixer gate_output_1_214(.a(output_2_214), .b(output_2_7), .y(output_1_214));
wire output_3_214, output_3_7, output_2_214;
mixer gate_output_2_214(.a(output_3_214), .b(output_3_7), .y(output_2_214));
wire output_4_214, output_4_7, output_3_214;
mixer gate_output_3_214(.a(output_4_214), .b(output_4_7), .y(output_3_214));
wire output_5_214, output_5_7, output_4_214;
mixer gate_output_4_214(.a(output_5_214), .b(output_5_7), .y(output_4_214));
wire output_6_214, output_6_7, output_5_214;
mixer gate_output_5_214(.a(output_6_214), .b(output_6_7), .y(output_5_214));
wire output_7_214, output_7_7, output_6_214;
mixer gate_output_6_214(.a(output_7_214), .b(output_7_7), .y(output_6_214));
wire output_8_214, output_8_7, output_7_214;
mixer gate_output_7_214(.a(output_8_214), .b(output_8_7), .y(output_7_214));
wire output_1_215, output_1_0, output_0_215;
mixer gate_output_0_215(.a(output_1_215), .b(output_1_0), .y(output_0_215));
wire output_2_215, output_2_0, output_1_215;
mixer gate_output_1_215(.a(output_2_215), .b(output_2_0), .y(output_1_215));
wire output_3_215, output_3_0, output_2_215;
mixer gate_output_2_215(.a(output_3_215), .b(output_3_0), .y(output_2_215));
wire output_4_215, output_4_0, output_3_215;
mixer gate_output_3_215(.a(output_4_215), .b(output_4_0), .y(output_3_215));
wire output_5_215, output_5_0, output_4_215;
mixer gate_output_4_215(.a(output_5_215), .b(output_5_0), .y(output_4_215));
wire output_6_215, output_6_0, output_5_215;
mixer gate_output_5_215(.a(output_6_215), .b(output_6_0), .y(output_5_215));
wire output_7_215, output_7_0, output_6_215;
mixer gate_output_6_215(.a(output_7_215), .b(output_7_0), .y(output_6_215));
wire output_8_215, output_8_0, output_7_215;
mixer gate_output_7_215(.a(output_8_215), .b(output_8_0), .y(output_7_215));
wire output_1_216, output_1_1, output_0_216;
mixer gate_output_0_216(.a(output_1_216), .b(output_1_1), .y(output_0_216));
wire output_2_216, output_2_1, output_1_216;
mixer gate_output_1_216(.a(output_2_216), .b(output_2_1), .y(output_1_216));
wire output_3_216, output_3_1, output_2_216;
mixer gate_output_2_216(.a(output_3_216), .b(output_3_1), .y(output_2_216));
wire output_4_216, output_4_1, output_3_216;
mixer gate_output_3_216(.a(output_4_216), .b(output_4_1), .y(output_3_216));
wire output_5_216, output_5_1, output_4_216;
mixer gate_output_4_216(.a(output_5_216), .b(output_5_1), .y(output_4_216));
wire output_6_216, output_6_1, output_5_216;
mixer gate_output_5_216(.a(output_6_216), .b(output_6_1), .y(output_5_216));
wire output_7_216, output_7_1, output_6_216;
mixer gate_output_6_216(.a(output_7_216), .b(output_7_1), .y(output_6_216));
wire output_8_216, output_8_1, output_7_216;
mixer gate_output_7_216(.a(output_8_216), .b(output_8_1), .y(output_7_216));
wire output_1_217, output_1_2, output_0_217;
mixer gate_output_0_217(.a(output_1_217), .b(output_1_2), .y(output_0_217));
wire output_2_217, output_2_2, output_1_217;
mixer gate_output_1_217(.a(output_2_217), .b(output_2_2), .y(output_1_217));
wire output_3_217, output_3_2, output_2_217;
mixer gate_output_2_217(.a(output_3_217), .b(output_3_2), .y(output_2_217));
wire output_4_217, output_4_2, output_3_217;
mixer gate_output_3_217(.a(output_4_217), .b(output_4_2), .y(output_3_217));
wire output_5_217, output_5_2, output_4_217;
mixer gate_output_4_217(.a(output_5_217), .b(output_5_2), .y(output_4_217));
wire output_6_217, output_6_2, output_5_217;
mixer gate_output_5_217(.a(output_6_217), .b(output_6_2), .y(output_5_217));
wire output_7_217, output_7_2, output_6_217;
mixer gate_output_6_217(.a(output_7_217), .b(output_7_2), .y(output_6_217));
wire output_8_217, output_8_2, output_7_217;
mixer gate_output_7_217(.a(output_8_217), .b(output_8_2), .y(output_7_217));
wire output_1_218, output_1_3, output_0_218;
mixer gate_output_0_218(.a(output_1_218), .b(output_1_3), .y(output_0_218));
wire output_2_218, output_2_3, output_1_218;
mixer gate_output_1_218(.a(output_2_218), .b(output_2_3), .y(output_1_218));
wire output_3_218, output_3_3, output_2_218;
mixer gate_output_2_218(.a(output_3_218), .b(output_3_3), .y(output_2_218));
wire output_4_218, output_4_3, output_3_218;
mixer gate_output_3_218(.a(output_4_218), .b(output_4_3), .y(output_3_218));
wire output_5_218, output_5_3, output_4_218;
mixer gate_output_4_218(.a(output_5_218), .b(output_5_3), .y(output_4_218));
wire output_6_218, output_6_3, output_5_218;
mixer gate_output_5_218(.a(output_6_218), .b(output_6_3), .y(output_5_218));
wire output_7_218, output_7_3, output_6_218;
mixer gate_output_6_218(.a(output_7_218), .b(output_7_3), .y(output_6_218));
wire output_8_218, output_8_3, output_7_218;
mixer gate_output_7_218(.a(output_8_218), .b(output_8_3), .y(output_7_218));
wire output_1_219, output_1_4, output_0_219;
mixer gate_output_0_219(.a(output_1_219), .b(output_1_4), .y(output_0_219));
wire output_2_219, output_2_4, output_1_219;
mixer gate_output_1_219(.a(output_2_219), .b(output_2_4), .y(output_1_219));
wire output_3_219, output_3_4, output_2_219;
mixer gate_output_2_219(.a(output_3_219), .b(output_3_4), .y(output_2_219));
wire output_4_219, output_4_4, output_3_219;
mixer gate_output_3_219(.a(output_4_219), .b(output_4_4), .y(output_3_219));
wire output_5_219, output_5_4, output_4_219;
mixer gate_output_4_219(.a(output_5_219), .b(output_5_4), .y(output_4_219));
wire output_6_219, output_6_4, output_5_219;
mixer gate_output_5_219(.a(output_6_219), .b(output_6_4), .y(output_5_219));
wire output_7_219, output_7_4, output_6_219;
mixer gate_output_6_219(.a(output_7_219), .b(output_7_4), .y(output_6_219));
wire output_8_219, output_8_4, output_7_219;
mixer gate_output_7_219(.a(output_8_219), .b(output_8_4), .y(output_7_219));
wire output_1_220, output_1_5, output_0_220;
mixer gate_output_0_220(.a(output_1_220), .b(output_1_5), .y(output_0_220));
wire output_2_220, output_2_5, output_1_220;
mixer gate_output_1_220(.a(output_2_220), .b(output_2_5), .y(output_1_220));
wire output_3_220, output_3_5, output_2_220;
mixer gate_output_2_220(.a(output_3_220), .b(output_3_5), .y(output_2_220));
wire output_4_220, output_4_5, output_3_220;
mixer gate_output_3_220(.a(output_4_220), .b(output_4_5), .y(output_3_220));
wire output_5_220, output_5_5, output_4_220;
mixer gate_output_4_220(.a(output_5_220), .b(output_5_5), .y(output_4_220));
wire output_6_220, output_6_5, output_5_220;
mixer gate_output_5_220(.a(output_6_220), .b(output_6_5), .y(output_5_220));
wire output_7_220, output_7_5, output_6_220;
mixer gate_output_6_220(.a(output_7_220), .b(output_7_5), .y(output_6_220));
wire output_8_220, output_8_5, output_7_220;
mixer gate_output_7_220(.a(output_8_220), .b(output_8_5), .y(output_7_220));
wire output_1_221, output_1_6, output_0_221;
mixer gate_output_0_221(.a(output_1_221), .b(output_1_6), .y(output_0_221));
wire output_2_221, output_2_6, output_1_221;
mixer gate_output_1_221(.a(output_2_221), .b(output_2_6), .y(output_1_221));
wire output_3_221, output_3_6, output_2_221;
mixer gate_output_2_221(.a(output_3_221), .b(output_3_6), .y(output_2_221));
wire output_4_221, output_4_6, output_3_221;
mixer gate_output_3_221(.a(output_4_221), .b(output_4_6), .y(output_3_221));
wire output_5_221, output_5_6, output_4_221;
mixer gate_output_4_221(.a(output_5_221), .b(output_5_6), .y(output_4_221));
wire output_6_221, output_6_6, output_5_221;
mixer gate_output_5_221(.a(output_6_221), .b(output_6_6), .y(output_5_221));
wire output_7_221, output_7_6, output_6_221;
mixer gate_output_6_221(.a(output_7_221), .b(output_7_6), .y(output_6_221));
wire output_8_221, output_8_6, output_7_221;
mixer gate_output_7_221(.a(output_8_221), .b(output_8_6), .y(output_7_221));
wire output_1_222, output_1_7, output_0_222;
mixer gate_output_0_222(.a(output_1_222), .b(output_1_7), .y(output_0_222));
wire output_2_222, output_2_7, output_1_222;
mixer gate_output_1_222(.a(output_2_222), .b(output_2_7), .y(output_1_222));
wire output_3_222, output_3_7, output_2_222;
mixer gate_output_2_222(.a(output_3_222), .b(output_3_7), .y(output_2_222));
wire output_4_222, output_4_7, output_3_222;
mixer gate_output_3_222(.a(output_4_222), .b(output_4_7), .y(output_3_222));
wire output_5_222, output_5_7, output_4_222;
mixer gate_output_4_222(.a(output_5_222), .b(output_5_7), .y(output_4_222));
wire output_6_222, output_6_7, output_5_222;
mixer gate_output_5_222(.a(output_6_222), .b(output_6_7), .y(output_5_222));
wire output_7_222, output_7_7, output_6_222;
mixer gate_output_6_222(.a(output_7_222), .b(output_7_7), .y(output_6_222));
wire output_8_222, output_8_7, output_7_222;
mixer gate_output_7_222(.a(output_8_222), .b(output_8_7), .y(output_7_222));
wire output_1_223, output_1_0, output_0_223;
mixer gate_output_0_223(.a(output_1_223), .b(output_1_0), .y(output_0_223));
wire output_2_223, output_2_0, output_1_223;
mixer gate_output_1_223(.a(output_2_223), .b(output_2_0), .y(output_1_223));
wire output_3_223, output_3_0, output_2_223;
mixer gate_output_2_223(.a(output_3_223), .b(output_3_0), .y(output_2_223));
wire output_4_223, output_4_0, output_3_223;
mixer gate_output_3_223(.a(output_4_223), .b(output_4_0), .y(output_3_223));
wire output_5_223, output_5_0, output_4_223;
mixer gate_output_4_223(.a(output_5_223), .b(output_5_0), .y(output_4_223));
wire output_6_223, output_6_0, output_5_223;
mixer gate_output_5_223(.a(output_6_223), .b(output_6_0), .y(output_5_223));
wire output_7_223, output_7_0, output_6_223;
mixer gate_output_6_223(.a(output_7_223), .b(output_7_0), .y(output_6_223));
wire output_8_223, output_8_0, output_7_223;
mixer gate_output_7_223(.a(output_8_223), .b(output_8_0), .y(output_7_223));
wire output_1_224, output_1_1, output_0_224;
mixer gate_output_0_224(.a(output_1_224), .b(output_1_1), .y(output_0_224));
wire output_2_224, output_2_1, output_1_224;
mixer gate_output_1_224(.a(output_2_224), .b(output_2_1), .y(output_1_224));
wire output_3_224, output_3_1, output_2_224;
mixer gate_output_2_224(.a(output_3_224), .b(output_3_1), .y(output_2_224));
wire output_4_224, output_4_1, output_3_224;
mixer gate_output_3_224(.a(output_4_224), .b(output_4_1), .y(output_3_224));
wire output_5_224, output_5_1, output_4_224;
mixer gate_output_4_224(.a(output_5_224), .b(output_5_1), .y(output_4_224));
wire output_6_224, output_6_1, output_5_224;
mixer gate_output_5_224(.a(output_6_224), .b(output_6_1), .y(output_5_224));
wire output_7_224, output_7_1, output_6_224;
mixer gate_output_6_224(.a(output_7_224), .b(output_7_1), .y(output_6_224));
wire output_8_224, output_8_1, output_7_224;
mixer gate_output_7_224(.a(output_8_224), .b(output_8_1), .y(output_7_224));
wire output_1_225, output_1_2, output_0_225;
mixer gate_output_0_225(.a(output_1_225), .b(output_1_2), .y(output_0_225));
wire output_2_225, output_2_2, output_1_225;
mixer gate_output_1_225(.a(output_2_225), .b(output_2_2), .y(output_1_225));
wire output_3_225, output_3_2, output_2_225;
mixer gate_output_2_225(.a(output_3_225), .b(output_3_2), .y(output_2_225));
wire output_4_225, output_4_2, output_3_225;
mixer gate_output_3_225(.a(output_4_225), .b(output_4_2), .y(output_3_225));
wire output_5_225, output_5_2, output_4_225;
mixer gate_output_4_225(.a(output_5_225), .b(output_5_2), .y(output_4_225));
wire output_6_225, output_6_2, output_5_225;
mixer gate_output_5_225(.a(output_6_225), .b(output_6_2), .y(output_5_225));
wire output_7_225, output_7_2, output_6_225;
mixer gate_output_6_225(.a(output_7_225), .b(output_7_2), .y(output_6_225));
wire output_8_225, output_8_2, output_7_225;
mixer gate_output_7_225(.a(output_8_225), .b(output_8_2), .y(output_7_225));
wire output_1_226, output_1_3, output_0_226;
mixer gate_output_0_226(.a(output_1_226), .b(output_1_3), .y(output_0_226));
wire output_2_226, output_2_3, output_1_226;
mixer gate_output_1_226(.a(output_2_226), .b(output_2_3), .y(output_1_226));
wire output_3_226, output_3_3, output_2_226;
mixer gate_output_2_226(.a(output_3_226), .b(output_3_3), .y(output_2_226));
wire output_4_226, output_4_3, output_3_226;
mixer gate_output_3_226(.a(output_4_226), .b(output_4_3), .y(output_3_226));
wire output_5_226, output_5_3, output_4_226;
mixer gate_output_4_226(.a(output_5_226), .b(output_5_3), .y(output_4_226));
wire output_6_226, output_6_3, output_5_226;
mixer gate_output_5_226(.a(output_6_226), .b(output_6_3), .y(output_5_226));
wire output_7_226, output_7_3, output_6_226;
mixer gate_output_6_226(.a(output_7_226), .b(output_7_3), .y(output_6_226));
wire output_8_226, output_8_3, output_7_226;
mixer gate_output_7_226(.a(output_8_226), .b(output_8_3), .y(output_7_226));
wire output_1_227, output_1_4, output_0_227;
mixer gate_output_0_227(.a(output_1_227), .b(output_1_4), .y(output_0_227));
wire output_2_227, output_2_4, output_1_227;
mixer gate_output_1_227(.a(output_2_227), .b(output_2_4), .y(output_1_227));
wire output_3_227, output_3_4, output_2_227;
mixer gate_output_2_227(.a(output_3_227), .b(output_3_4), .y(output_2_227));
wire output_4_227, output_4_4, output_3_227;
mixer gate_output_3_227(.a(output_4_227), .b(output_4_4), .y(output_3_227));
wire output_5_227, output_5_4, output_4_227;
mixer gate_output_4_227(.a(output_5_227), .b(output_5_4), .y(output_4_227));
wire output_6_227, output_6_4, output_5_227;
mixer gate_output_5_227(.a(output_6_227), .b(output_6_4), .y(output_5_227));
wire output_7_227, output_7_4, output_6_227;
mixer gate_output_6_227(.a(output_7_227), .b(output_7_4), .y(output_6_227));
wire output_8_227, output_8_4, output_7_227;
mixer gate_output_7_227(.a(output_8_227), .b(output_8_4), .y(output_7_227));
wire output_1_228, output_1_5, output_0_228;
mixer gate_output_0_228(.a(output_1_228), .b(output_1_5), .y(output_0_228));
wire output_2_228, output_2_5, output_1_228;
mixer gate_output_1_228(.a(output_2_228), .b(output_2_5), .y(output_1_228));
wire output_3_228, output_3_5, output_2_228;
mixer gate_output_2_228(.a(output_3_228), .b(output_3_5), .y(output_2_228));
wire output_4_228, output_4_5, output_3_228;
mixer gate_output_3_228(.a(output_4_228), .b(output_4_5), .y(output_3_228));
wire output_5_228, output_5_5, output_4_228;
mixer gate_output_4_228(.a(output_5_228), .b(output_5_5), .y(output_4_228));
wire output_6_228, output_6_5, output_5_228;
mixer gate_output_5_228(.a(output_6_228), .b(output_6_5), .y(output_5_228));
wire output_7_228, output_7_5, output_6_228;
mixer gate_output_6_228(.a(output_7_228), .b(output_7_5), .y(output_6_228));
wire output_8_228, output_8_5, output_7_228;
mixer gate_output_7_228(.a(output_8_228), .b(output_8_5), .y(output_7_228));
wire output_1_229, output_1_6, output_0_229;
mixer gate_output_0_229(.a(output_1_229), .b(output_1_6), .y(output_0_229));
wire output_2_229, output_2_6, output_1_229;
mixer gate_output_1_229(.a(output_2_229), .b(output_2_6), .y(output_1_229));
wire output_3_229, output_3_6, output_2_229;
mixer gate_output_2_229(.a(output_3_229), .b(output_3_6), .y(output_2_229));
wire output_4_229, output_4_6, output_3_229;
mixer gate_output_3_229(.a(output_4_229), .b(output_4_6), .y(output_3_229));
wire output_5_229, output_5_6, output_4_229;
mixer gate_output_4_229(.a(output_5_229), .b(output_5_6), .y(output_4_229));
wire output_6_229, output_6_6, output_5_229;
mixer gate_output_5_229(.a(output_6_229), .b(output_6_6), .y(output_5_229));
wire output_7_229, output_7_6, output_6_229;
mixer gate_output_6_229(.a(output_7_229), .b(output_7_6), .y(output_6_229));
wire output_8_229, output_8_6, output_7_229;
mixer gate_output_7_229(.a(output_8_229), .b(output_8_6), .y(output_7_229));
wire output_1_230, output_1_7, output_0_230;
mixer gate_output_0_230(.a(output_1_230), .b(output_1_7), .y(output_0_230));
wire output_2_230, output_2_7, output_1_230;
mixer gate_output_1_230(.a(output_2_230), .b(output_2_7), .y(output_1_230));
wire output_3_230, output_3_7, output_2_230;
mixer gate_output_2_230(.a(output_3_230), .b(output_3_7), .y(output_2_230));
wire output_4_230, output_4_7, output_3_230;
mixer gate_output_3_230(.a(output_4_230), .b(output_4_7), .y(output_3_230));
wire output_5_230, output_5_7, output_4_230;
mixer gate_output_4_230(.a(output_5_230), .b(output_5_7), .y(output_4_230));
wire output_6_230, output_6_7, output_5_230;
mixer gate_output_5_230(.a(output_6_230), .b(output_6_7), .y(output_5_230));
wire output_7_230, output_7_7, output_6_230;
mixer gate_output_6_230(.a(output_7_230), .b(output_7_7), .y(output_6_230));
wire output_8_230, output_8_7, output_7_230;
mixer gate_output_7_230(.a(output_8_230), .b(output_8_7), .y(output_7_230));
wire output_1_231, output_1_0, output_0_231;
mixer gate_output_0_231(.a(output_1_231), .b(output_1_0), .y(output_0_231));
wire output_2_231, output_2_0, output_1_231;
mixer gate_output_1_231(.a(output_2_231), .b(output_2_0), .y(output_1_231));
wire output_3_231, output_3_0, output_2_231;
mixer gate_output_2_231(.a(output_3_231), .b(output_3_0), .y(output_2_231));
wire output_4_231, output_4_0, output_3_231;
mixer gate_output_3_231(.a(output_4_231), .b(output_4_0), .y(output_3_231));
wire output_5_231, output_5_0, output_4_231;
mixer gate_output_4_231(.a(output_5_231), .b(output_5_0), .y(output_4_231));
wire output_6_231, output_6_0, output_5_231;
mixer gate_output_5_231(.a(output_6_231), .b(output_6_0), .y(output_5_231));
wire output_7_231, output_7_0, output_6_231;
mixer gate_output_6_231(.a(output_7_231), .b(output_7_0), .y(output_6_231));
wire output_8_231, output_8_0, output_7_231;
mixer gate_output_7_231(.a(output_8_231), .b(output_8_0), .y(output_7_231));
wire output_1_232, output_1_1, output_0_232;
mixer gate_output_0_232(.a(output_1_232), .b(output_1_1), .y(output_0_232));
wire output_2_232, output_2_1, output_1_232;
mixer gate_output_1_232(.a(output_2_232), .b(output_2_1), .y(output_1_232));
wire output_3_232, output_3_1, output_2_232;
mixer gate_output_2_232(.a(output_3_232), .b(output_3_1), .y(output_2_232));
wire output_4_232, output_4_1, output_3_232;
mixer gate_output_3_232(.a(output_4_232), .b(output_4_1), .y(output_3_232));
wire output_5_232, output_5_1, output_4_232;
mixer gate_output_4_232(.a(output_5_232), .b(output_5_1), .y(output_4_232));
wire output_6_232, output_6_1, output_5_232;
mixer gate_output_5_232(.a(output_6_232), .b(output_6_1), .y(output_5_232));
wire output_7_232, output_7_1, output_6_232;
mixer gate_output_6_232(.a(output_7_232), .b(output_7_1), .y(output_6_232));
wire output_8_232, output_8_1, output_7_232;
mixer gate_output_7_232(.a(output_8_232), .b(output_8_1), .y(output_7_232));
wire output_1_233, output_1_2, output_0_233;
mixer gate_output_0_233(.a(output_1_233), .b(output_1_2), .y(output_0_233));
wire output_2_233, output_2_2, output_1_233;
mixer gate_output_1_233(.a(output_2_233), .b(output_2_2), .y(output_1_233));
wire output_3_233, output_3_2, output_2_233;
mixer gate_output_2_233(.a(output_3_233), .b(output_3_2), .y(output_2_233));
wire output_4_233, output_4_2, output_3_233;
mixer gate_output_3_233(.a(output_4_233), .b(output_4_2), .y(output_3_233));
wire output_5_233, output_5_2, output_4_233;
mixer gate_output_4_233(.a(output_5_233), .b(output_5_2), .y(output_4_233));
wire output_6_233, output_6_2, output_5_233;
mixer gate_output_5_233(.a(output_6_233), .b(output_6_2), .y(output_5_233));
wire output_7_233, output_7_2, output_6_233;
mixer gate_output_6_233(.a(output_7_233), .b(output_7_2), .y(output_6_233));
wire output_8_233, output_8_2, output_7_233;
mixer gate_output_7_233(.a(output_8_233), .b(output_8_2), .y(output_7_233));
wire output_1_234, output_1_3, output_0_234;
mixer gate_output_0_234(.a(output_1_234), .b(output_1_3), .y(output_0_234));
wire output_2_234, output_2_3, output_1_234;
mixer gate_output_1_234(.a(output_2_234), .b(output_2_3), .y(output_1_234));
wire output_3_234, output_3_3, output_2_234;
mixer gate_output_2_234(.a(output_3_234), .b(output_3_3), .y(output_2_234));
wire output_4_234, output_4_3, output_3_234;
mixer gate_output_3_234(.a(output_4_234), .b(output_4_3), .y(output_3_234));
wire output_5_234, output_5_3, output_4_234;
mixer gate_output_4_234(.a(output_5_234), .b(output_5_3), .y(output_4_234));
wire output_6_234, output_6_3, output_5_234;
mixer gate_output_5_234(.a(output_6_234), .b(output_6_3), .y(output_5_234));
wire output_7_234, output_7_3, output_6_234;
mixer gate_output_6_234(.a(output_7_234), .b(output_7_3), .y(output_6_234));
wire output_8_234, output_8_3, output_7_234;
mixer gate_output_7_234(.a(output_8_234), .b(output_8_3), .y(output_7_234));
wire output_1_235, output_1_4, output_0_235;
mixer gate_output_0_235(.a(output_1_235), .b(output_1_4), .y(output_0_235));
wire output_2_235, output_2_4, output_1_235;
mixer gate_output_1_235(.a(output_2_235), .b(output_2_4), .y(output_1_235));
wire output_3_235, output_3_4, output_2_235;
mixer gate_output_2_235(.a(output_3_235), .b(output_3_4), .y(output_2_235));
wire output_4_235, output_4_4, output_3_235;
mixer gate_output_3_235(.a(output_4_235), .b(output_4_4), .y(output_3_235));
wire output_5_235, output_5_4, output_4_235;
mixer gate_output_4_235(.a(output_5_235), .b(output_5_4), .y(output_4_235));
wire output_6_235, output_6_4, output_5_235;
mixer gate_output_5_235(.a(output_6_235), .b(output_6_4), .y(output_5_235));
wire output_7_235, output_7_4, output_6_235;
mixer gate_output_6_235(.a(output_7_235), .b(output_7_4), .y(output_6_235));
wire output_8_235, output_8_4, output_7_235;
mixer gate_output_7_235(.a(output_8_235), .b(output_8_4), .y(output_7_235));
wire output_1_236, output_1_5, output_0_236;
mixer gate_output_0_236(.a(output_1_236), .b(output_1_5), .y(output_0_236));
wire output_2_236, output_2_5, output_1_236;
mixer gate_output_1_236(.a(output_2_236), .b(output_2_5), .y(output_1_236));
wire output_3_236, output_3_5, output_2_236;
mixer gate_output_2_236(.a(output_3_236), .b(output_3_5), .y(output_2_236));
wire output_4_236, output_4_5, output_3_236;
mixer gate_output_3_236(.a(output_4_236), .b(output_4_5), .y(output_3_236));
wire output_5_236, output_5_5, output_4_236;
mixer gate_output_4_236(.a(output_5_236), .b(output_5_5), .y(output_4_236));
wire output_6_236, output_6_5, output_5_236;
mixer gate_output_5_236(.a(output_6_236), .b(output_6_5), .y(output_5_236));
wire output_7_236, output_7_5, output_6_236;
mixer gate_output_6_236(.a(output_7_236), .b(output_7_5), .y(output_6_236));
wire output_8_236, output_8_5, output_7_236;
mixer gate_output_7_236(.a(output_8_236), .b(output_8_5), .y(output_7_236));
wire output_1_237, output_1_6, output_0_237;
mixer gate_output_0_237(.a(output_1_237), .b(output_1_6), .y(output_0_237));
wire output_2_237, output_2_6, output_1_237;
mixer gate_output_1_237(.a(output_2_237), .b(output_2_6), .y(output_1_237));
wire output_3_237, output_3_6, output_2_237;
mixer gate_output_2_237(.a(output_3_237), .b(output_3_6), .y(output_2_237));
wire output_4_237, output_4_6, output_3_237;
mixer gate_output_3_237(.a(output_4_237), .b(output_4_6), .y(output_3_237));
wire output_5_237, output_5_6, output_4_237;
mixer gate_output_4_237(.a(output_5_237), .b(output_5_6), .y(output_4_237));
wire output_6_237, output_6_6, output_5_237;
mixer gate_output_5_237(.a(output_6_237), .b(output_6_6), .y(output_5_237));
wire output_7_237, output_7_6, output_6_237;
mixer gate_output_6_237(.a(output_7_237), .b(output_7_6), .y(output_6_237));
wire output_8_237, output_8_6, output_7_237;
mixer gate_output_7_237(.a(output_8_237), .b(output_8_6), .y(output_7_237));
wire output_1_238, output_1_7, output_0_238;
mixer gate_output_0_238(.a(output_1_238), .b(output_1_7), .y(output_0_238));
wire output_2_238, output_2_7, output_1_238;
mixer gate_output_1_238(.a(output_2_238), .b(output_2_7), .y(output_1_238));
wire output_3_238, output_3_7, output_2_238;
mixer gate_output_2_238(.a(output_3_238), .b(output_3_7), .y(output_2_238));
wire output_4_238, output_4_7, output_3_238;
mixer gate_output_3_238(.a(output_4_238), .b(output_4_7), .y(output_3_238));
wire output_5_238, output_5_7, output_4_238;
mixer gate_output_4_238(.a(output_5_238), .b(output_5_7), .y(output_4_238));
wire output_6_238, output_6_7, output_5_238;
mixer gate_output_5_238(.a(output_6_238), .b(output_6_7), .y(output_5_238));
wire output_7_238, output_7_7, output_6_238;
mixer gate_output_6_238(.a(output_7_238), .b(output_7_7), .y(output_6_238));
wire output_8_238, output_8_7, output_7_238;
mixer gate_output_7_238(.a(output_8_238), .b(output_8_7), .y(output_7_238));
wire output_1_239, output_1_0, output_0_239;
mixer gate_output_0_239(.a(output_1_239), .b(output_1_0), .y(output_0_239));
wire output_2_239, output_2_0, output_1_239;
mixer gate_output_1_239(.a(output_2_239), .b(output_2_0), .y(output_1_239));
wire output_3_239, output_3_0, output_2_239;
mixer gate_output_2_239(.a(output_3_239), .b(output_3_0), .y(output_2_239));
wire output_4_239, output_4_0, output_3_239;
mixer gate_output_3_239(.a(output_4_239), .b(output_4_0), .y(output_3_239));
wire output_5_239, output_5_0, output_4_239;
mixer gate_output_4_239(.a(output_5_239), .b(output_5_0), .y(output_4_239));
wire output_6_239, output_6_0, output_5_239;
mixer gate_output_5_239(.a(output_6_239), .b(output_6_0), .y(output_5_239));
wire output_7_239, output_7_0, output_6_239;
mixer gate_output_6_239(.a(output_7_239), .b(output_7_0), .y(output_6_239));
wire output_8_239, output_8_0, output_7_239;
mixer gate_output_7_239(.a(output_8_239), .b(output_8_0), .y(output_7_239));
wire output_1_240, output_1_1, output_0_240;
mixer gate_output_0_240(.a(output_1_240), .b(output_1_1), .y(output_0_240));
wire output_2_240, output_2_1, output_1_240;
mixer gate_output_1_240(.a(output_2_240), .b(output_2_1), .y(output_1_240));
wire output_3_240, output_3_1, output_2_240;
mixer gate_output_2_240(.a(output_3_240), .b(output_3_1), .y(output_2_240));
wire output_4_240, output_4_1, output_3_240;
mixer gate_output_3_240(.a(output_4_240), .b(output_4_1), .y(output_3_240));
wire output_5_240, output_5_1, output_4_240;
mixer gate_output_4_240(.a(output_5_240), .b(output_5_1), .y(output_4_240));
wire output_6_240, output_6_1, output_5_240;
mixer gate_output_5_240(.a(output_6_240), .b(output_6_1), .y(output_5_240));
wire output_7_240, output_7_1, output_6_240;
mixer gate_output_6_240(.a(output_7_240), .b(output_7_1), .y(output_6_240));
wire output_8_240, output_8_1, output_7_240;
mixer gate_output_7_240(.a(output_8_240), .b(output_8_1), .y(output_7_240));
wire output_1_241, output_1_2, output_0_241;
mixer gate_output_0_241(.a(output_1_241), .b(output_1_2), .y(output_0_241));
wire output_2_241, output_2_2, output_1_241;
mixer gate_output_1_241(.a(output_2_241), .b(output_2_2), .y(output_1_241));
wire output_3_241, output_3_2, output_2_241;
mixer gate_output_2_241(.a(output_3_241), .b(output_3_2), .y(output_2_241));
wire output_4_241, output_4_2, output_3_241;
mixer gate_output_3_241(.a(output_4_241), .b(output_4_2), .y(output_3_241));
wire output_5_241, output_5_2, output_4_241;
mixer gate_output_4_241(.a(output_5_241), .b(output_5_2), .y(output_4_241));
wire output_6_241, output_6_2, output_5_241;
mixer gate_output_5_241(.a(output_6_241), .b(output_6_2), .y(output_5_241));
wire output_7_241, output_7_2, output_6_241;
mixer gate_output_6_241(.a(output_7_241), .b(output_7_2), .y(output_6_241));
wire output_8_241, output_8_2, output_7_241;
mixer gate_output_7_241(.a(output_8_241), .b(output_8_2), .y(output_7_241));
wire output_1_242, output_1_3, output_0_242;
mixer gate_output_0_242(.a(output_1_242), .b(output_1_3), .y(output_0_242));
wire output_2_242, output_2_3, output_1_242;
mixer gate_output_1_242(.a(output_2_242), .b(output_2_3), .y(output_1_242));
wire output_3_242, output_3_3, output_2_242;
mixer gate_output_2_242(.a(output_3_242), .b(output_3_3), .y(output_2_242));
wire output_4_242, output_4_3, output_3_242;
mixer gate_output_3_242(.a(output_4_242), .b(output_4_3), .y(output_3_242));
wire output_5_242, output_5_3, output_4_242;
mixer gate_output_4_242(.a(output_5_242), .b(output_5_3), .y(output_4_242));
wire output_6_242, output_6_3, output_5_242;
mixer gate_output_5_242(.a(output_6_242), .b(output_6_3), .y(output_5_242));
wire output_7_242, output_7_3, output_6_242;
mixer gate_output_6_242(.a(output_7_242), .b(output_7_3), .y(output_6_242));
wire output_8_242, output_8_3, output_7_242;
mixer gate_output_7_242(.a(output_8_242), .b(output_8_3), .y(output_7_242));
wire output_1_243, output_1_4, output_0_243;
mixer gate_output_0_243(.a(output_1_243), .b(output_1_4), .y(output_0_243));
wire output_2_243, output_2_4, output_1_243;
mixer gate_output_1_243(.a(output_2_243), .b(output_2_4), .y(output_1_243));
wire output_3_243, output_3_4, output_2_243;
mixer gate_output_2_243(.a(output_3_243), .b(output_3_4), .y(output_2_243));
wire output_4_243, output_4_4, output_3_243;
mixer gate_output_3_243(.a(output_4_243), .b(output_4_4), .y(output_3_243));
wire output_5_243, output_5_4, output_4_243;
mixer gate_output_4_243(.a(output_5_243), .b(output_5_4), .y(output_4_243));
wire output_6_243, output_6_4, output_5_243;
mixer gate_output_5_243(.a(output_6_243), .b(output_6_4), .y(output_5_243));
wire output_7_243, output_7_4, output_6_243;
mixer gate_output_6_243(.a(output_7_243), .b(output_7_4), .y(output_6_243));
wire output_8_243, output_8_4, output_7_243;
mixer gate_output_7_243(.a(output_8_243), .b(output_8_4), .y(output_7_243));
wire output_1_244, output_1_5, output_0_244;
mixer gate_output_0_244(.a(output_1_244), .b(output_1_5), .y(output_0_244));
wire output_2_244, output_2_5, output_1_244;
mixer gate_output_1_244(.a(output_2_244), .b(output_2_5), .y(output_1_244));
wire output_3_244, output_3_5, output_2_244;
mixer gate_output_2_244(.a(output_3_244), .b(output_3_5), .y(output_2_244));
wire output_4_244, output_4_5, output_3_244;
mixer gate_output_3_244(.a(output_4_244), .b(output_4_5), .y(output_3_244));
wire output_5_244, output_5_5, output_4_244;
mixer gate_output_4_244(.a(output_5_244), .b(output_5_5), .y(output_4_244));
wire output_6_244, output_6_5, output_5_244;
mixer gate_output_5_244(.a(output_6_244), .b(output_6_5), .y(output_5_244));
wire output_7_244, output_7_5, output_6_244;
mixer gate_output_6_244(.a(output_7_244), .b(output_7_5), .y(output_6_244));
wire output_8_244, output_8_5, output_7_244;
mixer gate_output_7_244(.a(output_8_244), .b(output_8_5), .y(output_7_244));
wire output_1_245, output_1_6, output_0_245;
mixer gate_output_0_245(.a(output_1_245), .b(output_1_6), .y(output_0_245));
wire output_2_245, output_2_6, output_1_245;
mixer gate_output_1_245(.a(output_2_245), .b(output_2_6), .y(output_1_245));
wire output_3_245, output_3_6, output_2_245;
mixer gate_output_2_245(.a(output_3_245), .b(output_3_6), .y(output_2_245));
wire output_4_245, output_4_6, output_3_245;
mixer gate_output_3_245(.a(output_4_245), .b(output_4_6), .y(output_3_245));
wire output_5_245, output_5_6, output_4_245;
mixer gate_output_4_245(.a(output_5_245), .b(output_5_6), .y(output_4_245));
wire output_6_245, output_6_6, output_5_245;
mixer gate_output_5_245(.a(output_6_245), .b(output_6_6), .y(output_5_245));
wire output_7_245, output_7_6, output_6_245;
mixer gate_output_6_245(.a(output_7_245), .b(output_7_6), .y(output_6_245));
wire output_8_245, output_8_6, output_7_245;
mixer gate_output_7_245(.a(output_8_245), .b(output_8_6), .y(output_7_245));
wire output_1_246, output_1_7, output_0_246;
mixer gate_output_0_246(.a(output_1_246), .b(output_1_7), .y(output_0_246));
wire output_2_246, output_2_7, output_1_246;
mixer gate_output_1_246(.a(output_2_246), .b(output_2_7), .y(output_1_246));
wire output_3_246, output_3_7, output_2_246;
mixer gate_output_2_246(.a(output_3_246), .b(output_3_7), .y(output_2_246));
wire output_4_246, output_4_7, output_3_246;
mixer gate_output_3_246(.a(output_4_246), .b(output_4_7), .y(output_3_246));
wire output_5_246, output_5_7, output_4_246;
mixer gate_output_4_246(.a(output_5_246), .b(output_5_7), .y(output_4_246));
wire output_6_246, output_6_7, output_5_246;
mixer gate_output_5_246(.a(output_6_246), .b(output_6_7), .y(output_5_246));
wire output_7_246, output_7_7, output_6_246;
mixer gate_output_6_246(.a(output_7_246), .b(output_7_7), .y(output_6_246));
wire output_8_246, output_8_7, output_7_246;
mixer gate_output_7_246(.a(output_8_246), .b(output_8_7), .y(output_7_246));
wire output_1_247, output_1_0, output_0_247;
mixer gate_output_0_247(.a(output_1_247), .b(output_1_0), .y(output_0_247));
wire output_2_247, output_2_0, output_1_247;
mixer gate_output_1_247(.a(output_2_247), .b(output_2_0), .y(output_1_247));
wire output_3_247, output_3_0, output_2_247;
mixer gate_output_2_247(.a(output_3_247), .b(output_3_0), .y(output_2_247));
wire output_4_247, output_4_0, output_3_247;
mixer gate_output_3_247(.a(output_4_247), .b(output_4_0), .y(output_3_247));
wire output_5_247, output_5_0, output_4_247;
mixer gate_output_4_247(.a(output_5_247), .b(output_5_0), .y(output_4_247));
wire output_6_247, output_6_0, output_5_247;
mixer gate_output_5_247(.a(output_6_247), .b(output_6_0), .y(output_5_247));
wire output_7_247, output_7_0, output_6_247;
mixer gate_output_6_247(.a(output_7_247), .b(output_7_0), .y(output_6_247));
wire output_8_247, output_8_0, output_7_247;
mixer gate_output_7_247(.a(output_8_247), .b(output_8_0), .y(output_7_247));
wire output_1_248, output_1_1, output_0_248;
mixer gate_output_0_248(.a(output_1_248), .b(output_1_1), .y(output_0_248));
wire output_2_248, output_2_1, output_1_248;
mixer gate_output_1_248(.a(output_2_248), .b(output_2_1), .y(output_1_248));
wire output_3_248, output_3_1, output_2_248;
mixer gate_output_2_248(.a(output_3_248), .b(output_3_1), .y(output_2_248));
wire output_4_248, output_4_1, output_3_248;
mixer gate_output_3_248(.a(output_4_248), .b(output_4_1), .y(output_3_248));
wire output_5_248, output_5_1, output_4_248;
mixer gate_output_4_248(.a(output_5_248), .b(output_5_1), .y(output_4_248));
wire output_6_248, output_6_1, output_5_248;
mixer gate_output_5_248(.a(output_6_248), .b(output_6_1), .y(output_5_248));
wire output_7_248, output_7_1, output_6_248;
mixer gate_output_6_248(.a(output_7_248), .b(output_7_1), .y(output_6_248));
wire output_8_248, output_8_1, output_7_248;
mixer gate_output_7_248(.a(output_8_248), .b(output_8_1), .y(output_7_248));
wire output_1_249, output_1_2, output_0_249;
mixer gate_output_0_249(.a(output_1_249), .b(output_1_2), .y(output_0_249));
wire output_2_249, output_2_2, output_1_249;
mixer gate_output_1_249(.a(output_2_249), .b(output_2_2), .y(output_1_249));
wire output_3_249, output_3_2, output_2_249;
mixer gate_output_2_249(.a(output_3_249), .b(output_3_2), .y(output_2_249));
wire output_4_249, output_4_2, output_3_249;
mixer gate_output_3_249(.a(output_4_249), .b(output_4_2), .y(output_3_249));
wire output_5_249, output_5_2, output_4_249;
mixer gate_output_4_249(.a(output_5_249), .b(output_5_2), .y(output_4_249));
wire output_6_249, output_6_2, output_5_249;
mixer gate_output_5_249(.a(output_6_249), .b(output_6_2), .y(output_5_249));
wire output_7_249, output_7_2, output_6_249;
mixer gate_output_6_249(.a(output_7_249), .b(output_7_2), .y(output_6_249));
wire output_8_249, output_8_2, output_7_249;
mixer gate_output_7_249(.a(output_8_249), .b(output_8_2), .y(output_7_249));
wire output_1_250, output_1_3, output_0_250;
mixer gate_output_0_250(.a(output_1_250), .b(output_1_3), .y(output_0_250));
wire output_2_250, output_2_3, output_1_250;
mixer gate_output_1_250(.a(output_2_250), .b(output_2_3), .y(output_1_250));
wire output_3_250, output_3_3, output_2_250;
mixer gate_output_2_250(.a(output_3_250), .b(output_3_3), .y(output_2_250));
wire output_4_250, output_4_3, output_3_250;
mixer gate_output_3_250(.a(output_4_250), .b(output_4_3), .y(output_3_250));
wire output_5_250, output_5_3, output_4_250;
mixer gate_output_4_250(.a(output_5_250), .b(output_5_3), .y(output_4_250));
wire output_6_250, output_6_3, output_5_250;
mixer gate_output_5_250(.a(output_6_250), .b(output_6_3), .y(output_5_250));
wire output_7_250, output_7_3, output_6_250;
mixer gate_output_6_250(.a(output_7_250), .b(output_7_3), .y(output_6_250));
wire output_8_250, output_8_3, output_7_250;
mixer gate_output_7_250(.a(output_8_250), .b(output_8_3), .y(output_7_250));
wire output_1_251, output_1_4, output_0_251;
mixer gate_output_0_251(.a(output_1_251), .b(output_1_4), .y(output_0_251));
wire output_2_251, output_2_4, output_1_251;
mixer gate_output_1_251(.a(output_2_251), .b(output_2_4), .y(output_1_251));
wire output_3_251, output_3_4, output_2_251;
mixer gate_output_2_251(.a(output_3_251), .b(output_3_4), .y(output_2_251));
wire output_4_251, output_4_4, output_3_251;
mixer gate_output_3_251(.a(output_4_251), .b(output_4_4), .y(output_3_251));
wire output_5_251, output_5_4, output_4_251;
mixer gate_output_4_251(.a(output_5_251), .b(output_5_4), .y(output_4_251));
wire output_6_251, output_6_4, output_5_251;
mixer gate_output_5_251(.a(output_6_251), .b(output_6_4), .y(output_5_251));
wire output_7_251, output_7_4, output_6_251;
mixer gate_output_6_251(.a(output_7_251), .b(output_7_4), .y(output_6_251));
wire output_8_251, output_8_4, output_7_251;
mixer gate_output_7_251(.a(output_8_251), .b(output_8_4), .y(output_7_251));
wire output_1_252, output_1_5, output_0_252;
mixer gate_output_0_252(.a(output_1_252), .b(output_1_5), .y(output_0_252));
wire output_2_252, output_2_5, output_1_252;
mixer gate_output_1_252(.a(output_2_252), .b(output_2_5), .y(output_1_252));
wire output_3_252, output_3_5, output_2_252;
mixer gate_output_2_252(.a(output_3_252), .b(output_3_5), .y(output_2_252));
wire output_4_252, output_4_5, output_3_252;
mixer gate_output_3_252(.a(output_4_252), .b(output_4_5), .y(output_3_252));
wire output_5_252, output_5_5, output_4_252;
mixer gate_output_4_252(.a(output_5_252), .b(output_5_5), .y(output_4_252));
wire output_6_252, output_6_5, output_5_252;
mixer gate_output_5_252(.a(output_6_252), .b(output_6_5), .y(output_5_252));
wire output_7_252, output_7_5, output_6_252;
mixer gate_output_6_252(.a(output_7_252), .b(output_7_5), .y(output_6_252));
wire output_8_252, output_8_5, output_7_252;
mixer gate_output_7_252(.a(output_8_252), .b(output_8_5), .y(output_7_252));
wire output_1_253, output_1_6, output_0_253;
mixer gate_output_0_253(.a(output_1_253), .b(output_1_6), .y(output_0_253));
wire output_2_253, output_2_6, output_1_253;
mixer gate_output_1_253(.a(output_2_253), .b(output_2_6), .y(output_1_253));
wire output_3_253, output_3_6, output_2_253;
mixer gate_output_2_253(.a(output_3_253), .b(output_3_6), .y(output_2_253));
wire output_4_253, output_4_6, output_3_253;
mixer gate_output_3_253(.a(output_4_253), .b(output_4_6), .y(output_3_253));
wire output_5_253, output_5_6, output_4_253;
mixer gate_output_4_253(.a(output_5_253), .b(output_5_6), .y(output_4_253));
wire output_6_253, output_6_6, output_5_253;
mixer gate_output_5_253(.a(output_6_253), .b(output_6_6), .y(output_5_253));
wire output_7_253, output_7_6, output_6_253;
mixer gate_output_6_253(.a(output_7_253), .b(output_7_6), .y(output_6_253));
wire output_8_253, output_8_6, output_7_253;
mixer gate_output_7_253(.a(output_8_253), .b(output_8_6), .y(output_7_253));
wire output_1_254, output_1_7, output_0_254;
mixer gate_output_0_254(.a(output_1_254), .b(output_1_7), .y(output_0_254));
wire output_2_254, output_2_7, output_1_254;
mixer gate_output_1_254(.a(output_2_254), .b(output_2_7), .y(output_1_254));
wire output_3_254, output_3_7, output_2_254;
mixer gate_output_2_254(.a(output_3_254), .b(output_3_7), .y(output_2_254));
wire output_4_254, output_4_7, output_3_254;
mixer gate_output_3_254(.a(output_4_254), .b(output_4_7), .y(output_3_254));
wire output_5_254, output_5_7, output_4_254;
mixer gate_output_4_254(.a(output_5_254), .b(output_5_7), .y(output_4_254));
wire output_6_254, output_6_7, output_5_254;
mixer gate_output_5_254(.a(output_6_254), .b(output_6_7), .y(output_5_254));
wire output_7_254, output_7_7, output_6_254;
mixer gate_output_6_254(.a(output_7_254), .b(output_7_7), .y(output_6_254));
wire output_8_254, output_8_7, output_7_254;
mixer gate_output_7_254(.a(output_8_254), .b(output_8_7), .y(output_7_254));
wire output_1_255, output_1_0, output_0_255;
mixer gate_output_0_255(.a(output_1_255), .b(output_1_0), .y(output_0_255));
wire output_2_255, output_2_0, output_1_255;
mixer gate_output_1_255(.a(output_2_255), .b(output_2_0), .y(output_1_255));
wire output_3_255, output_3_0, output_2_255;
mixer gate_output_2_255(.a(output_3_255), .b(output_3_0), .y(output_2_255));
wire output_4_255, output_4_0, output_3_255;
mixer gate_output_3_255(.a(output_4_255), .b(output_4_0), .y(output_3_255));
wire output_5_255, output_5_0, output_4_255;
mixer gate_output_4_255(.a(output_5_255), .b(output_5_0), .y(output_4_255));
wire output_6_255, output_6_0, output_5_255;
mixer gate_output_5_255(.a(output_6_255), .b(output_6_0), .y(output_5_255));
wire output_7_255, output_7_0, output_6_255;
mixer gate_output_6_255(.a(output_7_255), .b(output_7_0), .y(output_6_255));
wire output_8_255, output_8_0, output_7_255;
mixer gate_output_7_255(.a(output_8_255), .b(output_8_0), .y(output_7_255));
wire output_1_256, output_1_1, output_0_256;
mixer gate_output_0_256(.a(output_1_256), .b(output_1_1), .y(output_0_256));
wire output_2_256, output_2_1, output_1_256;
mixer gate_output_1_256(.a(output_2_256), .b(output_2_1), .y(output_1_256));
wire output_3_256, output_3_1, output_2_256;
mixer gate_output_2_256(.a(output_3_256), .b(output_3_1), .y(output_2_256));
wire output_4_256, output_4_1, output_3_256;
mixer gate_output_3_256(.a(output_4_256), .b(output_4_1), .y(output_3_256));
wire output_5_256, output_5_1, output_4_256;
mixer gate_output_4_256(.a(output_5_256), .b(output_5_1), .y(output_4_256));
wire output_6_256, output_6_1, output_5_256;
mixer gate_output_5_256(.a(output_6_256), .b(output_6_1), .y(output_5_256));
wire output_7_256, output_7_1, output_6_256;
mixer gate_output_6_256(.a(output_7_256), .b(output_7_1), .y(output_6_256));
wire output_8_256, output_8_1, output_7_256;
mixer gate_output_7_256(.a(output_8_256), .b(output_8_1), .y(output_7_256));
wire output_1_257, output_1_2, output_0_257;
mixer gate_output_0_257(.a(output_1_257), .b(output_1_2), .y(output_0_257));
wire output_2_257, output_2_2, output_1_257;
mixer gate_output_1_257(.a(output_2_257), .b(output_2_2), .y(output_1_257));
wire output_3_257, output_3_2, output_2_257;
mixer gate_output_2_257(.a(output_3_257), .b(output_3_2), .y(output_2_257));
wire output_4_257, output_4_2, output_3_257;
mixer gate_output_3_257(.a(output_4_257), .b(output_4_2), .y(output_3_257));
wire output_5_257, output_5_2, output_4_257;
mixer gate_output_4_257(.a(output_5_257), .b(output_5_2), .y(output_4_257));
wire output_6_257, output_6_2, output_5_257;
mixer gate_output_5_257(.a(output_6_257), .b(output_6_2), .y(output_5_257));
wire output_7_257, output_7_2, output_6_257;
mixer gate_output_6_257(.a(output_7_257), .b(output_7_2), .y(output_6_257));
wire output_8_257, output_8_2, output_7_257;
mixer gate_output_7_257(.a(output_8_257), .b(output_8_2), .y(output_7_257));
wire output_1_258, output_1_3, output_0_258;
mixer gate_output_0_258(.a(output_1_258), .b(output_1_3), .y(output_0_258));
wire output_2_258, output_2_3, output_1_258;
mixer gate_output_1_258(.a(output_2_258), .b(output_2_3), .y(output_1_258));
wire output_3_258, output_3_3, output_2_258;
mixer gate_output_2_258(.a(output_3_258), .b(output_3_3), .y(output_2_258));
wire output_4_258, output_4_3, output_3_258;
mixer gate_output_3_258(.a(output_4_258), .b(output_4_3), .y(output_3_258));
wire output_5_258, output_5_3, output_4_258;
mixer gate_output_4_258(.a(output_5_258), .b(output_5_3), .y(output_4_258));
wire output_6_258, output_6_3, output_5_258;
mixer gate_output_5_258(.a(output_6_258), .b(output_6_3), .y(output_5_258));
wire output_7_258, output_7_3, output_6_258;
mixer gate_output_6_258(.a(output_7_258), .b(output_7_3), .y(output_6_258));
wire output_8_258, output_8_3, output_7_258;
mixer gate_output_7_258(.a(output_8_258), .b(output_8_3), .y(output_7_258));
wire output_1_259, output_1_4, output_0_259;
mixer gate_output_0_259(.a(output_1_259), .b(output_1_4), .y(output_0_259));
wire output_2_259, output_2_4, output_1_259;
mixer gate_output_1_259(.a(output_2_259), .b(output_2_4), .y(output_1_259));
wire output_3_259, output_3_4, output_2_259;
mixer gate_output_2_259(.a(output_3_259), .b(output_3_4), .y(output_2_259));
wire output_4_259, output_4_4, output_3_259;
mixer gate_output_3_259(.a(output_4_259), .b(output_4_4), .y(output_3_259));
wire output_5_259, output_5_4, output_4_259;
mixer gate_output_4_259(.a(output_5_259), .b(output_5_4), .y(output_4_259));
wire output_6_259, output_6_4, output_5_259;
mixer gate_output_5_259(.a(output_6_259), .b(output_6_4), .y(output_5_259));
wire output_7_259, output_7_4, output_6_259;
mixer gate_output_6_259(.a(output_7_259), .b(output_7_4), .y(output_6_259));
wire output_8_259, output_8_4, output_7_259;
mixer gate_output_7_259(.a(output_8_259), .b(output_8_4), .y(output_7_259));
wire output_1_260, output_1_5, output_0_260;
mixer gate_output_0_260(.a(output_1_260), .b(output_1_5), .y(output_0_260));
wire output_2_260, output_2_5, output_1_260;
mixer gate_output_1_260(.a(output_2_260), .b(output_2_5), .y(output_1_260));
wire output_3_260, output_3_5, output_2_260;
mixer gate_output_2_260(.a(output_3_260), .b(output_3_5), .y(output_2_260));
wire output_4_260, output_4_5, output_3_260;
mixer gate_output_3_260(.a(output_4_260), .b(output_4_5), .y(output_3_260));
wire output_5_260, output_5_5, output_4_260;
mixer gate_output_4_260(.a(output_5_260), .b(output_5_5), .y(output_4_260));
wire output_6_260, output_6_5, output_5_260;
mixer gate_output_5_260(.a(output_6_260), .b(output_6_5), .y(output_5_260));
wire output_7_260, output_7_5, output_6_260;
mixer gate_output_6_260(.a(output_7_260), .b(output_7_5), .y(output_6_260));
wire output_8_260, output_8_5, output_7_260;
mixer gate_output_7_260(.a(output_8_260), .b(output_8_5), .y(output_7_260));
wire output_1_261, output_1_6, output_0_261;
mixer gate_output_0_261(.a(output_1_261), .b(output_1_6), .y(output_0_261));
wire output_2_261, output_2_6, output_1_261;
mixer gate_output_1_261(.a(output_2_261), .b(output_2_6), .y(output_1_261));
wire output_3_261, output_3_6, output_2_261;
mixer gate_output_2_261(.a(output_3_261), .b(output_3_6), .y(output_2_261));
wire output_4_261, output_4_6, output_3_261;
mixer gate_output_3_261(.a(output_4_261), .b(output_4_6), .y(output_3_261));
wire output_5_261, output_5_6, output_4_261;
mixer gate_output_4_261(.a(output_5_261), .b(output_5_6), .y(output_4_261));
wire output_6_261, output_6_6, output_5_261;
mixer gate_output_5_261(.a(output_6_261), .b(output_6_6), .y(output_5_261));
wire output_7_261, output_7_6, output_6_261;
mixer gate_output_6_261(.a(output_7_261), .b(output_7_6), .y(output_6_261));
wire output_8_261, output_8_6, output_7_261;
mixer gate_output_7_261(.a(output_8_261), .b(output_8_6), .y(output_7_261));
wire output_1_262, output_1_7, output_0_262;
mixer gate_output_0_262(.a(output_1_262), .b(output_1_7), .y(output_0_262));
wire output_2_262, output_2_7, output_1_262;
mixer gate_output_1_262(.a(output_2_262), .b(output_2_7), .y(output_1_262));
wire output_3_262, output_3_7, output_2_262;
mixer gate_output_2_262(.a(output_3_262), .b(output_3_7), .y(output_2_262));
wire output_4_262, output_4_7, output_3_262;
mixer gate_output_3_262(.a(output_4_262), .b(output_4_7), .y(output_3_262));
wire output_5_262, output_5_7, output_4_262;
mixer gate_output_4_262(.a(output_5_262), .b(output_5_7), .y(output_4_262));
wire output_6_262, output_6_7, output_5_262;
mixer gate_output_5_262(.a(output_6_262), .b(output_6_7), .y(output_5_262));
wire output_7_262, output_7_7, output_6_262;
mixer gate_output_6_262(.a(output_7_262), .b(output_7_7), .y(output_6_262));
wire output_8_262, output_8_7, output_7_262;
mixer gate_output_7_262(.a(output_8_262), .b(output_8_7), .y(output_7_262));
wire output_1_263, output_1_0, output_0_263;
mixer gate_output_0_263(.a(output_1_263), .b(output_1_0), .y(output_0_263));
wire output_2_263, output_2_0, output_1_263;
mixer gate_output_1_263(.a(output_2_263), .b(output_2_0), .y(output_1_263));
wire output_3_263, output_3_0, output_2_263;
mixer gate_output_2_263(.a(output_3_263), .b(output_3_0), .y(output_2_263));
wire output_4_263, output_4_0, output_3_263;
mixer gate_output_3_263(.a(output_4_263), .b(output_4_0), .y(output_3_263));
wire output_5_263, output_5_0, output_4_263;
mixer gate_output_4_263(.a(output_5_263), .b(output_5_0), .y(output_4_263));
wire output_6_263, output_6_0, output_5_263;
mixer gate_output_5_263(.a(output_6_263), .b(output_6_0), .y(output_5_263));
wire output_7_263, output_7_0, output_6_263;
mixer gate_output_6_263(.a(output_7_263), .b(output_7_0), .y(output_6_263));
wire output_8_263, output_8_0, output_7_263;
mixer gate_output_7_263(.a(output_8_263), .b(output_8_0), .y(output_7_263));
wire output_1_264, output_1_1, output_0_264;
mixer gate_output_0_264(.a(output_1_264), .b(output_1_1), .y(output_0_264));
wire output_2_264, output_2_1, output_1_264;
mixer gate_output_1_264(.a(output_2_264), .b(output_2_1), .y(output_1_264));
wire output_3_264, output_3_1, output_2_264;
mixer gate_output_2_264(.a(output_3_264), .b(output_3_1), .y(output_2_264));
wire output_4_264, output_4_1, output_3_264;
mixer gate_output_3_264(.a(output_4_264), .b(output_4_1), .y(output_3_264));
wire output_5_264, output_5_1, output_4_264;
mixer gate_output_4_264(.a(output_5_264), .b(output_5_1), .y(output_4_264));
wire output_6_264, output_6_1, output_5_264;
mixer gate_output_5_264(.a(output_6_264), .b(output_6_1), .y(output_5_264));
wire output_7_264, output_7_1, output_6_264;
mixer gate_output_6_264(.a(output_7_264), .b(output_7_1), .y(output_6_264));
wire output_8_264, output_8_1, output_7_264;
mixer gate_output_7_264(.a(output_8_264), .b(output_8_1), .y(output_7_264));
wire output_1_265, output_1_2, output_0_265;
mixer gate_output_0_265(.a(output_1_265), .b(output_1_2), .y(output_0_265));
wire output_2_265, output_2_2, output_1_265;
mixer gate_output_1_265(.a(output_2_265), .b(output_2_2), .y(output_1_265));
wire output_3_265, output_3_2, output_2_265;
mixer gate_output_2_265(.a(output_3_265), .b(output_3_2), .y(output_2_265));
wire output_4_265, output_4_2, output_3_265;
mixer gate_output_3_265(.a(output_4_265), .b(output_4_2), .y(output_3_265));
wire output_5_265, output_5_2, output_4_265;
mixer gate_output_4_265(.a(output_5_265), .b(output_5_2), .y(output_4_265));
wire output_6_265, output_6_2, output_5_265;
mixer gate_output_5_265(.a(output_6_265), .b(output_6_2), .y(output_5_265));
wire output_7_265, output_7_2, output_6_265;
mixer gate_output_6_265(.a(output_7_265), .b(output_7_2), .y(output_6_265));
wire output_8_265, output_8_2, output_7_265;
mixer gate_output_7_265(.a(output_8_265), .b(output_8_2), .y(output_7_265));
wire output_1_266, output_1_3, output_0_266;
mixer gate_output_0_266(.a(output_1_266), .b(output_1_3), .y(output_0_266));
wire output_2_266, output_2_3, output_1_266;
mixer gate_output_1_266(.a(output_2_266), .b(output_2_3), .y(output_1_266));
wire output_3_266, output_3_3, output_2_266;
mixer gate_output_2_266(.a(output_3_266), .b(output_3_3), .y(output_2_266));
wire output_4_266, output_4_3, output_3_266;
mixer gate_output_3_266(.a(output_4_266), .b(output_4_3), .y(output_3_266));
wire output_5_266, output_5_3, output_4_266;
mixer gate_output_4_266(.a(output_5_266), .b(output_5_3), .y(output_4_266));
wire output_6_266, output_6_3, output_5_266;
mixer gate_output_5_266(.a(output_6_266), .b(output_6_3), .y(output_5_266));
wire output_7_266, output_7_3, output_6_266;
mixer gate_output_6_266(.a(output_7_266), .b(output_7_3), .y(output_6_266));
wire output_8_266, output_8_3, output_7_266;
mixer gate_output_7_266(.a(output_8_266), .b(output_8_3), .y(output_7_266));
wire output_1_267, output_1_4, output_0_267;
mixer gate_output_0_267(.a(output_1_267), .b(output_1_4), .y(output_0_267));
wire output_2_267, output_2_4, output_1_267;
mixer gate_output_1_267(.a(output_2_267), .b(output_2_4), .y(output_1_267));
wire output_3_267, output_3_4, output_2_267;
mixer gate_output_2_267(.a(output_3_267), .b(output_3_4), .y(output_2_267));
wire output_4_267, output_4_4, output_3_267;
mixer gate_output_3_267(.a(output_4_267), .b(output_4_4), .y(output_3_267));
wire output_5_267, output_5_4, output_4_267;
mixer gate_output_4_267(.a(output_5_267), .b(output_5_4), .y(output_4_267));
wire output_6_267, output_6_4, output_5_267;
mixer gate_output_5_267(.a(output_6_267), .b(output_6_4), .y(output_5_267));
wire output_7_267, output_7_4, output_6_267;
mixer gate_output_6_267(.a(output_7_267), .b(output_7_4), .y(output_6_267));
wire output_8_267, output_8_4, output_7_267;
mixer gate_output_7_267(.a(output_8_267), .b(output_8_4), .y(output_7_267));
wire output_1_268, output_1_5, output_0_268;
mixer gate_output_0_268(.a(output_1_268), .b(output_1_5), .y(output_0_268));
wire output_2_268, output_2_5, output_1_268;
mixer gate_output_1_268(.a(output_2_268), .b(output_2_5), .y(output_1_268));
wire output_3_268, output_3_5, output_2_268;
mixer gate_output_2_268(.a(output_3_268), .b(output_3_5), .y(output_2_268));
wire output_4_268, output_4_5, output_3_268;
mixer gate_output_3_268(.a(output_4_268), .b(output_4_5), .y(output_3_268));
wire output_5_268, output_5_5, output_4_268;
mixer gate_output_4_268(.a(output_5_268), .b(output_5_5), .y(output_4_268));
wire output_6_268, output_6_5, output_5_268;
mixer gate_output_5_268(.a(output_6_268), .b(output_6_5), .y(output_5_268));
wire output_7_268, output_7_5, output_6_268;
mixer gate_output_6_268(.a(output_7_268), .b(output_7_5), .y(output_6_268));
wire output_8_268, output_8_5, output_7_268;
mixer gate_output_7_268(.a(output_8_268), .b(output_8_5), .y(output_7_268));
wire output_1_269, output_1_6, output_0_269;
mixer gate_output_0_269(.a(output_1_269), .b(output_1_6), .y(output_0_269));
wire output_2_269, output_2_6, output_1_269;
mixer gate_output_1_269(.a(output_2_269), .b(output_2_6), .y(output_1_269));
wire output_3_269, output_3_6, output_2_269;
mixer gate_output_2_269(.a(output_3_269), .b(output_3_6), .y(output_2_269));
wire output_4_269, output_4_6, output_3_269;
mixer gate_output_3_269(.a(output_4_269), .b(output_4_6), .y(output_3_269));
wire output_5_269, output_5_6, output_4_269;
mixer gate_output_4_269(.a(output_5_269), .b(output_5_6), .y(output_4_269));
wire output_6_269, output_6_6, output_5_269;
mixer gate_output_5_269(.a(output_6_269), .b(output_6_6), .y(output_5_269));
wire output_7_269, output_7_6, output_6_269;
mixer gate_output_6_269(.a(output_7_269), .b(output_7_6), .y(output_6_269));
wire output_8_269, output_8_6, output_7_269;
mixer gate_output_7_269(.a(output_8_269), .b(output_8_6), .y(output_7_269));
wire output_1_270, output_1_7, output_0_270;
mixer gate_output_0_270(.a(output_1_270), .b(output_1_7), .y(output_0_270));
wire output_2_270, output_2_7, output_1_270;
mixer gate_output_1_270(.a(output_2_270), .b(output_2_7), .y(output_1_270));
wire output_3_270, output_3_7, output_2_270;
mixer gate_output_2_270(.a(output_3_270), .b(output_3_7), .y(output_2_270));
wire output_4_270, output_4_7, output_3_270;
mixer gate_output_3_270(.a(output_4_270), .b(output_4_7), .y(output_3_270));
wire output_5_270, output_5_7, output_4_270;
mixer gate_output_4_270(.a(output_5_270), .b(output_5_7), .y(output_4_270));
wire output_6_270, output_6_7, output_5_270;
mixer gate_output_5_270(.a(output_6_270), .b(output_6_7), .y(output_5_270));
wire output_7_270, output_7_7, output_6_270;
mixer gate_output_6_270(.a(output_7_270), .b(output_7_7), .y(output_6_270));
wire output_8_270, output_8_7, output_7_270;
mixer gate_output_7_270(.a(output_8_270), .b(output_8_7), .y(output_7_270));
wire output_1_271, output_1_0, output_0_271;
mixer gate_output_0_271(.a(output_1_271), .b(output_1_0), .y(output_0_271));
wire output_2_271, output_2_0, output_1_271;
mixer gate_output_1_271(.a(output_2_271), .b(output_2_0), .y(output_1_271));
wire output_3_271, output_3_0, output_2_271;
mixer gate_output_2_271(.a(output_3_271), .b(output_3_0), .y(output_2_271));
wire output_4_271, output_4_0, output_3_271;
mixer gate_output_3_271(.a(output_4_271), .b(output_4_0), .y(output_3_271));
wire output_5_271, output_5_0, output_4_271;
mixer gate_output_4_271(.a(output_5_271), .b(output_5_0), .y(output_4_271));
wire output_6_271, output_6_0, output_5_271;
mixer gate_output_5_271(.a(output_6_271), .b(output_6_0), .y(output_5_271));
wire output_7_271, output_7_0, output_6_271;
mixer gate_output_6_271(.a(output_7_271), .b(output_7_0), .y(output_6_271));
wire output_8_271, output_8_0, output_7_271;
mixer gate_output_7_271(.a(output_8_271), .b(output_8_0), .y(output_7_271));
wire output_1_272, output_1_1, output_0_272;
mixer gate_output_0_272(.a(output_1_272), .b(output_1_1), .y(output_0_272));
wire output_2_272, output_2_1, output_1_272;
mixer gate_output_1_272(.a(output_2_272), .b(output_2_1), .y(output_1_272));
wire output_3_272, output_3_1, output_2_272;
mixer gate_output_2_272(.a(output_3_272), .b(output_3_1), .y(output_2_272));
wire output_4_272, output_4_1, output_3_272;
mixer gate_output_3_272(.a(output_4_272), .b(output_4_1), .y(output_3_272));
wire output_5_272, output_5_1, output_4_272;
mixer gate_output_4_272(.a(output_5_272), .b(output_5_1), .y(output_4_272));
wire output_6_272, output_6_1, output_5_272;
mixer gate_output_5_272(.a(output_6_272), .b(output_6_1), .y(output_5_272));
wire output_7_272, output_7_1, output_6_272;
mixer gate_output_6_272(.a(output_7_272), .b(output_7_1), .y(output_6_272));
wire output_8_272, output_8_1, output_7_272;
mixer gate_output_7_272(.a(output_8_272), .b(output_8_1), .y(output_7_272));
wire output_1_273, output_1_2, output_0_273;
mixer gate_output_0_273(.a(output_1_273), .b(output_1_2), .y(output_0_273));
wire output_2_273, output_2_2, output_1_273;
mixer gate_output_1_273(.a(output_2_273), .b(output_2_2), .y(output_1_273));
wire output_3_273, output_3_2, output_2_273;
mixer gate_output_2_273(.a(output_3_273), .b(output_3_2), .y(output_2_273));
wire output_4_273, output_4_2, output_3_273;
mixer gate_output_3_273(.a(output_4_273), .b(output_4_2), .y(output_3_273));
wire output_5_273, output_5_2, output_4_273;
mixer gate_output_4_273(.a(output_5_273), .b(output_5_2), .y(output_4_273));
wire output_6_273, output_6_2, output_5_273;
mixer gate_output_5_273(.a(output_6_273), .b(output_6_2), .y(output_5_273));
wire output_7_273, output_7_2, output_6_273;
mixer gate_output_6_273(.a(output_7_273), .b(output_7_2), .y(output_6_273));
wire output_8_273, output_8_2, output_7_273;
mixer gate_output_7_273(.a(output_8_273), .b(output_8_2), .y(output_7_273));
wire output_1_274, output_1_3, output_0_274;
mixer gate_output_0_274(.a(output_1_274), .b(output_1_3), .y(output_0_274));
wire output_2_274, output_2_3, output_1_274;
mixer gate_output_1_274(.a(output_2_274), .b(output_2_3), .y(output_1_274));
wire output_3_274, output_3_3, output_2_274;
mixer gate_output_2_274(.a(output_3_274), .b(output_3_3), .y(output_2_274));
wire output_4_274, output_4_3, output_3_274;
mixer gate_output_3_274(.a(output_4_274), .b(output_4_3), .y(output_3_274));
wire output_5_274, output_5_3, output_4_274;
mixer gate_output_4_274(.a(output_5_274), .b(output_5_3), .y(output_4_274));
wire output_6_274, output_6_3, output_5_274;
mixer gate_output_5_274(.a(output_6_274), .b(output_6_3), .y(output_5_274));
wire output_7_274, output_7_3, output_6_274;
mixer gate_output_6_274(.a(output_7_274), .b(output_7_3), .y(output_6_274));
wire output_8_274, output_8_3, output_7_274;
mixer gate_output_7_274(.a(output_8_274), .b(output_8_3), .y(output_7_274));
wire output_1_275, output_1_4, output_0_275;
mixer gate_output_0_275(.a(output_1_275), .b(output_1_4), .y(output_0_275));
wire output_2_275, output_2_4, output_1_275;
mixer gate_output_1_275(.a(output_2_275), .b(output_2_4), .y(output_1_275));
wire output_3_275, output_3_4, output_2_275;
mixer gate_output_2_275(.a(output_3_275), .b(output_3_4), .y(output_2_275));
wire output_4_275, output_4_4, output_3_275;
mixer gate_output_3_275(.a(output_4_275), .b(output_4_4), .y(output_3_275));
wire output_5_275, output_5_4, output_4_275;
mixer gate_output_4_275(.a(output_5_275), .b(output_5_4), .y(output_4_275));
wire output_6_275, output_6_4, output_5_275;
mixer gate_output_5_275(.a(output_6_275), .b(output_6_4), .y(output_5_275));
wire output_7_275, output_7_4, output_6_275;
mixer gate_output_6_275(.a(output_7_275), .b(output_7_4), .y(output_6_275));
wire output_8_275, output_8_4, output_7_275;
mixer gate_output_7_275(.a(output_8_275), .b(output_8_4), .y(output_7_275));
wire output_1_276, output_1_5, output_0_276;
mixer gate_output_0_276(.a(output_1_276), .b(output_1_5), .y(output_0_276));
wire output_2_276, output_2_5, output_1_276;
mixer gate_output_1_276(.a(output_2_276), .b(output_2_5), .y(output_1_276));
wire output_3_276, output_3_5, output_2_276;
mixer gate_output_2_276(.a(output_3_276), .b(output_3_5), .y(output_2_276));
wire output_4_276, output_4_5, output_3_276;
mixer gate_output_3_276(.a(output_4_276), .b(output_4_5), .y(output_3_276));
wire output_5_276, output_5_5, output_4_276;
mixer gate_output_4_276(.a(output_5_276), .b(output_5_5), .y(output_4_276));
wire output_6_276, output_6_5, output_5_276;
mixer gate_output_5_276(.a(output_6_276), .b(output_6_5), .y(output_5_276));
wire output_7_276, output_7_5, output_6_276;
mixer gate_output_6_276(.a(output_7_276), .b(output_7_5), .y(output_6_276));
wire output_8_276, output_8_5, output_7_276;
mixer gate_output_7_276(.a(output_8_276), .b(output_8_5), .y(output_7_276));
wire output_1_277, output_1_6, output_0_277;
mixer gate_output_0_277(.a(output_1_277), .b(output_1_6), .y(output_0_277));
wire output_2_277, output_2_6, output_1_277;
mixer gate_output_1_277(.a(output_2_277), .b(output_2_6), .y(output_1_277));
wire output_3_277, output_3_6, output_2_277;
mixer gate_output_2_277(.a(output_3_277), .b(output_3_6), .y(output_2_277));
wire output_4_277, output_4_6, output_3_277;
mixer gate_output_3_277(.a(output_4_277), .b(output_4_6), .y(output_3_277));
wire output_5_277, output_5_6, output_4_277;
mixer gate_output_4_277(.a(output_5_277), .b(output_5_6), .y(output_4_277));
wire output_6_277, output_6_6, output_5_277;
mixer gate_output_5_277(.a(output_6_277), .b(output_6_6), .y(output_5_277));
wire output_7_277, output_7_6, output_6_277;
mixer gate_output_6_277(.a(output_7_277), .b(output_7_6), .y(output_6_277));
wire output_8_277, output_8_6, output_7_277;
mixer gate_output_7_277(.a(output_8_277), .b(output_8_6), .y(output_7_277));
wire output_1_278, output_1_7, output_0_278;
mixer gate_output_0_278(.a(output_1_278), .b(output_1_7), .y(output_0_278));
wire output_2_278, output_2_7, output_1_278;
mixer gate_output_1_278(.a(output_2_278), .b(output_2_7), .y(output_1_278));
wire output_3_278, output_3_7, output_2_278;
mixer gate_output_2_278(.a(output_3_278), .b(output_3_7), .y(output_2_278));
wire output_4_278, output_4_7, output_3_278;
mixer gate_output_3_278(.a(output_4_278), .b(output_4_7), .y(output_3_278));
wire output_5_278, output_5_7, output_4_278;
mixer gate_output_4_278(.a(output_5_278), .b(output_5_7), .y(output_4_278));
wire output_6_278, output_6_7, output_5_278;
mixer gate_output_5_278(.a(output_6_278), .b(output_6_7), .y(output_5_278));
wire output_7_278, output_7_7, output_6_278;
mixer gate_output_6_278(.a(output_7_278), .b(output_7_7), .y(output_6_278));
wire output_8_278, output_8_7, output_7_278;
mixer gate_output_7_278(.a(output_8_278), .b(output_8_7), .y(output_7_278));
wire output_1_279, output_1_0, output_0_279;
mixer gate_output_0_279(.a(output_1_279), .b(output_1_0), .y(output_0_279));
wire output_2_279, output_2_0, output_1_279;
mixer gate_output_1_279(.a(output_2_279), .b(output_2_0), .y(output_1_279));
wire output_3_279, output_3_0, output_2_279;
mixer gate_output_2_279(.a(output_3_279), .b(output_3_0), .y(output_2_279));
wire output_4_279, output_4_0, output_3_279;
mixer gate_output_3_279(.a(output_4_279), .b(output_4_0), .y(output_3_279));
wire output_5_279, output_5_0, output_4_279;
mixer gate_output_4_279(.a(output_5_279), .b(output_5_0), .y(output_4_279));
wire output_6_279, output_6_0, output_5_279;
mixer gate_output_5_279(.a(output_6_279), .b(output_6_0), .y(output_5_279));
wire output_7_279, output_7_0, output_6_279;
mixer gate_output_6_279(.a(output_7_279), .b(output_7_0), .y(output_6_279));
wire output_8_279, output_8_0, output_7_279;
mixer gate_output_7_279(.a(output_8_279), .b(output_8_0), .y(output_7_279));
wire output_1_280, output_1_1, output_0_280;
mixer gate_output_0_280(.a(output_1_280), .b(output_1_1), .y(output_0_280));
wire output_2_280, output_2_1, output_1_280;
mixer gate_output_1_280(.a(output_2_280), .b(output_2_1), .y(output_1_280));
wire output_3_280, output_3_1, output_2_280;
mixer gate_output_2_280(.a(output_3_280), .b(output_3_1), .y(output_2_280));
wire output_4_280, output_4_1, output_3_280;
mixer gate_output_3_280(.a(output_4_280), .b(output_4_1), .y(output_3_280));
wire output_5_280, output_5_1, output_4_280;
mixer gate_output_4_280(.a(output_5_280), .b(output_5_1), .y(output_4_280));
wire output_6_280, output_6_1, output_5_280;
mixer gate_output_5_280(.a(output_6_280), .b(output_6_1), .y(output_5_280));
wire output_7_280, output_7_1, output_6_280;
mixer gate_output_6_280(.a(output_7_280), .b(output_7_1), .y(output_6_280));
wire output_8_280, output_8_1, output_7_280;
mixer gate_output_7_280(.a(output_8_280), .b(output_8_1), .y(output_7_280));
wire output_1_281, output_1_2, output_0_281;
mixer gate_output_0_281(.a(output_1_281), .b(output_1_2), .y(output_0_281));
wire output_2_281, output_2_2, output_1_281;
mixer gate_output_1_281(.a(output_2_281), .b(output_2_2), .y(output_1_281));
wire output_3_281, output_3_2, output_2_281;
mixer gate_output_2_281(.a(output_3_281), .b(output_3_2), .y(output_2_281));
wire output_4_281, output_4_2, output_3_281;
mixer gate_output_3_281(.a(output_4_281), .b(output_4_2), .y(output_3_281));
wire output_5_281, output_5_2, output_4_281;
mixer gate_output_4_281(.a(output_5_281), .b(output_5_2), .y(output_4_281));
wire output_6_281, output_6_2, output_5_281;
mixer gate_output_5_281(.a(output_6_281), .b(output_6_2), .y(output_5_281));
wire output_7_281, output_7_2, output_6_281;
mixer gate_output_6_281(.a(output_7_281), .b(output_7_2), .y(output_6_281));
wire output_8_281, output_8_2, output_7_281;
mixer gate_output_7_281(.a(output_8_281), .b(output_8_2), .y(output_7_281));
wire output_1_282, output_1_3, output_0_282;
mixer gate_output_0_282(.a(output_1_282), .b(output_1_3), .y(output_0_282));
wire output_2_282, output_2_3, output_1_282;
mixer gate_output_1_282(.a(output_2_282), .b(output_2_3), .y(output_1_282));
wire output_3_282, output_3_3, output_2_282;
mixer gate_output_2_282(.a(output_3_282), .b(output_3_3), .y(output_2_282));
wire output_4_282, output_4_3, output_3_282;
mixer gate_output_3_282(.a(output_4_282), .b(output_4_3), .y(output_3_282));
wire output_5_282, output_5_3, output_4_282;
mixer gate_output_4_282(.a(output_5_282), .b(output_5_3), .y(output_4_282));
wire output_6_282, output_6_3, output_5_282;
mixer gate_output_5_282(.a(output_6_282), .b(output_6_3), .y(output_5_282));
wire output_7_282, output_7_3, output_6_282;
mixer gate_output_6_282(.a(output_7_282), .b(output_7_3), .y(output_6_282));
wire output_8_282, output_8_3, output_7_282;
mixer gate_output_7_282(.a(output_8_282), .b(output_8_3), .y(output_7_282));
wire output_1_283, output_1_4, output_0_283;
mixer gate_output_0_283(.a(output_1_283), .b(output_1_4), .y(output_0_283));
wire output_2_283, output_2_4, output_1_283;
mixer gate_output_1_283(.a(output_2_283), .b(output_2_4), .y(output_1_283));
wire output_3_283, output_3_4, output_2_283;
mixer gate_output_2_283(.a(output_3_283), .b(output_3_4), .y(output_2_283));
wire output_4_283, output_4_4, output_3_283;
mixer gate_output_3_283(.a(output_4_283), .b(output_4_4), .y(output_3_283));
wire output_5_283, output_5_4, output_4_283;
mixer gate_output_4_283(.a(output_5_283), .b(output_5_4), .y(output_4_283));
wire output_6_283, output_6_4, output_5_283;
mixer gate_output_5_283(.a(output_6_283), .b(output_6_4), .y(output_5_283));
wire output_7_283, output_7_4, output_6_283;
mixer gate_output_6_283(.a(output_7_283), .b(output_7_4), .y(output_6_283));
wire output_8_283, output_8_4, output_7_283;
mixer gate_output_7_283(.a(output_8_283), .b(output_8_4), .y(output_7_283));
wire output_1_284, output_1_5, output_0_284;
mixer gate_output_0_284(.a(output_1_284), .b(output_1_5), .y(output_0_284));
wire output_2_284, output_2_5, output_1_284;
mixer gate_output_1_284(.a(output_2_284), .b(output_2_5), .y(output_1_284));
wire output_3_284, output_3_5, output_2_284;
mixer gate_output_2_284(.a(output_3_284), .b(output_3_5), .y(output_2_284));
wire output_4_284, output_4_5, output_3_284;
mixer gate_output_3_284(.a(output_4_284), .b(output_4_5), .y(output_3_284));
wire output_5_284, output_5_5, output_4_284;
mixer gate_output_4_284(.a(output_5_284), .b(output_5_5), .y(output_4_284));
wire output_6_284, output_6_5, output_5_284;
mixer gate_output_5_284(.a(output_6_284), .b(output_6_5), .y(output_5_284));
wire output_7_284, output_7_5, output_6_284;
mixer gate_output_6_284(.a(output_7_284), .b(output_7_5), .y(output_6_284));
wire output_8_284, output_8_5, output_7_284;
mixer gate_output_7_284(.a(output_8_284), .b(output_8_5), .y(output_7_284));
wire output_1_285, output_1_6, output_0_285;
mixer gate_output_0_285(.a(output_1_285), .b(output_1_6), .y(output_0_285));
wire output_2_285, output_2_6, output_1_285;
mixer gate_output_1_285(.a(output_2_285), .b(output_2_6), .y(output_1_285));
wire output_3_285, output_3_6, output_2_285;
mixer gate_output_2_285(.a(output_3_285), .b(output_3_6), .y(output_2_285));
wire output_4_285, output_4_6, output_3_285;
mixer gate_output_3_285(.a(output_4_285), .b(output_4_6), .y(output_3_285));
wire output_5_285, output_5_6, output_4_285;
mixer gate_output_4_285(.a(output_5_285), .b(output_5_6), .y(output_4_285));
wire output_6_285, output_6_6, output_5_285;
mixer gate_output_5_285(.a(output_6_285), .b(output_6_6), .y(output_5_285));
wire output_7_285, output_7_6, output_6_285;
mixer gate_output_6_285(.a(output_7_285), .b(output_7_6), .y(output_6_285));
wire output_8_285, output_8_6, output_7_285;
mixer gate_output_7_285(.a(output_8_285), .b(output_8_6), .y(output_7_285));
wire output_1_286, output_1_7, output_0_286;
mixer gate_output_0_286(.a(output_1_286), .b(output_1_7), .y(output_0_286));
wire output_2_286, output_2_7, output_1_286;
mixer gate_output_1_286(.a(output_2_286), .b(output_2_7), .y(output_1_286));
wire output_3_286, output_3_7, output_2_286;
mixer gate_output_2_286(.a(output_3_286), .b(output_3_7), .y(output_2_286));
wire output_4_286, output_4_7, output_3_286;
mixer gate_output_3_286(.a(output_4_286), .b(output_4_7), .y(output_3_286));
wire output_5_286, output_5_7, output_4_286;
mixer gate_output_4_286(.a(output_5_286), .b(output_5_7), .y(output_4_286));
wire output_6_286, output_6_7, output_5_286;
mixer gate_output_5_286(.a(output_6_286), .b(output_6_7), .y(output_5_286));
wire output_7_286, output_7_7, output_6_286;
mixer gate_output_6_286(.a(output_7_286), .b(output_7_7), .y(output_6_286));
wire output_8_286, output_8_7, output_7_286;
mixer gate_output_7_286(.a(output_8_286), .b(output_8_7), .y(output_7_286));
wire output_1_287, output_1_0, output_0_287;
mixer gate_output_0_287(.a(output_1_287), .b(output_1_0), .y(output_0_287));
wire output_2_287, output_2_0, output_1_287;
mixer gate_output_1_287(.a(output_2_287), .b(output_2_0), .y(output_1_287));
wire output_3_287, output_3_0, output_2_287;
mixer gate_output_2_287(.a(output_3_287), .b(output_3_0), .y(output_2_287));
wire output_4_287, output_4_0, output_3_287;
mixer gate_output_3_287(.a(output_4_287), .b(output_4_0), .y(output_3_287));
wire output_5_287, output_5_0, output_4_287;
mixer gate_output_4_287(.a(output_5_287), .b(output_5_0), .y(output_4_287));
wire output_6_287, output_6_0, output_5_287;
mixer gate_output_5_287(.a(output_6_287), .b(output_6_0), .y(output_5_287));
wire output_7_287, output_7_0, output_6_287;
mixer gate_output_6_287(.a(output_7_287), .b(output_7_0), .y(output_6_287));
wire output_8_287, output_8_0, output_7_287;
mixer gate_output_7_287(.a(output_8_287), .b(output_8_0), .y(output_7_287));
wire output_1_288, output_1_1, output_0_288;
mixer gate_output_0_288(.a(output_1_288), .b(output_1_1), .y(output_0_288));
wire output_2_288, output_2_1, output_1_288;
mixer gate_output_1_288(.a(output_2_288), .b(output_2_1), .y(output_1_288));
wire output_3_288, output_3_1, output_2_288;
mixer gate_output_2_288(.a(output_3_288), .b(output_3_1), .y(output_2_288));
wire output_4_288, output_4_1, output_3_288;
mixer gate_output_3_288(.a(output_4_288), .b(output_4_1), .y(output_3_288));
wire output_5_288, output_5_1, output_4_288;
mixer gate_output_4_288(.a(output_5_288), .b(output_5_1), .y(output_4_288));
wire output_6_288, output_6_1, output_5_288;
mixer gate_output_5_288(.a(output_6_288), .b(output_6_1), .y(output_5_288));
wire output_7_288, output_7_1, output_6_288;
mixer gate_output_6_288(.a(output_7_288), .b(output_7_1), .y(output_6_288));
wire output_8_288, output_8_1, output_7_288;
mixer gate_output_7_288(.a(output_8_288), .b(output_8_1), .y(output_7_288));
wire output_1_289, output_1_2, output_0_289;
mixer gate_output_0_289(.a(output_1_289), .b(output_1_2), .y(output_0_289));
wire output_2_289, output_2_2, output_1_289;
mixer gate_output_1_289(.a(output_2_289), .b(output_2_2), .y(output_1_289));
wire output_3_289, output_3_2, output_2_289;
mixer gate_output_2_289(.a(output_3_289), .b(output_3_2), .y(output_2_289));
wire output_4_289, output_4_2, output_3_289;
mixer gate_output_3_289(.a(output_4_289), .b(output_4_2), .y(output_3_289));
wire output_5_289, output_5_2, output_4_289;
mixer gate_output_4_289(.a(output_5_289), .b(output_5_2), .y(output_4_289));
wire output_6_289, output_6_2, output_5_289;
mixer gate_output_5_289(.a(output_6_289), .b(output_6_2), .y(output_5_289));
wire output_7_289, output_7_2, output_6_289;
mixer gate_output_6_289(.a(output_7_289), .b(output_7_2), .y(output_6_289));
wire output_8_289, output_8_2, output_7_289;
mixer gate_output_7_289(.a(output_8_289), .b(output_8_2), .y(output_7_289));
wire output_1_290, output_1_3, output_0_290;
mixer gate_output_0_290(.a(output_1_290), .b(output_1_3), .y(output_0_290));
wire output_2_290, output_2_3, output_1_290;
mixer gate_output_1_290(.a(output_2_290), .b(output_2_3), .y(output_1_290));
wire output_3_290, output_3_3, output_2_290;
mixer gate_output_2_290(.a(output_3_290), .b(output_3_3), .y(output_2_290));
wire output_4_290, output_4_3, output_3_290;
mixer gate_output_3_290(.a(output_4_290), .b(output_4_3), .y(output_3_290));
wire output_5_290, output_5_3, output_4_290;
mixer gate_output_4_290(.a(output_5_290), .b(output_5_3), .y(output_4_290));
wire output_6_290, output_6_3, output_5_290;
mixer gate_output_5_290(.a(output_6_290), .b(output_6_3), .y(output_5_290));
wire output_7_290, output_7_3, output_6_290;
mixer gate_output_6_290(.a(output_7_290), .b(output_7_3), .y(output_6_290));
wire output_8_290, output_8_3, output_7_290;
mixer gate_output_7_290(.a(output_8_290), .b(output_8_3), .y(output_7_290));
wire output_1_291, output_1_4, output_0_291;
mixer gate_output_0_291(.a(output_1_291), .b(output_1_4), .y(output_0_291));
wire output_2_291, output_2_4, output_1_291;
mixer gate_output_1_291(.a(output_2_291), .b(output_2_4), .y(output_1_291));
wire output_3_291, output_3_4, output_2_291;
mixer gate_output_2_291(.a(output_3_291), .b(output_3_4), .y(output_2_291));
wire output_4_291, output_4_4, output_3_291;
mixer gate_output_3_291(.a(output_4_291), .b(output_4_4), .y(output_3_291));
wire output_5_291, output_5_4, output_4_291;
mixer gate_output_4_291(.a(output_5_291), .b(output_5_4), .y(output_4_291));
wire output_6_291, output_6_4, output_5_291;
mixer gate_output_5_291(.a(output_6_291), .b(output_6_4), .y(output_5_291));
wire output_7_291, output_7_4, output_6_291;
mixer gate_output_6_291(.a(output_7_291), .b(output_7_4), .y(output_6_291));
wire output_8_291, output_8_4, output_7_291;
mixer gate_output_7_291(.a(output_8_291), .b(output_8_4), .y(output_7_291));
wire output_1_292, output_1_5, output_0_292;
mixer gate_output_0_292(.a(output_1_292), .b(output_1_5), .y(output_0_292));
wire output_2_292, output_2_5, output_1_292;
mixer gate_output_1_292(.a(output_2_292), .b(output_2_5), .y(output_1_292));
wire output_3_292, output_3_5, output_2_292;
mixer gate_output_2_292(.a(output_3_292), .b(output_3_5), .y(output_2_292));
wire output_4_292, output_4_5, output_3_292;
mixer gate_output_3_292(.a(output_4_292), .b(output_4_5), .y(output_3_292));
wire output_5_292, output_5_5, output_4_292;
mixer gate_output_4_292(.a(output_5_292), .b(output_5_5), .y(output_4_292));
wire output_6_292, output_6_5, output_5_292;
mixer gate_output_5_292(.a(output_6_292), .b(output_6_5), .y(output_5_292));
wire output_7_292, output_7_5, output_6_292;
mixer gate_output_6_292(.a(output_7_292), .b(output_7_5), .y(output_6_292));
wire output_8_292, output_8_5, output_7_292;
mixer gate_output_7_292(.a(output_8_292), .b(output_8_5), .y(output_7_292));
wire output_1_293, output_1_6, output_0_293;
mixer gate_output_0_293(.a(output_1_293), .b(output_1_6), .y(output_0_293));
wire output_2_293, output_2_6, output_1_293;
mixer gate_output_1_293(.a(output_2_293), .b(output_2_6), .y(output_1_293));
wire output_3_293, output_3_6, output_2_293;
mixer gate_output_2_293(.a(output_3_293), .b(output_3_6), .y(output_2_293));
wire output_4_293, output_4_6, output_3_293;
mixer gate_output_3_293(.a(output_4_293), .b(output_4_6), .y(output_3_293));
wire output_5_293, output_5_6, output_4_293;
mixer gate_output_4_293(.a(output_5_293), .b(output_5_6), .y(output_4_293));
wire output_6_293, output_6_6, output_5_293;
mixer gate_output_5_293(.a(output_6_293), .b(output_6_6), .y(output_5_293));
wire output_7_293, output_7_6, output_6_293;
mixer gate_output_6_293(.a(output_7_293), .b(output_7_6), .y(output_6_293));
wire output_8_293, output_8_6, output_7_293;
mixer gate_output_7_293(.a(output_8_293), .b(output_8_6), .y(output_7_293));
wire output_1_294, output_1_7, output_0_294;
mixer gate_output_0_294(.a(output_1_294), .b(output_1_7), .y(output_0_294));
wire output_2_294, output_2_7, output_1_294;
mixer gate_output_1_294(.a(output_2_294), .b(output_2_7), .y(output_1_294));
wire output_3_294, output_3_7, output_2_294;
mixer gate_output_2_294(.a(output_3_294), .b(output_3_7), .y(output_2_294));
wire output_4_294, output_4_7, output_3_294;
mixer gate_output_3_294(.a(output_4_294), .b(output_4_7), .y(output_3_294));
wire output_5_294, output_5_7, output_4_294;
mixer gate_output_4_294(.a(output_5_294), .b(output_5_7), .y(output_4_294));
wire output_6_294, output_6_7, output_5_294;
mixer gate_output_5_294(.a(output_6_294), .b(output_6_7), .y(output_5_294));
wire output_7_294, output_7_7, output_6_294;
mixer gate_output_6_294(.a(output_7_294), .b(output_7_7), .y(output_6_294));
wire output_8_294, output_8_7, output_7_294;
mixer gate_output_7_294(.a(output_8_294), .b(output_8_7), .y(output_7_294));
wire output_1_295, output_1_0, output_0_295;
mixer gate_output_0_295(.a(output_1_295), .b(output_1_0), .y(output_0_295));
wire output_2_295, output_2_0, output_1_295;
mixer gate_output_1_295(.a(output_2_295), .b(output_2_0), .y(output_1_295));
wire output_3_295, output_3_0, output_2_295;
mixer gate_output_2_295(.a(output_3_295), .b(output_3_0), .y(output_2_295));
wire output_4_295, output_4_0, output_3_295;
mixer gate_output_3_295(.a(output_4_295), .b(output_4_0), .y(output_3_295));
wire output_5_295, output_5_0, output_4_295;
mixer gate_output_4_295(.a(output_5_295), .b(output_5_0), .y(output_4_295));
wire output_6_295, output_6_0, output_5_295;
mixer gate_output_5_295(.a(output_6_295), .b(output_6_0), .y(output_5_295));
wire output_7_295, output_7_0, output_6_295;
mixer gate_output_6_295(.a(output_7_295), .b(output_7_0), .y(output_6_295));
wire output_8_295, output_8_0, output_7_295;
mixer gate_output_7_295(.a(output_8_295), .b(output_8_0), .y(output_7_295));
wire output_1_296, output_1_1, output_0_296;
mixer gate_output_0_296(.a(output_1_296), .b(output_1_1), .y(output_0_296));
wire output_2_296, output_2_1, output_1_296;
mixer gate_output_1_296(.a(output_2_296), .b(output_2_1), .y(output_1_296));
wire output_3_296, output_3_1, output_2_296;
mixer gate_output_2_296(.a(output_3_296), .b(output_3_1), .y(output_2_296));
wire output_4_296, output_4_1, output_3_296;
mixer gate_output_3_296(.a(output_4_296), .b(output_4_1), .y(output_3_296));
wire output_5_296, output_5_1, output_4_296;
mixer gate_output_4_296(.a(output_5_296), .b(output_5_1), .y(output_4_296));
wire output_6_296, output_6_1, output_5_296;
mixer gate_output_5_296(.a(output_6_296), .b(output_6_1), .y(output_5_296));
wire output_7_296, output_7_1, output_6_296;
mixer gate_output_6_296(.a(output_7_296), .b(output_7_1), .y(output_6_296));
wire output_8_296, output_8_1, output_7_296;
mixer gate_output_7_296(.a(output_8_296), .b(output_8_1), .y(output_7_296));
wire output_1_297, output_1_2, output_0_297;
mixer gate_output_0_297(.a(output_1_297), .b(output_1_2), .y(output_0_297));
wire output_2_297, output_2_2, output_1_297;
mixer gate_output_1_297(.a(output_2_297), .b(output_2_2), .y(output_1_297));
wire output_3_297, output_3_2, output_2_297;
mixer gate_output_2_297(.a(output_3_297), .b(output_3_2), .y(output_2_297));
wire output_4_297, output_4_2, output_3_297;
mixer gate_output_3_297(.a(output_4_297), .b(output_4_2), .y(output_3_297));
wire output_5_297, output_5_2, output_4_297;
mixer gate_output_4_297(.a(output_5_297), .b(output_5_2), .y(output_4_297));
wire output_6_297, output_6_2, output_5_297;
mixer gate_output_5_297(.a(output_6_297), .b(output_6_2), .y(output_5_297));
wire output_7_297, output_7_2, output_6_297;
mixer gate_output_6_297(.a(output_7_297), .b(output_7_2), .y(output_6_297));
wire output_8_297, output_8_2, output_7_297;
mixer gate_output_7_297(.a(output_8_297), .b(output_8_2), .y(output_7_297));
wire output_1_298, output_1_3, output_0_298;
mixer gate_output_0_298(.a(output_1_298), .b(output_1_3), .y(output_0_298));
wire output_2_298, output_2_3, output_1_298;
mixer gate_output_1_298(.a(output_2_298), .b(output_2_3), .y(output_1_298));
wire output_3_298, output_3_3, output_2_298;
mixer gate_output_2_298(.a(output_3_298), .b(output_3_3), .y(output_2_298));
wire output_4_298, output_4_3, output_3_298;
mixer gate_output_3_298(.a(output_4_298), .b(output_4_3), .y(output_3_298));
wire output_5_298, output_5_3, output_4_298;
mixer gate_output_4_298(.a(output_5_298), .b(output_5_3), .y(output_4_298));
wire output_6_298, output_6_3, output_5_298;
mixer gate_output_5_298(.a(output_6_298), .b(output_6_3), .y(output_5_298));
wire output_7_298, output_7_3, output_6_298;
mixer gate_output_6_298(.a(output_7_298), .b(output_7_3), .y(output_6_298));
wire output_8_298, output_8_3, output_7_298;
mixer gate_output_7_298(.a(output_8_298), .b(output_8_3), .y(output_7_298));
wire output_1_299, output_1_4, output_0_299;
mixer gate_output_0_299(.a(output_1_299), .b(output_1_4), .y(output_0_299));
wire output_2_299, output_2_4, output_1_299;
mixer gate_output_1_299(.a(output_2_299), .b(output_2_4), .y(output_1_299));
wire output_3_299, output_3_4, output_2_299;
mixer gate_output_2_299(.a(output_3_299), .b(output_3_4), .y(output_2_299));
wire output_4_299, output_4_4, output_3_299;
mixer gate_output_3_299(.a(output_4_299), .b(output_4_4), .y(output_3_299));
wire output_5_299, output_5_4, output_4_299;
mixer gate_output_4_299(.a(output_5_299), .b(output_5_4), .y(output_4_299));
wire output_6_299, output_6_4, output_5_299;
mixer gate_output_5_299(.a(output_6_299), .b(output_6_4), .y(output_5_299));
wire output_7_299, output_7_4, output_6_299;
mixer gate_output_6_299(.a(output_7_299), .b(output_7_4), .y(output_6_299));
wire output_8_299, output_8_4, output_7_299;
mixer gate_output_7_299(.a(output_8_299), .b(output_8_4), .y(output_7_299));
wire output_1_300, output_1_5, output_0_300;
mixer gate_output_0_300(.a(output_1_300), .b(output_1_5), .y(output_0_300));
wire output_2_300, output_2_5, output_1_300;
mixer gate_output_1_300(.a(output_2_300), .b(output_2_5), .y(output_1_300));
wire output_3_300, output_3_5, output_2_300;
mixer gate_output_2_300(.a(output_3_300), .b(output_3_5), .y(output_2_300));
wire output_4_300, output_4_5, output_3_300;
mixer gate_output_3_300(.a(output_4_300), .b(output_4_5), .y(output_3_300));
wire output_5_300, output_5_5, output_4_300;
mixer gate_output_4_300(.a(output_5_300), .b(output_5_5), .y(output_4_300));
wire output_6_300, output_6_5, output_5_300;
mixer gate_output_5_300(.a(output_6_300), .b(output_6_5), .y(output_5_300));
wire output_7_300, output_7_5, output_6_300;
mixer gate_output_6_300(.a(output_7_300), .b(output_7_5), .y(output_6_300));
wire output_8_300, output_8_5, output_7_300;
mixer gate_output_7_300(.a(output_8_300), .b(output_8_5), .y(output_7_300));
wire output_1_301, output_1_6, output_0_301;
mixer gate_output_0_301(.a(output_1_301), .b(output_1_6), .y(output_0_301));
wire output_2_301, output_2_6, output_1_301;
mixer gate_output_1_301(.a(output_2_301), .b(output_2_6), .y(output_1_301));
wire output_3_301, output_3_6, output_2_301;
mixer gate_output_2_301(.a(output_3_301), .b(output_3_6), .y(output_2_301));
wire output_4_301, output_4_6, output_3_301;
mixer gate_output_3_301(.a(output_4_301), .b(output_4_6), .y(output_3_301));
wire output_5_301, output_5_6, output_4_301;
mixer gate_output_4_301(.a(output_5_301), .b(output_5_6), .y(output_4_301));
wire output_6_301, output_6_6, output_5_301;
mixer gate_output_5_301(.a(output_6_301), .b(output_6_6), .y(output_5_301));
wire output_7_301, output_7_6, output_6_301;
mixer gate_output_6_301(.a(output_7_301), .b(output_7_6), .y(output_6_301));
wire output_8_301, output_8_6, output_7_301;
mixer gate_output_7_301(.a(output_8_301), .b(output_8_6), .y(output_7_301));
wire output_1_302, output_1_7, output_0_302;
mixer gate_output_0_302(.a(output_1_302), .b(output_1_7), .y(output_0_302));
wire output_2_302, output_2_7, output_1_302;
mixer gate_output_1_302(.a(output_2_302), .b(output_2_7), .y(output_1_302));
wire output_3_302, output_3_7, output_2_302;
mixer gate_output_2_302(.a(output_3_302), .b(output_3_7), .y(output_2_302));
wire output_4_302, output_4_7, output_3_302;
mixer gate_output_3_302(.a(output_4_302), .b(output_4_7), .y(output_3_302));
wire output_5_302, output_5_7, output_4_302;
mixer gate_output_4_302(.a(output_5_302), .b(output_5_7), .y(output_4_302));
wire output_6_302, output_6_7, output_5_302;
mixer gate_output_5_302(.a(output_6_302), .b(output_6_7), .y(output_5_302));
wire output_7_302, output_7_7, output_6_302;
mixer gate_output_6_302(.a(output_7_302), .b(output_7_7), .y(output_6_302));
wire output_8_302, output_8_7, output_7_302;
mixer gate_output_7_302(.a(output_8_302), .b(output_8_7), .y(output_7_302));
wire output_1_303, output_1_0, output_0_303;
mixer gate_output_0_303(.a(output_1_303), .b(output_1_0), .y(output_0_303));
wire output_2_303, output_2_0, output_1_303;
mixer gate_output_1_303(.a(output_2_303), .b(output_2_0), .y(output_1_303));
wire output_3_303, output_3_0, output_2_303;
mixer gate_output_2_303(.a(output_3_303), .b(output_3_0), .y(output_2_303));
wire output_4_303, output_4_0, output_3_303;
mixer gate_output_3_303(.a(output_4_303), .b(output_4_0), .y(output_3_303));
wire output_5_303, output_5_0, output_4_303;
mixer gate_output_4_303(.a(output_5_303), .b(output_5_0), .y(output_4_303));
wire output_6_303, output_6_0, output_5_303;
mixer gate_output_5_303(.a(output_6_303), .b(output_6_0), .y(output_5_303));
wire output_7_303, output_7_0, output_6_303;
mixer gate_output_6_303(.a(output_7_303), .b(output_7_0), .y(output_6_303));
wire output_8_303, output_8_0, output_7_303;
mixer gate_output_7_303(.a(output_8_303), .b(output_8_0), .y(output_7_303));
wire output_1_304, output_1_1, output_0_304;
mixer gate_output_0_304(.a(output_1_304), .b(output_1_1), .y(output_0_304));
wire output_2_304, output_2_1, output_1_304;
mixer gate_output_1_304(.a(output_2_304), .b(output_2_1), .y(output_1_304));
wire output_3_304, output_3_1, output_2_304;
mixer gate_output_2_304(.a(output_3_304), .b(output_3_1), .y(output_2_304));
wire output_4_304, output_4_1, output_3_304;
mixer gate_output_3_304(.a(output_4_304), .b(output_4_1), .y(output_3_304));
wire output_5_304, output_5_1, output_4_304;
mixer gate_output_4_304(.a(output_5_304), .b(output_5_1), .y(output_4_304));
wire output_6_304, output_6_1, output_5_304;
mixer gate_output_5_304(.a(output_6_304), .b(output_6_1), .y(output_5_304));
wire output_7_304, output_7_1, output_6_304;
mixer gate_output_6_304(.a(output_7_304), .b(output_7_1), .y(output_6_304));
wire output_8_304, output_8_1, output_7_304;
mixer gate_output_7_304(.a(output_8_304), .b(output_8_1), .y(output_7_304));
wire output_1_305, output_1_2, output_0_305;
mixer gate_output_0_305(.a(output_1_305), .b(output_1_2), .y(output_0_305));
wire output_2_305, output_2_2, output_1_305;
mixer gate_output_1_305(.a(output_2_305), .b(output_2_2), .y(output_1_305));
wire output_3_305, output_3_2, output_2_305;
mixer gate_output_2_305(.a(output_3_305), .b(output_3_2), .y(output_2_305));
wire output_4_305, output_4_2, output_3_305;
mixer gate_output_3_305(.a(output_4_305), .b(output_4_2), .y(output_3_305));
wire output_5_305, output_5_2, output_4_305;
mixer gate_output_4_305(.a(output_5_305), .b(output_5_2), .y(output_4_305));
wire output_6_305, output_6_2, output_5_305;
mixer gate_output_5_305(.a(output_6_305), .b(output_6_2), .y(output_5_305));
wire output_7_305, output_7_2, output_6_305;
mixer gate_output_6_305(.a(output_7_305), .b(output_7_2), .y(output_6_305));
wire output_8_305, output_8_2, output_7_305;
mixer gate_output_7_305(.a(output_8_305), .b(output_8_2), .y(output_7_305));
wire output_1_306, output_1_3, output_0_306;
mixer gate_output_0_306(.a(output_1_306), .b(output_1_3), .y(output_0_306));
wire output_2_306, output_2_3, output_1_306;
mixer gate_output_1_306(.a(output_2_306), .b(output_2_3), .y(output_1_306));
wire output_3_306, output_3_3, output_2_306;
mixer gate_output_2_306(.a(output_3_306), .b(output_3_3), .y(output_2_306));
wire output_4_306, output_4_3, output_3_306;
mixer gate_output_3_306(.a(output_4_306), .b(output_4_3), .y(output_3_306));
wire output_5_306, output_5_3, output_4_306;
mixer gate_output_4_306(.a(output_5_306), .b(output_5_3), .y(output_4_306));
wire output_6_306, output_6_3, output_5_306;
mixer gate_output_5_306(.a(output_6_306), .b(output_6_3), .y(output_5_306));
wire output_7_306, output_7_3, output_6_306;
mixer gate_output_6_306(.a(output_7_306), .b(output_7_3), .y(output_6_306));
wire output_8_306, output_8_3, output_7_306;
mixer gate_output_7_306(.a(output_8_306), .b(output_8_3), .y(output_7_306));
wire output_1_307, output_1_4, output_0_307;
mixer gate_output_0_307(.a(output_1_307), .b(output_1_4), .y(output_0_307));
wire output_2_307, output_2_4, output_1_307;
mixer gate_output_1_307(.a(output_2_307), .b(output_2_4), .y(output_1_307));
wire output_3_307, output_3_4, output_2_307;
mixer gate_output_2_307(.a(output_3_307), .b(output_3_4), .y(output_2_307));
wire output_4_307, output_4_4, output_3_307;
mixer gate_output_3_307(.a(output_4_307), .b(output_4_4), .y(output_3_307));
wire output_5_307, output_5_4, output_4_307;
mixer gate_output_4_307(.a(output_5_307), .b(output_5_4), .y(output_4_307));
wire output_6_307, output_6_4, output_5_307;
mixer gate_output_5_307(.a(output_6_307), .b(output_6_4), .y(output_5_307));
wire output_7_307, output_7_4, output_6_307;
mixer gate_output_6_307(.a(output_7_307), .b(output_7_4), .y(output_6_307));
wire output_8_307, output_8_4, output_7_307;
mixer gate_output_7_307(.a(output_8_307), .b(output_8_4), .y(output_7_307));
wire output_1_308, output_1_5, output_0_308;
mixer gate_output_0_308(.a(output_1_308), .b(output_1_5), .y(output_0_308));
wire output_2_308, output_2_5, output_1_308;
mixer gate_output_1_308(.a(output_2_308), .b(output_2_5), .y(output_1_308));
wire output_3_308, output_3_5, output_2_308;
mixer gate_output_2_308(.a(output_3_308), .b(output_3_5), .y(output_2_308));
wire output_4_308, output_4_5, output_3_308;
mixer gate_output_3_308(.a(output_4_308), .b(output_4_5), .y(output_3_308));
wire output_5_308, output_5_5, output_4_308;
mixer gate_output_4_308(.a(output_5_308), .b(output_5_5), .y(output_4_308));
wire output_6_308, output_6_5, output_5_308;
mixer gate_output_5_308(.a(output_6_308), .b(output_6_5), .y(output_5_308));
wire output_7_308, output_7_5, output_6_308;
mixer gate_output_6_308(.a(output_7_308), .b(output_7_5), .y(output_6_308));
wire output_8_308, output_8_5, output_7_308;
mixer gate_output_7_308(.a(output_8_308), .b(output_8_5), .y(output_7_308));
wire output_1_309, output_1_6, output_0_309;
mixer gate_output_0_309(.a(output_1_309), .b(output_1_6), .y(output_0_309));
wire output_2_309, output_2_6, output_1_309;
mixer gate_output_1_309(.a(output_2_309), .b(output_2_6), .y(output_1_309));
wire output_3_309, output_3_6, output_2_309;
mixer gate_output_2_309(.a(output_3_309), .b(output_3_6), .y(output_2_309));
wire output_4_309, output_4_6, output_3_309;
mixer gate_output_3_309(.a(output_4_309), .b(output_4_6), .y(output_3_309));
wire output_5_309, output_5_6, output_4_309;
mixer gate_output_4_309(.a(output_5_309), .b(output_5_6), .y(output_4_309));
wire output_6_309, output_6_6, output_5_309;
mixer gate_output_5_309(.a(output_6_309), .b(output_6_6), .y(output_5_309));
wire output_7_309, output_7_6, output_6_309;
mixer gate_output_6_309(.a(output_7_309), .b(output_7_6), .y(output_6_309));
wire output_8_309, output_8_6, output_7_309;
mixer gate_output_7_309(.a(output_8_309), .b(output_8_6), .y(output_7_309));
wire output_1_310, output_1_7, output_0_310;
mixer gate_output_0_310(.a(output_1_310), .b(output_1_7), .y(output_0_310));
wire output_2_310, output_2_7, output_1_310;
mixer gate_output_1_310(.a(output_2_310), .b(output_2_7), .y(output_1_310));
wire output_3_310, output_3_7, output_2_310;
mixer gate_output_2_310(.a(output_3_310), .b(output_3_7), .y(output_2_310));
wire output_4_310, output_4_7, output_3_310;
mixer gate_output_3_310(.a(output_4_310), .b(output_4_7), .y(output_3_310));
wire output_5_310, output_5_7, output_4_310;
mixer gate_output_4_310(.a(output_5_310), .b(output_5_7), .y(output_4_310));
wire output_6_310, output_6_7, output_5_310;
mixer gate_output_5_310(.a(output_6_310), .b(output_6_7), .y(output_5_310));
wire output_7_310, output_7_7, output_6_310;
mixer gate_output_6_310(.a(output_7_310), .b(output_7_7), .y(output_6_310));
wire output_8_310, output_8_7, output_7_310;
mixer gate_output_7_310(.a(output_8_310), .b(output_8_7), .y(output_7_310));
wire output_1_311, output_1_0, output_0_311;
mixer gate_output_0_311(.a(output_1_311), .b(output_1_0), .y(output_0_311));
wire output_2_311, output_2_0, output_1_311;
mixer gate_output_1_311(.a(output_2_311), .b(output_2_0), .y(output_1_311));
wire output_3_311, output_3_0, output_2_311;
mixer gate_output_2_311(.a(output_3_311), .b(output_3_0), .y(output_2_311));
wire output_4_311, output_4_0, output_3_311;
mixer gate_output_3_311(.a(output_4_311), .b(output_4_0), .y(output_3_311));
wire output_5_311, output_5_0, output_4_311;
mixer gate_output_4_311(.a(output_5_311), .b(output_5_0), .y(output_4_311));
wire output_6_311, output_6_0, output_5_311;
mixer gate_output_5_311(.a(output_6_311), .b(output_6_0), .y(output_5_311));
wire output_7_311, output_7_0, output_6_311;
mixer gate_output_6_311(.a(output_7_311), .b(output_7_0), .y(output_6_311));
wire output_8_311, output_8_0, output_7_311;
mixer gate_output_7_311(.a(output_8_311), .b(output_8_0), .y(output_7_311));
wire output_1_312, output_1_1, output_0_312;
mixer gate_output_0_312(.a(output_1_312), .b(output_1_1), .y(output_0_312));
wire output_2_312, output_2_1, output_1_312;
mixer gate_output_1_312(.a(output_2_312), .b(output_2_1), .y(output_1_312));
wire output_3_312, output_3_1, output_2_312;
mixer gate_output_2_312(.a(output_3_312), .b(output_3_1), .y(output_2_312));
wire output_4_312, output_4_1, output_3_312;
mixer gate_output_3_312(.a(output_4_312), .b(output_4_1), .y(output_3_312));
wire output_5_312, output_5_1, output_4_312;
mixer gate_output_4_312(.a(output_5_312), .b(output_5_1), .y(output_4_312));
wire output_6_312, output_6_1, output_5_312;
mixer gate_output_5_312(.a(output_6_312), .b(output_6_1), .y(output_5_312));
wire output_7_312, output_7_1, output_6_312;
mixer gate_output_6_312(.a(output_7_312), .b(output_7_1), .y(output_6_312));
wire output_8_312, output_8_1, output_7_312;
mixer gate_output_7_312(.a(output_8_312), .b(output_8_1), .y(output_7_312));
wire output_1_313, output_1_2, output_0_313;
mixer gate_output_0_313(.a(output_1_313), .b(output_1_2), .y(output_0_313));
wire output_2_313, output_2_2, output_1_313;
mixer gate_output_1_313(.a(output_2_313), .b(output_2_2), .y(output_1_313));
wire output_3_313, output_3_2, output_2_313;
mixer gate_output_2_313(.a(output_3_313), .b(output_3_2), .y(output_2_313));
wire output_4_313, output_4_2, output_3_313;
mixer gate_output_3_313(.a(output_4_313), .b(output_4_2), .y(output_3_313));
wire output_5_313, output_5_2, output_4_313;
mixer gate_output_4_313(.a(output_5_313), .b(output_5_2), .y(output_4_313));
wire output_6_313, output_6_2, output_5_313;
mixer gate_output_5_313(.a(output_6_313), .b(output_6_2), .y(output_5_313));
wire output_7_313, output_7_2, output_6_313;
mixer gate_output_6_313(.a(output_7_313), .b(output_7_2), .y(output_6_313));
wire output_8_313, output_8_2, output_7_313;
mixer gate_output_7_313(.a(output_8_313), .b(output_8_2), .y(output_7_313));
wire output_1_314, output_1_3, output_0_314;
mixer gate_output_0_314(.a(output_1_314), .b(output_1_3), .y(output_0_314));
wire output_2_314, output_2_3, output_1_314;
mixer gate_output_1_314(.a(output_2_314), .b(output_2_3), .y(output_1_314));
wire output_3_314, output_3_3, output_2_314;
mixer gate_output_2_314(.a(output_3_314), .b(output_3_3), .y(output_2_314));
wire output_4_314, output_4_3, output_3_314;
mixer gate_output_3_314(.a(output_4_314), .b(output_4_3), .y(output_3_314));
wire output_5_314, output_5_3, output_4_314;
mixer gate_output_4_314(.a(output_5_314), .b(output_5_3), .y(output_4_314));
wire output_6_314, output_6_3, output_5_314;
mixer gate_output_5_314(.a(output_6_314), .b(output_6_3), .y(output_5_314));
wire output_7_314, output_7_3, output_6_314;
mixer gate_output_6_314(.a(output_7_314), .b(output_7_3), .y(output_6_314));
wire output_8_314, output_8_3, output_7_314;
mixer gate_output_7_314(.a(output_8_314), .b(output_8_3), .y(output_7_314));
wire output_1_315, output_1_4, output_0_315;
mixer gate_output_0_315(.a(output_1_315), .b(output_1_4), .y(output_0_315));
wire output_2_315, output_2_4, output_1_315;
mixer gate_output_1_315(.a(output_2_315), .b(output_2_4), .y(output_1_315));
wire output_3_315, output_3_4, output_2_315;
mixer gate_output_2_315(.a(output_3_315), .b(output_3_4), .y(output_2_315));
wire output_4_315, output_4_4, output_3_315;
mixer gate_output_3_315(.a(output_4_315), .b(output_4_4), .y(output_3_315));
wire output_5_315, output_5_4, output_4_315;
mixer gate_output_4_315(.a(output_5_315), .b(output_5_4), .y(output_4_315));
wire output_6_315, output_6_4, output_5_315;
mixer gate_output_5_315(.a(output_6_315), .b(output_6_4), .y(output_5_315));
wire output_7_315, output_7_4, output_6_315;
mixer gate_output_6_315(.a(output_7_315), .b(output_7_4), .y(output_6_315));
wire output_8_315, output_8_4, output_7_315;
mixer gate_output_7_315(.a(output_8_315), .b(output_8_4), .y(output_7_315));
wire output_1_316, output_1_5, output_0_316;
mixer gate_output_0_316(.a(output_1_316), .b(output_1_5), .y(output_0_316));
wire output_2_316, output_2_5, output_1_316;
mixer gate_output_1_316(.a(output_2_316), .b(output_2_5), .y(output_1_316));
wire output_3_316, output_3_5, output_2_316;
mixer gate_output_2_316(.a(output_3_316), .b(output_3_5), .y(output_2_316));
wire output_4_316, output_4_5, output_3_316;
mixer gate_output_3_316(.a(output_4_316), .b(output_4_5), .y(output_3_316));
wire output_5_316, output_5_5, output_4_316;
mixer gate_output_4_316(.a(output_5_316), .b(output_5_5), .y(output_4_316));
wire output_6_316, output_6_5, output_5_316;
mixer gate_output_5_316(.a(output_6_316), .b(output_6_5), .y(output_5_316));
wire output_7_316, output_7_5, output_6_316;
mixer gate_output_6_316(.a(output_7_316), .b(output_7_5), .y(output_6_316));
wire output_8_316, output_8_5, output_7_316;
mixer gate_output_7_316(.a(output_8_316), .b(output_8_5), .y(output_7_316));
wire output_1_317, output_1_6, output_0_317;
mixer gate_output_0_317(.a(output_1_317), .b(output_1_6), .y(output_0_317));
wire output_2_317, output_2_6, output_1_317;
mixer gate_output_1_317(.a(output_2_317), .b(output_2_6), .y(output_1_317));
wire output_3_317, output_3_6, output_2_317;
mixer gate_output_2_317(.a(output_3_317), .b(output_3_6), .y(output_2_317));
wire output_4_317, output_4_6, output_3_317;
mixer gate_output_3_317(.a(output_4_317), .b(output_4_6), .y(output_3_317));
wire output_5_317, output_5_6, output_4_317;
mixer gate_output_4_317(.a(output_5_317), .b(output_5_6), .y(output_4_317));
wire output_6_317, output_6_6, output_5_317;
mixer gate_output_5_317(.a(output_6_317), .b(output_6_6), .y(output_5_317));
wire output_7_317, output_7_6, output_6_317;
mixer gate_output_6_317(.a(output_7_317), .b(output_7_6), .y(output_6_317));
wire output_8_317, output_8_6, output_7_317;
mixer gate_output_7_317(.a(output_8_317), .b(output_8_6), .y(output_7_317));
wire output_1_318, output_1_7, output_0_318;
mixer gate_output_0_318(.a(output_1_318), .b(output_1_7), .y(output_0_318));
wire output_2_318, output_2_7, output_1_318;
mixer gate_output_1_318(.a(output_2_318), .b(output_2_7), .y(output_1_318));
wire output_3_318, output_3_7, output_2_318;
mixer gate_output_2_318(.a(output_3_318), .b(output_3_7), .y(output_2_318));
wire output_4_318, output_4_7, output_3_318;
mixer gate_output_3_318(.a(output_4_318), .b(output_4_7), .y(output_3_318));
wire output_5_318, output_5_7, output_4_318;
mixer gate_output_4_318(.a(output_5_318), .b(output_5_7), .y(output_4_318));
wire output_6_318, output_6_7, output_5_318;
mixer gate_output_5_318(.a(output_6_318), .b(output_6_7), .y(output_5_318));
wire output_7_318, output_7_7, output_6_318;
mixer gate_output_6_318(.a(output_7_318), .b(output_7_7), .y(output_6_318));
wire output_8_318, output_8_7, output_7_318;
mixer gate_output_7_318(.a(output_8_318), .b(output_8_7), .y(output_7_318));
wire output_1_319, output_1_0, output_0_319;
mixer gate_output_0_319(.a(output_1_319), .b(output_1_0), .y(output_0_319));
wire output_2_319, output_2_0, output_1_319;
mixer gate_output_1_319(.a(output_2_319), .b(output_2_0), .y(output_1_319));
wire output_3_319, output_3_0, output_2_319;
mixer gate_output_2_319(.a(output_3_319), .b(output_3_0), .y(output_2_319));
wire output_4_319, output_4_0, output_3_319;
mixer gate_output_3_319(.a(output_4_319), .b(output_4_0), .y(output_3_319));
wire output_5_319, output_5_0, output_4_319;
mixer gate_output_4_319(.a(output_5_319), .b(output_5_0), .y(output_4_319));
wire output_6_319, output_6_0, output_5_319;
mixer gate_output_5_319(.a(output_6_319), .b(output_6_0), .y(output_5_319));
wire output_7_319, output_7_0, output_6_319;
mixer gate_output_6_319(.a(output_7_319), .b(output_7_0), .y(output_6_319));
wire output_8_319, output_8_0, output_7_319;
mixer gate_output_7_319(.a(output_8_319), .b(output_8_0), .y(output_7_319));
wire output_1_320, output_1_1, output_0_320;
mixer gate_output_0_320(.a(output_1_320), .b(output_1_1), .y(output_0_320));
wire output_2_320, output_2_1, output_1_320;
mixer gate_output_1_320(.a(output_2_320), .b(output_2_1), .y(output_1_320));
wire output_3_320, output_3_1, output_2_320;
mixer gate_output_2_320(.a(output_3_320), .b(output_3_1), .y(output_2_320));
wire output_4_320, output_4_1, output_3_320;
mixer gate_output_3_320(.a(output_4_320), .b(output_4_1), .y(output_3_320));
wire output_5_320, output_5_1, output_4_320;
mixer gate_output_4_320(.a(output_5_320), .b(output_5_1), .y(output_4_320));
wire output_6_320, output_6_1, output_5_320;
mixer gate_output_5_320(.a(output_6_320), .b(output_6_1), .y(output_5_320));
wire output_7_320, output_7_1, output_6_320;
mixer gate_output_6_320(.a(output_7_320), .b(output_7_1), .y(output_6_320));
wire output_8_320, output_8_1, output_7_320;
mixer gate_output_7_320(.a(output_8_320), .b(output_8_1), .y(output_7_320));
wire output_1_321, output_1_2, output_0_321;
mixer gate_output_0_321(.a(output_1_321), .b(output_1_2), .y(output_0_321));
wire output_2_321, output_2_2, output_1_321;
mixer gate_output_1_321(.a(output_2_321), .b(output_2_2), .y(output_1_321));
wire output_3_321, output_3_2, output_2_321;
mixer gate_output_2_321(.a(output_3_321), .b(output_3_2), .y(output_2_321));
wire output_4_321, output_4_2, output_3_321;
mixer gate_output_3_321(.a(output_4_321), .b(output_4_2), .y(output_3_321));
wire output_5_321, output_5_2, output_4_321;
mixer gate_output_4_321(.a(output_5_321), .b(output_5_2), .y(output_4_321));
wire output_6_321, output_6_2, output_5_321;
mixer gate_output_5_321(.a(output_6_321), .b(output_6_2), .y(output_5_321));
wire output_7_321, output_7_2, output_6_321;
mixer gate_output_6_321(.a(output_7_321), .b(output_7_2), .y(output_6_321));
wire output_8_321, output_8_2, output_7_321;
mixer gate_output_7_321(.a(output_8_321), .b(output_8_2), .y(output_7_321));
wire output_1_322, output_1_3, output_0_322;
mixer gate_output_0_322(.a(output_1_322), .b(output_1_3), .y(output_0_322));
wire output_2_322, output_2_3, output_1_322;
mixer gate_output_1_322(.a(output_2_322), .b(output_2_3), .y(output_1_322));
wire output_3_322, output_3_3, output_2_322;
mixer gate_output_2_322(.a(output_3_322), .b(output_3_3), .y(output_2_322));
wire output_4_322, output_4_3, output_3_322;
mixer gate_output_3_322(.a(output_4_322), .b(output_4_3), .y(output_3_322));
wire output_5_322, output_5_3, output_4_322;
mixer gate_output_4_322(.a(output_5_322), .b(output_5_3), .y(output_4_322));
wire output_6_322, output_6_3, output_5_322;
mixer gate_output_5_322(.a(output_6_322), .b(output_6_3), .y(output_5_322));
wire output_7_322, output_7_3, output_6_322;
mixer gate_output_6_322(.a(output_7_322), .b(output_7_3), .y(output_6_322));
wire output_8_322, output_8_3, output_7_322;
mixer gate_output_7_322(.a(output_8_322), .b(output_8_3), .y(output_7_322));
wire output_1_323, output_1_4, output_0_323;
mixer gate_output_0_323(.a(output_1_323), .b(output_1_4), .y(output_0_323));
wire output_2_323, output_2_4, output_1_323;
mixer gate_output_1_323(.a(output_2_323), .b(output_2_4), .y(output_1_323));
wire output_3_323, output_3_4, output_2_323;
mixer gate_output_2_323(.a(output_3_323), .b(output_3_4), .y(output_2_323));
wire output_4_323, output_4_4, output_3_323;
mixer gate_output_3_323(.a(output_4_323), .b(output_4_4), .y(output_3_323));
wire output_5_323, output_5_4, output_4_323;
mixer gate_output_4_323(.a(output_5_323), .b(output_5_4), .y(output_4_323));
wire output_6_323, output_6_4, output_5_323;
mixer gate_output_5_323(.a(output_6_323), .b(output_6_4), .y(output_5_323));
wire output_7_323, output_7_4, output_6_323;
mixer gate_output_6_323(.a(output_7_323), .b(output_7_4), .y(output_6_323));
wire output_8_323, output_8_4, output_7_323;
mixer gate_output_7_323(.a(output_8_323), .b(output_8_4), .y(output_7_323));
wire output_1_324, output_1_5, output_0_324;
mixer gate_output_0_324(.a(output_1_324), .b(output_1_5), .y(output_0_324));
wire output_2_324, output_2_5, output_1_324;
mixer gate_output_1_324(.a(output_2_324), .b(output_2_5), .y(output_1_324));
wire output_3_324, output_3_5, output_2_324;
mixer gate_output_2_324(.a(output_3_324), .b(output_3_5), .y(output_2_324));
wire output_4_324, output_4_5, output_3_324;
mixer gate_output_3_324(.a(output_4_324), .b(output_4_5), .y(output_3_324));
wire output_5_324, output_5_5, output_4_324;
mixer gate_output_4_324(.a(output_5_324), .b(output_5_5), .y(output_4_324));
wire output_6_324, output_6_5, output_5_324;
mixer gate_output_5_324(.a(output_6_324), .b(output_6_5), .y(output_5_324));
wire output_7_324, output_7_5, output_6_324;
mixer gate_output_6_324(.a(output_7_324), .b(output_7_5), .y(output_6_324));
wire output_8_324, output_8_5, output_7_324;
mixer gate_output_7_324(.a(output_8_324), .b(output_8_5), .y(output_7_324));
wire output_1_325, output_1_6, output_0_325;
mixer gate_output_0_325(.a(output_1_325), .b(output_1_6), .y(output_0_325));
wire output_2_325, output_2_6, output_1_325;
mixer gate_output_1_325(.a(output_2_325), .b(output_2_6), .y(output_1_325));
wire output_3_325, output_3_6, output_2_325;
mixer gate_output_2_325(.a(output_3_325), .b(output_3_6), .y(output_2_325));
wire output_4_325, output_4_6, output_3_325;
mixer gate_output_3_325(.a(output_4_325), .b(output_4_6), .y(output_3_325));
wire output_5_325, output_5_6, output_4_325;
mixer gate_output_4_325(.a(output_5_325), .b(output_5_6), .y(output_4_325));
wire output_6_325, output_6_6, output_5_325;
mixer gate_output_5_325(.a(output_6_325), .b(output_6_6), .y(output_5_325));
wire output_7_325, output_7_6, output_6_325;
mixer gate_output_6_325(.a(output_7_325), .b(output_7_6), .y(output_6_325));
wire output_8_325, output_8_6, output_7_325;
mixer gate_output_7_325(.a(output_8_325), .b(output_8_6), .y(output_7_325));
wire output_1_326, output_1_7, output_0_326;
mixer gate_output_0_326(.a(output_1_326), .b(output_1_7), .y(output_0_326));
wire output_2_326, output_2_7, output_1_326;
mixer gate_output_1_326(.a(output_2_326), .b(output_2_7), .y(output_1_326));
wire output_3_326, output_3_7, output_2_326;
mixer gate_output_2_326(.a(output_3_326), .b(output_3_7), .y(output_2_326));
wire output_4_326, output_4_7, output_3_326;
mixer gate_output_3_326(.a(output_4_326), .b(output_4_7), .y(output_3_326));
wire output_5_326, output_5_7, output_4_326;
mixer gate_output_4_326(.a(output_5_326), .b(output_5_7), .y(output_4_326));
wire output_6_326, output_6_7, output_5_326;
mixer gate_output_5_326(.a(output_6_326), .b(output_6_7), .y(output_5_326));
wire output_7_326, output_7_7, output_6_326;
mixer gate_output_6_326(.a(output_7_326), .b(output_7_7), .y(output_6_326));
wire output_8_326, output_8_7, output_7_326;
mixer gate_output_7_326(.a(output_8_326), .b(output_8_7), .y(output_7_326));
wire output_1_327, output_1_0, output_0_327;
mixer gate_output_0_327(.a(output_1_327), .b(output_1_0), .y(output_0_327));
wire output_2_327, output_2_0, output_1_327;
mixer gate_output_1_327(.a(output_2_327), .b(output_2_0), .y(output_1_327));
wire output_3_327, output_3_0, output_2_327;
mixer gate_output_2_327(.a(output_3_327), .b(output_3_0), .y(output_2_327));
wire output_4_327, output_4_0, output_3_327;
mixer gate_output_3_327(.a(output_4_327), .b(output_4_0), .y(output_3_327));
wire output_5_327, output_5_0, output_4_327;
mixer gate_output_4_327(.a(output_5_327), .b(output_5_0), .y(output_4_327));
wire output_6_327, output_6_0, output_5_327;
mixer gate_output_5_327(.a(output_6_327), .b(output_6_0), .y(output_5_327));
wire output_7_327, output_7_0, output_6_327;
mixer gate_output_6_327(.a(output_7_327), .b(output_7_0), .y(output_6_327));
wire output_8_327, output_8_0, output_7_327;
mixer gate_output_7_327(.a(output_8_327), .b(output_8_0), .y(output_7_327));
wire output_1_328, output_1_1, output_0_328;
mixer gate_output_0_328(.a(output_1_328), .b(output_1_1), .y(output_0_328));
wire output_2_328, output_2_1, output_1_328;
mixer gate_output_1_328(.a(output_2_328), .b(output_2_1), .y(output_1_328));
wire output_3_328, output_3_1, output_2_328;
mixer gate_output_2_328(.a(output_3_328), .b(output_3_1), .y(output_2_328));
wire output_4_328, output_4_1, output_3_328;
mixer gate_output_3_328(.a(output_4_328), .b(output_4_1), .y(output_3_328));
wire output_5_328, output_5_1, output_4_328;
mixer gate_output_4_328(.a(output_5_328), .b(output_5_1), .y(output_4_328));
wire output_6_328, output_6_1, output_5_328;
mixer gate_output_5_328(.a(output_6_328), .b(output_6_1), .y(output_5_328));
wire output_7_328, output_7_1, output_6_328;
mixer gate_output_6_328(.a(output_7_328), .b(output_7_1), .y(output_6_328));
wire output_8_328, output_8_1, output_7_328;
mixer gate_output_7_328(.a(output_8_328), .b(output_8_1), .y(output_7_328));
wire output_1_329, output_1_2, output_0_329;
mixer gate_output_0_329(.a(output_1_329), .b(output_1_2), .y(output_0_329));
wire output_2_329, output_2_2, output_1_329;
mixer gate_output_1_329(.a(output_2_329), .b(output_2_2), .y(output_1_329));
wire output_3_329, output_3_2, output_2_329;
mixer gate_output_2_329(.a(output_3_329), .b(output_3_2), .y(output_2_329));
wire output_4_329, output_4_2, output_3_329;
mixer gate_output_3_329(.a(output_4_329), .b(output_4_2), .y(output_3_329));
wire output_5_329, output_5_2, output_4_329;
mixer gate_output_4_329(.a(output_5_329), .b(output_5_2), .y(output_4_329));
wire output_6_329, output_6_2, output_5_329;
mixer gate_output_5_329(.a(output_6_329), .b(output_6_2), .y(output_5_329));
wire output_7_329, output_7_2, output_6_329;
mixer gate_output_6_329(.a(output_7_329), .b(output_7_2), .y(output_6_329));
wire output_8_329, output_8_2, output_7_329;
mixer gate_output_7_329(.a(output_8_329), .b(output_8_2), .y(output_7_329));
wire output_1_330, output_1_3, output_0_330;
mixer gate_output_0_330(.a(output_1_330), .b(output_1_3), .y(output_0_330));
wire output_2_330, output_2_3, output_1_330;
mixer gate_output_1_330(.a(output_2_330), .b(output_2_3), .y(output_1_330));
wire output_3_330, output_3_3, output_2_330;
mixer gate_output_2_330(.a(output_3_330), .b(output_3_3), .y(output_2_330));
wire output_4_330, output_4_3, output_3_330;
mixer gate_output_3_330(.a(output_4_330), .b(output_4_3), .y(output_3_330));
wire output_5_330, output_5_3, output_4_330;
mixer gate_output_4_330(.a(output_5_330), .b(output_5_3), .y(output_4_330));
wire output_6_330, output_6_3, output_5_330;
mixer gate_output_5_330(.a(output_6_330), .b(output_6_3), .y(output_5_330));
wire output_7_330, output_7_3, output_6_330;
mixer gate_output_6_330(.a(output_7_330), .b(output_7_3), .y(output_6_330));
wire output_8_330, output_8_3, output_7_330;
mixer gate_output_7_330(.a(output_8_330), .b(output_8_3), .y(output_7_330));
wire output_1_331, output_1_4, output_0_331;
mixer gate_output_0_331(.a(output_1_331), .b(output_1_4), .y(output_0_331));
wire output_2_331, output_2_4, output_1_331;
mixer gate_output_1_331(.a(output_2_331), .b(output_2_4), .y(output_1_331));
wire output_3_331, output_3_4, output_2_331;
mixer gate_output_2_331(.a(output_3_331), .b(output_3_4), .y(output_2_331));
wire output_4_331, output_4_4, output_3_331;
mixer gate_output_3_331(.a(output_4_331), .b(output_4_4), .y(output_3_331));
wire output_5_331, output_5_4, output_4_331;
mixer gate_output_4_331(.a(output_5_331), .b(output_5_4), .y(output_4_331));
wire output_6_331, output_6_4, output_5_331;
mixer gate_output_5_331(.a(output_6_331), .b(output_6_4), .y(output_5_331));
wire output_7_331, output_7_4, output_6_331;
mixer gate_output_6_331(.a(output_7_331), .b(output_7_4), .y(output_6_331));
wire output_8_331, output_8_4, output_7_331;
mixer gate_output_7_331(.a(output_8_331), .b(output_8_4), .y(output_7_331));
wire output_1_332, output_1_5, output_0_332;
mixer gate_output_0_332(.a(output_1_332), .b(output_1_5), .y(output_0_332));
wire output_2_332, output_2_5, output_1_332;
mixer gate_output_1_332(.a(output_2_332), .b(output_2_5), .y(output_1_332));
wire output_3_332, output_3_5, output_2_332;
mixer gate_output_2_332(.a(output_3_332), .b(output_3_5), .y(output_2_332));
wire output_4_332, output_4_5, output_3_332;
mixer gate_output_3_332(.a(output_4_332), .b(output_4_5), .y(output_3_332));
wire output_5_332, output_5_5, output_4_332;
mixer gate_output_4_332(.a(output_5_332), .b(output_5_5), .y(output_4_332));
wire output_6_332, output_6_5, output_5_332;
mixer gate_output_5_332(.a(output_6_332), .b(output_6_5), .y(output_5_332));
wire output_7_332, output_7_5, output_6_332;
mixer gate_output_6_332(.a(output_7_332), .b(output_7_5), .y(output_6_332));
wire output_8_332, output_8_5, output_7_332;
mixer gate_output_7_332(.a(output_8_332), .b(output_8_5), .y(output_7_332));
wire output_1_333, output_1_6, output_0_333;
mixer gate_output_0_333(.a(output_1_333), .b(output_1_6), .y(output_0_333));
wire output_2_333, output_2_6, output_1_333;
mixer gate_output_1_333(.a(output_2_333), .b(output_2_6), .y(output_1_333));
wire output_3_333, output_3_6, output_2_333;
mixer gate_output_2_333(.a(output_3_333), .b(output_3_6), .y(output_2_333));
wire output_4_333, output_4_6, output_3_333;
mixer gate_output_3_333(.a(output_4_333), .b(output_4_6), .y(output_3_333));
wire output_5_333, output_5_6, output_4_333;
mixer gate_output_4_333(.a(output_5_333), .b(output_5_6), .y(output_4_333));
wire output_6_333, output_6_6, output_5_333;
mixer gate_output_5_333(.a(output_6_333), .b(output_6_6), .y(output_5_333));
wire output_7_333, output_7_6, output_6_333;
mixer gate_output_6_333(.a(output_7_333), .b(output_7_6), .y(output_6_333));
wire output_8_333, output_8_6, output_7_333;
mixer gate_output_7_333(.a(output_8_333), .b(output_8_6), .y(output_7_333));
wire output_1_334, output_1_7, output_0_334;
mixer gate_output_0_334(.a(output_1_334), .b(output_1_7), .y(output_0_334));
wire output_2_334, output_2_7, output_1_334;
mixer gate_output_1_334(.a(output_2_334), .b(output_2_7), .y(output_1_334));
wire output_3_334, output_3_7, output_2_334;
mixer gate_output_2_334(.a(output_3_334), .b(output_3_7), .y(output_2_334));
wire output_4_334, output_4_7, output_3_334;
mixer gate_output_3_334(.a(output_4_334), .b(output_4_7), .y(output_3_334));
wire output_5_334, output_5_7, output_4_334;
mixer gate_output_4_334(.a(output_5_334), .b(output_5_7), .y(output_4_334));
wire output_6_334, output_6_7, output_5_334;
mixer gate_output_5_334(.a(output_6_334), .b(output_6_7), .y(output_5_334));
wire output_7_334, output_7_7, output_6_334;
mixer gate_output_6_334(.a(output_7_334), .b(output_7_7), .y(output_6_334));
wire output_8_334, output_8_7, output_7_334;
mixer gate_output_7_334(.a(output_8_334), .b(output_8_7), .y(output_7_334));
wire output_1_335, output_1_0, output_0_335;
mixer gate_output_0_335(.a(output_1_335), .b(output_1_0), .y(output_0_335));
wire output_2_335, output_2_0, output_1_335;
mixer gate_output_1_335(.a(output_2_335), .b(output_2_0), .y(output_1_335));
wire output_3_335, output_3_0, output_2_335;
mixer gate_output_2_335(.a(output_3_335), .b(output_3_0), .y(output_2_335));
wire output_4_335, output_4_0, output_3_335;
mixer gate_output_3_335(.a(output_4_335), .b(output_4_0), .y(output_3_335));
wire output_5_335, output_5_0, output_4_335;
mixer gate_output_4_335(.a(output_5_335), .b(output_5_0), .y(output_4_335));
wire output_6_335, output_6_0, output_5_335;
mixer gate_output_5_335(.a(output_6_335), .b(output_6_0), .y(output_5_335));
wire output_7_335, output_7_0, output_6_335;
mixer gate_output_6_335(.a(output_7_335), .b(output_7_0), .y(output_6_335));
wire output_8_335, output_8_0, output_7_335;
mixer gate_output_7_335(.a(output_8_335), .b(output_8_0), .y(output_7_335));
wire output_1_336, output_1_1, output_0_336;
mixer gate_output_0_336(.a(output_1_336), .b(output_1_1), .y(output_0_336));
wire output_2_336, output_2_1, output_1_336;
mixer gate_output_1_336(.a(output_2_336), .b(output_2_1), .y(output_1_336));
wire output_3_336, output_3_1, output_2_336;
mixer gate_output_2_336(.a(output_3_336), .b(output_3_1), .y(output_2_336));
wire output_4_336, output_4_1, output_3_336;
mixer gate_output_3_336(.a(output_4_336), .b(output_4_1), .y(output_3_336));
wire output_5_336, output_5_1, output_4_336;
mixer gate_output_4_336(.a(output_5_336), .b(output_5_1), .y(output_4_336));
wire output_6_336, output_6_1, output_5_336;
mixer gate_output_5_336(.a(output_6_336), .b(output_6_1), .y(output_5_336));
wire output_7_336, output_7_1, output_6_336;
mixer gate_output_6_336(.a(output_7_336), .b(output_7_1), .y(output_6_336));
wire output_8_336, output_8_1, output_7_336;
mixer gate_output_7_336(.a(output_8_336), .b(output_8_1), .y(output_7_336));
wire output_1_337, output_1_2, output_0_337;
mixer gate_output_0_337(.a(output_1_337), .b(output_1_2), .y(output_0_337));
wire output_2_337, output_2_2, output_1_337;
mixer gate_output_1_337(.a(output_2_337), .b(output_2_2), .y(output_1_337));
wire output_3_337, output_3_2, output_2_337;
mixer gate_output_2_337(.a(output_3_337), .b(output_3_2), .y(output_2_337));
wire output_4_337, output_4_2, output_3_337;
mixer gate_output_3_337(.a(output_4_337), .b(output_4_2), .y(output_3_337));
wire output_5_337, output_5_2, output_4_337;
mixer gate_output_4_337(.a(output_5_337), .b(output_5_2), .y(output_4_337));
wire output_6_337, output_6_2, output_5_337;
mixer gate_output_5_337(.a(output_6_337), .b(output_6_2), .y(output_5_337));
wire output_7_337, output_7_2, output_6_337;
mixer gate_output_6_337(.a(output_7_337), .b(output_7_2), .y(output_6_337));
wire output_8_337, output_8_2, output_7_337;
mixer gate_output_7_337(.a(output_8_337), .b(output_8_2), .y(output_7_337));
wire output_1_338, output_1_3, output_0_338;
mixer gate_output_0_338(.a(output_1_338), .b(output_1_3), .y(output_0_338));
wire output_2_338, output_2_3, output_1_338;
mixer gate_output_1_338(.a(output_2_338), .b(output_2_3), .y(output_1_338));
wire output_3_338, output_3_3, output_2_338;
mixer gate_output_2_338(.a(output_3_338), .b(output_3_3), .y(output_2_338));
wire output_4_338, output_4_3, output_3_338;
mixer gate_output_3_338(.a(output_4_338), .b(output_4_3), .y(output_3_338));
wire output_5_338, output_5_3, output_4_338;
mixer gate_output_4_338(.a(output_5_338), .b(output_5_3), .y(output_4_338));
wire output_6_338, output_6_3, output_5_338;
mixer gate_output_5_338(.a(output_6_338), .b(output_6_3), .y(output_5_338));
wire output_7_338, output_7_3, output_6_338;
mixer gate_output_6_338(.a(output_7_338), .b(output_7_3), .y(output_6_338));
wire output_8_338, output_8_3, output_7_338;
mixer gate_output_7_338(.a(output_8_338), .b(output_8_3), .y(output_7_338));
wire output_1_339, output_1_4, output_0_339;
mixer gate_output_0_339(.a(output_1_339), .b(output_1_4), .y(output_0_339));
wire output_2_339, output_2_4, output_1_339;
mixer gate_output_1_339(.a(output_2_339), .b(output_2_4), .y(output_1_339));
wire output_3_339, output_3_4, output_2_339;
mixer gate_output_2_339(.a(output_3_339), .b(output_3_4), .y(output_2_339));
wire output_4_339, output_4_4, output_3_339;
mixer gate_output_3_339(.a(output_4_339), .b(output_4_4), .y(output_3_339));
wire output_5_339, output_5_4, output_4_339;
mixer gate_output_4_339(.a(output_5_339), .b(output_5_4), .y(output_4_339));
wire output_6_339, output_6_4, output_5_339;
mixer gate_output_5_339(.a(output_6_339), .b(output_6_4), .y(output_5_339));
wire output_7_339, output_7_4, output_6_339;
mixer gate_output_6_339(.a(output_7_339), .b(output_7_4), .y(output_6_339));
wire output_8_339, output_8_4, output_7_339;
mixer gate_output_7_339(.a(output_8_339), .b(output_8_4), .y(output_7_339));
wire output_1_340, output_1_5, output_0_340;
mixer gate_output_0_340(.a(output_1_340), .b(output_1_5), .y(output_0_340));
wire output_2_340, output_2_5, output_1_340;
mixer gate_output_1_340(.a(output_2_340), .b(output_2_5), .y(output_1_340));
wire output_3_340, output_3_5, output_2_340;
mixer gate_output_2_340(.a(output_3_340), .b(output_3_5), .y(output_2_340));
wire output_4_340, output_4_5, output_3_340;
mixer gate_output_3_340(.a(output_4_340), .b(output_4_5), .y(output_3_340));
wire output_5_340, output_5_5, output_4_340;
mixer gate_output_4_340(.a(output_5_340), .b(output_5_5), .y(output_4_340));
wire output_6_340, output_6_5, output_5_340;
mixer gate_output_5_340(.a(output_6_340), .b(output_6_5), .y(output_5_340));
wire output_7_340, output_7_5, output_6_340;
mixer gate_output_6_340(.a(output_7_340), .b(output_7_5), .y(output_6_340));
wire output_8_340, output_8_5, output_7_340;
mixer gate_output_7_340(.a(output_8_340), .b(output_8_5), .y(output_7_340));
wire output_1_341, output_1_6, output_0_341;
mixer gate_output_0_341(.a(output_1_341), .b(output_1_6), .y(output_0_341));
wire output_2_341, output_2_6, output_1_341;
mixer gate_output_1_341(.a(output_2_341), .b(output_2_6), .y(output_1_341));
wire output_3_341, output_3_6, output_2_341;
mixer gate_output_2_341(.a(output_3_341), .b(output_3_6), .y(output_2_341));
wire output_4_341, output_4_6, output_3_341;
mixer gate_output_3_341(.a(output_4_341), .b(output_4_6), .y(output_3_341));
wire output_5_341, output_5_6, output_4_341;
mixer gate_output_4_341(.a(output_5_341), .b(output_5_6), .y(output_4_341));
wire output_6_341, output_6_6, output_5_341;
mixer gate_output_5_341(.a(output_6_341), .b(output_6_6), .y(output_5_341));
wire output_7_341, output_7_6, output_6_341;
mixer gate_output_6_341(.a(output_7_341), .b(output_7_6), .y(output_6_341));
wire output_8_341, output_8_6, output_7_341;
mixer gate_output_7_341(.a(output_8_341), .b(output_8_6), .y(output_7_341));
wire output_1_342, output_1_7, output_0_342;
mixer gate_output_0_342(.a(output_1_342), .b(output_1_7), .y(output_0_342));
wire output_2_342, output_2_7, output_1_342;
mixer gate_output_1_342(.a(output_2_342), .b(output_2_7), .y(output_1_342));
wire output_3_342, output_3_7, output_2_342;
mixer gate_output_2_342(.a(output_3_342), .b(output_3_7), .y(output_2_342));
wire output_4_342, output_4_7, output_3_342;
mixer gate_output_3_342(.a(output_4_342), .b(output_4_7), .y(output_3_342));
wire output_5_342, output_5_7, output_4_342;
mixer gate_output_4_342(.a(output_5_342), .b(output_5_7), .y(output_4_342));
wire output_6_342, output_6_7, output_5_342;
mixer gate_output_5_342(.a(output_6_342), .b(output_6_7), .y(output_5_342));
wire output_7_342, output_7_7, output_6_342;
mixer gate_output_6_342(.a(output_7_342), .b(output_7_7), .y(output_6_342));
wire output_8_342, output_8_7, output_7_342;
mixer gate_output_7_342(.a(output_8_342), .b(output_8_7), .y(output_7_342));
wire output_1_343, output_1_0, output_0_343;
mixer gate_output_0_343(.a(output_1_343), .b(output_1_0), .y(output_0_343));
wire output_2_343, output_2_0, output_1_343;
mixer gate_output_1_343(.a(output_2_343), .b(output_2_0), .y(output_1_343));
wire output_3_343, output_3_0, output_2_343;
mixer gate_output_2_343(.a(output_3_343), .b(output_3_0), .y(output_2_343));
wire output_4_343, output_4_0, output_3_343;
mixer gate_output_3_343(.a(output_4_343), .b(output_4_0), .y(output_3_343));
wire output_5_343, output_5_0, output_4_343;
mixer gate_output_4_343(.a(output_5_343), .b(output_5_0), .y(output_4_343));
wire output_6_343, output_6_0, output_5_343;
mixer gate_output_5_343(.a(output_6_343), .b(output_6_0), .y(output_5_343));
wire output_7_343, output_7_0, output_6_343;
mixer gate_output_6_343(.a(output_7_343), .b(output_7_0), .y(output_6_343));
wire output_8_343, output_8_0, output_7_343;
mixer gate_output_7_343(.a(output_8_343), .b(output_8_0), .y(output_7_343));
wire output_1_344, output_1_1, output_0_344;
mixer gate_output_0_344(.a(output_1_344), .b(output_1_1), .y(output_0_344));
wire output_2_344, output_2_1, output_1_344;
mixer gate_output_1_344(.a(output_2_344), .b(output_2_1), .y(output_1_344));
wire output_3_344, output_3_1, output_2_344;
mixer gate_output_2_344(.a(output_3_344), .b(output_3_1), .y(output_2_344));
wire output_4_344, output_4_1, output_3_344;
mixer gate_output_3_344(.a(output_4_344), .b(output_4_1), .y(output_3_344));
wire output_5_344, output_5_1, output_4_344;
mixer gate_output_4_344(.a(output_5_344), .b(output_5_1), .y(output_4_344));
wire output_6_344, output_6_1, output_5_344;
mixer gate_output_5_344(.a(output_6_344), .b(output_6_1), .y(output_5_344));
wire output_7_344, output_7_1, output_6_344;
mixer gate_output_6_344(.a(output_7_344), .b(output_7_1), .y(output_6_344));
wire output_8_344, output_8_1, output_7_344;
mixer gate_output_7_344(.a(output_8_344), .b(output_8_1), .y(output_7_344));
wire output_1_345, output_1_2, output_0_345;
mixer gate_output_0_345(.a(output_1_345), .b(output_1_2), .y(output_0_345));
wire output_2_345, output_2_2, output_1_345;
mixer gate_output_1_345(.a(output_2_345), .b(output_2_2), .y(output_1_345));
wire output_3_345, output_3_2, output_2_345;
mixer gate_output_2_345(.a(output_3_345), .b(output_3_2), .y(output_2_345));
wire output_4_345, output_4_2, output_3_345;
mixer gate_output_3_345(.a(output_4_345), .b(output_4_2), .y(output_3_345));
wire output_5_345, output_5_2, output_4_345;
mixer gate_output_4_345(.a(output_5_345), .b(output_5_2), .y(output_4_345));
wire output_6_345, output_6_2, output_5_345;
mixer gate_output_5_345(.a(output_6_345), .b(output_6_2), .y(output_5_345));
wire output_7_345, output_7_2, output_6_345;
mixer gate_output_6_345(.a(output_7_345), .b(output_7_2), .y(output_6_345));
wire output_8_345, output_8_2, output_7_345;
mixer gate_output_7_345(.a(output_8_345), .b(output_8_2), .y(output_7_345));
wire output_1_346, output_1_3, output_0_346;
mixer gate_output_0_346(.a(output_1_346), .b(output_1_3), .y(output_0_346));
wire output_2_346, output_2_3, output_1_346;
mixer gate_output_1_346(.a(output_2_346), .b(output_2_3), .y(output_1_346));
wire output_3_346, output_3_3, output_2_346;
mixer gate_output_2_346(.a(output_3_346), .b(output_3_3), .y(output_2_346));
wire output_4_346, output_4_3, output_3_346;
mixer gate_output_3_346(.a(output_4_346), .b(output_4_3), .y(output_3_346));
wire output_5_346, output_5_3, output_4_346;
mixer gate_output_4_346(.a(output_5_346), .b(output_5_3), .y(output_4_346));
wire output_6_346, output_6_3, output_5_346;
mixer gate_output_5_346(.a(output_6_346), .b(output_6_3), .y(output_5_346));
wire output_7_346, output_7_3, output_6_346;
mixer gate_output_6_346(.a(output_7_346), .b(output_7_3), .y(output_6_346));
wire output_8_346, output_8_3, output_7_346;
mixer gate_output_7_346(.a(output_8_346), .b(output_8_3), .y(output_7_346));
wire output_1_347, output_1_4, output_0_347;
mixer gate_output_0_347(.a(output_1_347), .b(output_1_4), .y(output_0_347));
wire output_2_347, output_2_4, output_1_347;
mixer gate_output_1_347(.a(output_2_347), .b(output_2_4), .y(output_1_347));
wire output_3_347, output_3_4, output_2_347;
mixer gate_output_2_347(.a(output_3_347), .b(output_3_4), .y(output_2_347));
wire output_4_347, output_4_4, output_3_347;
mixer gate_output_3_347(.a(output_4_347), .b(output_4_4), .y(output_3_347));
wire output_5_347, output_5_4, output_4_347;
mixer gate_output_4_347(.a(output_5_347), .b(output_5_4), .y(output_4_347));
wire output_6_347, output_6_4, output_5_347;
mixer gate_output_5_347(.a(output_6_347), .b(output_6_4), .y(output_5_347));
wire output_7_347, output_7_4, output_6_347;
mixer gate_output_6_347(.a(output_7_347), .b(output_7_4), .y(output_6_347));
wire output_8_347, output_8_4, output_7_347;
mixer gate_output_7_347(.a(output_8_347), .b(output_8_4), .y(output_7_347));
wire output_1_348, output_1_5, output_0_348;
mixer gate_output_0_348(.a(output_1_348), .b(output_1_5), .y(output_0_348));
wire output_2_348, output_2_5, output_1_348;
mixer gate_output_1_348(.a(output_2_348), .b(output_2_5), .y(output_1_348));
wire output_3_348, output_3_5, output_2_348;
mixer gate_output_2_348(.a(output_3_348), .b(output_3_5), .y(output_2_348));
wire output_4_348, output_4_5, output_3_348;
mixer gate_output_3_348(.a(output_4_348), .b(output_4_5), .y(output_3_348));
wire output_5_348, output_5_5, output_4_348;
mixer gate_output_4_348(.a(output_5_348), .b(output_5_5), .y(output_4_348));
wire output_6_348, output_6_5, output_5_348;
mixer gate_output_5_348(.a(output_6_348), .b(output_6_5), .y(output_5_348));
wire output_7_348, output_7_5, output_6_348;
mixer gate_output_6_348(.a(output_7_348), .b(output_7_5), .y(output_6_348));
wire output_8_348, output_8_5, output_7_348;
mixer gate_output_7_348(.a(output_8_348), .b(output_8_5), .y(output_7_348));
wire output_1_349, output_1_6, output_0_349;
mixer gate_output_0_349(.a(output_1_349), .b(output_1_6), .y(output_0_349));
wire output_2_349, output_2_6, output_1_349;
mixer gate_output_1_349(.a(output_2_349), .b(output_2_6), .y(output_1_349));
wire output_3_349, output_3_6, output_2_349;
mixer gate_output_2_349(.a(output_3_349), .b(output_3_6), .y(output_2_349));
wire output_4_349, output_4_6, output_3_349;
mixer gate_output_3_349(.a(output_4_349), .b(output_4_6), .y(output_3_349));
wire output_5_349, output_5_6, output_4_349;
mixer gate_output_4_349(.a(output_5_349), .b(output_5_6), .y(output_4_349));
wire output_6_349, output_6_6, output_5_349;
mixer gate_output_5_349(.a(output_6_349), .b(output_6_6), .y(output_5_349));
wire output_7_349, output_7_6, output_6_349;
mixer gate_output_6_349(.a(output_7_349), .b(output_7_6), .y(output_6_349));
wire output_8_349, output_8_6, output_7_349;
mixer gate_output_7_349(.a(output_8_349), .b(output_8_6), .y(output_7_349));
wire output_1_350, output_1_7, output_0_350;
mixer gate_output_0_350(.a(output_1_350), .b(output_1_7), .y(output_0_350));
wire output_2_350, output_2_7, output_1_350;
mixer gate_output_1_350(.a(output_2_350), .b(output_2_7), .y(output_1_350));
wire output_3_350, output_3_7, output_2_350;
mixer gate_output_2_350(.a(output_3_350), .b(output_3_7), .y(output_2_350));
wire output_4_350, output_4_7, output_3_350;
mixer gate_output_3_350(.a(output_4_350), .b(output_4_7), .y(output_3_350));
wire output_5_350, output_5_7, output_4_350;
mixer gate_output_4_350(.a(output_5_350), .b(output_5_7), .y(output_4_350));
wire output_6_350, output_6_7, output_5_350;
mixer gate_output_5_350(.a(output_6_350), .b(output_6_7), .y(output_5_350));
wire output_7_350, output_7_7, output_6_350;
mixer gate_output_6_350(.a(output_7_350), .b(output_7_7), .y(output_6_350));
wire output_8_350, output_8_7, output_7_350;
mixer gate_output_7_350(.a(output_8_350), .b(output_8_7), .y(output_7_350));
wire output_1_351, output_1_0, output_0_351;
mixer gate_output_0_351(.a(output_1_351), .b(output_1_0), .y(output_0_351));
wire output_2_351, output_2_0, output_1_351;
mixer gate_output_1_351(.a(output_2_351), .b(output_2_0), .y(output_1_351));
wire output_3_351, output_3_0, output_2_351;
mixer gate_output_2_351(.a(output_3_351), .b(output_3_0), .y(output_2_351));
wire output_4_351, output_4_0, output_3_351;
mixer gate_output_3_351(.a(output_4_351), .b(output_4_0), .y(output_3_351));
wire output_5_351, output_5_0, output_4_351;
mixer gate_output_4_351(.a(output_5_351), .b(output_5_0), .y(output_4_351));
wire output_6_351, output_6_0, output_5_351;
mixer gate_output_5_351(.a(output_6_351), .b(output_6_0), .y(output_5_351));
wire output_7_351, output_7_0, output_6_351;
mixer gate_output_6_351(.a(output_7_351), .b(output_7_0), .y(output_6_351));
wire output_8_351, output_8_0, output_7_351;
mixer gate_output_7_351(.a(output_8_351), .b(output_8_0), .y(output_7_351));
wire output_1_352, output_1_1, output_0_352;
mixer gate_output_0_352(.a(output_1_352), .b(output_1_1), .y(output_0_352));
wire output_2_352, output_2_1, output_1_352;
mixer gate_output_1_352(.a(output_2_352), .b(output_2_1), .y(output_1_352));
wire output_3_352, output_3_1, output_2_352;
mixer gate_output_2_352(.a(output_3_352), .b(output_3_1), .y(output_2_352));
wire output_4_352, output_4_1, output_3_352;
mixer gate_output_3_352(.a(output_4_352), .b(output_4_1), .y(output_3_352));
wire output_5_352, output_5_1, output_4_352;
mixer gate_output_4_352(.a(output_5_352), .b(output_5_1), .y(output_4_352));
wire output_6_352, output_6_1, output_5_352;
mixer gate_output_5_352(.a(output_6_352), .b(output_6_1), .y(output_5_352));
wire output_7_352, output_7_1, output_6_352;
mixer gate_output_6_352(.a(output_7_352), .b(output_7_1), .y(output_6_352));
wire output_8_352, output_8_1, output_7_352;
mixer gate_output_7_352(.a(output_8_352), .b(output_8_1), .y(output_7_352));
wire output_1_353, output_1_2, output_0_353;
mixer gate_output_0_353(.a(output_1_353), .b(output_1_2), .y(output_0_353));
wire output_2_353, output_2_2, output_1_353;
mixer gate_output_1_353(.a(output_2_353), .b(output_2_2), .y(output_1_353));
wire output_3_353, output_3_2, output_2_353;
mixer gate_output_2_353(.a(output_3_353), .b(output_3_2), .y(output_2_353));
wire output_4_353, output_4_2, output_3_353;
mixer gate_output_3_353(.a(output_4_353), .b(output_4_2), .y(output_3_353));
wire output_5_353, output_5_2, output_4_353;
mixer gate_output_4_353(.a(output_5_353), .b(output_5_2), .y(output_4_353));
wire output_6_353, output_6_2, output_5_353;
mixer gate_output_5_353(.a(output_6_353), .b(output_6_2), .y(output_5_353));
wire output_7_353, output_7_2, output_6_353;
mixer gate_output_6_353(.a(output_7_353), .b(output_7_2), .y(output_6_353));
wire output_8_353, output_8_2, output_7_353;
mixer gate_output_7_353(.a(output_8_353), .b(output_8_2), .y(output_7_353));
wire output_1_354, output_1_3, output_0_354;
mixer gate_output_0_354(.a(output_1_354), .b(output_1_3), .y(output_0_354));
wire output_2_354, output_2_3, output_1_354;
mixer gate_output_1_354(.a(output_2_354), .b(output_2_3), .y(output_1_354));
wire output_3_354, output_3_3, output_2_354;
mixer gate_output_2_354(.a(output_3_354), .b(output_3_3), .y(output_2_354));
wire output_4_354, output_4_3, output_3_354;
mixer gate_output_3_354(.a(output_4_354), .b(output_4_3), .y(output_3_354));
wire output_5_354, output_5_3, output_4_354;
mixer gate_output_4_354(.a(output_5_354), .b(output_5_3), .y(output_4_354));
wire output_6_354, output_6_3, output_5_354;
mixer gate_output_5_354(.a(output_6_354), .b(output_6_3), .y(output_5_354));
wire output_7_354, output_7_3, output_6_354;
mixer gate_output_6_354(.a(output_7_354), .b(output_7_3), .y(output_6_354));
wire output_8_354, output_8_3, output_7_354;
mixer gate_output_7_354(.a(output_8_354), .b(output_8_3), .y(output_7_354));
wire output_1_355, output_1_4, output_0_355;
mixer gate_output_0_355(.a(output_1_355), .b(output_1_4), .y(output_0_355));
wire output_2_355, output_2_4, output_1_355;
mixer gate_output_1_355(.a(output_2_355), .b(output_2_4), .y(output_1_355));
wire output_3_355, output_3_4, output_2_355;
mixer gate_output_2_355(.a(output_3_355), .b(output_3_4), .y(output_2_355));
wire output_4_355, output_4_4, output_3_355;
mixer gate_output_3_355(.a(output_4_355), .b(output_4_4), .y(output_3_355));
wire output_5_355, output_5_4, output_4_355;
mixer gate_output_4_355(.a(output_5_355), .b(output_5_4), .y(output_4_355));
wire output_6_355, output_6_4, output_5_355;
mixer gate_output_5_355(.a(output_6_355), .b(output_6_4), .y(output_5_355));
wire output_7_355, output_7_4, output_6_355;
mixer gate_output_6_355(.a(output_7_355), .b(output_7_4), .y(output_6_355));
wire output_8_355, output_8_4, output_7_355;
mixer gate_output_7_355(.a(output_8_355), .b(output_8_4), .y(output_7_355));
wire output_1_356, output_1_5, output_0_356;
mixer gate_output_0_356(.a(output_1_356), .b(output_1_5), .y(output_0_356));
wire output_2_356, output_2_5, output_1_356;
mixer gate_output_1_356(.a(output_2_356), .b(output_2_5), .y(output_1_356));
wire output_3_356, output_3_5, output_2_356;
mixer gate_output_2_356(.a(output_3_356), .b(output_3_5), .y(output_2_356));
wire output_4_356, output_4_5, output_3_356;
mixer gate_output_3_356(.a(output_4_356), .b(output_4_5), .y(output_3_356));
wire output_5_356, output_5_5, output_4_356;
mixer gate_output_4_356(.a(output_5_356), .b(output_5_5), .y(output_4_356));
wire output_6_356, output_6_5, output_5_356;
mixer gate_output_5_356(.a(output_6_356), .b(output_6_5), .y(output_5_356));
wire output_7_356, output_7_5, output_6_356;
mixer gate_output_6_356(.a(output_7_356), .b(output_7_5), .y(output_6_356));
wire output_8_356, output_8_5, output_7_356;
mixer gate_output_7_356(.a(output_8_356), .b(output_8_5), .y(output_7_356));
wire output_1_357, output_1_6, output_0_357;
mixer gate_output_0_357(.a(output_1_357), .b(output_1_6), .y(output_0_357));
wire output_2_357, output_2_6, output_1_357;
mixer gate_output_1_357(.a(output_2_357), .b(output_2_6), .y(output_1_357));
wire output_3_357, output_3_6, output_2_357;
mixer gate_output_2_357(.a(output_3_357), .b(output_3_6), .y(output_2_357));
wire output_4_357, output_4_6, output_3_357;
mixer gate_output_3_357(.a(output_4_357), .b(output_4_6), .y(output_3_357));
wire output_5_357, output_5_6, output_4_357;
mixer gate_output_4_357(.a(output_5_357), .b(output_5_6), .y(output_4_357));
wire output_6_357, output_6_6, output_5_357;
mixer gate_output_5_357(.a(output_6_357), .b(output_6_6), .y(output_5_357));
wire output_7_357, output_7_6, output_6_357;
mixer gate_output_6_357(.a(output_7_357), .b(output_7_6), .y(output_6_357));
wire output_8_357, output_8_6, output_7_357;
mixer gate_output_7_357(.a(output_8_357), .b(output_8_6), .y(output_7_357));
wire output_1_358, output_1_7, output_0_358;
mixer gate_output_0_358(.a(output_1_358), .b(output_1_7), .y(output_0_358));
wire output_2_358, output_2_7, output_1_358;
mixer gate_output_1_358(.a(output_2_358), .b(output_2_7), .y(output_1_358));
wire output_3_358, output_3_7, output_2_358;
mixer gate_output_2_358(.a(output_3_358), .b(output_3_7), .y(output_2_358));
wire output_4_358, output_4_7, output_3_358;
mixer gate_output_3_358(.a(output_4_358), .b(output_4_7), .y(output_3_358));
wire output_5_358, output_5_7, output_4_358;
mixer gate_output_4_358(.a(output_5_358), .b(output_5_7), .y(output_4_358));
wire output_6_358, output_6_7, output_5_358;
mixer gate_output_5_358(.a(output_6_358), .b(output_6_7), .y(output_5_358));
wire output_7_358, output_7_7, output_6_358;
mixer gate_output_6_358(.a(output_7_358), .b(output_7_7), .y(output_6_358));
wire output_8_358, output_8_7, output_7_358;
mixer gate_output_7_358(.a(output_8_358), .b(output_8_7), .y(output_7_358));
wire output_1_359, output_1_0, output_0_359;
mixer gate_output_0_359(.a(output_1_359), .b(output_1_0), .y(output_0_359));
wire output_2_359, output_2_0, output_1_359;
mixer gate_output_1_359(.a(output_2_359), .b(output_2_0), .y(output_1_359));
wire output_3_359, output_3_0, output_2_359;
mixer gate_output_2_359(.a(output_3_359), .b(output_3_0), .y(output_2_359));
wire output_4_359, output_4_0, output_3_359;
mixer gate_output_3_359(.a(output_4_359), .b(output_4_0), .y(output_3_359));
wire output_5_359, output_5_0, output_4_359;
mixer gate_output_4_359(.a(output_5_359), .b(output_5_0), .y(output_4_359));
wire output_6_359, output_6_0, output_5_359;
mixer gate_output_5_359(.a(output_6_359), .b(output_6_0), .y(output_5_359));
wire output_7_359, output_7_0, output_6_359;
mixer gate_output_6_359(.a(output_7_359), .b(output_7_0), .y(output_6_359));
wire output_8_359, output_8_0, output_7_359;
mixer gate_output_7_359(.a(output_8_359), .b(output_8_0), .y(output_7_359));
wire output_1_360, output_1_1, output_0_360;
mixer gate_output_0_360(.a(output_1_360), .b(output_1_1), .y(output_0_360));
wire output_2_360, output_2_1, output_1_360;
mixer gate_output_1_360(.a(output_2_360), .b(output_2_1), .y(output_1_360));
wire output_3_360, output_3_1, output_2_360;
mixer gate_output_2_360(.a(output_3_360), .b(output_3_1), .y(output_2_360));
wire output_4_360, output_4_1, output_3_360;
mixer gate_output_3_360(.a(output_4_360), .b(output_4_1), .y(output_3_360));
wire output_5_360, output_5_1, output_4_360;
mixer gate_output_4_360(.a(output_5_360), .b(output_5_1), .y(output_4_360));
wire output_6_360, output_6_1, output_5_360;
mixer gate_output_5_360(.a(output_6_360), .b(output_6_1), .y(output_5_360));
wire output_7_360, output_7_1, output_6_360;
mixer gate_output_6_360(.a(output_7_360), .b(output_7_1), .y(output_6_360));
wire output_8_360, output_8_1, output_7_360;
mixer gate_output_7_360(.a(output_8_360), .b(output_8_1), .y(output_7_360));
wire output_1_361, output_1_2, output_0_361;
mixer gate_output_0_361(.a(output_1_361), .b(output_1_2), .y(output_0_361));
wire output_2_361, output_2_2, output_1_361;
mixer gate_output_1_361(.a(output_2_361), .b(output_2_2), .y(output_1_361));
wire output_3_361, output_3_2, output_2_361;
mixer gate_output_2_361(.a(output_3_361), .b(output_3_2), .y(output_2_361));
wire output_4_361, output_4_2, output_3_361;
mixer gate_output_3_361(.a(output_4_361), .b(output_4_2), .y(output_3_361));
wire output_5_361, output_5_2, output_4_361;
mixer gate_output_4_361(.a(output_5_361), .b(output_5_2), .y(output_4_361));
wire output_6_361, output_6_2, output_5_361;
mixer gate_output_5_361(.a(output_6_361), .b(output_6_2), .y(output_5_361));
wire output_7_361, output_7_2, output_6_361;
mixer gate_output_6_361(.a(output_7_361), .b(output_7_2), .y(output_6_361));
wire output_8_361, output_8_2, output_7_361;
mixer gate_output_7_361(.a(output_8_361), .b(output_8_2), .y(output_7_361));
wire output_1_362, output_1_3, output_0_362;
mixer gate_output_0_362(.a(output_1_362), .b(output_1_3), .y(output_0_362));
wire output_2_362, output_2_3, output_1_362;
mixer gate_output_1_362(.a(output_2_362), .b(output_2_3), .y(output_1_362));
wire output_3_362, output_3_3, output_2_362;
mixer gate_output_2_362(.a(output_3_362), .b(output_3_3), .y(output_2_362));
wire output_4_362, output_4_3, output_3_362;
mixer gate_output_3_362(.a(output_4_362), .b(output_4_3), .y(output_3_362));
wire output_5_362, output_5_3, output_4_362;
mixer gate_output_4_362(.a(output_5_362), .b(output_5_3), .y(output_4_362));
wire output_6_362, output_6_3, output_5_362;
mixer gate_output_5_362(.a(output_6_362), .b(output_6_3), .y(output_5_362));
wire output_7_362, output_7_3, output_6_362;
mixer gate_output_6_362(.a(output_7_362), .b(output_7_3), .y(output_6_362));
wire output_8_362, output_8_3, output_7_362;
mixer gate_output_7_362(.a(output_8_362), .b(output_8_3), .y(output_7_362));
wire output_1_363, output_1_4, output_0_363;
mixer gate_output_0_363(.a(output_1_363), .b(output_1_4), .y(output_0_363));
wire output_2_363, output_2_4, output_1_363;
mixer gate_output_1_363(.a(output_2_363), .b(output_2_4), .y(output_1_363));
wire output_3_363, output_3_4, output_2_363;
mixer gate_output_2_363(.a(output_3_363), .b(output_3_4), .y(output_2_363));
wire output_4_363, output_4_4, output_3_363;
mixer gate_output_3_363(.a(output_4_363), .b(output_4_4), .y(output_3_363));
wire output_5_363, output_5_4, output_4_363;
mixer gate_output_4_363(.a(output_5_363), .b(output_5_4), .y(output_4_363));
wire output_6_363, output_6_4, output_5_363;
mixer gate_output_5_363(.a(output_6_363), .b(output_6_4), .y(output_5_363));
wire output_7_363, output_7_4, output_6_363;
mixer gate_output_6_363(.a(output_7_363), .b(output_7_4), .y(output_6_363));
wire output_8_363, output_8_4, output_7_363;
mixer gate_output_7_363(.a(output_8_363), .b(output_8_4), .y(output_7_363));
wire output_1_364, output_1_5, output_0_364;
mixer gate_output_0_364(.a(output_1_364), .b(output_1_5), .y(output_0_364));
wire output_2_364, output_2_5, output_1_364;
mixer gate_output_1_364(.a(output_2_364), .b(output_2_5), .y(output_1_364));
wire output_3_364, output_3_5, output_2_364;
mixer gate_output_2_364(.a(output_3_364), .b(output_3_5), .y(output_2_364));
wire output_4_364, output_4_5, output_3_364;
mixer gate_output_3_364(.a(output_4_364), .b(output_4_5), .y(output_3_364));
wire output_5_364, output_5_5, output_4_364;
mixer gate_output_4_364(.a(output_5_364), .b(output_5_5), .y(output_4_364));
wire output_6_364, output_6_5, output_5_364;
mixer gate_output_5_364(.a(output_6_364), .b(output_6_5), .y(output_5_364));
wire output_7_364, output_7_5, output_6_364;
mixer gate_output_6_364(.a(output_7_364), .b(output_7_5), .y(output_6_364));
wire output_8_364, output_8_5, output_7_364;
mixer gate_output_7_364(.a(output_8_364), .b(output_8_5), .y(output_7_364));
wire output_1_365, output_1_6, output_0_365;
mixer gate_output_0_365(.a(output_1_365), .b(output_1_6), .y(output_0_365));
wire output_2_365, output_2_6, output_1_365;
mixer gate_output_1_365(.a(output_2_365), .b(output_2_6), .y(output_1_365));
wire output_3_365, output_3_6, output_2_365;
mixer gate_output_2_365(.a(output_3_365), .b(output_3_6), .y(output_2_365));
wire output_4_365, output_4_6, output_3_365;
mixer gate_output_3_365(.a(output_4_365), .b(output_4_6), .y(output_3_365));
wire output_5_365, output_5_6, output_4_365;
mixer gate_output_4_365(.a(output_5_365), .b(output_5_6), .y(output_4_365));
wire output_6_365, output_6_6, output_5_365;
mixer gate_output_5_365(.a(output_6_365), .b(output_6_6), .y(output_5_365));
wire output_7_365, output_7_6, output_6_365;
mixer gate_output_6_365(.a(output_7_365), .b(output_7_6), .y(output_6_365));
wire output_8_365, output_8_6, output_7_365;
mixer gate_output_7_365(.a(output_8_365), .b(output_8_6), .y(output_7_365));
wire output_1_366, output_1_7, output_0_366;
mixer gate_output_0_366(.a(output_1_366), .b(output_1_7), .y(output_0_366));
wire output_2_366, output_2_7, output_1_366;
mixer gate_output_1_366(.a(output_2_366), .b(output_2_7), .y(output_1_366));
wire output_3_366, output_3_7, output_2_366;
mixer gate_output_2_366(.a(output_3_366), .b(output_3_7), .y(output_2_366));
wire output_4_366, output_4_7, output_3_366;
mixer gate_output_3_366(.a(output_4_366), .b(output_4_7), .y(output_3_366));
wire output_5_366, output_5_7, output_4_366;
mixer gate_output_4_366(.a(output_5_366), .b(output_5_7), .y(output_4_366));
wire output_6_366, output_6_7, output_5_366;
mixer gate_output_5_366(.a(output_6_366), .b(output_6_7), .y(output_5_366));
wire output_7_366, output_7_7, output_6_366;
mixer gate_output_6_366(.a(output_7_366), .b(output_7_7), .y(output_6_366));
wire output_8_366, output_8_7, output_7_366;
mixer gate_output_7_366(.a(output_8_366), .b(output_8_7), .y(output_7_366));
wire output_1_367, output_1_0, output_0_367;
mixer gate_output_0_367(.a(output_1_367), .b(output_1_0), .y(output_0_367));
wire output_2_367, output_2_0, output_1_367;
mixer gate_output_1_367(.a(output_2_367), .b(output_2_0), .y(output_1_367));
wire output_3_367, output_3_0, output_2_367;
mixer gate_output_2_367(.a(output_3_367), .b(output_3_0), .y(output_2_367));
wire output_4_367, output_4_0, output_3_367;
mixer gate_output_3_367(.a(output_4_367), .b(output_4_0), .y(output_3_367));
wire output_5_367, output_5_0, output_4_367;
mixer gate_output_4_367(.a(output_5_367), .b(output_5_0), .y(output_4_367));
wire output_6_367, output_6_0, output_5_367;
mixer gate_output_5_367(.a(output_6_367), .b(output_6_0), .y(output_5_367));
wire output_7_367, output_7_0, output_6_367;
mixer gate_output_6_367(.a(output_7_367), .b(output_7_0), .y(output_6_367));
wire output_8_367, output_8_0, output_7_367;
mixer gate_output_7_367(.a(output_8_367), .b(output_8_0), .y(output_7_367));
wire output_1_368, output_1_1, output_0_368;
mixer gate_output_0_368(.a(output_1_368), .b(output_1_1), .y(output_0_368));
wire output_2_368, output_2_1, output_1_368;
mixer gate_output_1_368(.a(output_2_368), .b(output_2_1), .y(output_1_368));
wire output_3_368, output_3_1, output_2_368;
mixer gate_output_2_368(.a(output_3_368), .b(output_3_1), .y(output_2_368));
wire output_4_368, output_4_1, output_3_368;
mixer gate_output_3_368(.a(output_4_368), .b(output_4_1), .y(output_3_368));
wire output_5_368, output_5_1, output_4_368;
mixer gate_output_4_368(.a(output_5_368), .b(output_5_1), .y(output_4_368));
wire output_6_368, output_6_1, output_5_368;
mixer gate_output_5_368(.a(output_6_368), .b(output_6_1), .y(output_5_368));
wire output_7_368, output_7_1, output_6_368;
mixer gate_output_6_368(.a(output_7_368), .b(output_7_1), .y(output_6_368));
wire output_8_368, output_8_1, output_7_368;
mixer gate_output_7_368(.a(output_8_368), .b(output_8_1), .y(output_7_368));
wire output_1_369, output_1_2, output_0_369;
mixer gate_output_0_369(.a(output_1_369), .b(output_1_2), .y(output_0_369));
wire output_2_369, output_2_2, output_1_369;
mixer gate_output_1_369(.a(output_2_369), .b(output_2_2), .y(output_1_369));
wire output_3_369, output_3_2, output_2_369;
mixer gate_output_2_369(.a(output_3_369), .b(output_3_2), .y(output_2_369));
wire output_4_369, output_4_2, output_3_369;
mixer gate_output_3_369(.a(output_4_369), .b(output_4_2), .y(output_3_369));
wire output_5_369, output_5_2, output_4_369;
mixer gate_output_4_369(.a(output_5_369), .b(output_5_2), .y(output_4_369));
wire output_6_369, output_6_2, output_5_369;
mixer gate_output_5_369(.a(output_6_369), .b(output_6_2), .y(output_5_369));
wire output_7_369, output_7_2, output_6_369;
mixer gate_output_6_369(.a(output_7_369), .b(output_7_2), .y(output_6_369));
wire output_8_369, output_8_2, output_7_369;
mixer gate_output_7_369(.a(output_8_369), .b(output_8_2), .y(output_7_369));
wire output_1_370, output_1_3, output_0_370;
mixer gate_output_0_370(.a(output_1_370), .b(output_1_3), .y(output_0_370));
wire output_2_370, output_2_3, output_1_370;
mixer gate_output_1_370(.a(output_2_370), .b(output_2_3), .y(output_1_370));
wire output_3_370, output_3_3, output_2_370;
mixer gate_output_2_370(.a(output_3_370), .b(output_3_3), .y(output_2_370));
wire output_4_370, output_4_3, output_3_370;
mixer gate_output_3_370(.a(output_4_370), .b(output_4_3), .y(output_3_370));
wire output_5_370, output_5_3, output_4_370;
mixer gate_output_4_370(.a(output_5_370), .b(output_5_3), .y(output_4_370));
wire output_6_370, output_6_3, output_5_370;
mixer gate_output_5_370(.a(output_6_370), .b(output_6_3), .y(output_5_370));
wire output_7_370, output_7_3, output_6_370;
mixer gate_output_6_370(.a(output_7_370), .b(output_7_3), .y(output_6_370));
wire output_8_370, output_8_3, output_7_370;
mixer gate_output_7_370(.a(output_8_370), .b(output_8_3), .y(output_7_370));
wire output_1_371, output_1_4, output_0_371;
mixer gate_output_0_371(.a(output_1_371), .b(output_1_4), .y(output_0_371));
wire output_2_371, output_2_4, output_1_371;
mixer gate_output_1_371(.a(output_2_371), .b(output_2_4), .y(output_1_371));
wire output_3_371, output_3_4, output_2_371;
mixer gate_output_2_371(.a(output_3_371), .b(output_3_4), .y(output_2_371));
wire output_4_371, output_4_4, output_3_371;
mixer gate_output_3_371(.a(output_4_371), .b(output_4_4), .y(output_3_371));
wire output_5_371, output_5_4, output_4_371;
mixer gate_output_4_371(.a(output_5_371), .b(output_5_4), .y(output_4_371));
wire output_6_371, output_6_4, output_5_371;
mixer gate_output_5_371(.a(output_6_371), .b(output_6_4), .y(output_5_371));
wire output_7_371, output_7_4, output_6_371;
mixer gate_output_6_371(.a(output_7_371), .b(output_7_4), .y(output_6_371));
wire output_8_371, output_8_4, output_7_371;
mixer gate_output_7_371(.a(output_8_371), .b(output_8_4), .y(output_7_371));
wire output_1_372, output_1_5, output_0_372;
mixer gate_output_0_372(.a(output_1_372), .b(output_1_5), .y(output_0_372));
wire output_2_372, output_2_5, output_1_372;
mixer gate_output_1_372(.a(output_2_372), .b(output_2_5), .y(output_1_372));
wire output_3_372, output_3_5, output_2_372;
mixer gate_output_2_372(.a(output_3_372), .b(output_3_5), .y(output_2_372));
wire output_4_372, output_4_5, output_3_372;
mixer gate_output_3_372(.a(output_4_372), .b(output_4_5), .y(output_3_372));
wire output_5_372, output_5_5, output_4_372;
mixer gate_output_4_372(.a(output_5_372), .b(output_5_5), .y(output_4_372));
wire output_6_372, output_6_5, output_5_372;
mixer gate_output_5_372(.a(output_6_372), .b(output_6_5), .y(output_5_372));
wire output_7_372, output_7_5, output_6_372;
mixer gate_output_6_372(.a(output_7_372), .b(output_7_5), .y(output_6_372));
wire output_8_372, output_8_5, output_7_372;
mixer gate_output_7_372(.a(output_8_372), .b(output_8_5), .y(output_7_372));
wire output_1_373, output_1_6, output_0_373;
mixer gate_output_0_373(.a(output_1_373), .b(output_1_6), .y(output_0_373));
wire output_2_373, output_2_6, output_1_373;
mixer gate_output_1_373(.a(output_2_373), .b(output_2_6), .y(output_1_373));
wire output_3_373, output_3_6, output_2_373;
mixer gate_output_2_373(.a(output_3_373), .b(output_3_6), .y(output_2_373));
wire output_4_373, output_4_6, output_3_373;
mixer gate_output_3_373(.a(output_4_373), .b(output_4_6), .y(output_3_373));
wire output_5_373, output_5_6, output_4_373;
mixer gate_output_4_373(.a(output_5_373), .b(output_5_6), .y(output_4_373));
wire output_6_373, output_6_6, output_5_373;
mixer gate_output_5_373(.a(output_6_373), .b(output_6_6), .y(output_5_373));
wire output_7_373, output_7_6, output_6_373;
mixer gate_output_6_373(.a(output_7_373), .b(output_7_6), .y(output_6_373));
wire output_8_373, output_8_6, output_7_373;
mixer gate_output_7_373(.a(output_8_373), .b(output_8_6), .y(output_7_373));
wire output_1_374, output_1_7, output_0_374;
mixer gate_output_0_374(.a(output_1_374), .b(output_1_7), .y(output_0_374));
wire output_2_374, output_2_7, output_1_374;
mixer gate_output_1_374(.a(output_2_374), .b(output_2_7), .y(output_1_374));
wire output_3_374, output_3_7, output_2_374;
mixer gate_output_2_374(.a(output_3_374), .b(output_3_7), .y(output_2_374));
wire output_4_374, output_4_7, output_3_374;
mixer gate_output_3_374(.a(output_4_374), .b(output_4_7), .y(output_3_374));
wire output_5_374, output_5_7, output_4_374;
mixer gate_output_4_374(.a(output_5_374), .b(output_5_7), .y(output_4_374));
wire output_6_374, output_6_7, output_5_374;
mixer gate_output_5_374(.a(output_6_374), .b(output_6_7), .y(output_5_374));
wire output_7_374, output_7_7, output_6_374;
mixer gate_output_6_374(.a(output_7_374), .b(output_7_7), .y(output_6_374));
wire output_8_374, output_8_7, output_7_374;
mixer gate_output_7_374(.a(output_8_374), .b(output_8_7), .y(output_7_374));
wire output_1_375, output_1_0, output_0_375;
mixer gate_output_0_375(.a(output_1_375), .b(output_1_0), .y(output_0_375));
wire output_2_375, output_2_0, output_1_375;
mixer gate_output_1_375(.a(output_2_375), .b(output_2_0), .y(output_1_375));
wire output_3_375, output_3_0, output_2_375;
mixer gate_output_2_375(.a(output_3_375), .b(output_3_0), .y(output_2_375));
wire output_4_375, output_4_0, output_3_375;
mixer gate_output_3_375(.a(output_4_375), .b(output_4_0), .y(output_3_375));
wire output_5_375, output_5_0, output_4_375;
mixer gate_output_4_375(.a(output_5_375), .b(output_5_0), .y(output_4_375));
wire output_6_375, output_6_0, output_5_375;
mixer gate_output_5_375(.a(output_6_375), .b(output_6_0), .y(output_5_375));
wire output_7_375, output_7_0, output_6_375;
mixer gate_output_6_375(.a(output_7_375), .b(output_7_0), .y(output_6_375));
wire output_8_375, output_8_0, output_7_375;
mixer gate_output_7_375(.a(output_8_375), .b(output_8_0), .y(output_7_375));
wire output_1_376, output_1_1, output_0_376;
mixer gate_output_0_376(.a(output_1_376), .b(output_1_1), .y(output_0_376));
wire output_2_376, output_2_1, output_1_376;
mixer gate_output_1_376(.a(output_2_376), .b(output_2_1), .y(output_1_376));
wire output_3_376, output_3_1, output_2_376;
mixer gate_output_2_376(.a(output_3_376), .b(output_3_1), .y(output_2_376));
wire output_4_376, output_4_1, output_3_376;
mixer gate_output_3_376(.a(output_4_376), .b(output_4_1), .y(output_3_376));
wire output_5_376, output_5_1, output_4_376;
mixer gate_output_4_376(.a(output_5_376), .b(output_5_1), .y(output_4_376));
wire output_6_376, output_6_1, output_5_376;
mixer gate_output_5_376(.a(output_6_376), .b(output_6_1), .y(output_5_376));
wire output_7_376, output_7_1, output_6_376;
mixer gate_output_6_376(.a(output_7_376), .b(output_7_1), .y(output_6_376));
wire output_8_376, output_8_1, output_7_376;
mixer gate_output_7_376(.a(output_8_376), .b(output_8_1), .y(output_7_376));
wire output_1_377, output_1_2, output_0_377;
mixer gate_output_0_377(.a(output_1_377), .b(output_1_2), .y(output_0_377));
wire output_2_377, output_2_2, output_1_377;
mixer gate_output_1_377(.a(output_2_377), .b(output_2_2), .y(output_1_377));
wire output_3_377, output_3_2, output_2_377;
mixer gate_output_2_377(.a(output_3_377), .b(output_3_2), .y(output_2_377));
wire output_4_377, output_4_2, output_3_377;
mixer gate_output_3_377(.a(output_4_377), .b(output_4_2), .y(output_3_377));
wire output_5_377, output_5_2, output_4_377;
mixer gate_output_4_377(.a(output_5_377), .b(output_5_2), .y(output_4_377));
wire output_6_377, output_6_2, output_5_377;
mixer gate_output_5_377(.a(output_6_377), .b(output_6_2), .y(output_5_377));
wire output_7_377, output_7_2, output_6_377;
mixer gate_output_6_377(.a(output_7_377), .b(output_7_2), .y(output_6_377));
wire output_8_377, output_8_2, output_7_377;
mixer gate_output_7_377(.a(output_8_377), .b(output_8_2), .y(output_7_377));
wire output_1_378, output_1_3, output_0_378;
mixer gate_output_0_378(.a(output_1_378), .b(output_1_3), .y(output_0_378));
wire output_2_378, output_2_3, output_1_378;
mixer gate_output_1_378(.a(output_2_378), .b(output_2_3), .y(output_1_378));
wire output_3_378, output_3_3, output_2_378;
mixer gate_output_2_378(.a(output_3_378), .b(output_3_3), .y(output_2_378));
wire output_4_378, output_4_3, output_3_378;
mixer gate_output_3_378(.a(output_4_378), .b(output_4_3), .y(output_3_378));
wire output_5_378, output_5_3, output_4_378;
mixer gate_output_4_378(.a(output_5_378), .b(output_5_3), .y(output_4_378));
wire output_6_378, output_6_3, output_5_378;
mixer gate_output_5_378(.a(output_6_378), .b(output_6_3), .y(output_5_378));
wire output_7_378, output_7_3, output_6_378;
mixer gate_output_6_378(.a(output_7_378), .b(output_7_3), .y(output_6_378));
wire output_8_378, output_8_3, output_7_378;
mixer gate_output_7_378(.a(output_8_378), .b(output_8_3), .y(output_7_378));
wire output_1_379, output_1_4, output_0_379;
mixer gate_output_0_379(.a(output_1_379), .b(output_1_4), .y(output_0_379));
wire output_2_379, output_2_4, output_1_379;
mixer gate_output_1_379(.a(output_2_379), .b(output_2_4), .y(output_1_379));
wire output_3_379, output_3_4, output_2_379;
mixer gate_output_2_379(.a(output_3_379), .b(output_3_4), .y(output_2_379));
wire output_4_379, output_4_4, output_3_379;
mixer gate_output_3_379(.a(output_4_379), .b(output_4_4), .y(output_3_379));
wire output_5_379, output_5_4, output_4_379;
mixer gate_output_4_379(.a(output_5_379), .b(output_5_4), .y(output_4_379));
wire output_6_379, output_6_4, output_5_379;
mixer gate_output_5_379(.a(output_6_379), .b(output_6_4), .y(output_5_379));
wire output_7_379, output_7_4, output_6_379;
mixer gate_output_6_379(.a(output_7_379), .b(output_7_4), .y(output_6_379));
wire output_8_379, output_8_4, output_7_379;
mixer gate_output_7_379(.a(output_8_379), .b(output_8_4), .y(output_7_379));
wire output_1_380, output_1_5, output_0_380;
mixer gate_output_0_380(.a(output_1_380), .b(output_1_5), .y(output_0_380));
wire output_2_380, output_2_5, output_1_380;
mixer gate_output_1_380(.a(output_2_380), .b(output_2_5), .y(output_1_380));
wire output_3_380, output_3_5, output_2_380;
mixer gate_output_2_380(.a(output_3_380), .b(output_3_5), .y(output_2_380));
wire output_4_380, output_4_5, output_3_380;
mixer gate_output_3_380(.a(output_4_380), .b(output_4_5), .y(output_3_380));
wire output_5_380, output_5_5, output_4_380;
mixer gate_output_4_380(.a(output_5_380), .b(output_5_5), .y(output_4_380));
wire output_6_380, output_6_5, output_5_380;
mixer gate_output_5_380(.a(output_6_380), .b(output_6_5), .y(output_5_380));
wire output_7_380, output_7_5, output_6_380;
mixer gate_output_6_380(.a(output_7_380), .b(output_7_5), .y(output_6_380));
wire output_8_380, output_8_5, output_7_380;
mixer gate_output_7_380(.a(output_8_380), .b(output_8_5), .y(output_7_380));
wire output_1_381, output_1_6, output_0_381;
mixer gate_output_0_381(.a(output_1_381), .b(output_1_6), .y(output_0_381));
wire output_2_381, output_2_6, output_1_381;
mixer gate_output_1_381(.a(output_2_381), .b(output_2_6), .y(output_1_381));
wire output_3_381, output_3_6, output_2_381;
mixer gate_output_2_381(.a(output_3_381), .b(output_3_6), .y(output_2_381));
wire output_4_381, output_4_6, output_3_381;
mixer gate_output_3_381(.a(output_4_381), .b(output_4_6), .y(output_3_381));
wire output_5_381, output_5_6, output_4_381;
mixer gate_output_4_381(.a(output_5_381), .b(output_5_6), .y(output_4_381));
wire output_6_381, output_6_6, output_5_381;
mixer gate_output_5_381(.a(output_6_381), .b(output_6_6), .y(output_5_381));
wire output_7_381, output_7_6, output_6_381;
mixer gate_output_6_381(.a(output_7_381), .b(output_7_6), .y(output_6_381));
wire output_8_381, output_8_6, output_7_381;
mixer gate_output_7_381(.a(output_8_381), .b(output_8_6), .y(output_7_381));
wire output_1_382, output_1_7, output_0_382;
mixer gate_output_0_382(.a(output_1_382), .b(output_1_7), .y(output_0_382));
wire output_2_382, output_2_7, output_1_382;
mixer gate_output_1_382(.a(output_2_382), .b(output_2_7), .y(output_1_382));
wire output_3_382, output_3_7, output_2_382;
mixer gate_output_2_382(.a(output_3_382), .b(output_3_7), .y(output_2_382));
wire output_4_382, output_4_7, output_3_382;
mixer gate_output_3_382(.a(output_4_382), .b(output_4_7), .y(output_3_382));
wire output_5_382, output_5_7, output_4_382;
mixer gate_output_4_382(.a(output_5_382), .b(output_5_7), .y(output_4_382));
wire output_6_382, output_6_7, output_5_382;
mixer gate_output_5_382(.a(output_6_382), .b(output_6_7), .y(output_5_382));
wire output_7_382, output_7_7, output_6_382;
mixer gate_output_6_382(.a(output_7_382), .b(output_7_7), .y(output_6_382));
wire output_8_382, output_8_7, output_7_382;
mixer gate_output_7_382(.a(output_8_382), .b(output_8_7), .y(output_7_382));
wire output_1_383, output_1_0, output_0_383;
mixer gate_output_0_383(.a(output_1_383), .b(output_1_0), .y(output_0_383));
wire output_2_383, output_2_0, output_1_383;
mixer gate_output_1_383(.a(output_2_383), .b(output_2_0), .y(output_1_383));
wire output_3_383, output_3_0, output_2_383;
mixer gate_output_2_383(.a(output_3_383), .b(output_3_0), .y(output_2_383));
wire output_4_383, output_4_0, output_3_383;
mixer gate_output_3_383(.a(output_4_383), .b(output_4_0), .y(output_3_383));
wire output_5_383, output_5_0, output_4_383;
mixer gate_output_4_383(.a(output_5_383), .b(output_5_0), .y(output_4_383));
wire output_6_383, output_6_0, output_5_383;
mixer gate_output_5_383(.a(output_6_383), .b(output_6_0), .y(output_5_383));
wire output_7_383, output_7_0, output_6_383;
mixer gate_output_6_383(.a(output_7_383), .b(output_7_0), .y(output_6_383));
wire output_8_383, output_8_0, output_7_383;
mixer gate_output_7_383(.a(output_8_383), .b(output_8_0), .y(output_7_383));
wire output_1_384, output_1_1, output_0_384;
mixer gate_output_0_384(.a(output_1_384), .b(output_1_1), .y(output_0_384));
wire output_2_384, output_2_1, output_1_384;
mixer gate_output_1_384(.a(output_2_384), .b(output_2_1), .y(output_1_384));
wire output_3_384, output_3_1, output_2_384;
mixer gate_output_2_384(.a(output_3_384), .b(output_3_1), .y(output_2_384));
wire output_4_384, output_4_1, output_3_384;
mixer gate_output_3_384(.a(output_4_384), .b(output_4_1), .y(output_3_384));
wire output_5_384, output_5_1, output_4_384;
mixer gate_output_4_384(.a(output_5_384), .b(output_5_1), .y(output_4_384));
wire output_6_384, output_6_1, output_5_384;
mixer gate_output_5_384(.a(output_6_384), .b(output_6_1), .y(output_5_384));
wire output_7_384, output_7_1, output_6_384;
mixer gate_output_6_384(.a(output_7_384), .b(output_7_1), .y(output_6_384));
wire output_8_384, output_8_1, output_7_384;
mixer gate_output_7_384(.a(output_8_384), .b(output_8_1), .y(output_7_384));
wire output_1_385, output_1_2, output_0_385;
mixer gate_output_0_385(.a(output_1_385), .b(output_1_2), .y(output_0_385));
wire output_2_385, output_2_2, output_1_385;
mixer gate_output_1_385(.a(output_2_385), .b(output_2_2), .y(output_1_385));
wire output_3_385, output_3_2, output_2_385;
mixer gate_output_2_385(.a(output_3_385), .b(output_3_2), .y(output_2_385));
wire output_4_385, output_4_2, output_3_385;
mixer gate_output_3_385(.a(output_4_385), .b(output_4_2), .y(output_3_385));
wire output_5_385, output_5_2, output_4_385;
mixer gate_output_4_385(.a(output_5_385), .b(output_5_2), .y(output_4_385));
wire output_6_385, output_6_2, output_5_385;
mixer gate_output_5_385(.a(output_6_385), .b(output_6_2), .y(output_5_385));
wire output_7_385, output_7_2, output_6_385;
mixer gate_output_6_385(.a(output_7_385), .b(output_7_2), .y(output_6_385));
wire output_8_385, output_8_2, output_7_385;
mixer gate_output_7_385(.a(output_8_385), .b(output_8_2), .y(output_7_385));
wire output_1_386, output_1_3, output_0_386;
mixer gate_output_0_386(.a(output_1_386), .b(output_1_3), .y(output_0_386));
wire output_2_386, output_2_3, output_1_386;
mixer gate_output_1_386(.a(output_2_386), .b(output_2_3), .y(output_1_386));
wire output_3_386, output_3_3, output_2_386;
mixer gate_output_2_386(.a(output_3_386), .b(output_3_3), .y(output_2_386));
wire output_4_386, output_4_3, output_3_386;
mixer gate_output_3_386(.a(output_4_386), .b(output_4_3), .y(output_3_386));
wire output_5_386, output_5_3, output_4_386;
mixer gate_output_4_386(.a(output_5_386), .b(output_5_3), .y(output_4_386));
wire output_6_386, output_6_3, output_5_386;
mixer gate_output_5_386(.a(output_6_386), .b(output_6_3), .y(output_5_386));
wire output_7_386, output_7_3, output_6_386;
mixer gate_output_6_386(.a(output_7_386), .b(output_7_3), .y(output_6_386));
wire output_8_386, output_8_3, output_7_386;
mixer gate_output_7_386(.a(output_8_386), .b(output_8_3), .y(output_7_386));
wire output_1_387, output_1_4, output_0_387;
mixer gate_output_0_387(.a(output_1_387), .b(output_1_4), .y(output_0_387));
wire output_2_387, output_2_4, output_1_387;
mixer gate_output_1_387(.a(output_2_387), .b(output_2_4), .y(output_1_387));
wire output_3_387, output_3_4, output_2_387;
mixer gate_output_2_387(.a(output_3_387), .b(output_3_4), .y(output_2_387));
wire output_4_387, output_4_4, output_3_387;
mixer gate_output_3_387(.a(output_4_387), .b(output_4_4), .y(output_3_387));
wire output_5_387, output_5_4, output_4_387;
mixer gate_output_4_387(.a(output_5_387), .b(output_5_4), .y(output_4_387));
wire output_6_387, output_6_4, output_5_387;
mixer gate_output_5_387(.a(output_6_387), .b(output_6_4), .y(output_5_387));
wire output_7_387, output_7_4, output_6_387;
mixer gate_output_6_387(.a(output_7_387), .b(output_7_4), .y(output_6_387));
wire output_8_387, output_8_4, output_7_387;
mixer gate_output_7_387(.a(output_8_387), .b(output_8_4), .y(output_7_387));
wire output_1_388, output_1_5, output_0_388;
mixer gate_output_0_388(.a(output_1_388), .b(output_1_5), .y(output_0_388));
wire output_2_388, output_2_5, output_1_388;
mixer gate_output_1_388(.a(output_2_388), .b(output_2_5), .y(output_1_388));
wire output_3_388, output_3_5, output_2_388;
mixer gate_output_2_388(.a(output_3_388), .b(output_3_5), .y(output_2_388));
wire output_4_388, output_4_5, output_3_388;
mixer gate_output_3_388(.a(output_4_388), .b(output_4_5), .y(output_3_388));
wire output_5_388, output_5_5, output_4_388;
mixer gate_output_4_388(.a(output_5_388), .b(output_5_5), .y(output_4_388));
wire output_6_388, output_6_5, output_5_388;
mixer gate_output_5_388(.a(output_6_388), .b(output_6_5), .y(output_5_388));
wire output_7_388, output_7_5, output_6_388;
mixer gate_output_6_388(.a(output_7_388), .b(output_7_5), .y(output_6_388));
wire output_8_388, output_8_5, output_7_388;
mixer gate_output_7_388(.a(output_8_388), .b(output_8_5), .y(output_7_388));
wire output_1_389, output_1_6, output_0_389;
mixer gate_output_0_389(.a(output_1_389), .b(output_1_6), .y(output_0_389));
wire output_2_389, output_2_6, output_1_389;
mixer gate_output_1_389(.a(output_2_389), .b(output_2_6), .y(output_1_389));
wire output_3_389, output_3_6, output_2_389;
mixer gate_output_2_389(.a(output_3_389), .b(output_3_6), .y(output_2_389));
wire output_4_389, output_4_6, output_3_389;
mixer gate_output_3_389(.a(output_4_389), .b(output_4_6), .y(output_3_389));
wire output_5_389, output_5_6, output_4_389;
mixer gate_output_4_389(.a(output_5_389), .b(output_5_6), .y(output_4_389));
wire output_6_389, output_6_6, output_5_389;
mixer gate_output_5_389(.a(output_6_389), .b(output_6_6), .y(output_5_389));
wire output_7_389, output_7_6, output_6_389;
mixer gate_output_6_389(.a(output_7_389), .b(output_7_6), .y(output_6_389));
wire output_8_389, output_8_6, output_7_389;
mixer gate_output_7_389(.a(output_8_389), .b(output_8_6), .y(output_7_389));
wire output_1_390, output_1_7, output_0_390;
mixer gate_output_0_390(.a(output_1_390), .b(output_1_7), .y(output_0_390));
wire output_2_390, output_2_7, output_1_390;
mixer gate_output_1_390(.a(output_2_390), .b(output_2_7), .y(output_1_390));
wire output_3_390, output_3_7, output_2_390;
mixer gate_output_2_390(.a(output_3_390), .b(output_3_7), .y(output_2_390));
wire output_4_390, output_4_7, output_3_390;
mixer gate_output_3_390(.a(output_4_390), .b(output_4_7), .y(output_3_390));
wire output_5_390, output_5_7, output_4_390;
mixer gate_output_4_390(.a(output_5_390), .b(output_5_7), .y(output_4_390));
wire output_6_390, output_6_7, output_5_390;
mixer gate_output_5_390(.a(output_6_390), .b(output_6_7), .y(output_5_390));
wire output_7_390, output_7_7, output_6_390;
mixer gate_output_6_390(.a(output_7_390), .b(output_7_7), .y(output_6_390));
wire output_8_390, output_8_7, output_7_390;
mixer gate_output_7_390(.a(output_8_390), .b(output_8_7), .y(output_7_390));
wire output_1_391, output_1_0, output_0_391;
mixer gate_output_0_391(.a(output_1_391), .b(output_1_0), .y(output_0_391));
wire output_2_391, output_2_0, output_1_391;
mixer gate_output_1_391(.a(output_2_391), .b(output_2_0), .y(output_1_391));
wire output_3_391, output_3_0, output_2_391;
mixer gate_output_2_391(.a(output_3_391), .b(output_3_0), .y(output_2_391));
wire output_4_391, output_4_0, output_3_391;
mixer gate_output_3_391(.a(output_4_391), .b(output_4_0), .y(output_3_391));
wire output_5_391, output_5_0, output_4_391;
mixer gate_output_4_391(.a(output_5_391), .b(output_5_0), .y(output_4_391));
wire output_6_391, output_6_0, output_5_391;
mixer gate_output_5_391(.a(output_6_391), .b(output_6_0), .y(output_5_391));
wire output_7_391, output_7_0, output_6_391;
mixer gate_output_6_391(.a(output_7_391), .b(output_7_0), .y(output_6_391));
wire output_8_391, output_8_0, output_7_391;
mixer gate_output_7_391(.a(output_8_391), .b(output_8_0), .y(output_7_391));
wire output_1_392, output_1_1, output_0_392;
mixer gate_output_0_392(.a(output_1_392), .b(output_1_1), .y(output_0_392));
wire output_2_392, output_2_1, output_1_392;
mixer gate_output_1_392(.a(output_2_392), .b(output_2_1), .y(output_1_392));
wire output_3_392, output_3_1, output_2_392;
mixer gate_output_2_392(.a(output_3_392), .b(output_3_1), .y(output_2_392));
wire output_4_392, output_4_1, output_3_392;
mixer gate_output_3_392(.a(output_4_392), .b(output_4_1), .y(output_3_392));
wire output_5_392, output_5_1, output_4_392;
mixer gate_output_4_392(.a(output_5_392), .b(output_5_1), .y(output_4_392));
wire output_6_392, output_6_1, output_5_392;
mixer gate_output_5_392(.a(output_6_392), .b(output_6_1), .y(output_5_392));
wire output_7_392, output_7_1, output_6_392;
mixer gate_output_6_392(.a(output_7_392), .b(output_7_1), .y(output_6_392));
wire output_8_392, output_8_1, output_7_392;
mixer gate_output_7_392(.a(output_8_392), .b(output_8_1), .y(output_7_392));
wire output_1_393, output_1_2, output_0_393;
mixer gate_output_0_393(.a(output_1_393), .b(output_1_2), .y(output_0_393));
wire output_2_393, output_2_2, output_1_393;
mixer gate_output_1_393(.a(output_2_393), .b(output_2_2), .y(output_1_393));
wire output_3_393, output_3_2, output_2_393;
mixer gate_output_2_393(.a(output_3_393), .b(output_3_2), .y(output_2_393));
wire output_4_393, output_4_2, output_3_393;
mixer gate_output_3_393(.a(output_4_393), .b(output_4_2), .y(output_3_393));
wire output_5_393, output_5_2, output_4_393;
mixer gate_output_4_393(.a(output_5_393), .b(output_5_2), .y(output_4_393));
wire output_6_393, output_6_2, output_5_393;
mixer gate_output_5_393(.a(output_6_393), .b(output_6_2), .y(output_5_393));
wire output_7_393, output_7_2, output_6_393;
mixer gate_output_6_393(.a(output_7_393), .b(output_7_2), .y(output_6_393));
wire output_8_393, output_8_2, output_7_393;
mixer gate_output_7_393(.a(output_8_393), .b(output_8_2), .y(output_7_393));
wire output_1_394, output_1_3, output_0_394;
mixer gate_output_0_394(.a(output_1_394), .b(output_1_3), .y(output_0_394));
wire output_2_394, output_2_3, output_1_394;
mixer gate_output_1_394(.a(output_2_394), .b(output_2_3), .y(output_1_394));
wire output_3_394, output_3_3, output_2_394;
mixer gate_output_2_394(.a(output_3_394), .b(output_3_3), .y(output_2_394));
wire output_4_394, output_4_3, output_3_394;
mixer gate_output_3_394(.a(output_4_394), .b(output_4_3), .y(output_3_394));
wire output_5_394, output_5_3, output_4_394;
mixer gate_output_4_394(.a(output_5_394), .b(output_5_3), .y(output_4_394));
wire output_6_394, output_6_3, output_5_394;
mixer gate_output_5_394(.a(output_6_394), .b(output_6_3), .y(output_5_394));
wire output_7_394, output_7_3, output_6_394;
mixer gate_output_6_394(.a(output_7_394), .b(output_7_3), .y(output_6_394));
wire output_8_394, output_8_3, output_7_394;
mixer gate_output_7_394(.a(output_8_394), .b(output_8_3), .y(output_7_394));
wire output_1_395, output_1_4, output_0_395;
mixer gate_output_0_395(.a(output_1_395), .b(output_1_4), .y(output_0_395));
wire output_2_395, output_2_4, output_1_395;
mixer gate_output_1_395(.a(output_2_395), .b(output_2_4), .y(output_1_395));
wire output_3_395, output_3_4, output_2_395;
mixer gate_output_2_395(.a(output_3_395), .b(output_3_4), .y(output_2_395));
wire output_4_395, output_4_4, output_3_395;
mixer gate_output_3_395(.a(output_4_395), .b(output_4_4), .y(output_3_395));
wire output_5_395, output_5_4, output_4_395;
mixer gate_output_4_395(.a(output_5_395), .b(output_5_4), .y(output_4_395));
wire output_6_395, output_6_4, output_5_395;
mixer gate_output_5_395(.a(output_6_395), .b(output_6_4), .y(output_5_395));
wire output_7_395, output_7_4, output_6_395;
mixer gate_output_6_395(.a(output_7_395), .b(output_7_4), .y(output_6_395));
wire output_8_395, output_8_4, output_7_395;
mixer gate_output_7_395(.a(output_8_395), .b(output_8_4), .y(output_7_395));
wire output_1_396, output_1_5, output_0_396;
mixer gate_output_0_396(.a(output_1_396), .b(output_1_5), .y(output_0_396));
wire output_2_396, output_2_5, output_1_396;
mixer gate_output_1_396(.a(output_2_396), .b(output_2_5), .y(output_1_396));
wire output_3_396, output_3_5, output_2_396;
mixer gate_output_2_396(.a(output_3_396), .b(output_3_5), .y(output_2_396));
wire output_4_396, output_4_5, output_3_396;
mixer gate_output_3_396(.a(output_4_396), .b(output_4_5), .y(output_3_396));
wire output_5_396, output_5_5, output_4_396;
mixer gate_output_4_396(.a(output_5_396), .b(output_5_5), .y(output_4_396));
wire output_6_396, output_6_5, output_5_396;
mixer gate_output_5_396(.a(output_6_396), .b(output_6_5), .y(output_5_396));
wire output_7_396, output_7_5, output_6_396;
mixer gate_output_6_396(.a(output_7_396), .b(output_7_5), .y(output_6_396));
wire output_8_396, output_8_5, output_7_396;
mixer gate_output_7_396(.a(output_8_396), .b(output_8_5), .y(output_7_396));
wire output_1_397, output_1_6, output_0_397;
mixer gate_output_0_397(.a(output_1_397), .b(output_1_6), .y(output_0_397));
wire output_2_397, output_2_6, output_1_397;
mixer gate_output_1_397(.a(output_2_397), .b(output_2_6), .y(output_1_397));
wire output_3_397, output_3_6, output_2_397;
mixer gate_output_2_397(.a(output_3_397), .b(output_3_6), .y(output_2_397));
wire output_4_397, output_4_6, output_3_397;
mixer gate_output_3_397(.a(output_4_397), .b(output_4_6), .y(output_3_397));
wire output_5_397, output_5_6, output_4_397;
mixer gate_output_4_397(.a(output_5_397), .b(output_5_6), .y(output_4_397));
wire output_6_397, output_6_6, output_5_397;
mixer gate_output_5_397(.a(output_6_397), .b(output_6_6), .y(output_5_397));
wire output_7_397, output_7_6, output_6_397;
mixer gate_output_6_397(.a(output_7_397), .b(output_7_6), .y(output_6_397));
wire output_8_397, output_8_6, output_7_397;
mixer gate_output_7_397(.a(output_8_397), .b(output_8_6), .y(output_7_397));
wire output_1_398, output_1_7, output_0_398;
mixer gate_output_0_398(.a(output_1_398), .b(output_1_7), .y(output_0_398));
wire output_2_398, output_2_7, output_1_398;
mixer gate_output_1_398(.a(output_2_398), .b(output_2_7), .y(output_1_398));
wire output_3_398, output_3_7, output_2_398;
mixer gate_output_2_398(.a(output_3_398), .b(output_3_7), .y(output_2_398));
wire output_4_398, output_4_7, output_3_398;
mixer gate_output_3_398(.a(output_4_398), .b(output_4_7), .y(output_3_398));
wire output_5_398, output_5_7, output_4_398;
mixer gate_output_4_398(.a(output_5_398), .b(output_5_7), .y(output_4_398));
wire output_6_398, output_6_7, output_5_398;
mixer gate_output_5_398(.a(output_6_398), .b(output_6_7), .y(output_5_398));
wire output_7_398, output_7_7, output_6_398;
mixer gate_output_6_398(.a(output_7_398), .b(output_7_7), .y(output_6_398));
wire output_8_398, output_8_7, output_7_398;
mixer gate_output_7_398(.a(output_8_398), .b(output_8_7), .y(output_7_398));
wire output_1_399, output_1_0, output_0_399;
mixer gate_output_0_399(.a(output_1_399), .b(output_1_0), .y(output_0_399));
wire output_2_399, output_2_0, output_1_399;
mixer gate_output_1_399(.a(output_2_399), .b(output_2_0), .y(output_1_399));
wire output_3_399, output_3_0, output_2_399;
mixer gate_output_2_399(.a(output_3_399), .b(output_3_0), .y(output_2_399));
wire output_4_399, output_4_0, output_3_399;
mixer gate_output_3_399(.a(output_4_399), .b(output_4_0), .y(output_3_399));
wire output_5_399, output_5_0, output_4_399;
mixer gate_output_4_399(.a(output_5_399), .b(output_5_0), .y(output_4_399));
wire output_6_399, output_6_0, output_5_399;
mixer gate_output_5_399(.a(output_6_399), .b(output_6_0), .y(output_5_399));
wire output_7_399, output_7_0, output_6_399;
mixer gate_output_6_399(.a(output_7_399), .b(output_7_0), .y(output_6_399));
wire output_8_399, output_8_0, output_7_399;
mixer gate_output_7_399(.a(output_8_399), .b(output_8_0), .y(output_7_399));
wire output_1_400, output_1_1, output_0_400;
mixer gate_output_0_400(.a(output_1_400), .b(output_1_1), .y(output_0_400));
wire output_2_400, output_2_1, output_1_400;
mixer gate_output_1_400(.a(output_2_400), .b(output_2_1), .y(output_1_400));
wire output_3_400, output_3_1, output_2_400;
mixer gate_output_2_400(.a(output_3_400), .b(output_3_1), .y(output_2_400));
wire output_4_400, output_4_1, output_3_400;
mixer gate_output_3_400(.a(output_4_400), .b(output_4_1), .y(output_3_400));
wire output_5_400, output_5_1, output_4_400;
mixer gate_output_4_400(.a(output_5_400), .b(output_5_1), .y(output_4_400));
wire output_6_400, output_6_1, output_5_400;
mixer gate_output_5_400(.a(output_6_400), .b(output_6_1), .y(output_5_400));
wire output_7_400, output_7_1, output_6_400;
mixer gate_output_6_400(.a(output_7_400), .b(output_7_1), .y(output_6_400));
wire output_8_400, output_8_1, output_7_400;
mixer gate_output_7_400(.a(output_8_400), .b(output_8_1), .y(output_7_400));
wire output_1_401, output_1_2, output_0_401;
mixer gate_output_0_401(.a(output_1_401), .b(output_1_2), .y(output_0_401));
wire output_2_401, output_2_2, output_1_401;
mixer gate_output_1_401(.a(output_2_401), .b(output_2_2), .y(output_1_401));
wire output_3_401, output_3_2, output_2_401;
mixer gate_output_2_401(.a(output_3_401), .b(output_3_2), .y(output_2_401));
wire output_4_401, output_4_2, output_3_401;
mixer gate_output_3_401(.a(output_4_401), .b(output_4_2), .y(output_3_401));
wire output_5_401, output_5_2, output_4_401;
mixer gate_output_4_401(.a(output_5_401), .b(output_5_2), .y(output_4_401));
wire output_6_401, output_6_2, output_5_401;
mixer gate_output_5_401(.a(output_6_401), .b(output_6_2), .y(output_5_401));
wire output_7_401, output_7_2, output_6_401;
mixer gate_output_6_401(.a(output_7_401), .b(output_7_2), .y(output_6_401));
wire output_8_401, output_8_2, output_7_401;
mixer gate_output_7_401(.a(output_8_401), .b(output_8_2), .y(output_7_401));
wire output_1_402, output_1_3, output_0_402;
mixer gate_output_0_402(.a(output_1_402), .b(output_1_3), .y(output_0_402));
wire output_2_402, output_2_3, output_1_402;
mixer gate_output_1_402(.a(output_2_402), .b(output_2_3), .y(output_1_402));
wire output_3_402, output_3_3, output_2_402;
mixer gate_output_2_402(.a(output_3_402), .b(output_3_3), .y(output_2_402));
wire output_4_402, output_4_3, output_3_402;
mixer gate_output_3_402(.a(output_4_402), .b(output_4_3), .y(output_3_402));
wire output_5_402, output_5_3, output_4_402;
mixer gate_output_4_402(.a(output_5_402), .b(output_5_3), .y(output_4_402));
wire output_6_402, output_6_3, output_5_402;
mixer gate_output_5_402(.a(output_6_402), .b(output_6_3), .y(output_5_402));
wire output_7_402, output_7_3, output_6_402;
mixer gate_output_6_402(.a(output_7_402), .b(output_7_3), .y(output_6_402));
wire output_8_402, output_8_3, output_7_402;
mixer gate_output_7_402(.a(output_8_402), .b(output_8_3), .y(output_7_402));
wire output_1_403, output_1_4, output_0_403;
mixer gate_output_0_403(.a(output_1_403), .b(output_1_4), .y(output_0_403));
wire output_2_403, output_2_4, output_1_403;
mixer gate_output_1_403(.a(output_2_403), .b(output_2_4), .y(output_1_403));
wire output_3_403, output_3_4, output_2_403;
mixer gate_output_2_403(.a(output_3_403), .b(output_3_4), .y(output_2_403));
wire output_4_403, output_4_4, output_3_403;
mixer gate_output_3_403(.a(output_4_403), .b(output_4_4), .y(output_3_403));
wire output_5_403, output_5_4, output_4_403;
mixer gate_output_4_403(.a(output_5_403), .b(output_5_4), .y(output_4_403));
wire output_6_403, output_6_4, output_5_403;
mixer gate_output_5_403(.a(output_6_403), .b(output_6_4), .y(output_5_403));
wire output_7_403, output_7_4, output_6_403;
mixer gate_output_6_403(.a(output_7_403), .b(output_7_4), .y(output_6_403));
wire output_8_403, output_8_4, output_7_403;
mixer gate_output_7_403(.a(output_8_403), .b(output_8_4), .y(output_7_403));
wire output_1_404, output_1_5, output_0_404;
mixer gate_output_0_404(.a(output_1_404), .b(output_1_5), .y(output_0_404));
wire output_2_404, output_2_5, output_1_404;
mixer gate_output_1_404(.a(output_2_404), .b(output_2_5), .y(output_1_404));
wire output_3_404, output_3_5, output_2_404;
mixer gate_output_2_404(.a(output_3_404), .b(output_3_5), .y(output_2_404));
wire output_4_404, output_4_5, output_3_404;
mixer gate_output_3_404(.a(output_4_404), .b(output_4_5), .y(output_3_404));
wire output_5_404, output_5_5, output_4_404;
mixer gate_output_4_404(.a(output_5_404), .b(output_5_5), .y(output_4_404));
wire output_6_404, output_6_5, output_5_404;
mixer gate_output_5_404(.a(output_6_404), .b(output_6_5), .y(output_5_404));
wire output_7_404, output_7_5, output_6_404;
mixer gate_output_6_404(.a(output_7_404), .b(output_7_5), .y(output_6_404));
wire output_8_404, output_8_5, output_7_404;
mixer gate_output_7_404(.a(output_8_404), .b(output_8_5), .y(output_7_404));
wire output_1_405, output_1_6, output_0_405;
mixer gate_output_0_405(.a(output_1_405), .b(output_1_6), .y(output_0_405));
wire output_2_405, output_2_6, output_1_405;
mixer gate_output_1_405(.a(output_2_405), .b(output_2_6), .y(output_1_405));
wire output_3_405, output_3_6, output_2_405;
mixer gate_output_2_405(.a(output_3_405), .b(output_3_6), .y(output_2_405));
wire output_4_405, output_4_6, output_3_405;
mixer gate_output_3_405(.a(output_4_405), .b(output_4_6), .y(output_3_405));
wire output_5_405, output_5_6, output_4_405;
mixer gate_output_4_405(.a(output_5_405), .b(output_5_6), .y(output_4_405));
wire output_6_405, output_6_6, output_5_405;
mixer gate_output_5_405(.a(output_6_405), .b(output_6_6), .y(output_5_405));
wire output_7_405, output_7_6, output_6_405;
mixer gate_output_6_405(.a(output_7_405), .b(output_7_6), .y(output_6_405));
wire output_8_405, output_8_6, output_7_405;
mixer gate_output_7_405(.a(output_8_405), .b(output_8_6), .y(output_7_405));
wire output_1_406, output_1_7, output_0_406;
mixer gate_output_0_406(.a(output_1_406), .b(output_1_7), .y(output_0_406));
wire output_2_406, output_2_7, output_1_406;
mixer gate_output_1_406(.a(output_2_406), .b(output_2_7), .y(output_1_406));
wire output_3_406, output_3_7, output_2_406;
mixer gate_output_2_406(.a(output_3_406), .b(output_3_7), .y(output_2_406));
wire output_4_406, output_4_7, output_3_406;
mixer gate_output_3_406(.a(output_4_406), .b(output_4_7), .y(output_3_406));
wire output_5_406, output_5_7, output_4_406;
mixer gate_output_4_406(.a(output_5_406), .b(output_5_7), .y(output_4_406));
wire output_6_406, output_6_7, output_5_406;
mixer gate_output_5_406(.a(output_6_406), .b(output_6_7), .y(output_5_406));
wire output_7_406, output_7_7, output_6_406;
mixer gate_output_6_406(.a(output_7_406), .b(output_7_7), .y(output_6_406));
wire output_8_406, output_8_7, output_7_406;
mixer gate_output_7_406(.a(output_8_406), .b(output_8_7), .y(output_7_406));
wire output_1_407, output_1_0, output_0_407;
mixer gate_output_0_407(.a(output_1_407), .b(output_1_0), .y(output_0_407));
wire output_2_407, output_2_0, output_1_407;
mixer gate_output_1_407(.a(output_2_407), .b(output_2_0), .y(output_1_407));
wire output_3_407, output_3_0, output_2_407;
mixer gate_output_2_407(.a(output_3_407), .b(output_3_0), .y(output_2_407));
wire output_4_407, output_4_0, output_3_407;
mixer gate_output_3_407(.a(output_4_407), .b(output_4_0), .y(output_3_407));
wire output_5_407, output_5_0, output_4_407;
mixer gate_output_4_407(.a(output_5_407), .b(output_5_0), .y(output_4_407));
wire output_6_407, output_6_0, output_5_407;
mixer gate_output_5_407(.a(output_6_407), .b(output_6_0), .y(output_5_407));
wire output_7_407, output_7_0, output_6_407;
mixer gate_output_6_407(.a(output_7_407), .b(output_7_0), .y(output_6_407));
wire output_8_407, output_8_0, output_7_407;
mixer gate_output_7_407(.a(output_8_407), .b(output_8_0), .y(output_7_407));
wire output_1_408, output_1_1, output_0_408;
mixer gate_output_0_408(.a(output_1_408), .b(output_1_1), .y(output_0_408));
wire output_2_408, output_2_1, output_1_408;
mixer gate_output_1_408(.a(output_2_408), .b(output_2_1), .y(output_1_408));
wire output_3_408, output_3_1, output_2_408;
mixer gate_output_2_408(.a(output_3_408), .b(output_3_1), .y(output_2_408));
wire output_4_408, output_4_1, output_3_408;
mixer gate_output_3_408(.a(output_4_408), .b(output_4_1), .y(output_3_408));
wire output_5_408, output_5_1, output_4_408;
mixer gate_output_4_408(.a(output_5_408), .b(output_5_1), .y(output_4_408));
wire output_6_408, output_6_1, output_5_408;
mixer gate_output_5_408(.a(output_6_408), .b(output_6_1), .y(output_5_408));
wire output_7_408, output_7_1, output_6_408;
mixer gate_output_6_408(.a(output_7_408), .b(output_7_1), .y(output_6_408));
wire output_8_408, output_8_1, output_7_408;
mixer gate_output_7_408(.a(output_8_408), .b(output_8_1), .y(output_7_408));
wire output_1_409, output_1_2, output_0_409;
mixer gate_output_0_409(.a(output_1_409), .b(output_1_2), .y(output_0_409));
wire output_2_409, output_2_2, output_1_409;
mixer gate_output_1_409(.a(output_2_409), .b(output_2_2), .y(output_1_409));
wire output_3_409, output_3_2, output_2_409;
mixer gate_output_2_409(.a(output_3_409), .b(output_3_2), .y(output_2_409));
wire output_4_409, output_4_2, output_3_409;
mixer gate_output_3_409(.a(output_4_409), .b(output_4_2), .y(output_3_409));
wire output_5_409, output_5_2, output_4_409;
mixer gate_output_4_409(.a(output_5_409), .b(output_5_2), .y(output_4_409));
wire output_6_409, output_6_2, output_5_409;
mixer gate_output_5_409(.a(output_6_409), .b(output_6_2), .y(output_5_409));
wire output_7_409, output_7_2, output_6_409;
mixer gate_output_6_409(.a(output_7_409), .b(output_7_2), .y(output_6_409));
wire output_8_409, output_8_2, output_7_409;
mixer gate_output_7_409(.a(output_8_409), .b(output_8_2), .y(output_7_409));
wire output_1_410, output_1_3, output_0_410;
mixer gate_output_0_410(.a(output_1_410), .b(output_1_3), .y(output_0_410));
wire output_2_410, output_2_3, output_1_410;
mixer gate_output_1_410(.a(output_2_410), .b(output_2_3), .y(output_1_410));
wire output_3_410, output_3_3, output_2_410;
mixer gate_output_2_410(.a(output_3_410), .b(output_3_3), .y(output_2_410));
wire output_4_410, output_4_3, output_3_410;
mixer gate_output_3_410(.a(output_4_410), .b(output_4_3), .y(output_3_410));
wire output_5_410, output_5_3, output_4_410;
mixer gate_output_4_410(.a(output_5_410), .b(output_5_3), .y(output_4_410));
wire output_6_410, output_6_3, output_5_410;
mixer gate_output_5_410(.a(output_6_410), .b(output_6_3), .y(output_5_410));
wire output_7_410, output_7_3, output_6_410;
mixer gate_output_6_410(.a(output_7_410), .b(output_7_3), .y(output_6_410));
wire output_8_410, output_8_3, output_7_410;
mixer gate_output_7_410(.a(output_8_410), .b(output_8_3), .y(output_7_410));
wire output_1_411, output_1_4, output_0_411;
mixer gate_output_0_411(.a(output_1_411), .b(output_1_4), .y(output_0_411));
wire output_2_411, output_2_4, output_1_411;
mixer gate_output_1_411(.a(output_2_411), .b(output_2_4), .y(output_1_411));
wire output_3_411, output_3_4, output_2_411;
mixer gate_output_2_411(.a(output_3_411), .b(output_3_4), .y(output_2_411));
wire output_4_411, output_4_4, output_3_411;
mixer gate_output_3_411(.a(output_4_411), .b(output_4_4), .y(output_3_411));
wire output_5_411, output_5_4, output_4_411;
mixer gate_output_4_411(.a(output_5_411), .b(output_5_4), .y(output_4_411));
wire output_6_411, output_6_4, output_5_411;
mixer gate_output_5_411(.a(output_6_411), .b(output_6_4), .y(output_5_411));
wire output_7_411, output_7_4, output_6_411;
mixer gate_output_6_411(.a(output_7_411), .b(output_7_4), .y(output_6_411));
wire output_8_411, output_8_4, output_7_411;
mixer gate_output_7_411(.a(output_8_411), .b(output_8_4), .y(output_7_411));
wire output_1_412, output_1_5, output_0_412;
mixer gate_output_0_412(.a(output_1_412), .b(output_1_5), .y(output_0_412));
wire output_2_412, output_2_5, output_1_412;
mixer gate_output_1_412(.a(output_2_412), .b(output_2_5), .y(output_1_412));
wire output_3_412, output_3_5, output_2_412;
mixer gate_output_2_412(.a(output_3_412), .b(output_3_5), .y(output_2_412));
wire output_4_412, output_4_5, output_3_412;
mixer gate_output_3_412(.a(output_4_412), .b(output_4_5), .y(output_3_412));
wire output_5_412, output_5_5, output_4_412;
mixer gate_output_4_412(.a(output_5_412), .b(output_5_5), .y(output_4_412));
wire output_6_412, output_6_5, output_5_412;
mixer gate_output_5_412(.a(output_6_412), .b(output_6_5), .y(output_5_412));
wire output_7_412, output_7_5, output_6_412;
mixer gate_output_6_412(.a(output_7_412), .b(output_7_5), .y(output_6_412));
wire output_8_412, output_8_5, output_7_412;
mixer gate_output_7_412(.a(output_8_412), .b(output_8_5), .y(output_7_412));
wire output_1_413, output_1_6, output_0_413;
mixer gate_output_0_413(.a(output_1_413), .b(output_1_6), .y(output_0_413));
wire output_2_413, output_2_6, output_1_413;
mixer gate_output_1_413(.a(output_2_413), .b(output_2_6), .y(output_1_413));
wire output_3_413, output_3_6, output_2_413;
mixer gate_output_2_413(.a(output_3_413), .b(output_3_6), .y(output_2_413));
wire output_4_413, output_4_6, output_3_413;
mixer gate_output_3_413(.a(output_4_413), .b(output_4_6), .y(output_3_413));
wire output_5_413, output_5_6, output_4_413;
mixer gate_output_4_413(.a(output_5_413), .b(output_5_6), .y(output_4_413));
wire output_6_413, output_6_6, output_5_413;
mixer gate_output_5_413(.a(output_6_413), .b(output_6_6), .y(output_5_413));
wire output_7_413, output_7_6, output_6_413;
mixer gate_output_6_413(.a(output_7_413), .b(output_7_6), .y(output_6_413));
wire output_8_413, output_8_6, output_7_413;
mixer gate_output_7_413(.a(output_8_413), .b(output_8_6), .y(output_7_413));
wire output_1_414, output_1_7, output_0_414;
mixer gate_output_0_414(.a(output_1_414), .b(output_1_7), .y(output_0_414));
wire output_2_414, output_2_7, output_1_414;
mixer gate_output_1_414(.a(output_2_414), .b(output_2_7), .y(output_1_414));
wire output_3_414, output_3_7, output_2_414;
mixer gate_output_2_414(.a(output_3_414), .b(output_3_7), .y(output_2_414));
wire output_4_414, output_4_7, output_3_414;
mixer gate_output_3_414(.a(output_4_414), .b(output_4_7), .y(output_3_414));
wire output_5_414, output_5_7, output_4_414;
mixer gate_output_4_414(.a(output_5_414), .b(output_5_7), .y(output_4_414));
wire output_6_414, output_6_7, output_5_414;
mixer gate_output_5_414(.a(output_6_414), .b(output_6_7), .y(output_5_414));
wire output_7_414, output_7_7, output_6_414;
mixer gate_output_6_414(.a(output_7_414), .b(output_7_7), .y(output_6_414));
wire output_8_414, output_8_7, output_7_414;
mixer gate_output_7_414(.a(output_8_414), .b(output_8_7), .y(output_7_414));
wire output_1_415, output_1_0, output_0_415;
mixer gate_output_0_415(.a(output_1_415), .b(output_1_0), .y(output_0_415));
wire output_2_415, output_2_0, output_1_415;
mixer gate_output_1_415(.a(output_2_415), .b(output_2_0), .y(output_1_415));
wire output_3_415, output_3_0, output_2_415;
mixer gate_output_2_415(.a(output_3_415), .b(output_3_0), .y(output_2_415));
wire output_4_415, output_4_0, output_3_415;
mixer gate_output_3_415(.a(output_4_415), .b(output_4_0), .y(output_3_415));
wire output_5_415, output_5_0, output_4_415;
mixer gate_output_4_415(.a(output_5_415), .b(output_5_0), .y(output_4_415));
wire output_6_415, output_6_0, output_5_415;
mixer gate_output_5_415(.a(output_6_415), .b(output_6_0), .y(output_5_415));
wire output_7_415, output_7_0, output_6_415;
mixer gate_output_6_415(.a(output_7_415), .b(output_7_0), .y(output_6_415));
wire output_8_415, output_8_0, output_7_415;
mixer gate_output_7_415(.a(output_8_415), .b(output_8_0), .y(output_7_415));
wire output_1_416, output_1_1, output_0_416;
mixer gate_output_0_416(.a(output_1_416), .b(output_1_1), .y(output_0_416));
wire output_2_416, output_2_1, output_1_416;
mixer gate_output_1_416(.a(output_2_416), .b(output_2_1), .y(output_1_416));
wire output_3_416, output_3_1, output_2_416;
mixer gate_output_2_416(.a(output_3_416), .b(output_3_1), .y(output_2_416));
wire output_4_416, output_4_1, output_3_416;
mixer gate_output_3_416(.a(output_4_416), .b(output_4_1), .y(output_3_416));
wire output_5_416, output_5_1, output_4_416;
mixer gate_output_4_416(.a(output_5_416), .b(output_5_1), .y(output_4_416));
wire output_6_416, output_6_1, output_5_416;
mixer gate_output_5_416(.a(output_6_416), .b(output_6_1), .y(output_5_416));
wire output_7_416, output_7_1, output_6_416;
mixer gate_output_6_416(.a(output_7_416), .b(output_7_1), .y(output_6_416));
wire output_8_416, output_8_1, output_7_416;
mixer gate_output_7_416(.a(output_8_416), .b(output_8_1), .y(output_7_416));
wire output_1_417, output_1_2, output_0_417;
mixer gate_output_0_417(.a(output_1_417), .b(output_1_2), .y(output_0_417));
wire output_2_417, output_2_2, output_1_417;
mixer gate_output_1_417(.a(output_2_417), .b(output_2_2), .y(output_1_417));
wire output_3_417, output_3_2, output_2_417;
mixer gate_output_2_417(.a(output_3_417), .b(output_3_2), .y(output_2_417));
wire output_4_417, output_4_2, output_3_417;
mixer gate_output_3_417(.a(output_4_417), .b(output_4_2), .y(output_3_417));
wire output_5_417, output_5_2, output_4_417;
mixer gate_output_4_417(.a(output_5_417), .b(output_5_2), .y(output_4_417));
wire output_6_417, output_6_2, output_5_417;
mixer gate_output_5_417(.a(output_6_417), .b(output_6_2), .y(output_5_417));
wire output_7_417, output_7_2, output_6_417;
mixer gate_output_6_417(.a(output_7_417), .b(output_7_2), .y(output_6_417));
wire output_8_417, output_8_2, output_7_417;
mixer gate_output_7_417(.a(output_8_417), .b(output_8_2), .y(output_7_417));
wire output_1_418, output_1_3, output_0_418;
mixer gate_output_0_418(.a(output_1_418), .b(output_1_3), .y(output_0_418));
wire output_2_418, output_2_3, output_1_418;
mixer gate_output_1_418(.a(output_2_418), .b(output_2_3), .y(output_1_418));
wire output_3_418, output_3_3, output_2_418;
mixer gate_output_2_418(.a(output_3_418), .b(output_3_3), .y(output_2_418));
wire output_4_418, output_4_3, output_3_418;
mixer gate_output_3_418(.a(output_4_418), .b(output_4_3), .y(output_3_418));
wire output_5_418, output_5_3, output_4_418;
mixer gate_output_4_418(.a(output_5_418), .b(output_5_3), .y(output_4_418));
wire output_6_418, output_6_3, output_5_418;
mixer gate_output_5_418(.a(output_6_418), .b(output_6_3), .y(output_5_418));
wire output_7_418, output_7_3, output_6_418;
mixer gate_output_6_418(.a(output_7_418), .b(output_7_3), .y(output_6_418));
wire output_8_418, output_8_3, output_7_418;
mixer gate_output_7_418(.a(output_8_418), .b(output_8_3), .y(output_7_418));
wire output_1_419, output_1_4, output_0_419;
mixer gate_output_0_419(.a(output_1_419), .b(output_1_4), .y(output_0_419));
wire output_2_419, output_2_4, output_1_419;
mixer gate_output_1_419(.a(output_2_419), .b(output_2_4), .y(output_1_419));
wire output_3_419, output_3_4, output_2_419;
mixer gate_output_2_419(.a(output_3_419), .b(output_3_4), .y(output_2_419));
wire output_4_419, output_4_4, output_3_419;
mixer gate_output_3_419(.a(output_4_419), .b(output_4_4), .y(output_3_419));
wire output_5_419, output_5_4, output_4_419;
mixer gate_output_4_419(.a(output_5_419), .b(output_5_4), .y(output_4_419));
wire output_6_419, output_6_4, output_5_419;
mixer gate_output_5_419(.a(output_6_419), .b(output_6_4), .y(output_5_419));
wire output_7_419, output_7_4, output_6_419;
mixer gate_output_6_419(.a(output_7_419), .b(output_7_4), .y(output_6_419));
wire output_8_419, output_8_4, output_7_419;
mixer gate_output_7_419(.a(output_8_419), .b(output_8_4), .y(output_7_419));
wire output_1_420, output_1_5, output_0_420;
mixer gate_output_0_420(.a(output_1_420), .b(output_1_5), .y(output_0_420));
wire output_2_420, output_2_5, output_1_420;
mixer gate_output_1_420(.a(output_2_420), .b(output_2_5), .y(output_1_420));
wire output_3_420, output_3_5, output_2_420;
mixer gate_output_2_420(.a(output_3_420), .b(output_3_5), .y(output_2_420));
wire output_4_420, output_4_5, output_3_420;
mixer gate_output_3_420(.a(output_4_420), .b(output_4_5), .y(output_3_420));
wire output_5_420, output_5_5, output_4_420;
mixer gate_output_4_420(.a(output_5_420), .b(output_5_5), .y(output_4_420));
wire output_6_420, output_6_5, output_5_420;
mixer gate_output_5_420(.a(output_6_420), .b(output_6_5), .y(output_5_420));
wire output_7_420, output_7_5, output_6_420;
mixer gate_output_6_420(.a(output_7_420), .b(output_7_5), .y(output_6_420));
wire output_8_420, output_8_5, output_7_420;
mixer gate_output_7_420(.a(output_8_420), .b(output_8_5), .y(output_7_420));
wire output_1_421, output_1_6, output_0_421;
mixer gate_output_0_421(.a(output_1_421), .b(output_1_6), .y(output_0_421));
wire output_2_421, output_2_6, output_1_421;
mixer gate_output_1_421(.a(output_2_421), .b(output_2_6), .y(output_1_421));
wire output_3_421, output_3_6, output_2_421;
mixer gate_output_2_421(.a(output_3_421), .b(output_3_6), .y(output_2_421));
wire output_4_421, output_4_6, output_3_421;
mixer gate_output_3_421(.a(output_4_421), .b(output_4_6), .y(output_3_421));
wire output_5_421, output_5_6, output_4_421;
mixer gate_output_4_421(.a(output_5_421), .b(output_5_6), .y(output_4_421));
wire output_6_421, output_6_6, output_5_421;
mixer gate_output_5_421(.a(output_6_421), .b(output_6_6), .y(output_5_421));
wire output_7_421, output_7_6, output_6_421;
mixer gate_output_6_421(.a(output_7_421), .b(output_7_6), .y(output_6_421));
wire output_8_421, output_8_6, output_7_421;
mixer gate_output_7_421(.a(output_8_421), .b(output_8_6), .y(output_7_421));
wire output_1_422, output_1_7, output_0_422;
mixer gate_output_0_422(.a(output_1_422), .b(output_1_7), .y(output_0_422));
wire output_2_422, output_2_7, output_1_422;
mixer gate_output_1_422(.a(output_2_422), .b(output_2_7), .y(output_1_422));
wire output_3_422, output_3_7, output_2_422;
mixer gate_output_2_422(.a(output_3_422), .b(output_3_7), .y(output_2_422));
wire output_4_422, output_4_7, output_3_422;
mixer gate_output_3_422(.a(output_4_422), .b(output_4_7), .y(output_3_422));
wire output_5_422, output_5_7, output_4_422;
mixer gate_output_4_422(.a(output_5_422), .b(output_5_7), .y(output_4_422));
wire output_6_422, output_6_7, output_5_422;
mixer gate_output_5_422(.a(output_6_422), .b(output_6_7), .y(output_5_422));
wire output_7_422, output_7_7, output_6_422;
mixer gate_output_6_422(.a(output_7_422), .b(output_7_7), .y(output_6_422));
wire output_8_422, output_8_7, output_7_422;
mixer gate_output_7_422(.a(output_8_422), .b(output_8_7), .y(output_7_422));
wire output_1_423, output_1_0, output_0_423;
mixer gate_output_0_423(.a(output_1_423), .b(output_1_0), .y(output_0_423));
wire output_2_423, output_2_0, output_1_423;
mixer gate_output_1_423(.a(output_2_423), .b(output_2_0), .y(output_1_423));
wire output_3_423, output_3_0, output_2_423;
mixer gate_output_2_423(.a(output_3_423), .b(output_3_0), .y(output_2_423));
wire output_4_423, output_4_0, output_3_423;
mixer gate_output_3_423(.a(output_4_423), .b(output_4_0), .y(output_3_423));
wire output_5_423, output_5_0, output_4_423;
mixer gate_output_4_423(.a(output_5_423), .b(output_5_0), .y(output_4_423));
wire output_6_423, output_6_0, output_5_423;
mixer gate_output_5_423(.a(output_6_423), .b(output_6_0), .y(output_5_423));
wire output_7_423, output_7_0, output_6_423;
mixer gate_output_6_423(.a(output_7_423), .b(output_7_0), .y(output_6_423));
wire output_8_423, output_8_0, output_7_423;
mixer gate_output_7_423(.a(output_8_423), .b(output_8_0), .y(output_7_423));
wire output_1_424, output_1_1, output_0_424;
mixer gate_output_0_424(.a(output_1_424), .b(output_1_1), .y(output_0_424));
wire output_2_424, output_2_1, output_1_424;
mixer gate_output_1_424(.a(output_2_424), .b(output_2_1), .y(output_1_424));
wire output_3_424, output_3_1, output_2_424;
mixer gate_output_2_424(.a(output_3_424), .b(output_3_1), .y(output_2_424));
wire output_4_424, output_4_1, output_3_424;
mixer gate_output_3_424(.a(output_4_424), .b(output_4_1), .y(output_3_424));
wire output_5_424, output_5_1, output_4_424;
mixer gate_output_4_424(.a(output_5_424), .b(output_5_1), .y(output_4_424));
wire output_6_424, output_6_1, output_5_424;
mixer gate_output_5_424(.a(output_6_424), .b(output_6_1), .y(output_5_424));
wire output_7_424, output_7_1, output_6_424;
mixer gate_output_6_424(.a(output_7_424), .b(output_7_1), .y(output_6_424));
wire output_8_424, output_8_1, output_7_424;
mixer gate_output_7_424(.a(output_8_424), .b(output_8_1), .y(output_7_424));
wire output_1_425, output_1_2, output_0_425;
mixer gate_output_0_425(.a(output_1_425), .b(output_1_2), .y(output_0_425));
wire output_2_425, output_2_2, output_1_425;
mixer gate_output_1_425(.a(output_2_425), .b(output_2_2), .y(output_1_425));
wire output_3_425, output_3_2, output_2_425;
mixer gate_output_2_425(.a(output_3_425), .b(output_3_2), .y(output_2_425));
wire output_4_425, output_4_2, output_3_425;
mixer gate_output_3_425(.a(output_4_425), .b(output_4_2), .y(output_3_425));
wire output_5_425, output_5_2, output_4_425;
mixer gate_output_4_425(.a(output_5_425), .b(output_5_2), .y(output_4_425));
wire output_6_425, output_6_2, output_5_425;
mixer gate_output_5_425(.a(output_6_425), .b(output_6_2), .y(output_5_425));
wire output_7_425, output_7_2, output_6_425;
mixer gate_output_6_425(.a(output_7_425), .b(output_7_2), .y(output_6_425));
wire output_8_425, output_8_2, output_7_425;
mixer gate_output_7_425(.a(output_8_425), .b(output_8_2), .y(output_7_425));
wire output_1_426, output_1_3, output_0_426;
mixer gate_output_0_426(.a(output_1_426), .b(output_1_3), .y(output_0_426));
wire output_2_426, output_2_3, output_1_426;
mixer gate_output_1_426(.a(output_2_426), .b(output_2_3), .y(output_1_426));
wire output_3_426, output_3_3, output_2_426;
mixer gate_output_2_426(.a(output_3_426), .b(output_3_3), .y(output_2_426));
wire output_4_426, output_4_3, output_3_426;
mixer gate_output_3_426(.a(output_4_426), .b(output_4_3), .y(output_3_426));
wire output_5_426, output_5_3, output_4_426;
mixer gate_output_4_426(.a(output_5_426), .b(output_5_3), .y(output_4_426));
wire output_6_426, output_6_3, output_5_426;
mixer gate_output_5_426(.a(output_6_426), .b(output_6_3), .y(output_5_426));
wire output_7_426, output_7_3, output_6_426;
mixer gate_output_6_426(.a(output_7_426), .b(output_7_3), .y(output_6_426));
wire output_8_426, output_8_3, output_7_426;
mixer gate_output_7_426(.a(output_8_426), .b(output_8_3), .y(output_7_426));
wire output_1_427, output_1_4, output_0_427;
mixer gate_output_0_427(.a(output_1_427), .b(output_1_4), .y(output_0_427));
wire output_2_427, output_2_4, output_1_427;
mixer gate_output_1_427(.a(output_2_427), .b(output_2_4), .y(output_1_427));
wire output_3_427, output_3_4, output_2_427;
mixer gate_output_2_427(.a(output_3_427), .b(output_3_4), .y(output_2_427));
wire output_4_427, output_4_4, output_3_427;
mixer gate_output_3_427(.a(output_4_427), .b(output_4_4), .y(output_3_427));
wire output_5_427, output_5_4, output_4_427;
mixer gate_output_4_427(.a(output_5_427), .b(output_5_4), .y(output_4_427));
wire output_6_427, output_6_4, output_5_427;
mixer gate_output_5_427(.a(output_6_427), .b(output_6_4), .y(output_5_427));
wire output_7_427, output_7_4, output_6_427;
mixer gate_output_6_427(.a(output_7_427), .b(output_7_4), .y(output_6_427));
wire output_8_427, output_8_4, output_7_427;
mixer gate_output_7_427(.a(output_8_427), .b(output_8_4), .y(output_7_427));
wire output_1_428, output_1_5, output_0_428;
mixer gate_output_0_428(.a(output_1_428), .b(output_1_5), .y(output_0_428));
wire output_2_428, output_2_5, output_1_428;
mixer gate_output_1_428(.a(output_2_428), .b(output_2_5), .y(output_1_428));
wire output_3_428, output_3_5, output_2_428;
mixer gate_output_2_428(.a(output_3_428), .b(output_3_5), .y(output_2_428));
wire output_4_428, output_4_5, output_3_428;
mixer gate_output_3_428(.a(output_4_428), .b(output_4_5), .y(output_3_428));
wire output_5_428, output_5_5, output_4_428;
mixer gate_output_4_428(.a(output_5_428), .b(output_5_5), .y(output_4_428));
wire output_6_428, output_6_5, output_5_428;
mixer gate_output_5_428(.a(output_6_428), .b(output_6_5), .y(output_5_428));
wire output_7_428, output_7_5, output_6_428;
mixer gate_output_6_428(.a(output_7_428), .b(output_7_5), .y(output_6_428));
wire output_8_428, output_8_5, output_7_428;
mixer gate_output_7_428(.a(output_8_428), .b(output_8_5), .y(output_7_428));
wire output_1_429, output_1_6, output_0_429;
mixer gate_output_0_429(.a(output_1_429), .b(output_1_6), .y(output_0_429));
wire output_2_429, output_2_6, output_1_429;
mixer gate_output_1_429(.a(output_2_429), .b(output_2_6), .y(output_1_429));
wire output_3_429, output_3_6, output_2_429;
mixer gate_output_2_429(.a(output_3_429), .b(output_3_6), .y(output_2_429));
wire output_4_429, output_4_6, output_3_429;
mixer gate_output_3_429(.a(output_4_429), .b(output_4_6), .y(output_3_429));
wire output_5_429, output_5_6, output_4_429;
mixer gate_output_4_429(.a(output_5_429), .b(output_5_6), .y(output_4_429));
wire output_6_429, output_6_6, output_5_429;
mixer gate_output_5_429(.a(output_6_429), .b(output_6_6), .y(output_5_429));
wire output_7_429, output_7_6, output_6_429;
mixer gate_output_6_429(.a(output_7_429), .b(output_7_6), .y(output_6_429));
wire output_8_429, output_8_6, output_7_429;
mixer gate_output_7_429(.a(output_8_429), .b(output_8_6), .y(output_7_429));
wire output_1_430, output_1_7, output_0_430;
mixer gate_output_0_430(.a(output_1_430), .b(output_1_7), .y(output_0_430));
wire output_2_430, output_2_7, output_1_430;
mixer gate_output_1_430(.a(output_2_430), .b(output_2_7), .y(output_1_430));
wire output_3_430, output_3_7, output_2_430;
mixer gate_output_2_430(.a(output_3_430), .b(output_3_7), .y(output_2_430));
wire output_4_430, output_4_7, output_3_430;
mixer gate_output_3_430(.a(output_4_430), .b(output_4_7), .y(output_3_430));
wire output_5_430, output_5_7, output_4_430;
mixer gate_output_4_430(.a(output_5_430), .b(output_5_7), .y(output_4_430));
wire output_6_430, output_6_7, output_5_430;
mixer gate_output_5_430(.a(output_6_430), .b(output_6_7), .y(output_5_430));
wire output_7_430, output_7_7, output_6_430;
mixer gate_output_6_430(.a(output_7_430), .b(output_7_7), .y(output_6_430));
wire output_8_430, output_8_7, output_7_430;
mixer gate_output_7_430(.a(output_8_430), .b(output_8_7), .y(output_7_430));
wire output_1_431, output_1_0, output_0_431;
mixer gate_output_0_431(.a(output_1_431), .b(output_1_0), .y(output_0_431));
wire output_2_431, output_2_0, output_1_431;
mixer gate_output_1_431(.a(output_2_431), .b(output_2_0), .y(output_1_431));
wire output_3_431, output_3_0, output_2_431;
mixer gate_output_2_431(.a(output_3_431), .b(output_3_0), .y(output_2_431));
wire output_4_431, output_4_0, output_3_431;
mixer gate_output_3_431(.a(output_4_431), .b(output_4_0), .y(output_3_431));
wire output_5_431, output_5_0, output_4_431;
mixer gate_output_4_431(.a(output_5_431), .b(output_5_0), .y(output_4_431));
wire output_6_431, output_6_0, output_5_431;
mixer gate_output_5_431(.a(output_6_431), .b(output_6_0), .y(output_5_431));
wire output_7_431, output_7_0, output_6_431;
mixer gate_output_6_431(.a(output_7_431), .b(output_7_0), .y(output_6_431));
wire output_8_431, output_8_0, output_7_431;
mixer gate_output_7_431(.a(output_8_431), .b(output_8_0), .y(output_7_431));
wire output_1_432, output_1_1, output_0_432;
mixer gate_output_0_432(.a(output_1_432), .b(output_1_1), .y(output_0_432));
wire output_2_432, output_2_1, output_1_432;
mixer gate_output_1_432(.a(output_2_432), .b(output_2_1), .y(output_1_432));
wire output_3_432, output_3_1, output_2_432;
mixer gate_output_2_432(.a(output_3_432), .b(output_3_1), .y(output_2_432));
wire output_4_432, output_4_1, output_3_432;
mixer gate_output_3_432(.a(output_4_432), .b(output_4_1), .y(output_3_432));
wire output_5_432, output_5_1, output_4_432;
mixer gate_output_4_432(.a(output_5_432), .b(output_5_1), .y(output_4_432));
wire output_6_432, output_6_1, output_5_432;
mixer gate_output_5_432(.a(output_6_432), .b(output_6_1), .y(output_5_432));
wire output_7_432, output_7_1, output_6_432;
mixer gate_output_6_432(.a(output_7_432), .b(output_7_1), .y(output_6_432));
wire output_8_432, output_8_1, output_7_432;
mixer gate_output_7_432(.a(output_8_432), .b(output_8_1), .y(output_7_432));
wire output_1_433, output_1_2, output_0_433;
mixer gate_output_0_433(.a(output_1_433), .b(output_1_2), .y(output_0_433));
wire output_2_433, output_2_2, output_1_433;
mixer gate_output_1_433(.a(output_2_433), .b(output_2_2), .y(output_1_433));
wire output_3_433, output_3_2, output_2_433;
mixer gate_output_2_433(.a(output_3_433), .b(output_3_2), .y(output_2_433));
wire output_4_433, output_4_2, output_3_433;
mixer gate_output_3_433(.a(output_4_433), .b(output_4_2), .y(output_3_433));
wire output_5_433, output_5_2, output_4_433;
mixer gate_output_4_433(.a(output_5_433), .b(output_5_2), .y(output_4_433));
wire output_6_433, output_6_2, output_5_433;
mixer gate_output_5_433(.a(output_6_433), .b(output_6_2), .y(output_5_433));
wire output_7_433, output_7_2, output_6_433;
mixer gate_output_6_433(.a(output_7_433), .b(output_7_2), .y(output_6_433));
wire output_8_433, output_8_2, output_7_433;
mixer gate_output_7_433(.a(output_8_433), .b(output_8_2), .y(output_7_433));
wire output_1_434, output_1_3, output_0_434;
mixer gate_output_0_434(.a(output_1_434), .b(output_1_3), .y(output_0_434));
wire output_2_434, output_2_3, output_1_434;
mixer gate_output_1_434(.a(output_2_434), .b(output_2_3), .y(output_1_434));
wire output_3_434, output_3_3, output_2_434;
mixer gate_output_2_434(.a(output_3_434), .b(output_3_3), .y(output_2_434));
wire output_4_434, output_4_3, output_3_434;
mixer gate_output_3_434(.a(output_4_434), .b(output_4_3), .y(output_3_434));
wire output_5_434, output_5_3, output_4_434;
mixer gate_output_4_434(.a(output_5_434), .b(output_5_3), .y(output_4_434));
wire output_6_434, output_6_3, output_5_434;
mixer gate_output_5_434(.a(output_6_434), .b(output_6_3), .y(output_5_434));
wire output_7_434, output_7_3, output_6_434;
mixer gate_output_6_434(.a(output_7_434), .b(output_7_3), .y(output_6_434));
wire output_8_434, output_8_3, output_7_434;
mixer gate_output_7_434(.a(output_8_434), .b(output_8_3), .y(output_7_434));
wire output_1_435, output_1_4, output_0_435;
mixer gate_output_0_435(.a(output_1_435), .b(output_1_4), .y(output_0_435));
wire output_2_435, output_2_4, output_1_435;
mixer gate_output_1_435(.a(output_2_435), .b(output_2_4), .y(output_1_435));
wire output_3_435, output_3_4, output_2_435;
mixer gate_output_2_435(.a(output_3_435), .b(output_3_4), .y(output_2_435));
wire output_4_435, output_4_4, output_3_435;
mixer gate_output_3_435(.a(output_4_435), .b(output_4_4), .y(output_3_435));
wire output_5_435, output_5_4, output_4_435;
mixer gate_output_4_435(.a(output_5_435), .b(output_5_4), .y(output_4_435));
wire output_6_435, output_6_4, output_5_435;
mixer gate_output_5_435(.a(output_6_435), .b(output_6_4), .y(output_5_435));
wire output_7_435, output_7_4, output_6_435;
mixer gate_output_6_435(.a(output_7_435), .b(output_7_4), .y(output_6_435));
wire output_8_435, output_8_4, output_7_435;
mixer gate_output_7_435(.a(output_8_435), .b(output_8_4), .y(output_7_435));
wire output_1_436, output_1_5, output_0_436;
mixer gate_output_0_436(.a(output_1_436), .b(output_1_5), .y(output_0_436));
wire output_2_436, output_2_5, output_1_436;
mixer gate_output_1_436(.a(output_2_436), .b(output_2_5), .y(output_1_436));
wire output_3_436, output_3_5, output_2_436;
mixer gate_output_2_436(.a(output_3_436), .b(output_3_5), .y(output_2_436));
wire output_4_436, output_4_5, output_3_436;
mixer gate_output_3_436(.a(output_4_436), .b(output_4_5), .y(output_3_436));
wire output_5_436, output_5_5, output_4_436;
mixer gate_output_4_436(.a(output_5_436), .b(output_5_5), .y(output_4_436));
wire output_6_436, output_6_5, output_5_436;
mixer gate_output_5_436(.a(output_6_436), .b(output_6_5), .y(output_5_436));
wire output_7_436, output_7_5, output_6_436;
mixer gate_output_6_436(.a(output_7_436), .b(output_7_5), .y(output_6_436));
wire output_8_436, output_8_5, output_7_436;
mixer gate_output_7_436(.a(output_8_436), .b(output_8_5), .y(output_7_436));
wire output_1_437, output_1_6, output_0_437;
mixer gate_output_0_437(.a(output_1_437), .b(output_1_6), .y(output_0_437));
wire output_2_437, output_2_6, output_1_437;
mixer gate_output_1_437(.a(output_2_437), .b(output_2_6), .y(output_1_437));
wire output_3_437, output_3_6, output_2_437;
mixer gate_output_2_437(.a(output_3_437), .b(output_3_6), .y(output_2_437));
wire output_4_437, output_4_6, output_3_437;
mixer gate_output_3_437(.a(output_4_437), .b(output_4_6), .y(output_3_437));
wire output_5_437, output_5_6, output_4_437;
mixer gate_output_4_437(.a(output_5_437), .b(output_5_6), .y(output_4_437));
wire output_6_437, output_6_6, output_5_437;
mixer gate_output_5_437(.a(output_6_437), .b(output_6_6), .y(output_5_437));
wire output_7_437, output_7_6, output_6_437;
mixer gate_output_6_437(.a(output_7_437), .b(output_7_6), .y(output_6_437));
wire output_8_437, output_8_6, output_7_437;
mixer gate_output_7_437(.a(output_8_437), .b(output_8_6), .y(output_7_437));
wire output_1_438, output_1_7, output_0_438;
mixer gate_output_0_438(.a(output_1_438), .b(output_1_7), .y(output_0_438));
wire output_2_438, output_2_7, output_1_438;
mixer gate_output_1_438(.a(output_2_438), .b(output_2_7), .y(output_1_438));
wire output_3_438, output_3_7, output_2_438;
mixer gate_output_2_438(.a(output_3_438), .b(output_3_7), .y(output_2_438));
wire output_4_438, output_4_7, output_3_438;
mixer gate_output_3_438(.a(output_4_438), .b(output_4_7), .y(output_3_438));
wire output_5_438, output_5_7, output_4_438;
mixer gate_output_4_438(.a(output_5_438), .b(output_5_7), .y(output_4_438));
wire output_6_438, output_6_7, output_5_438;
mixer gate_output_5_438(.a(output_6_438), .b(output_6_7), .y(output_5_438));
wire output_7_438, output_7_7, output_6_438;
mixer gate_output_6_438(.a(output_7_438), .b(output_7_7), .y(output_6_438));
wire output_8_438, output_8_7, output_7_438;
mixer gate_output_7_438(.a(output_8_438), .b(output_8_7), .y(output_7_438));
wire output_1_439, output_1_0, output_0_439;
mixer gate_output_0_439(.a(output_1_439), .b(output_1_0), .y(output_0_439));
wire output_2_439, output_2_0, output_1_439;
mixer gate_output_1_439(.a(output_2_439), .b(output_2_0), .y(output_1_439));
wire output_3_439, output_3_0, output_2_439;
mixer gate_output_2_439(.a(output_3_439), .b(output_3_0), .y(output_2_439));
wire output_4_439, output_4_0, output_3_439;
mixer gate_output_3_439(.a(output_4_439), .b(output_4_0), .y(output_3_439));
wire output_5_439, output_5_0, output_4_439;
mixer gate_output_4_439(.a(output_5_439), .b(output_5_0), .y(output_4_439));
wire output_6_439, output_6_0, output_5_439;
mixer gate_output_5_439(.a(output_6_439), .b(output_6_0), .y(output_5_439));
wire output_7_439, output_7_0, output_6_439;
mixer gate_output_6_439(.a(output_7_439), .b(output_7_0), .y(output_6_439));
wire output_8_439, output_8_0, output_7_439;
mixer gate_output_7_439(.a(output_8_439), .b(output_8_0), .y(output_7_439));
wire output_1_440, output_1_1, output_0_440;
mixer gate_output_0_440(.a(output_1_440), .b(output_1_1), .y(output_0_440));
wire output_2_440, output_2_1, output_1_440;
mixer gate_output_1_440(.a(output_2_440), .b(output_2_1), .y(output_1_440));
wire output_3_440, output_3_1, output_2_440;
mixer gate_output_2_440(.a(output_3_440), .b(output_3_1), .y(output_2_440));
wire output_4_440, output_4_1, output_3_440;
mixer gate_output_3_440(.a(output_4_440), .b(output_4_1), .y(output_3_440));
wire output_5_440, output_5_1, output_4_440;
mixer gate_output_4_440(.a(output_5_440), .b(output_5_1), .y(output_4_440));
wire output_6_440, output_6_1, output_5_440;
mixer gate_output_5_440(.a(output_6_440), .b(output_6_1), .y(output_5_440));
wire output_7_440, output_7_1, output_6_440;
mixer gate_output_6_440(.a(output_7_440), .b(output_7_1), .y(output_6_440));
wire output_8_440, output_8_1, output_7_440;
mixer gate_output_7_440(.a(output_8_440), .b(output_8_1), .y(output_7_440));
wire output_1_441, output_1_2, output_0_441;
mixer gate_output_0_441(.a(output_1_441), .b(output_1_2), .y(output_0_441));
wire output_2_441, output_2_2, output_1_441;
mixer gate_output_1_441(.a(output_2_441), .b(output_2_2), .y(output_1_441));
wire output_3_441, output_3_2, output_2_441;
mixer gate_output_2_441(.a(output_3_441), .b(output_3_2), .y(output_2_441));
wire output_4_441, output_4_2, output_3_441;
mixer gate_output_3_441(.a(output_4_441), .b(output_4_2), .y(output_3_441));
wire output_5_441, output_5_2, output_4_441;
mixer gate_output_4_441(.a(output_5_441), .b(output_5_2), .y(output_4_441));
wire output_6_441, output_6_2, output_5_441;
mixer gate_output_5_441(.a(output_6_441), .b(output_6_2), .y(output_5_441));
wire output_7_441, output_7_2, output_6_441;
mixer gate_output_6_441(.a(output_7_441), .b(output_7_2), .y(output_6_441));
wire output_8_441, output_8_2, output_7_441;
mixer gate_output_7_441(.a(output_8_441), .b(output_8_2), .y(output_7_441));
wire output_1_442, output_1_3, output_0_442;
mixer gate_output_0_442(.a(output_1_442), .b(output_1_3), .y(output_0_442));
wire output_2_442, output_2_3, output_1_442;
mixer gate_output_1_442(.a(output_2_442), .b(output_2_3), .y(output_1_442));
wire output_3_442, output_3_3, output_2_442;
mixer gate_output_2_442(.a(output_3_442), .b(output_3_3), .y(output_2_442));
wire output_4_442, output_4_3, output_3_442;
mixer gate_output_3_442(.a(output_4_442), .b(output_4_3), .y(output_3_442));
wire output_5_442, output_5_3, output_4_442;
mixer gate_output_4_442(.a(output_5_442), .b(output_5_3), .y(output_4_442));
wire output_6_442, output_6_3, output_5_442;
mixer gate_output_5_442(.a(output_6_442), .b(output_6_3), .y(output_5_442));
wire output_7_442, output_7_3, output_6_442;
mixer gate_output_6_442(.a(output_7_442), .b(output_7_3), .y(output_6_442));
wire output_8_442, output_8_3, output_7_442;
mixer gate_output_7_442(.a(output_8_442), .b(output_8_3), .y(output_7_442));
wire output_1_443, output_1_4, output_0_443;
mixer gate_output_0_443(.a(output_1_443), .b(output_1_4), .y(output_0_443));
wire output_2_443, output_2_4, output_1_443;
mixer gate_output_1_443(.a(output_2_443), .b(output_2_4), .y(output_1_443));
wire output_3_443, output_3_4, output_2_443;
mixer gate_output_2_443(.a(output_3_443), .b(output_3_4), .y(output_2_443));
wire output_4_443, output_4_4, output_3_443;
mixer gate_output_3_443(.a(output_4_443), .b(output_4_4), .y(output_3_443));
wire output_5_443, output_5_4, output_4_443;
mixer gate_output_4_443(.a(output_5_443), .b(output_5_4), .y(output_4_443));
wire output_6_443, output_6_4, output_5_443;
mixer gate_output_5_443(.a(output_6_443), .b(output_6_4), .y(output_5_443));
wire output_7_443, output_7_4, output_6_443;
mixer gate_output_6_443(.a(output_7_443), .b(output_7_4), .y(output_6_443));
wire output_8_443, output_8_4, output_7_443;
mixer gate_output_7_443(.a(output_8_443), .b(output_8_4), .y(output_7_443));
wire output_1_444, output_1_5, output_0_444;
mixer gate_output_0_444(.a(output_1_444), .b(output_1_5), .y(output_0_444));
wire output_2_444, output_2_5, output_1_444;
mixer gate_output_1_444(.a(output_2_444), .b(output_2_5), .y(output_1_444));
wire output_3_444, output_3_5, output_2_444;
mixer gate_output_2_444(.a(output_3_444), .b(output_3_5), .y(output_2_444));
wire output_4_444, output_4_5, output_3_444;
mixer gate_output_3_444(.a(output_4_444), .b(output_4_5), .y(output_3_444));
wire output_5_444, output_5_5, output_4_444;
mixer gate_output_4_444(.a(output_5_444), .b(output_5_5), .y(output_4_444));
wire output_6_444, output_6_5, output_5_444;
mixer gate_output_5_444(.a(output_6_444), .b(output_6_5), .y(output_5_444));
wire output_7_444, output_7_5, output_6_444;
mixer gate_output_6_444(.a(output_7_444), .b(output_7_5), .y(output_6_444));
wire output_8_444, output_8_5, output_7_444;
mixer gate_output_7_444(.a(output_8_444), .b(output_8_5), .y(output_7_444));
wire output_1_445, output_1_6, output_0_445;
mixer gate_output_0_445(.a(output_1_445), .b(output_1_6), .y(output_0_445));
wire output_2_445, output_2_6, output_1_445;
mixer gate_output_1_445(.a(output_2_445), .b(output_2_6), .y(output_1_445));
wire output_3_445, output_3_6, output_2_445;
mixer gate_output_2_445(.a(output_3_445), .b(output_3_6), .y(output_2_445));
wire output_4_445, output_4_6, output_3_445;
mixer gate_output_3_445(.a(output_4_445), .b(output_4_6), .y(output_3_445));
wire output_5_445, output_5_6, output_4_445;
mixer gate_output_4_445(.a(output_5_445), .b(output_5_6), .y(output_4_445));
wire output_6_445, output_6_6, output_5_445;
mixer gate_output_5_445(.a(output_6_445), .b(output_6_6), .y(output_5_445));
wire output_7_445, output_7_6, output_6_445;
mixer gate_output_6_445(.a(output_7_445), .b(output_7_6), .y(output_6_445));
wire output_8_445, output_8_6, output_7_445;
mixer gate_output_7_445(.a(output_8_445), .b(output_8_6), .y(output_7_445));
wire output_1_446, output_1_7, output_0_446;
mixer gate_output_0_446(.a(output_1_446), .b(output_1_7), .y(output_0_446));
wire output_2_446, output_2_7, output_1_446;
mixer gate_output_1_446(.a(output_2_446), .b(output_2_7), .y(output_1_446));
wire output_3_446, output_3_7, output_2_446;
mixer gate_output_2_446(.a(output_3_446), .b(output_3_7), .y(output_2_446));
wire output_4_446, output_4_7, output_3_446;
mixer gate_output_3_446(.a(output_4_446), .b(output_4_7), .y(output_3_446));
wire output_5_446, output_5_7, output_4_446;
mixer gate_output_4_446(.a(output_5_446), .b(output_5_7), .y(output_4_446));
wire output_6_446, output_6_7, output_5_446;
mixer gate_output_5_446(.a(output_6_446), .b(output_6_7), .y(output_5_446));
wire output_7_446, output_7_7, output_6_446;
mixer gate_output_6_446(.a(output_7_446), .b(output_7_7), .y(output_6_446));
wire output_8_446, output_8_7, output_7_446;
mixer gate_output_7_446(.a(output_8_446), .b(output_8_7), .y(output_7_446));
wire output_1_447, output_1_0, output_0_447;
mixer gate_output_0_447(.a(output_1_447), .b(output_1_0), .y(output_0_447));
wire output_2_447, output_2_0, output_1_447;
mixer gate_output_1_447(.a(output_2_447), .b(output_2_0), .y(output_1_447));
wire output_3_447, output_3_0, output_2_447;
mixer gate_output_2_447(.a(output_3_447), .b(output_3_0), .y(output_2_447));
wire output_4_447, output_4_0, output_3_447;
mixer gate_output_3_447(.a(output_4_447), .b(output_4_0), .y(output_3_447));
wire output_5_447, output_5_0, output_4_447;
mixer gate_output_4_447(.a(output_5_447), .b(output_5_0), .y(output_4_447));
wire output_6_447, output_6_0, output_5_447;
mixer gate_output_5_447(.a(output_6_447), .b(output_6_0), .y(output_5_447));
wire output_7_447, output_7_0, output_6_447;
mixer gate_output_6_447(.a(output_7_447), .b(output_7_0), .y(output_6_447));
wire output_8_447, output_8_0, output_7_447;
mixer gate_output_7_447(.a(output_8_447), .b(output_8_0), .y(output_7_447));
wire output_1_448, output_1_1, output_0_448;
mixer gate_output_0_448(.a(output_1_448), .b(output_1_1), .y(output_0_448));
wire output_2_448, output_2_1, output_1_448;
mixer gate_output_1_448(.a(output_2_448), .b(output_2_1), .y(output_1_448));
wire output_3_448, output_3_1, output_2_448;
mixer gate_output_2_448(.a(output_3_448), .b(output_3_1), .y(output_2_448));
wire output_4_448, output_4_1, output_3_448;
mixer gate_output_3_448(.a(output_4_448), .b(output_4_1), .y(output_3_448));
wire output_5_448, output_5_1, output_4_448;
mixer gate_output_4_448(.a(output_5_448), .b(output_5_1), .y(output_4_448));
wire output_6_448, output_6_1, output_5_448;
mixer gate_output_5_448(.a(output_6_448), .b(output_6_1), .y(output_5_448));
wire output_7_448, output_7_1, output_6_448;
mixer gate_output_6_448(.a(output_7_448), .b(output_7_1), .y(output_6_448));
wire output_8_448, output_8_1, output_7_448;
mixer gate_output_7_448(.a(output_8_448), .b(output_8_1), .y(output_7_448));
wire output_1_449, output_1_2, output_0_449;
mixer gate_output_0_449(.a(output_1_449), .b(output_1_2), .y(output_0_449));
wire output_2_449, output_2_2, output_1_449;
mixer gate_output_1_449(.a(output_2_449), .b(output_2_2), .y(output_1_449));
wire output_3_449, output_3_2, output_2_449;
mixer gate_output_2_449(.a(output_3_449), .b(output_3_2), .y(output_2_449));
wire output_4_449, output_4_2, output_3_449;
mixer gate_output_3_449(.a(output_4_449), .b(output_4_2), .y(output_3_449));
wire output_5_449, output_5_2, output_4_449;
mixer gate_output_4_449(.a(output_5_449), .b(output_5_2), .y(output_4_449));
wire output_6_449, output_6_2, output_5_449;
mixer gate_output_5_449(.a(output_6_449), .b(output_6_2), .y(output_5_449));
wire output_7_449, output_7_2, output_6_449;
mixer gate_output_6_449(.a(output_7_449), .b(output_7_2), .y(output_6_449));
wire output_8_449, output_8_2, output_7_449;
mixer gate_output_7_449(.a(output_8_449), .b(output_8_2), .y(output_7_449));
wire output_1_450, output_1_3, output_0_450;
mixer gate_output_0_450(.a(output_1_450), .b(output_1_3), .y(output_0_450));
wire output_2_450, output_2_3, output_1_450;
mixer gate_output_1_450(.a(output_2_450), .b(output_2_3), .y(output_1_450));
wire output_3_450, output_3_3, output_2_450;
mixer gate_output_2_450(.a(output_3_450), .b(output_3_3), .y(output_2_450));
wire output_4_450, output_4_3, output_3_450;
mixer gate_output_3_450(.a(output_4_450), .b(output_4_3), .y(output_3_450));
wire output_5_450, output_5_3, output_4_450;
mixer gate_output_4_450(.a(output_5_450), .b(output_5_3), .y(output_4_450));
wire output_6_450, output_6_3, output_5_450;
mixer gate_output_5_450(.a(output_6_450), .b(output_6_3), .y(output_5_450));
wire output_7_450, output_7_3, output_6_450;
mixer gate_output_6_450(.a(output_7_450), .b(output_7_3), .y(output_6_450));
wire output_8_450, output_8_3, output_7_450;
mixer gate_output_7_450(.a(output_8_450), .b(output_8_3), .y(output_7_450));
wire output_1_451, output_1_4, output_0_451;
mixer gate_output_0_451(.a(output_1_451), .b(output_1_4), .y(output_0_451));
wire output_2_451, output_2_4, output_1_451;
mixer gate_output_1_451(.a(output_2_451), .b(output_2_4), .y(output_1_451));
wire output_3_451, output_3_4, output_2_451;
mixer gate_output_2_451(.a(output_3_451), .b(output_3_4), .y(output_2_451));
wire output_4_451, output_4_4, output_3_451;
mixer gate_output_3_451(.a(output_4_451), .b(output_4_4), .y(output_3_451));
wire output_5_451, output_5_4, output_4_451;
mixer gate_output_4_451(.a(output_5_451), .b(output_5_4), .y(output_4_451));
wire output_6_451, output_6_4, output_5_451;
mixer gate_output_5_451(.a(output_6_451), .b(output_6_4), .y(output_5_451));
wire output_7_451, output_7_4, output_6_451;
mixer gate_output_6_451(.a(output_7_451), .b(output_7_4), .y(output_6_451));
wire output_8_451, output_8_4, output_7_451;
mixer gate_output_7_451(.a(output_8_451), .b(output_8_4), .y(output_7_451));
wire output_1_452, output_1_5, output_0_452;
mixer gate_output_0_452(.a(output_1_452), .b(output_1_5), .y(output_0_452));
wire output_2_452, output_2_5, output_1_452;
mixer gate_output_1_452(.a(output_2_452), .b(output_2_5), .y(output_1_452));
wire output_3_452, output_3_5, output_2_452;
mixer gate_output_2_452(.a(output_3_452), .b(output_3_5), .y(output_2_452));
wire output_4_452, output_4_5, output_3_452;
mixer gate_output_3_452(.a(output_4_452), .b(output_4_5), .y(output_3_452));
wire output_5_452, output_5_5, output_4_452;
mixer gate_output_4_452(.a(output_5_452), .b(output_5_5), .y(output_4_452));
wire output_6_452, output_6_5, output_5_452;
mixer gate_output_5_452(.a(output_6_452), .b(output_6_5), .y(output_5_452));
wire output_7_452, output_7_5, output_6_452;
mixer gate_output_6_452(.a(output_7_452), .b(output_7_5), .y(output_6_452));
wire output_8_452, output_8_5, output_7_452;
mixer gate_output_7_452(.a(output_8_452), .b(output_8_5), .y(output_7_452));
wire output_1_453, output_1_6, output_0_453;
mixer gate_output_0_453(.a(output_1_453), .b(output_1_6), .y(output_0_453));
wire output_2_453, output_2_6, output_1_453;
mixer gate_output_1_453(.a(output_2_453), .b(output_2_6), .y(output_1_453));
wire output_3_453, output_3_6, output_2_453;
mixer gate_output_2_453(.a(output_3_453), .b(output_3_6), .y(output_2_453));
wire output_4_453, output_4_6, output_3_453;
mixer gate_output_3_453(.a(output_4_453), .b(output_4_6), .y(output_3_453));
wire output_5_453, output_5_6, output_4_453;
mixer gate_output_4_453(.a(output_5_453), .b(output_5_6), .y(output_4_453));
wire output_6_453, output_6_6, output_5_453;
mixer gate_output_5_453(.a(output_6_453), .b(output_6_6), .y(output_5_453));
wire output_7_453, output_7_6, output_6_453;
mixer gate_output_6_453(.a(output_7_453), .b(output_7_6), .y(output_6_453));
wire output_8_453, output_8_6, output_7_453;
mixer gate_output_7_453(.a(output_8_453), .b(output_8_6), .y(output_7_453));
wire output_1_454, output_1_7, output_0_454;
mixer gate_output_0_454(.a(output_1_454), .b(output_1_7), .y(output_0_454));
wire output_2_454, output_2_7, output_1_454;
mixer gate_output_1_454(.a(output_2_454), .b(output_2_7), .y(output_1_454));
wire output_3_454, output_3_7, output_2_454;
mixer gate_output_2_454(.a(output_3_454), .b(output_3_7), .y(output_2_454));
wire output_4_454, output_4_7, output_3_454;
mixer gate_output_3_454(.a(output_4_454), .b(output_4_7), .y(output_3_454));
wire output_5_454, output_5_7, output_4_454;
mixer gate_output_4_454(.a(output_5_454), .b(output_5_7), .y(output_4_454));
wire output_6_454, output_6_7, output_5_454;
mixer gate_output_5_454(.a(output_6_454), .b(output_6_7), .y(output_5_454));
wire output_7_454, output_7_7, output_6_454;
mixer gate_output_6_454(.a(output_7_454), .b(output_7_7), .y(output_6_454));
wire output_8_454, output_8_7, output_7_454;
mixer gate_output_7_454(.a(output_8_454), .b(output_8_7), .y(output_7_454));
wire output_1_455, output_1_0, output_0_455;
mixer gate_output_0_455(.a(output_1_455), .b(output_1_0), .y(output_0_455));
wire output_2_455, output_2_0, output_1_455;
mixer gate_output_1_455(.a(output_2_455), .b(output_2_0), .y(output_1_455));
wire output_3_455, output_3_0, output_2_455;
mixer gate_output_2_455(.a(output_3_455), .b(output_3_0), .y(output_2_455));
wire output_4_455, output_4_0, output_3_455;
mixer gate_output_3_455(.a(output_4_455), .b(output_4_0), .y(output_3_455));
wire output_5_455, output_5_0, output_4_455;
mixer gate_output_4_455(.a(output_5_455), .b(output_5_0), .y(output_4_455));
wire output_6_455, output_6_0, output_5_455;
mixer gate_output_5_455(.a(output_6_455), .b(output_6_0), .y(output_5_455));
wire output_7_455, output_7_0, output_6_455;
mixer gate_output_6_455(.a(output_7_455), .b(output_7_0), .y(output_6_455));
wire output_8_455, output_8_0, output_7_455;
mixer gate_output_7_455(.a(output_8_455), .b(output_8_0), .y(output_7_455));
wire output_1_456, output_1_1, output_0_456;
mixer gate_output_0_456(.a(output_1_456), .b(output_1_1), .y(output_0_456));
wire output_2_456, output_2_1, output_1_456;
mixer gate_output_1_456(.a(output_2_456), .b(output_2_1), .y(output_1_456));
wire output_3_456, output_3_1, output_2_456;
mixer gate_output_2_456(.a(output_3_456), .b(output_3_1), .y(output_2_456));
wire output_4_456, output_4_1, output_3_456;
mixer gate_output_3_456(.a(output_4_456), .b(output_4_1), .y(output_3_456));
wire output_5_456, output_5_1, output_4_456;
mixer gate_output_4_456(.a(output_5_456), .b(output_5_1), .y(output_4_456));
wire output_6_456, output_6_1, output_5_456;
mixer gate_output_5_456(.a(output_6_456), .b(output_6_1), .y(output_5_456));
wire output_7_456, output_7_1, output_6_456;
mixer gate_output_6_456(.a(output_7_456), .b(output_7_1), .y(output_6_456));
wire output_8_456, output_8_1, output_7_456;
mixer gate_output_7_456(.a(output_8_456), .b(output_8_1), .y(output_7_456));
wire output_1_457, output_1_2, output_0_457;
mixer gate_output_0_457(.a(output_1_457), .b(output_1_2), .y(output_0_457));
wire output_2_457, output_2_2, output_1_457;
mixer gate_output_1_457(.a(output_2_457), .b(output_2_2), .y(output_1_457));
wire output_3_457, output_3_2, output_2_457;
mixer gate_output_2_457(.a(output_3_457), .b(output_3_2), .y(output_2_457));
wire output_4_457, output_4_2, output_3_457;
mixer gate_output_3_457(.a(output_4_457), .b(output_4_2), .y(output_3_457));
wire output_5_457, output_5_2, output_4_457;
mixer gate_output_4_457(.a(output_5_457), .b(output_5_2), .y(output_4_457));
wire output_6_457, output_6_2, output_5_457;
mixer gate_output_5_457(.a(output_6_457), .b(output_6_2), .y(output_5_457));
wire output_7_457, output_7_2, output_6_457;
mixer gate_output_6_457(.a(output_7_457), .b(output_7_2), .y(output_6_457));
wire output_8_457, output_8_2, output_7_457;
mixer gate_output_7_457(.a(output_8_457), .b(output_8_2), .y(output_7_457));
wire output_1_458, output_1_3, output_0_458;
mixer gate_output_0_458(.a(output_1_458), .b(output_1_3), .y(output_0_458));
wire output_2_458, output_2_3, output_1_458;
mixer gate_output_1_458(.a(output_2_458), .b(output_2_3), .y(output_1_458));
wire output_3_458, output_3_3, output_2_458;
mixer gate_output_2_458(.a(output_3_458), .b(output_3_3), .y(output_2_458));
wire output_4_458, output_4_3, output_3_458;
mixer gate_output_3_458(.a(output_4_458), .b(output_4_3), .y(output_3_458));
wire output_5_458, output_5_3, output_4_458;
mixer gate_output_4_458(.a(output_5_458), .b(output_5_3), .y(output_4_458));
wire output_6_458, output_6_3, output_5_458;
mixer gate_output_5_458(.a(output_6_458), .b(output_6_3), .y(output_5_458));
wire output_7_458, output_7_3, output_6_458;
mixer gate_output_6_458(.a(output_7_458), .b(output_7_3), .y(output_6_458));
wire output_8_458, output_8_3, output_7_458;
mixer gate_output_7_458(.a(output_8_458), .b(output_8_3), .y(output_7_458));
wire output_1_459, output_1_4, output_0_459;
mixer gate_output_0_459(.a(output_1_459), .b(output_1_4), .y(output_0_459));
wire output_2_459, output_2_4, output_1_459;
mixer gate_output_1_459(.a(output_2_459), .b(output_2_4), .y(output_1_459));
wire output_3_459, output_3_4, output_2_459;
mixer gate_output_2_459(.a(output_3_459), .b(output_3_4), .y(output_2_459));
wire output_4_459, output_4_4, output_3_459;
mixer gate_output_3_459(.a(output_4_459), .b(output_4_4), .y(output_3_459));
wire output_5_459, output_5_4, output_4_459;
mixer gate_output_4_459(.a(output_5_459), .b(output_5_4), .y(output_4_459));
wire output_6_459, output_6_4, output_5_459;
mixer gate_output_5_459(.a(output_6_459), .b(output_6_4), .y(output_5_459));
wire output_7_459, output_7_4, output_6_459;
mixer gate_output_6_459(.a(output_7_459), .b(output_7_4), .y(output_6_459));
wire output_8_459, output_8_4, output_7_459;
mixer gate_output_7_459(.a(output_8_459), .b(output_8_4), .y(output_7_459));
wire output_1_460, output_1_5, output_0_460;
mixer gate_output_0_460(.a(output_1_460), .b(output_1_5), .y(output_0_460));
wire output_2_460, output_2_5, output_1_460;
mixer gate_output_1_460(.a(output_2_460), .b(output_2_5), .y(output_1_460));
wire output_3_460, output_3_5, output_2_460;
mixer gate_output_2_460(.a(output_3_460), .b(output_3_5), .y(output_2_460));
wire output_4_460, output_4_5, output_3_460;
mixer gate_output_3_460(.a(output_4_460), .b(output_4_5), .y(output_3_460));
wire output_5_460, output_5_5, output_4_460;
mixer gate_output_4_460(.a(output_5_460), .b(output_5_5), .y(output_4_460));
wire output_6_460, output_6_5, output_5_460;
mixer gate_output_5_460(.a(output_6_460), .b(output_6_5), .y(output_5_460));
wire output_7_460, output_7_5, output_6_460;
mixer gate_output_6_460(.a(output_7_460), .b(output_7_5), .y(output_6_460));
wire output_8_460, output_8_5, output_7_460;
mixer gate_output_7_460(.a(output_8_460), .b(output_8_5), .y(output_7_460));
wire output_1_461, output_1_6, output_0_461;
mixer gate_output_0_461(.a(output_1_461), .b(output_1_6), .y(output_0_461));
wire output_2_461, output_2_6, output_1_461;
mixer gate_output_1_461(.a(output_2_461), .b(output_2_6), .y(output_1_461));
wire output_3_461, output_3_6, output_2_461;
mixer gate_output_2_461(.a(output_3_461), .b(output_3_6), .y(output_2_461));
wire output_4_461, output_4_6, output_3_461;
mixer gate_output_3_461(.a(output_4_461), .b(output_4_6), .y(output_3_461));
wire output_5_461, output_5_6, output_4_461;
mixer gate_output_4_461(.a(output_5_461), .b(output_5_6), .y(output_4_461));
wire output_6_461, output_6_6, output_5_461;
mixer gate_output_5_461(.a(output_6_461), .b(output_6_6), .y(output_5_461));
wire output_7_461, output_7_6, output_6_461;
mixer gate_output_6_461(.a(output_7_461), .b(output_7_6), .y(output_6_461));
wire output_8_461, output_8_6, output_7_461;
mixer gate_output_7_461(.a(output_8_461), .b(output_8_6), .y(output_7_461));
wire output_1_462, output_1_7, output_0_462;
mixer gate_output_0_462(.a(output_1_462), .b(output_1_7), .y(output_0_462));
wire output_2_462, output_2_7, output_1_462;
mixer gate_output_1_462(.a(output_2_462), .b(output_2_7), .y(output_1_462));
wire output_3_462, output_3_7, output_2_462;
mixer gate_output_2_462(.a(output_3_462), .b(output_3_7), .y(output_2_462));
wire output_4_462, output_4_7, output_3_462;
mixer gate_output_3_462(.a(output_4_462), .b(output_4_7), .y(output_3_462));
wire output_5_462, output_5_7, output_4_462;
mixer gate_output_4_462(.a(output_5_462), .b(output_5_7), .y(output_4_462));
wire output_6_462, output_6_7, output_5_462;
mixer gate_output_5_462(.a(output_6_462), .b(output_6_7), .y(output_5_462));
wire output_7_462, output_7_7, output_6_462;
mixer gate_output_6_462(.a(output_7_462), .b(output_7_7), .y(output_6_462));
wire output_8_462, output_8_7, output_7_462;
mixer gate_output_7_462(.a(output_8_462), .b(output_8_7), .y(output_7_462));
wire output_1_463, output_1_0, output_0_463;
mixer gate_output_0_463(.a(output_1_463), .b(output_1_0), .y(output_0_463));
wire output_2_463, output_2_0, output_1_463;
mixer gate_output_1_463(.a(output_2_463), .b(output_2_0), .y(output_1_463));
wire output_3_463, output_3_0, output_2_463;
mixer gate_output_2_463(.a(output_3_463), .b(output_3_0), .y(output_2_463));
wire output_4_463, output_4_0, output_3_463;
mixer gate_output_3_463(.a(output_4_463), .b(output_4_0), .y(output_3_463));
wire output_5_463, output_5_0, output_4_463;
mixer gate_output_4_463(.a(output_5_463), .b(output_5_0), .y(output_4_463));
wire output_6_463, output_6_0, output_5_463;
mixer gate_output_5_463(.a(output_6_463), .b(output_6_0), .y(output_5_463));
wire output_7_463, output_7_0, output_6_463;
mixer gate_output_6_463(.a(output_7_463), .b(output_7_0), .y(output_6_463));
wire output_8_463, output_8_0, output_7_463;
mixer gate_output_7_463(.a(output_8_463), .b(output_8_0), .y(output_7_463));
wire output_1_464, output_1_1, output_0_464;
mixer gate_output_0_464(.a(output_1_464), .b(output_1_1), .y(output_0_464));
wire output_2_464, output_2_1, output_1_464;
mixer gate_output_1_464(.a(output_2_464), .b(output_2_1), .y(output_1_464));
wire output_3_464, output_3_1, output_2_464;
mixer gate_output_2_464(.a(output_3_464), .b(output_3_1), .y(output_2_464));
wire output_4_464, output_4_1, output_3_464;
mixer gate_output_3_464(.a(output_4_464), .b(output_4_1), .y(output_3_464));
wire output_5_464, output_5_1, output_4_464;
mixer gate_output_4_464(.a(output_5_464), .b(output_5_1), .y(output_4_464));
wire output_6_464, output_6_1, output_5_464;
mixer gate_output_5_464(.a(output_6_464), .b(output_6_1), .y(output_5_464));
wire output_7_464, output_7_1, output_6_464;
mixer gate_output_6_464(.a(output_7_464), .b(output_7_1), .y(output_6_464));
wire output_8_464, output_8_1, output_7_464;
mixer gate_output_7_464(.a(output_8_464), .b(output_8_1), .y(output_7_464));
wire output_1_465, output_1_2, output_0_465;
mixer gate_output_0_465(.a(output_1_465), .b(output_1_2), .y(output_0_465));
wire output_2_465, output_2_2, output_1_465;
mixer gate_output_1_465(.a(output_2_465), .b(output_2_2), .y(output_1_465));
wire output_3_465, output_3_2, output_2_465;
mixer gate_output_2_465(.a(output_3_465), .b(output_3_2), .y(output_2_465));
wire output_4_465, output_4_2, output_3_465;
mixer gate_output_3_465(.a(output_4_465), .b(output_4_2), .y(output_3_465));
wire output_5_465, output_5_2, output_4_465;
mixer gate_output_4_465(.a(output_5_465), .b(output_5_2), .y(output_4_465));
wire output_6_465, output_6_2, output_5_465;
mixer gate_output_5_465(.a(output_6_465), .b(output_6_2), .y(output_5_465));
wire output_7_465, output_7_2, output_6_465;
mixer gate_output_6_465(.a(output_7_465), .b(output_7_2), .y(output_6_465));
wire output_8_465, output_8_2, output_7_465;
mixer gate_output_7_465(.a(output_8_465), .b(output_8_2), .y(output_7_465));
wire output_1_466, output_1_3, output_0_466;
mixer gate_output_0_466(.a(output_1_466), .b(output_1_3), .y(output_0_466));
wire output_2_466, output_2_3, output_1_466;
mixer gate_output_1_466(.a(output_2_466), .b(output_2_3), .y(output_1_466));
wire output_3_466, output_3_3, output_2_466;
mixer gate_output_2_466(.a(output_3_466), .b(output_3_3), .y(output_2_466));
wire output_4_466, output_4_3, output_3_466;
mixer gate_output_3_466(.a(output_4_466), .b(output_4_3), .y(output_3_466));
wire output_5_466, output_5_3, output_4_466;
mixer gate_output_4_466(.a(output_5_466), .b(output_5_3), .y(output_4_466));
wire output_6_466, output_6_3, output_5_466;
mixer gate_output_5_466(.a(output_6_466), .b(output_6_3), .y(output_5_466));
wire output_7_466, output_7_3, output_6_466;
mixer gate_output_6_466(.a(output_7_466), .b(output_7_3), .y(output_6_466));
wire output_8_466, output_8_3, output_7_466;
mixer gate_output_7_466(.a(output_8_466), .b(output_8_3), .y(output_7_466));
wire output_1_467, output_1_4, output_0_467;
mixer gate_output_0_467(.a(output_1_467), .b(output_1_4), .y(output_0_467));
wire output_2_467, output_2_4, output_1_467;
mixer gate_output_1_467(.a(output_2_467), .b(output_2_4), .y(output_1_467));
wire output_3_467, output_3_4, output_2_467;
mixer gate_output_2_467(.a(output_3_467), .b(output_3_4), .y(output_2_467));
wire output_4_467, output_4_4, output_3_467;
mixer gate_output_3_467(.a(output_4_467), .b(output_4_4), .y(output_3_467));
wire output_5_467, output_5_4, output_4_467;
mixer gate_output_4_467(.a(output_5_467), .b(output_5_4), .y(output_4_467));
wire output_6_467, output_6_4, output_5_467;
mixer gate_output_5_467(.a(output_6_467), .b(output_6_4), .y(output_5_467));
wire output_7_467, output_7_4, output_6_467;
mixer gate_output_6_467(.a(output_7_467), .b(output_7_4), .y(output_6_467));
wire output_8_467, output_8_4, output_7_467;
mixer gate_output_7_467(.a(output_8_467), .b(output_8_4), .y(output_7_467));
wire output_1_468, output_1_5, output_0_468;
mixer gate_output_0_468(.a(output_1_468), .b(output_1_5), .y(output_0_468));
wire output_2_468, output_2_5, output_1_468;
mixer gate_output_1_468(.a(output_2_468), .b(output_2_5), .y(output_1_468));
wire output_3_468, output_3_5, output_2_468;
mixer gate_output_2_468(.a(output_3_468), .b(output_3_5), .y(output_2_468));
wire output_4_468, output_4_5, output_3_468;
mixer gate_output_3_468(.a(output_4_468), .b(output_4_5), .y(output_3_468));
wire output_5_468, output_5_5, output_4_468;
mixer gate_output_4_468(.a(output_5_468), .b(output_5_5), .y(output_4_468));
wire output_6_468, output_6_5, output_5_468;
mixer gate_output_5_468(.a(output_6_468), .b(output_6_5), .y(output_5_468));
wire output_7_468, output_7_5, output_6_468;
mixer gate_output_6_468(.a(output_7_468), .b(output_7_5), .y(output_6_468));
wire output_8_468, output_8_5, output_7_468;
mixer gate_output_7_468(.a(output_8_468), .b(output_8_5), .y(output_7_468));
wire output_1_469, output_1_6, output_0_469;
mixer gate_output_0_469(.a(output_1_469), .b(output_1_6), .y(output_0_469));
wire output_2_469, output_2_6, output_1_469;
mixer gate_output_1_469(.a(output_2_469), .b(output_2_6), .y(output_1_469));
wire output_3_469, output_3_6, output_2_469;
mixer gate_output_2_469(.a(output_3_469), .b(output_3_6), .y(output_2_469));
wire output_4_469, output_4_6, output_3_469;
mixer gate_output_3_469(.a(output_4_469), .b(output_4_6), .y(output_3_469));
wire output_5_469, output_5_6, output_4_469;
mixer gate_output_4_469(.a(output_5_469), .b(output_5_6), .y(output_4_469));
wire output_6_469, output_6_6, output_5_469;
mixer gate_output_5_469(.a(output_6_469), .b(output_6_6), .y(output_5_469));
wire output_7_469, output_7_6, output_6_469;
mixer gate_output_6_469(.a(output_7_469), .b(output_7_6), .y(output_6_469));
wire output_8_469, output_8_6, output_7_469;
mixer gate_output_7_469(.a(output_8_469), .b(output_8_6), .y(output_7_469));
wire output_1_470, output_1_7, output_0_470;
mixer gate_output_0_470(.a(output_1_470), .b(output_1_7), .y(output_0_470));
wire output_2_470, output_2_7, output_1_470;
mixer gate_output_1_470(.a(output_2_470), .b(output_2_7), .y(output_1_470));
wire output_3_470, output_3_7, output_2_470;
mixer gate_output_2_470(.a(output_3_470), .b(output_3_7), .y(output_2_470));
wire output_4_470, output_4_7, output_3_470;
mixer gate_output_3_470(.a(output_4_470), .b(output_4_7), .y(output_3_470));
wire output_5_470, output_5_7, output_4_470;
mixer gate_output_4_470(.a(output_5_470), .b(output_5_7), .y(output_4_470));
wire output_6_470, output_6_7, output_5_470;
mixer gate_output_5_470(.a(output_6_470), .b(output_6_7), .y(output_5_470));
wire output_7_470, output_7_7, output_6_470;
mixer gate_output_6_470(.a(output_7_470), .b(output_7_7), .y(output_6_470));
wire output_8_470, output_8_7, output_7_470;
mixer gate_output_7_470(.a(output_8_470), .b(output_8_7), .y(output_7_470));
wire output_1_471, output_1_0, output_0_471;
mixer gate_output_0_471(.a(output_1_471), .b(output_1_0), .y(output_0_471));
wire output_2_471, output_2_0, output_1_471;
mixer gate_output_1_471(.a(output_2_471), .b(output_2_0), .y(output_1_471));
wire output_3_471, output_3_0, output_2_471;
mixer gate_output_2_471(.a(output_3_471), .b(output_3_0), .y(output_2_471));
wire output_4_471, output_4_0, output_3_471;
mixer gate_output_3_471(.a(output_4_471), .b(output_4_0), .y(output_3_471));
wire output_5_471, output_5_0, output_4_471;
mixer gate_output_4_471(.a(output_5_471), .b(output_5_0), .y(output_4_471));
wire output_6_471, output_6_0, output_5_471;
mixer gate_output_5_471(.a(output_6_471), .b(output_6_0), .y(output_5_471));
wire output_7_471, output_7_0, output_6_471;
mixer gate_output_6_471(.a(output_7_471), .b(output_7_0), .y(output_6_471));
wire output_8_471, output_8_0, output_7_471;
mixer gate_output_7_471(.a(output_8_471), .b(output_8_0), .y(output_7_471));
wire output_1_472, output_1_1, output_0_472;
mixer gate_output_0_472(.a(output_1_472), .b(output_1_1), .y(output_0_472));
wire output_2_472, output_2_1, output_1_472;
mixer gate_output_1_472(.a(output_2_472), .b(output_2_1), .y(output_1_472));
wire output_3_472, output_3_1, output_2_472;
mixer gate_output_2_472(.a(output_3_472), .b(output_3_1), .y(output_2_472));
wire output_4_472, output_4_1, output_3_472;
mixer gate_output_3_472(.a(output_4_472), .b(output_4_1), .y(output_3_472));
wire output_5_472, output_5_1, output_4_472;
mixer gate_output_4_472(.a(output_5_472), .b(output_5_1), .y(output_4_472));
wire output_6_472, output_6_1, output_5_472;
mixer gate_output_5_472(.a(output_6_472), .b(output_6_1), .y(output_5_472));
wire output_7_472, output_7_1, output_6_472;
mixer gate_output_6_472(.a(output_7_472), .b(output_7_1), .y(output_6_472));
wire output_8_472, output_8_1, output_7_472;
mixer gate_output_7_472(.a(output_8_472), .b(output_8_1), .y(output_7_472));
wire output_1_473, output_1_2, output_0_473;
mixer gate_output_0_473(.a(output_1_473), .b(output_1_2), .y(output_0_473));
wire output_2_473, output_2_2, output_1_473;
mixer gate_output_1_473(.a(output_2_473), .b(output_2_2), .y(output_1_473));
wire output_3_473, output_3_2, output_2_473;
mixer gate_output_2_473(.a(output_3_473), .b(output_3_2), .y(output_2_473));
wire output_4_473, output_4_2, output_3_473;
mixer gate_output_3_473(.a(output_4_473), .b(output_4_2), .y(output_3_473));
wire output_5_473, output_5_2, output_4_473;
mixer gate_output_4_473(.a(output_5_473), .b(output_5_2), .y(output_4_473));
wire output_6_473, output_6_2, output_5_473;
mixer gate_output_5_473(.a(output_6_473), .b(output_6_2), .y(output_5_473));
wire output_7_473, output_7_2, output_6_473;
mixer gate_output_6_473(.a(output_7_473), .b(output_7_2), .y(output_6_473));
wire output_8_473, output_8_2, output_7_473;
mixer gate_output_7_473(.a(output_8_473), .b(output_8_2), .y(output_7_473));
wire output_1_474, output_1_3, output_0_474;
mixer gate_output_0_474(.a(output_1_474), .b(output_1_3), .y(output_0_474));
wire output_2_474, output_2_3, output_1_474;
mixer gate_output_1_474(.a(output_2_474), .b(output_2_3), .y(output_1_474));
wire output_3_474, output_3_3, output_2_474;
mixer gate_output_2_474(.a(output_3_474), .b(output_3_3), .y(output_2_474));
wire output_4_474, output_4_3, output_3_474;
mixer gate_output_3_474(.a(output_4_474), .b(output_4_3), .y(output_3_474));
wire output_5_474, output_5_3, output_4_474;
mixer gate_output_4_474(.a(output_5_474), .b(output_5_3), .y(output_4_474));
wire output_6_474, output_6_3, output_5_474;
mixer gate_output_5_474(.a(output_6_474), .b(output_6_3), .y(output_5_474));
wire output_7_474, output_7_3, output_6_474;
mixer gate_output_6_474(.a(output_7_474), .b(output_7_3), .y(output_6_474));
wire output_8_474, output_8_3, output_7_474;
mixer gate_output_7_474(.a(output_8_474), .b(output_8_3), .y(output_7_474));
wire output_1_475, output_1_4, output_0_475;
mixer gate_output_0_475(.a(output_1_475), .b(output_1_4), .y(output_0_475));
wire output_2_475, output_2_4, output_1_475;
mixer gate_output_1_475(.a(output_2_475), .b(output_2_4), .y(output_1_475));
wire output_3_475, output_3_4, output_2_475;
mixer gate_output_2_475(.a(output_3_475), .b(output_3_4), .y(output_2_475));
wire output_4_475, output_4_4, output_3_475;
mixer gate_output_3_475(.a(output_4_475), .b(output_4_4), .y(output_3_475));
wire output_5_475, output_5_4, output_4_475;
mixer gate_output_4_475(.a(output_5_475), .b(output_5_4), .y(output_4_475));
wire output_6_475, output_6_4, output_5_475;
mixer gate_output_5_475(.a(output_6_475), .b(output_6_4), .y(output_5_475));
wire output_7_475, output_7_4, output_6_475;
mixer gate_output_6_475(.a(output_7_475), .b(output_7_4), .y(output_6_475));
wire output_8_475, output_8_4, output_7_475;
mixer gate_output_7_475(.a(output_8_475), .b(output_8_4), .y(output_7_475));
wire output_1_476, output_1_5, output_0_476;
mixer gate_output_0_476(.a(output_1_476), .b(output_1_5), .y(output_0_476));
wire output_2_476, output_2_5, output_1_476;
mixer gate_output_1_476(.a(output_2_476), .b(output_2_5), .y(output_1_476));
wire output_3_476, output_3_5, output_2_476;
mixer gate_output_2_476(.a(output_3_476), .b(output_3_5), .y(output_2_476));
wire output_4_476, output_4_5, output_3_476;
mixer gate_output_3_476(.a(output_4_476), .b(output_4_5), .y(output_3_476));
wire output_5_476, output_5_5, output_4_476;
mixer gate_output_4_476(.a(output_5_476), .b(output_5_5), .y(output_4_476));
wire output_6_476, output_6_5, output_5_476;
mixer gate_output_5_476(.a(output_6_476), .b(output_6_5), .y(output_5_476));
wire output_7_476, output_7_5, output_6_476;
mixer gate_output_6_476(.a(output_7_476), .b(output_7_5), .y(output_6_476));
wire output_8_476, output_8_5, output_7_476;
mixer gate_output_7_476(.a(output_8_476), .b(output_8_5), .y(output_7_476));
wire output_1_477, output_1_6, output_0_477;
mixer gate_output_0_477(.a(output_1_477), .b(output_1_6), .y(output_0_477));
wire output_2_477, output_2_6, output_1_477;
mixer gate_output_1_477(.a(output_2_477), .b(output_2_6), .y(output_1_477));
wire output_3_477, output_3_6, output_2_477;
mixer gate_output_2_477(.a(output_3_477), .b(output_3_6), .y(output_2_477));
wire output_4_477, output_4_6, output_3_477;
mixer gate_output_3_477(.a(output_4_477), .b(output_4_6), .y(output_3_477));
wire output_5_477, output_5_6, output_4_477;
mixer gate_output_4_477(.a(output_5_477), .b(output_5_6), .y(output_4_477));
wire output_6_477, output_6_6, output_5_477;
mixer gate_output_5_477(.a(output_6_477), .b(output_6_6), .y(output_5_477));
wire output_7_477, output_7_6, output_6_477;
mixer gate_output_6_477(.a(output_7_477), .b(output_7_6), .y(output_6_477));
wire output_8_477, output_8_6, output_7_477;
mixer gate_output_7_477(.a(output_8_477), .b(output_8_6), .y(output_7_477));
wire output_1_478, output_1_7, output_0_478;
mixer gate_output_0_478(.a(output_1_478), .b(output_1_7), .y(output_0_478));
wire output_2_478, output_2_7, output_1_478;
mixer gate_output_1_478(.a(output_2_478), .b(output_2_7), .y(output_1_478));
wire output_3_478, output_3_7, output_2_478;
mixer gate_output_2_478(.a(output_3_478), .b(output_3_7), .y(output_2_478));
wire output_4_478, output_4_7, output_3_478;
mixer gate_output_3_478(.a(output_4_478), .b(output_4_7), .y(output_3_478));
wire output_5_478, output_5_7, output_4_478;
mixer gate_output_4_478(.a(output_5_478), .b(output_5_7), .y(output_4_478));
wire output_6_478, output_6_7, output_5_478;
mixer gate_output_5_478(.a(output_6_478), .b(output_6_7), .y(output_5_478));
wire output_7_478, output_7_7, output_6_478;
mixer gate_output_6_478(.a(output_7_478), .b(output_7_7), .y(output_6_478));
wire output_8_478, output_8_7, output_7_478;
mixer gate_output_7_478(.a(output_8_478), .b(output_8_7), .y(output_7_478));
wire output_1_479, output_1_0, output_0_479;
mixer gate_output_0_479(.a(output_1_479), .b(output_1_0), .y(output_0_479));
wire output_2_479, output_2_0, output_1_479;
mixer gate_output_1_479(.a(output_2_479), .b(output_2_0), .y(output_1_479));
wire output_3_479, output_3_0, output_2_479;
mixer gate_output_2_479(.a(output_3_479), .b(output_3_0), .y(output_2_479));
wire output_4_479, output_4_0, output_3_479;
mixer gate_output_3_479(.a(output_4_479), .b(output_4_0), .y(output_3_479));
wire output_5_479, output_5_0, output_4_479;
mixer gate_output_4_479(.a(output_5_479), .b(output_5_0), .y(output_4_479));
wire output_6_479, output_6_0, output_5_479;
mixer gate_output_5_479(.a(output_6_479), .b(output_6_0), .y(output_5_479));
wire output_7_479, output_7_0, output_6_479;
mixer gate_output_6_479(.a(output_7_479), .b(output_7_0), .y(output_6_479));
wire output_8_479, output_8_0, output_7_479;
mixer gate_output_7_479(.a(output_8_479), .b(output_8_0), .y(output_7_479));
wire output_1_480, output_1_1, output_0_480;
mixer gate_output_0_480(.a(output_1_480), .b(output_1_1), .y(output_0_480));
wire output_2_480, output_2_1, output_1_480;
mixer gate_output_1_480(.a(output_2_480), .b(output_2_1), .y(output_1_480));
wire output_3_480, output_3_1, output_2_480;
mixer gate_output_2_480(.a(output_3_480), .b(output_3_1), .y(output_2_480));
wire output_4_480, output_4_1, output_3_480;
mixer gate_output_3_480(.a(output_4_480), .b(output_4_1), .y(output_3_480));
wire output_5_480, output_5_1, output_4_480;
mixer gate_output_4_480(.a(output_5_480), .b(output_5_1), .y(output_4_480));
wire output_6_480, output_6_1, output_5_480;
mixer gate_output_5_480(.a(output_6_480), .b(output_6_1), .y(output_5_480));
wire output_7_480, output_7_1, output_6_480;
mixer gate_output_6_480(.a(output_7_480), .b(output_7_1), .y(output_6_480));
wire output_8_480, output_8_1, output_7_480;
mixer gate_output_7_480(.a(output_8_480), .b(output_8_1), .y(output_7_480));
wire output_1_481, output_1_2, output_0_481;
mixer gate_output_0_481(.a(output_1_481), .b(output_1_2), .y(output_0_481));
wire output_2_481, output_2_2, output_1_481;
mixer gate_output_1_481(.a(output_2_481), .b(output_2_2), .y(output_1_481));
wire output_3_481, output_3_2, output_2_481;
mixer gate_output_2_481(.a(output_3_481), .b(output_3_2), .y(output_2_481));
wire output_4_481, output_4_2, output_3_481;
mixer gate_output_3_481(.a(output_4_481), .b(output_4_2), .y(output_3_481));
wire output_5_481, output_5_2, output_4_481;
mixer gate_output_4_481(.a(output_5_481), .b(output_5_2), .y(output_4_481));
wire output_6_481, output_6_2, output_5_481;
mixer gate_output_5_481(.a(output_6_481), .b(output_6_2), .y(output_5_481));
wire output_7_481, output_7_2, output_6_481;
mixer gate_output_6_481(.a(output_7_481), .b(output_7_2), .y(output_6_481));
wire output_8_481, output_8_2, output_7_481;
mixer gate_output_7_481(.a(output_8_481), .b(output_8_2), .y(output_7_481));
wire output_1_482, output_1_3, output_0_482;
mixer gate_output_0_482(.a(output_1_482), .b(output_1_3), .y(output_0_482));
wire output_2_482, output_2_3, output_1_482;
mixer gate_output_1_482(.a(output_2_482), .b(output_2_3), .y(output_1_482));
wire output_3_482, output_3_3, output_2_482;
mixer gate_output_2_482(.a(output_3_482), .b(output_3_3), .y(output_2_482));
wire output_4_482, output_4_3, output_3_482;
mixer gate_output_3_482(.a(output_4_482), .b(output_4_3), .y(output_3_482));
wire output_5_482, output_5_3, output_4_482;
mixer gate_output_4_482(.a(output_5_482), .b(output_5_3), .y(output_4_482));
wire output_6_482, output_6_3, output_5_482;
mixer gate_output_5_482(.a(output_6_482), .b(output_6_3), .y(output_5_482));
wire output_7_482, output_7_3, output_6_482;
mixer gate_output_6_482(.a(output_7_482), .b(output_7_3), .y(output_6_482));
wire output_8_482, output_8_3, output_7_482;
mixer gate_output_7_482(.a(output_8_482), .b(output_8_3), .y(output_7_482));
wire output_1_483, output_1_4, output_0_483;
mixer gate_output_0_483(.a(output_1_483), .b(output_1_4), .y(output_0_483));
wire output_2_483, output_2_4, output_1_483;
mixer gate_output_1_483(.a(output_2_483), .b(output_2_4), .y(output_1_483));
wire output_3_483, output_3_4, output_2_483;
mixer gate_output_2_483(.a(output_3_483), .b(output_3_4), .y(output_2_483));
wire output_4_483, output_4_4, output_3_483;
mixer gate_output_3_483(.a(output_4_483), .b(output_4_4), .y(output_3_483));
wire output_5_483, output_5_4, output_4_483;
mixer gate_output_4_483(.a(output_5_483), .b(output_5_4), .y(output_4_483));
wire output_6_483, output_6_4, output_5_483;
mixer gate_output_5_483(.a(output_6_483), .b(output_6_4), .y(output_5_483));
wire output_7_483, output_7_4, output_6_483;
mixer gate_output_6_483(.a(output_7_483), .b(output_7_4), .y(output_6_483));
wire output_8_483, output_8_4, output_7_483;
mixer gate_output_7_483(.a(output_8_483), .b(output_8_4), .y(output_7_483));
wire output_1_484, output_1_5, output_0_484;
mixer gate_output_0_484(.a(output_1_484), .b(output_1_5), .y(output_0_484));
wire output_2_484, output_2_5, output_1_484;
mixer gate_output_1_484(.a(output_2_484), .b(output_2_5), .y(output_1_484));
wire output_3_484, output_3_5, output_2_484;
mixer gate_output_2_484(.a(output_3_484), .b(output_3_5), .y(output_2_484));
wire output_4_484, output_4_5, output_3_484;
mixer gate_output_3_484(.a(output_4_484), .b(output_4_5), .y(output_3_484));
wire output_5_484, output_5_5, output_4_484;
mixer gate_output_4_484(.a(output_5_484), .b(output_5_5), .y(output_4_484));
wire output_6_484, output_6_5, output_5_484;
mixer gate_output_5_484(.a(output_6_484), .b(output_6_5), .y(output_5_484));
wire output_7_484, output_7_5, output_6_484;
mixer gate_output_6_484(.a(output_7_484), .b(output_7_5), .y(output_6_484));
wire output_8_484, output_8_5, output_7_484;
mixer gate_output_7_484(.a(output_8_484), .b(output_8_5), .y(output_7_484));
wire output_1_485, output_1_6, output_0_485;
mixer gate_output_0_485(.a(output_1_485), .b(output_1_6), .y(output_0_485));
wire output_2_485, output_2_6, output_1_485;
mixer gate_output_1_485(.a(output_2_485), .b(output_2_6), .y(output_1_485));
wire output_3_485, output_3_6, output_2_485;
mixer gate_output_2_485(.a(output_3_485), .b(output_3_6), .y(output_2_485));
wire output_4_485, output_4_6, output_3_485;
mixer gate_output_3_485(.a(output_4_485), .b(output_4_6), .y(output_3_485));
wire output_5_485, output_5_6, output_4_485;
mixer gate_output_4_485(.a(output_5_485), .b(output_5_6), .y(output_4_485));
wire output_6_485, output_6_6, output_5_485;
mixer gate_output_5_485(.a(output_6_485), .b(output_6_6), .y(output_5_485));
wire output_7_485, output_7_6, output_6_485;
mixer gate_output_6_485(.a(output_7_485), .b(output_7_6), .y(output_6_485));
wire output_8_485, output_8_6, output_7_485;
mixer gate_output_7_485(.a(output_8_485), .b(output_8_6), .y(output_7_485));
wire output_1_486, output_1_7, output_0_486;
mixer gate_output_0_486(.a(output_1_486), .b(output_1_7), .y(output_0_486));
wire output_2_486, output_2_7, output_1_486;
mixer gate_output_1_486(.a(output_2_486), .b(output_2_7), .y(output_1_486));
wire output_3_486, output_3_7, output_2_486;
mixer gate_output_2_486(.a(output_3_486), .b(output_3_7), .y(output_2_486));
wire output_4_486, output_4_7, output_3_486;
mixer gate_output_3_486(.a(output_4_486), .b(output_4_7), .y(output_3_486));
wire output_5_486, output_5_7, output_4_486;
mixer gate_output_4_486(.a(output_5_486), .b(output_5_7), .y(output_4_486));
wire output_6_486, output_6_7, output_5_486;
mixer gate_output_5_486(.a(output_6_486), .b(output_6_7), .y(output_5_486));
wire output_7_486, output_7_7, output_6_486;
mixer gate_output_6_486(.a(output_7_486), .b(output_7_7), .y(output_6_486));
wire output_8_486, output_8_7, output_7_486;
mixer gate_output_7_486(.a(output_8_486), .b(output_8_7), .y(output_7_486));
wire output_1_487, output_1_0, output_0_487;
mixer gate_output_0_487(.a(output_1_487), .b(output_1_0), .y(output_0_487));
wire output_2_487, output_2_0, output_1_487;
mixer gate_output_1_487(.a(output_2_487), .b(output_2_0), .y(output_1_487));
wire output_3_487, output_3_0, output_2_487;
mixer gate_output_2_487(.a(output_3_487), .b(output_3_0), .y(output_2_487));
wire output_4_487, output_4_0, output_3_487;
mixer gate_output_3_487(.a(output_4_487), .b(output_4_0), .y(output_3_487));
wire output_5_487, output_5_0, output_4_487;
mixer gate_output_4_487(.a(output_5_487), .b(output_5_0), .y(output_4_487));
wire output_6_487, output_6_0, output_5_487;
mixer gate_output_5_487(.a(output_6_487), .b(output_6_0), .y(output_5_487));
wire output_7_487, output_7_0, output_6_487;
mixer gate_output_6_487(.a(output_7_487), .b(output_7_0), .y(output_6_487));
wire output_8_487, output_8_0, output_7_487;
mixer gate_output_7_487(.a(output_8_487), .b(output_8_0), .y(output_7_487));
wire output_1_488, output_1_1, output_0_488;
mixer gate_output_0_488(.a(output_1_488), .b(output_1_1), .y(output_0_488));
wire output_2_488, output_2_1, output_1_488;
mixer gate_output_1_488(.a(output_2_488), .b(output_2_1), .y(output_1_488));
wire output_3_488, output_3_1, output_2_488;
mixer gate_output_2_488(.a(output_3_488), .b(output_3_1), .y(output_2_488));
wire output_4_488, output_4_1, output_3_488;
mixer gate_output_3_488(.a(output_4_488), .b(output_4_1), .y(output_3_488));
wire output_5_488, output_5_1, output_4_488;
mixer gate_output_4_488(.a(output_5_488), .b(output_5_1), .y(output_4_488));
wire output_6_488, output_6_1, output_5_488;
mixer gate_output_5_488(.a(output_6_488), .b(output_6_1), .y(output_5_488));
wire output_7_488, output_7_1, output_6_488;
mixer gate_output_6_488(.a(output_7_488), .b(output_7_1), .y(output_6_488));
wire output_8_488, output_8_1, output_7_488;
mixer gate_output_7_488(.a(output_8_488), .b(output_8_1), .y(output_7_488));
wire output_1_489, output_1_2, output_0_489;
mixer gate_output_0_489(.a(output_1_489), .b(output_1_2), .y(output_0_489));
wire output_2_489, output_2_2, output_1_489;
mixer gate_output_1_489(.a(output_2_489), .b(output_2_2), .y(output_1_489));
wire output_3_489, output_3_2, output_2_489;
mixer gate_output_2_489(.a(output_3_489), .b(output_3_2), .y(output_2_489));
wire output_4_489, output_4_2, output_3_489;
mixer gate_output_3_489(.a(output_4_489), .b(output_4_2), .y(output_3_489));
wire output_5_489, output_5_2, output_4_489;
mixer gate_output_4_489(.a(output_5_489), .b(output_5_2), .y(output_4_489));
wire output_6_489, output_6_2, output_5_489;
mixer gate_output_5_489(.a(output_6_489), .b(output_6_2), .y(output_5_489));
wire output_7_489, output_7_2, output_6_489;
mixer gate_output_6_489(.a(output_7_489), .b(output_7_2), .y(output_6_489));
wire output_8_489, output_8_2, output_7_489;
mixer gate_output_7_489(.a(output_8_489), .b(output_8_2), .y(output_7_489));
wire output_1_490, output_1_3, output_0_490;
mixer gate_output_0_490(.a(output_1_490), .b(output_1_3), .y(output_0_490));
wire output_2_490, output_2_3, output_1_490;
mixer gate_output_1_490(.a(output_2_490), .b(output_2_3), .y(output_1_490));
wire output_3_490, output_3_3, output_2_490;
mixer gate_output_2_490(.a(output_3_490), .b(output_3_3), .y(output_2_490));
wire output_4_490, output_4_3, output_3_490;
mixer gate_output_3_490(.a(output_4_490), .b(output_4_3), .y(output_3_490));
wire output_5_490, output_5_3, output_4_490;
mixer gate_output_4_490(.a(output_5_490), .b(output_5_3), .y(output_4_490));
wire output_6_490, output_6_3, output_5_490;
mixer gate_output_5_490(.a(output_6_490), .b(output_6_3), .y(output_5_490));
wire output_7_490, output_7_3, output_6_490;
mixer gate_output_6_490(.a(output_7_490), .b(output_7_3), .y(output_6_490));
wire output_8_490, output_8_3, output_7_490;
mixer gate_output_7_490(.a(output_8_490), .b(output_8_3), .y(output_7_490));
wire output_1_491, output_1_4, output_0_491;
mixer gate_output_0_491(.a(output_1_491), .b(output_1_4), .y(output_0_491));
wire output_2_491, output_2_4, output_1_491;
mixer gate_output_1_491(.a(output_2_491), .b(output_2_4), .y(output_1_491));
wire output_3_491, output_3_4, output_2_491;
mixer gate_output_2_491(.a(output_3_491), .b(output_3_4), .y(output_2_491));
wire output_4_491, output_4_4, output_3_491;
mixer gate_output_3_491(.a(output_4_491), .b(output_4_4), .y(output_3_491));
wire output_5_491, output_5_4, output_4_491;
mixer gate_output_4_491(.a(output_5_491), .b(output_5_4), .y(output_4_491));
wire output_6_491, output_6_4, output_5_491;
mixer gate_output_5_491(.a(output_6_491), .b(output_6_4), .y(output_5_491));
wire output_7_491, output_7_4, output_6_491;
mixer gate_output_6_491(.a(output_7_491), .b(output_7_4), .y(output_6_491));
wire output_8_491, output_8_4, output_7_491;
mixer gate_output_7_491(.a(output_8_491), .b(output_8_4), .y(output_7_491));
wire output_1_492, output_1_5, output_0_492;
mixer gate_output_0_492(.a(output_1_492), .b(output_1_5), .y(output_0_492));
wire output_2_492, output_2_5, output_1_492;
mixer gate_output_1_492(.a(output_2_492), .b(output_2_5), .y(output_1_492));
wire output_3_492, output_3_5, output_2_492;
mixer gate_output_2_492(.a(output_3_492), .b(output_3_5), .y(output_2_492));
wire output_4_492, output_4_5, output_3_492;
mixer gate_output_3_492(.a(output_4_492), .b(output_4_5), .y(output_3_492));
wire output_5_492, output_5_5, output_4_492;
mixer gate_output_4_492(.a(output_5_492), .b(output_5_5), .y(output_4_492));
wire output_6_492, output_6_5, output_5_492;
mixer gate_output_5_492(.a(output_6_492), .b(output_6_5), .y(output_5_492));
wire output_7_492, output_7_5, output_6_492;
mixer gate_output_6_492(.a(output_7_492), .b(output_7_5), .y(output_6_492));
wire output_8_492, output_8_5, output_7_492;
mixer gate_output_7_492(.a(output_8_492), .b(output_8_5), .y(output_7_492));
wire output_1_493, output_1_6, output_0_493;
mixer gate_output_0_493(.a(output_1_493), .b(output_1_6), .y(output_0_493));
wire output_2_493, output_2_6, output_1_493;
mixer gate_output_1_493(.a(output_2_493), .b(output_2_6), .y(output_1_493));
wire output_3_493, output_3_6, output_2_493;
mixer gate_output_2_493(.a(output_3_493), .b(output_3_6), .y(output_2_493));
wire output_4_493, output_4_6, output_3_493;
mixer gate_output_3_493(.a(output_4_493), .b(output_4_6), .y(output_3_493));
wire output_5_493, output_5_6, output_4_493;
mixer gate_output_4_493(.a(output_5_493), .b(output_5_6), .y(output_4_493));
wire output_6_493, output_6_6, output_5_493;
mixer gate_output_5_493(.a(output_6_493), .b(output_6_6), .y(output_5_493));
wire output_7_493, output_7_6, output_6_493;
mixer gate_output_6_493(.a(output_7_493), .b(output_7_6), .y(output_6_493));
wire output_8_493, output_8_6, output_7_493;
mixer gate_output_7_493(.a(output_8_493), .b(output_8_6), .y(output_7_493));
wire output_1_494, output_1_7, output_0_494;
mixer gate_output_0_494(.a(output_1_494), .b(output_1_7), .y(output_0_494));
wire output_2_494, output_2_7, output_1_494;
mixer gate_output_1_494(.a(output_2_494), .b(output_2_7), .y(output_1_494));
wire output_3_494, output_3_7, output_2_494;
mixer gate_output_2_494(.a(output_3_494), .b(output_3_7), .y(output_2_494));
wire output_4_494, output_4_7, output_3_494;
mixer gate_output_3_494(.a(output_4_494), .b(output_4_7), .y(output_3_494));
wire output_5_494, output_5_7, output_4_494;
mixer gate_output_4_494(.a(output_5_494), .b(output_5_7), .y(output_4_494));
wire output_6_494, output_6_7, output_5_494;
mixer gate_output_5_494(.a(output_6_494), .b(output_6_7), .y(output_5_494));
wire output_7_494, output_7_7, output_6_494;
mixer gate_output_6_494(.a(output_7_494), .b(output_7_7), .y(output_6_494));
wire output_8_494, output_8_7, output_7_494;
mixer gate_output_7_494(.a(output_8_494), .b(output_8_7), .y(output_7_494));
wire output_1_495, output_1_0, output_0_495;
mixer gate_output_0_495(.a(output_1_495), .b(output_1_0), .y(output_0_495));
wire output_2_495, output_2_0, output_1_495;
mixer gate_output_1_495(.a(output_2_495), .b(output_2_0), .y(output_1_495));
wire output_3_495, output_3_0, output_2_495;
mixer gate_output_2_495(.a(output_3_495), .b(output_3_0), .y(output_2_495));
wire output_4_495, output_4_0, output_3_495;
mixer gate_output_3_495(.a(output_4_495), .b(output_4_0), .y(output_3_495));
wire output_5_495, output_5_0, output_4_495;
mixer gate_output_4_495(.a(output_5_495), .b(output_5_0), .y(output_4_495));
wire output_6_495, output_6_0, output_5_495;
mixer gate_output_5_495(.a(output_6_495), .b(output_6_0), .y(output_5_495));
wire output_7_495, output_7_0, output_6_495;
mixer gate_output_6_495(.a(output_7_495), .b(output_7_0), .y(output_6_495));
wire output_8_495, output_8_0, output_7_495;
mixer gate_output_7_495(.a(output_8_495), .b(output_8_0), .y(output_7_495));
wire output_1_496, output_1_1, output_0_496;
mixer gate_output_0_496(.a(output_1_496), .b(output_1_1), .y(output_0_496));
wire output_2_496, output_2_1, output_1_496;
mixer gate_output_1_496(.a(output_2_496), .b(output_2_1), .y(output_1_496));
wire output_3_496, output_3_1, output_2_496;
mixer gate_output_2_496(.a(output_3_496), .b(output_3_1), .y(output_2_496));
wire output_4_496, output_4_1, output_3_496;
mixer gate_output_3_496(.a(output_4_496), .b(output_4_1), .y(output_3_496));
wire output_5_496, output_5_1, output_4_496;
mixer gate_output_4_496(.a(output_5_496), .b(output_5_1), .y(output_4_496));
wire output_6_496, output_6_1, output_5_496;
mixer gate_output_5_496(.a(output_6_496), .b(output_6_1), .y(output_5_496));
wire output_7_496, output_7_1, output_6_496;
mixer gate_output_6_496(.a(output_7_496), .b(output_7_1), .y(output_6_496));
wire output_8_496, output_8_1, output_7_496;
mixer gate_output_7_496(.a(output_8_496), .b(output_8_1), .y(output_7_496));
wire output_1_497, output_1_2, output_0_497;
mixer gate_output_0_497(.a(output_1_497), .b(output_1_2), .y(output_0_497));
wire output_2_497, output_2_2, output_1_497;
mixer gate_output_1_497(.a(output_2_497), .b(output_2_2), .y(output_1_497));
wire output_3_497, output_3_2, output_2_497;
mixer gate_output_2_497(.a(output_3_497), .b(output_3_2), .y(output_2_497));
wire output_4_497, output_4_2, output_3_497;
mixer gate_output_3_497(.a(output_4_497), .b(output_4_2), .y(output_3_497));
wire output_5_497, output_5_2, output_4_497;
mixer gate_output_4_497(.a(output_5_497), .b(output_5_2), .y(output_4_497));
wire output_6_497, output_6_2, output_5_497;
mixer gate_output_5_497(.a(output_6_497), .b(output_6_2), .y(output_5_497));
wire output_7_497, output_7_2, output_6_497;
mixer gate_output_6_497(.a(output_7_497), .b(output_7_2), .y(output_6_497));
wire output_8_497, output_8_2, output_7_497;
mixer gate_output_7_497(.a(output_8_497), .b(output_8_2), .y(output_7_497));
wire output_1_498, output_1_3, output_0_498;
mixer gate_output_0_498(.a(output_1_498), .b(output_1_3), .y(output_0_498));
wire output_2_498, output_2_3, output_1_498;
mixer gate_output_1_498(.a(output_2_498), .b(output_2_3), .y(output_1_498));
wire output_3_498, output_3_3, output_2_498;
mixer gate_output_2_498(.a(output_3_498), .b(output_3_3), .y(output_2_498));
wire output_4_498, output_4_3, output_3_498;
mixer gate_output_3_498(.a(output_4_498), .b(output_4_3), .y(output_3_498));
wire output_5_498, output_5_3, output_4_498;
mixer gate_output_4_498(.a(output_5_498), .b(output_5_3), .y(output_4_498));
wire output_6_498, output_6_3, output_5_498;
mixer gate_output_5_498(.a(output_6_498), .b(output_6_3), .y(output_5_498));
wire output_7_498, output_7_3, output_6_498;
mixer gate_output_6_498(.a(output_7_498), .b(output_7_3), .y(output_6_498));
wire output_8_498, output_8_3, output_7_498;
mixer gate_output_7_498(.a(output_8_498), .b(output_8_3), .y(output_7_498));
wire output_1_499, output_1_4, output_0_499;
mixer gate_output_0_499(.a(output_1_499), .b(output_1_4), .y(output_0_499));
wire output_2_499, output_2_4, output_1_499;
mixer gate_output_1_499(.a(output_2_499), .b(output_2_4), .y(output_1_499));
wire output_3_499, output_3_4, output_2_499;
mixer gate_output_2_499(.a(output_3_499), .b(output_3_4), .y(output_2_499));
wire output_4_499, output_4_4, output_3_499;
mixer gate_output_3_499(.a(output_4_499), .b(output_4_4), .y(output_3_499));
wire output_5_499, output_5_4, output_4_499;
mixer gate_output_4_499(.a(output_5_499), .b(output_5_4), .y(output_4_499));
wire output_6_499, output_6_4, output_5_499;
mixer gate_output_5_499(.a(output_6_499), .b(output_6_4), .y(output_5_499));
wire output_7_499, output_7_4, output_6_499;
mixer gate_output_6_499(.a(output_7_499), .b(output_7_4), .y(output_6_499));
wire output_8_499, output_8_4, output_7_499;
mixer gate_output_7_499(.a(output_8_499), .b(output_8_4), .y(output_7_499));
wire output_1_500, output_1_5, output_0_500;
mixer gate_output_0_500(.a(output_1_500), .b(output_1_5), .y(output_0_500));
wire output_2_500, output_2_5, output_1_500;
mixer gate_output_1_500(.a(output_2_500), .b(output_2_5), .y(output_1_500));
wire output_3_500, output_3_5, output_2_500;
mixer gate_output_2_500(.a(output_3_500), .b(output_3_5), .y(output_2_500));
wire output_4_500, output_4_5, output_3_500;
mixer gate_output_3_500(.a(output_4_500), .b(output_4_5), .y(output_3_500));
wire output_5_500, output_5_5, output_4_500;
mixer gate_output_4_500(.a(output_5_500), .b(output_5_5), .y(output_4_500));
wire output_6_500, output_6_5, output_5_500;
mixer gate_output_5_500(.a(output_6_500), .b(output_6_5), .y(output_5_500));
wire output_7_500, output_7_5, output_6_500;
mixer gate_output_6_500(.a(output_7_500), .b(output_7_5), .y(output_6_500));
wire output_8_500, output_8_5, output_7_500;
mixer gate_output_7_500(.a(output_8_500), .b(output_8_5), .y(output_7_500));
wire output_1_501, output_1_6, output_0_501;
mixer gate_output_0_501(.a(output_1_501), .b(output_1_6), .y(output_0_501));
wire output_2_501, output_2_6, output_1_501;
mixer gate_output_1_501(.a(output_2_501), .b(output_2_6), .y(output_1_501));
wire output_3_501, output_3_6, output_2_501;
mixer gate_output_2_501(.a(output_3_501), .b(output_3_6), .y(output_2_501));
wire output_4_501, output_4_6, output_3_501;
mixer gate_output_3_501(.a(output_4_501), .b(output_4_6), .y(output_3_501));
wire output_5_501, output_5_6, output_4_501;
mixer gate_output_4_501(.a(output_5_501), .b(output_5_6), .y(output_4_501));
wire output_6_501, output_6_6, output_5_501;
mixer gate_output_5_501(.a(output_6_501), .b(output_6_6), .y(output_5_501));
wire output_7_501, output_7_6, output_6_501;
mixer gate_output_6_501(.a(output_7_501), .b(output_7_6), .y(output_6_501));
wire output_8_501, output_8_6, output_7_501;
mixer gate_output_7_501(.a(output_8_501), .b(output_8_6), .y(output_7_501));
wire output_1_502, output_1_7, output_0_502;
mixer gate_output_0_502(.a(output_1_502), .b(output_1_7), .y(output_0_502));
wire output_2_502, output_2_7, output_1_502;
mixer gate_output_1_502(.a(output_2_502), .b(output_2_7), .y(output_1_502));
wire output_3_502, output_3_7, output_2_502;
mixer gate_output_2_502(.a(output_3_502), .b(output_3_7), .y(output_2_502));
wire output_4_502, output_4_7, output_3_502;
mixer gate_output_3_502(.a(output_4_502), .b(output_4_7), .y(output_3_502));
wire output_5_502, output_5_7, output_4_502;
mixer gate_output_4_502(.a(output_5_502), .b(output_5_7), .y(output_4_502));
wire output_6_502, output_6_7, output_5_502;
mixer gate_output_5_502(.a(output_6_502), .b(output_6_7), .y(output_5_502));
wire output_7_502, output_7_7, output_6_502;
mixer gate_output_6_502(.a(output_7_502), .b(output_7_7), .y(output_6_502));
wire output_8_502, output_8_7, output_7_502;
mixer gate_output_7_502(.a(output_8_502), .b(output_8_7), .y(output_7_502));
wire output_1_503, output_1_0, output_0_503;
mixer gate_output_0_503(.a(output_1_503), .b(output_1_0), .y(output_0_503));
wire output_2_503, output_2_0, output_1_503;
mixer gate_output_1_503(.a(output_2_503), .b(output_2_0), .y(output_1_503));
wire output_3_503, output_3_0, output_2_503;
mixer gate_output_2_503(.a(output_3_503), .b(output_3_0), .y(output_2_503));
wire output_4_503, output_4_0, output_3_503;
mixer gate_output_3_503(.a(output_4_503), .b(output_4_0), .y(output_3_503));
wire output_5_503, output_5_0, output_4_503;
mixer gate_output_4_503(.a(output_5_503), .b(output_5_0), .y(output_4_503));
wire output_6_503, output_6_0, output_5_503;
mixer gate_output_5_503(.a(output_6_503), .b(output_6_0), .y(output_5_503));
wire output_7_503, output_7_0, output_6_503;
mixer gate_output_6_503(.a(output_7_503), .b(output_7_0), .y(output_6_503));
wire output_8_503, output_8_0, output_7_503;
mixer gate_output_7_503(.a(output_8_503), .b(output_8_0), .y(output_7_503));
wire output_1_504, output_1_1, output_0_504;
mixer gate_output_0_504(.a(output_1_504), .b(output_1_1), .y(output_0_504));
wire output_2_504, output_2_1, output_1_504;
mixer gate_output_1_504(.a(output_2_504), .b(output_2_1), .y(output_1_504));
wire output_3_504, output_3_1, output_2_504;
mixer gate_output_2_504(.a(output_3_504), .b(output_3_1), .y(output_2_504));
wire output_4_504, output_4_1, output_3_504;
mixer gate_output_3_504(.a(output_4_504), .b(output_4_1), .y(output_3_504));
wire output_5_504, output_5_1, output_4_504;
mixer gate_output_4_504(.a(output_5_504), .b(output_5_1), .y(output_4_504));
wire output_6_504, output_6_1, output_5_504;
mixer gate_output_5_504(.a(output_6_504), .b(output_6_1), .y(output_5_504));
wire output_7_504, output_7_1, output_6_504;
mixer gate_output_6_504(.a(output_7_504), .b(output_7_1), .y(output_6_504));
wire output_8_504, output_8_1, output_7_504;
mixer gate_output_7_504(.a(output_8_504), .b(output_8_1), .y(output_7_504));
wire output_1_505, output_1_2, output_0_505;
mixer gate_output_0_505(.a(output_1_505), .b(output_1_2), .y(output_0_505));
wire output_2_505, output_2_2, output_1_505;
mixer gate_output_1_505(.a(output_2_505), .b(output_2_2), .y(output_1_505));
wire output_3_505, output_3_2, output_2_505;
mixer gate_output_2_505(.a(output_3_505), .b(output_3_2), .y(output_2_505));
wire output_4_505, output_4_2, output_3_505;
mixer gate_output_3_505(.a(output_4_505), .b(output_4_2), .y(output_3_505));
wire output_5_505, output_5_2, output_4_505;
mixer gate_output_4_505(.a(output_5_505), .b(output_5_2), .y(output_4_505));
wire output_6_505, output_6_2, output_5_505;
mixer gate_output_5_505(.a(output_6_505), .b(output_6_2), .y(output_5_505));
wire output_7_505, output_7_2, output_6_505;
mixer gate_output_6_505(.a(output_7_505), .b(output_7_2), .y(output_6_505));
wire output_8_505, output_8_2, output_7_505;
mixer gate_output_7_505(.a(output_8_505), .b(output_8_2), .y(output_7_505));
wire output_1_506, output_1_3, output_0_506;
mixer gate_output_0_506(.a(output_1_506), .b(output_1_3), .y(output_0_506));
wire output_2_506, output_2_3, output_1_506;
mixer gate_output_1_506(.a(output_2_506), .b(output_2_3), .y(output_1_506));
wire output_3_506, output_3_3, output_2_506;
mixer gate_output_2_506(.a(output_3_506), .b(output_3_3), .y(output_2_506));
wire output_4_506, output_4_3, output_3_506;
mixer gate_output_3_506(.a(output_4_506), .b(output_4_3), .y(output_3_506));
wire output_5_506, output_5_3, output_4_506;
mixer gate_output_4_506(.a(output_5_506), .b(output_5_3), .y(output_4_506));
wire output_6_506, output_6_3, output_5_506;
mixer gate_output_5_506(.a(output_6_506), .b(output_6_3), .y(output_5_506));
wire output_7_506, output_7_3, output_6_506;
mixer gate_output_6_506(.a(output_7_506), .b(output_7_3), .y(output_6_506));
wire output_8_506, output_8_3, output_7_506;
mixer gate_output_7_506(.a(output_8_506), .b(output_8_3), .y(output_7_506));
wire output_1_507, output_1_4, output_0_507;
mixer gate_output_0_507(.a(output_1_507), .b(output_1_4), .y(output_0_507));
wire output_2_507, output_2_4, output_1_507;
mixer gate_output_1_507(.a(output_2_507), .b(output_2_4), .y(output_1_507));
wire output_3_507, output_3_4, output_2_507;
mixer gate_output_2_507(.a(output_3_507), .b(output_3_4), .y(output_2_507));
wire output_4_507, output_4_4, output_3_507;
mixer gate_output_3_507(.a(output_4_507), .b(output_4_4), .y(output_3_507));
wire output_5_507, output_5_4, output_4_507;
mixer gate_output_4_507(.a(output_5_507), .b(output_5_4), .y(output_4_507));
wire output_6_507, output_6_4, output_5_507;
mixer gate_output_5_507(.a(output_6_507), .b(output_6_4), .y(output_5_507));
wire output_7_507, output_7_4, output_6_507;
mixer gate_output_6_507(.a(output_7_507), .b(output_7_4), .y(output_6_507));
wire output_8_507, output_8_4, output_7_507;
mixer gate_output_7_507(.a(output_8_507), .b(output_8_4), .y(output_7_507));
wire output_1_508, output_1_5, output_0_508;
mixer gate_output_0_508(.a(output_1_508), .b(output_1_5), .y(output_0_508));
wire output_2_508, output_2_5, output_1_508;
mixer gate_output_1_508(.a(output_2_508), .b(output_2_5), .y(output_1_508));
wire output_3_508, output_3_5, output_2_508;
mixer gate_output_2_508(.a(output_3_508), .b(output_3_5), .y(output_2_508));
wire output_4_508, output_4_5, output_3_508;
mixer gate_output_3_508(.a(output_4_508), .b(output_4_5), .y(output_3_508));
wire output_5_508, output_5_5, output_4_508;
mixer gate_output_4_508(.a(output_5_508), .b(output_5_5), .y(output_4_508));
wire output_6_508, output_6_5, output_5_508;
mixer gate_output_5_508(.a(output_6_508), .b(output_6_5), .y(output_5_508));
wire output_7_508, output_7_5, output_6_508;
mixer gate_output_6_508(.a(output_7_508), .b(output_7_5), .y(output_6_508));
wire output_8_508, output_8_5, output_7_508;
mixer gate_output_7_508(.a(output_8_508), .b(output_8_5), .y(output_7_508));
wire output_1_509, output_1_6, output_0_509;
mixer gate_output_0_509(.a(output_1_509), .b(output_1_6), .y(output_0_509));
wire output_2_509, output_2_6, output_1_509;
mixer gate_output_1_509(.a(output_2_509), .b(output_2_6), .y(output_1_509));
wire output_3_509, output_3_6, output_2_509;
mixer gate_output_2_509(.a(output_3_509), .b(output_3_6), .y(output_2_509));
wire output_4_509, output_4_6, output_3_509;
mixer gate_output_3_509(.a(output_4_509), .b(output_4_6), .y(output_3_509));
wire output_5_509, output_5_6, output_4_509;
mixer gate_output_4_509(.a(output_5_509), .b(output_5_6), .y(output_4_509));
wire output_6_509, output_6_6, output_5_509;
mixer gate_output_5_509(.a(output_6_509), .b(output_6_6), .y(output_5_509));
wire output_7_509, output_7_6, output_6_509;
mixer gate_output_6_509(.a(output_7_509), .b(output_7_6), .y(output_6_509));
wire output_8_509, output_8_6, output_7_509;
mixer gate_output_7_509(.a(output_8_509), .b(output_8_6), .y(output_7_509));
wire output_1_510, output_1_7, output_0_510;
mixer gate_output_0_510(.a(output_1_510), .b(output_1_7), .y(output_0_510));
wire output_2_510, output_2_7, output_1_510;
mixer gate_output_1_510(.a(output_2_510), .b(output_2_7), .y(output_1_510));
wire output_3_510, output_3_7, output_2_510;
mixer gate_output_2_510(.a(output_3_510), .b(output_3_7), .y(output_2_510));
wire output_4_510, output_4_7, output_3_510;
mixer gate_output_3_510(.a(output_4_510), .b(output_4_7), .y(output_3_510));
wire output_5_510, output_5_7, output_4_510;
mixer gate_output_4_510(.a(output_5_510), .b(output_5_7), .y(output_4_510));
wire output_6_510, output_6_7, output_5_510;
mixer gate_output_5_510(.a(output_6_510), .b(output_6_7), .y(output_5_510));
wire output_7_510, output_7_7, output_6_510;
mixer gate_output_6_510(.a(output_7_510), .b(output_7_7), .y(output_6_510));
wire output_8_510, output_8_7, output_7_510;
mixer gate_output_7_510(.a(output_8_510), .b(output_8_7), .y(output_7_510));
wire output_1_511, output_1_0, output_0_511;
mixer gate_output_0_511(.a(output_1_511), .b(output_1_0), .y(output_0_511));
wire output_2_511, output_2_0, output_1_511;
mixer gate_output_1_511(.a(output_2_511), .b(output_2_0), .y(output_1_511));
wire output_3_511, output_3_0, output_2_511;
mixer gate_output_2_511(.a(output_3_511), .b(output_3_0), .y(output_2_511));
wire output_4_511, output_4_0, output_3_511;
mixer gate_output_3_511(.a(output_4_511), .b(output_4_0), .y(output_3_511));
wire output_5_511, output_5_0, output_4_511;
mixer gate_output_4_511(.a(output_5_511), .b(output_5_0), .y(output_4_511));
wire output_6_511, output_6_0, output_5_511;
mixer gate_output_5_511(.a(output_6_511), .b(output_6_0), .y(output_5_511));
wire output_7_511, output_7_0, output_6_511;
mixer gate_output_6_511(.a(output_7_511), .b(output_7_0), .y(output_6_511));
wire output_8_511, output_8_0, output_7_511;
mixer gate_output_7_511(.a(output_8_511), .b(output_8_0), .y(output_7_511));
assign output_0 = output_0_0;
wire output_0_512;
assign output_0_512 = input_0;
assign output_1 = output_1_0;
wire output_1_512;
assign output_1_512 = input_1;
assign output_2 = output_2_0;
wire output_2_512;
assign output_2_512 = input_2;
assign output_3 = output_3_0;
wire output_3_512;
assign output_3_512 = input_3;
assign output_4 = output_4_0;
wire output_4_512;
assign output_4_512 = input_4;
assign output_5 = output_5_0;
wire output_5_512;
assign output_5_512 = input_5;
assign output_6 = output_6_0;
wire output_6_512;
assign output_6_512 = input_6;
assign output_7 = output_7_0;
wire output_7_512;
assign output_7_512 = input_7;
endmodule
