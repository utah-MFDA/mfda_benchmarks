module fanout2_braid_16_16 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,output output_8,output output_9,output output_10,output output_11,output output_12,output output_13,output output_14,output output_15,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_9_0, output_9_1, output_8_0;
mixer gate_output_8_0(.a(output_9_0), .b(output_9_1), .y(output_8_0));
wire output_10_0, output_10_1, output_9_0;
mixer gate_output_9_0(.a(output_10_0), .b(output_10_1), .y(output_9_0));
wire output_11_0, output_11_1, output_10_0;
mixer gate_output_10_0(.a(output_11_0), .b(output_11_1), .y(output_10_0));
wire output_12_0, output_12_1, output_11_0;
mixer gate_output_11_0(.a(output_12_0), .b(output_12_1), .y(output_11_0));
wire output_13_0, output_13_1, output_12_0;
mixer gate_output_12_0(.a(output_13_0), .b(output_13_1), .y(output_12_0));
wire output_14_0, output_14_1, output_13_0;
mixer gate_output_13_0(.a(output_14_0), .b(output_14_1), .y(output_13_0));
wire output_15_0, output_15_1, output_14_0;
mixer gate_output_14_0(.a(output_15_0), .b(output_15_1), .y(output_14_0));
wire output_16_0, output_16_1, output_15_0;
mixer gate_output_15_0(.a(output_16_0), .b(output_16_1), .y(output_15_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_9_1, output_9_2, output_8_1;
mixer gate_output_8_1(.a(output_9_1), .b(output_9_2), .y(output_8_1));
wire output_10_1, output_10_2, output_9_1;
mixer gate_output_9_1(.a(output_10_1), .b(output_10_2), .y(output_9_1));
wire output_11_1, output_11_2, output_10_1;
mixer gate_output_10_1(.a(output_11_1), .b(output_11_2), .y(output_10_1));
wire output_12_1, output_12_2, output_11_1;
mixer gate_output_11_1(.a(output_12_1), .b(output_12_2), .y(output_11_1));
wire output_13_1, output_13_2, output_12_1;
mixer gate_output_12_1(.a(output_13_1), .b(output_13_2), .y(output_12_1));
wire output_14_1, output_14_2, output_13_1;
mixer gate_output_13_1(.a(output_14_1), .b(output_14_2), .y(output_13_1));
wire output_15_1, output_15_2, output_14_1;
mixer gate_output_14_1(.a(output_15_1), .b(output_15_2), .y(output_14_1));
wire output_16_1, output_16_2, output_15_1;
mixer gate_output_15_1(.a(output_16_1), .b(output_16_2), .y(output_15_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_9_2, output_9_3, output_8_2;
mixer gate_output_8_2(.a(output_9_2), .b(output_9_3), .y(output_8_2));
wire output_10_2, output_10_3, output_9_2;
mixer gate_output_9_2(.a(output_10_2), .b(output_10_3), .y(output_9_2));
wire output_11_2, output_11_3, output_10_2;
mixer gate_output_10_2(.a(output_11_2), .b(output_11_3), .y(output_10_2));
wire output_12_2, output_12_3, output_11_2;
mixer gate_output_11_2(.a(output_12_2), .b(output_12_3), .y(output_11_2));
wire output_13_2, output_13_3, output_12_2;
mixer gate_output_12_2(.a(output_13_2), .b(output_13_3), .y(output_12_2));
wire output_14_2, output_14_3, output_13_2;
mixer gate_output_13_2(.a(output_14_2), .b(output_14_3), .y(output_13_2));
wire output_15_2, output_15_3, output_14_2;
mixer gate_output_14_2(.a(output_15_2), .b(output_15_3), .y(output_14_2));
wire output_16_2, output_16_3, output_15_2;
mixer gate_output_15_2(.a(output_16_2), .b(output_16_3), .y(output_15_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_9_3, output_9_4, output_8_3;
mixer gate_output_8_3(.a(output_9_3), .b(output_9_4), .y(output_8_3));
wire output_10_3, output_10_4, output_9_3;
mixer gate_output_9_3(.a(output_10_3), .b(output_10_4), .y(output_9_3));
wire output_11_3, output_11_4, output_10_3;
mixer gate_output_10_3(.a(output_11_3), .b(output_11_4), .y(output_10_3));
wire output_12_3, output_12_4, output_11_3;
mixer gate_output_11_3(.a(output_12_3), .b(output_12_4), .y(output_11_3));
wire output_13_3, output_13_4, output_12_3;
mixer gate_output_12_3(.a(output_13_3), .b(output_13_4), .y(output_12_3));
wire output_14_3, output_14_4, output_13_3;
mixer gate_output_13_3(.a(output_14_3), .b(output_14_4), .y(output_13_3));
wire output_15_3, output_15_4, output_14_3;
mixer gate_output_14_3(.a(output_15_3), .b(output_15_4), .y(output_14_3));
wire output_16_3, output_16_4, output_15_3;
mixer gate_output_15_3(.a(output_16_3), .b(output_16_4), .y(output_15_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_9_4, output_9_5, output_8_4;
mixer gate_output_8_4(.a(output_9_4), .b(output_9_5), .y(output_8_4));
wire output_10_4, output_10_5, output_9_4;
mixer gate_output_9_4(.a(output_10_4), .b(output_10_5), .y(output_9_4));
wire output_11_4, output_11_5, output_10_4;
mixer gate_output_10_4(.a(output_11_4), .b(output_11_5), .y(output_10_4));
wire output_12_4, output_12_5, output_11_4;
mixer gate_output_11_4(.a(output_12_4), .b(output_12_5), .y(output_11_4));
wire output_13_4, output_13_5, output_12_4;
mixer gate_output_12_4(.a(output_13_4), .b(output_13_5), .y(output_12_4));
wire output_14_4, output_14_5, output_13_4;
mixer gate_output_13_4(.a(output_14_4), .b(output_14_5), .y(output_13_4));
wire output_15_4, output_15_5, output_14_4;
mixer gate_output_14_4(.a(output_15_4), .b(output_15_5), .y(output_14_4));
wire output_16_4, output_16_5, output_15_4;
mixer gate_output_15_4(.a(output_16_4), .b(output_16_5), .y(output_15_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_9_5, output_9_6, output_8_5;
mixer gate_output_8_5(.a(output_9_5), .b(output_9_6), .y(output_8_5));
wire output_10_5, output_10_6, output_9_5;
mixer gate_output_9_5(.a(output_10_5), .b(output_10_6), .y(output_9_5));
wire output_11_5, output_11_6, output_10_5;
mixer gate_output_10_5(.a(output_11_5), .b(output_11_6), .y(output_10_5));
wire output_12_5, output_12_6, output_11_5;
mixer gate_output_11_5(.a(output_12_5), .b(output_12_6), .y(output_11_5));
wire output_13_5, output_13_6, output_12_5;
mixer gate_output_12_5(.a(output_13_5), .b(output_13_6), .y(output_12_5));
wire output_14_5, output_14_6, output_13_5;
mixer gate_output_13_5(.a(output_14_5), .b(output_14_6), .y(output_13_5));
wire output_15_5, output_15_6, output_14_5;
mixer gate_output_14_5(.a(output_15_5), .b(output_15_6), .y(output_14_5));
wire output_16_5, output_16_6, output_15_5;
mixer gate_output_15_5(.a(output_16_5), .b(output_16_6), .y(output_15_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_9_6, output_9_7, output_8_6;
mixer gate_output_8_6(.a(output_9_6), .b(output_9_7), .y(output_8_6));
wire output_10_6, output_10_7, output_9_6;
mixer gate_output_9_6(.a(output_10_6), .b(output_10_7), .y(output_9_6));
wire output_11_6, output_11_7, output_10_6;
mixer gate_output_10_6(.a(output_11_6), .b(output_11_7), .y(output_10_6));
wire output_12_6, output_12_7, output_11_6;
mixer gate_output_11_6(.a(output_12_6), .b(output_12_7), .y(output_11_6));
wire output_13_6, output_13_7, output_12_6;
mixer gate_output_12_6(.a(output_13_6), .b(output_13_7), .y(output_12_6));
wire output_14_6, output_14_7, output_13_6;
mixer gate_output_13_6(.a(output_14_6), .b(output_14_7), .y(output_13_6));
wire output_15_6, output_15_7, output_14_6;
mixer gate_output_14_6(.a(output_15_6), .b(output_15_7), .y(output_14_6));
wire output_16_6, output_16_7, output_15_6;
mixer gate_output_15_6(.a(output_16_6), .b(output_16_7), .y(output_15_6));
wire output_1_7, output_1_8, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_8), .y(output_0_7));
wire output_2_7, output_2_8, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_8), .y(output_1_7));
wire output_3_7, output_3_8, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_8), .y(output_2_7));
wire output_4_7, output_4_8, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_8), .y(output_3_7));
wire output_5_7, output_5_8, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_8), .y(output_4_7));
wire output_6_7, output_6_8, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_8), .y(output_5_7));
wire output_7_7, output_7_8, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_8), .y(output_6_7));
wire output_8_7, output_8_8, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_8), .y(output_7_7));
wire output_9_7, output_9_8, output_8_7;
mixer gate_output_8_7(.a(output_9_7), .b(output_9_8), .y(output_8_7));
wire output_10_7, output_10_8, output_9_7;
mixer gate_output_9_7(.a(output_10_7), .b(output_10_8), .y(output_9_7));
wire output_11_7, output_11_8, output_10_7;
mixer gate_output_10_7(.a(output_11_7), .b(output_11_8), .y(output_10_7));
wire output_12_7, output_12_8, output_11_7;
mixer gate_output_11_7(.a(output_12_7), .b(output_12_8), .y(output_11_7));
wire output_13_7, output_13_8, output_12_7;
mixer gate_output_12_7(.a(output_13_7), .b(output_13_8), .y(output_12_7));
wire output_14_7, output_14_8, output_13_7;
mixer gate_output_13_7(.a(output_14_7), .b(output_14_8), .y(output_13_7));
wire output_15_7, output_15_8, output_14_7;
mixer gate_output_14_7(.a(output_15_7), .b(output_15_8), .y(output_14_7));
wire output_16_7, output_16_8, output_15_7;
mixer gate_output_15_7(.a(output_16_7), .b(output_16_8), .y(output_15_7));
wire output_1_8, output_1_9, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_9), .y(output_0_8));
wire output_2_8, output_2_9, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_9), .y(output_1_8));
wire output_3_8, output_3_9, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_9), .y(output_2_8));
wire output_4_8, output_4_9, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_9), .y(output_3_8));
wire output_5_8, output_5_9, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_9), .y(output_4_8));
wire output_6_8, output_6_9, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_9), .y(output_5_8));
wire output_7_8, output_7_9, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_9), .y(output_6_8));
wire output_8_8, output_8_9, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_9), .y(output_7_8));
wire output_9_8, output_9_9, output_8_8;
mixer gate_output_8_8(.a(output_9_8), .b(output_9_9), .y(output_8_8));
wire output_10_8, output_10_9, output_9_8;
mixer gate_output_9_8(.a(output_10_8), .b(output_10_9), .y(output_9_8));
wire output_11_8, output_11_9, output_10_8;
mixer gate_output_10_8(.a(output_11_8), .b(output_11_9), .y(output_10_8));
wire output_12_8, output_12_9, output_11_8;
mixer gate_output_11_8(.a(output_12_8), .b(output_12_9), .y(output_11_8));
wire output_13_8, output_13_9, output_12_8;
mixer gate_output_12_8(.a(output_13_8), .b(output_13_9), .y(output_12_8));
wire output_14_8, output_14_9, output_13_8;
mixer gate_output_13_8(.a(output_14_8), .b(output_14_9), .y(output_13_8));
wire output_15_8, output_15_9, output_14_8;
mixer gate_output_14_8(.a(output_15_8), .b(output_15_9), .y(output_14_8));
wire output_16_8, output_16_9, output_15_8;
mixer gate_output_15_8(.a(output_16_8), .b(output_16_9), .y(output_15_8));
wire output_1_9, output_1_10, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_10), .y(output_0_9));
wire output_2_9, output_2_10, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_10), .y(output_1_9));
wire output_3_9, output_3_10, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_10), .y(output_2_9));
wire output_4_9, output_4_10, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_10), .y(output_3_9));
wire output_5_9, output_5_10, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_10), .y(output_4_9));
wire output_6_9, output_6_10, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_10), .y(output_5_9));
wire output_7_9, output_7_10, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_10), .y(output_6_9));
wire output_8_9, output_8_10, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_10), .y(output_7_9));
wire output_9_9, output_9_10, output_8_9;
mixer gate_output_8_9(.a(output_9_9), .b(output_9_10), .y(output_8_9));
wire output_10_9, output_10_10, output_9_9;
mixer gate_output_9_9(.a(output_10_9), .b(output_10_10), .y(output_9_9));
wire output_11_9, output_11_10, output_10_9;
mixer gate_output_10_9(.a(output_11_9), .b(output_11_10), .y(output_10_9));
wire output_12_9, output_12_10, output_11_9;
mixer gate_output_11_9(.a(output_12_9), .b(output_12_10), .y(output_11_9));
wire output_13_9, output_13_10, output_12_9;
mixer gate_output_12_9(.a(output_13_9), .b(output_13_10), .y(output_12_9));
wire output_14_9, output_14_10, output_13_9;
mixer gate_output_13_9(.a(output_14_9), .b(output_14_10), .y(output_13_9));
wire output_15_9, output_15_10, output_14_9;
mixer gate_output_14_9(.a(output_15_9), .b(output_15_10), .y(output_14_9));
wire output_16_9, output_16_10, output_15_9;
mixer gate_output_15_9(.a(output_16_9), .b(output_16_10), .y(output_15_9));
wire output_1_10, output_1_11, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_11), .y(output_0_10));
wire output_2_10, output_2_11, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_11), .y(output_1_10));
wire output_3_10, output_3_11, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_11), .y(output_2_10));
wire output_4_10, output_4_11, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_11), .y(output_3_10));
wire output_5_10, output_5_11, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_11), .y(output_4_10));
wire output_6_10, output_6_11, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_11), .y(output_5_10));
wire output_7_10, output_7_11, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_11), .y(output_6_10));
wire output_8_10, output_8_11, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_11), .y(output_7_10));
wire output_9_10, output_9_11, output_8_10;
mixer gate_output_8_10(.a(output_9_10), .b(output_9_11), .y(output_8_10));
wire output_10_10, output_10_11, output_9_10;
mixer gate_output_9_10(.a(output_10_10), .b(output_10_11), .y(output_9_10));
wire output_11_10, output_11_11, output_10_10;
mixer gate_output_10_10(.a(output_11_10), .b(output_11_11), .y(output_10_10));
wire output_12_10, output_12_11, output_11_10;
mixer gate_output_11_10(.a(output_12_10), .b(output_12_11), .y(output_11_10));
wire output_13_10, output_13_11, output_12_10;
mixer gate_output_12_10(.a(output_13_10), .b(output_13_11), .y(output_12_10));
wire output_14_10, output_14_11, output_13_10;
mixer gate_output_13_10(.a(output_14_10), .b(output_14_11), .y(output_13_10));
wire output_15_10, output_15_11, output_14_10;
mixer gate_output_14_10(.a(output_15_10), .b(output_15_11), .y(output_14_10));
wire output_16_10, output_16_11, output_15_10;
mixer gate_output_15_10(.a(output_16_10), .b(output_16_11), .y(output_15_10));
wire output_1_11, output_1_12, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_12), .y(output_0_11));
wire output_2_11, output_2_12, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_12), .y(output_1_11));
wire output_3_11, output_3_12, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_12), .y(output_2_11));
wire output_4_11, output_4_12, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_12), .y(output_3_11));
wire output_5_11, output_5_12, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_12), .y(output_4_11));
wire output_6_11, output_6_12, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_12), .y(output_5_11));
wire output_7_11, output_7_12, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_12), .y(output_6_11));
wire output_8_11, output_8_12, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_12), .y(output_7_11));
wire output_9_11, output_9_12, output_8_11;
mixer gate_output_8_11(.a(output_9_11), .b(output_9_12), .y(output_8_11));
wire output_10_11, output_10_12, output_9_11;
mixer gate_output_9_11(.a(output_10_11), .b(output_10_12), .y(output_9_11));
wire output_11_11, output_11_12, output_10_11;
mixer gate_output_10_11(.a(output_11_11), .b(output_11_12), .y(output_10_11));
wire output_12_11, output_12_12, output_11_11;
mixer gate_output_11_11(.a(output_12_11), .b(output_12_12), .y(output_11_11));
wire output_13_11, output_13_12, output_12_11;
mixer gate_output_12_11(.a(output_13_11), .b(output_13_12), .y(output_12_11));
wire output_14_11, output_14_12, output_13_11;
mixer gate_output_13_11(.a(output_14_11), .b(output_14_12), .y(output_13_11));
wire output_15_11, output_15_12, output_14_11;
mixer gate_output_14_11(.a(output_15_11), .b(output_15_12), .y(output_14_11));
wire output_16_11, output_16_12, output_15_11;
mixer gate_output_15_11(.a(output_16_11), .b(output_16_12), .y(output_15_11));
wire output_1_12, output_1_13, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_13), .y(output_0_12));
wire output_2_12, output_2_13, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_13), .y(output_1_12));
wire output_3_12, output_3_13, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_13), .y(output_2_12));
wire output_4_12, output_4_13, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_13), .y(output_3_12));
wire output_5_12, output_5_13, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_13), .y(output_4_12));
wire output_6_12, output_6_13, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_13), .y(output_5_12));
wire output_7_12, output_7_13, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_13), .y(output_6_12));
wire output_8_12, output_8_13, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_13), .y(output_7_12));
wire output_9_12, output_9_13, output_8_12;
mixer gate_output_8_12(.a(output_9_12), .b(output_9_13), .y(output_8_12));
wire output_10_12, output_10_13, output_9_12;
mixer gate_output_9_12(.a(output_10_12), .b(output_10_13), .y(output_9_12));
wire output_11_12, output_11_13, output_10_12;
mixer gate_output_10_12(.a(output_11_12), .b(output_11_13), .y(output_10_12));
wire output_12_12, output_12_13, output_11_12;
mixer gate_output_11_12(.a(output_12_12), .b(output_12_13), .y(output_11_12));
wire output_13_12, output_13_13, output_12_12;
mixer gate_output_12_12(.a(output_13_12), .b(output_13_13), .y(output_12_12));
wire output_14_12, output_14_13, output_13_12;
mixer gate_output_13_12(.a(output_14_12), .b(output_14_13), .y(output_13_12));
wire output_15_12, output_15_13, output_14_12;
mixer gate_output_14_12(.a(output_15_12), .b(output_15_13), .y(output_14_12));
wire output_16_12, output_16_13, output_15_12;
mixer gate_output_15_12(.a(output_16_12), .b(output_16_13), .y(output_15_12));
wire output_1_13, output_1_14, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_14), .y(output_0_13));
wire output_2_13, output_2_14, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_14), .y(output_1_13));
wire output_3_13, output_3_14, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_14), .y(output_2_13));
wire output_4_13, output_4_14, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_14), .y(output_3_13));
wire output_5_13, output_5_14, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_14), .y(output_4_13));
wire output_6_13, output_6_14, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_14), .y(output_5_13));
wire output_7_13, output_7_14, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_14), .y(output_6_13));
wire output_8_13, output_8_14, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_14), .y(output_7_13));
wire output_9_13, output_9_14, output_8_13;
mixer gate_output_8_13(.a(output_9_13), .b(output_9_14), .y(output_8_13));
wire output_10_13, output_10_14, output_9_13;
mixer gate_output_9_13(.a(output_10_13), .b(output_10_14), .y(output_9_13));
wire output_11_13, output_11_14, output_10_13;
mixer gate_output_10_13(.a(output_11_13), .b(output_11_14), .y(output_10_13));
wire output_12_13, output_12_14, output_11_13;
mixer gate_output_11_13(.a(output_12_13), .b(output_12_14), .y(output_11_13));
wire output_13_13, output_13_14, output_12_13;
mixer gate_output_12_13(.a(output_13_13), .b(output_13_14), .y(output_12_13));
wire output_14_13, output_14_14, output_13_13;
mixer gate_output_13_13(.a(output_14_13), .b(output_14_14), .y(output_13_13));
wire output_15_13, output_15_14, output_14_13;
mixer gate_output_14_13(.a(output_15_13), .b(output_15_14), .y(output_14_13));
wire output_16_13, output_16_14, output_15_13;
mixer gate_output_15_13(.a(output_16_13), .b(output_16_14), .y(output_15_13));
wire output_1_14, output_1_15, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_15), .y(output_0_14));
wire output_2_14, output_2_15, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_15), .y(output_1_14));
wire output_3_14, output_3_15, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_15), .y(output_2_14));
wire output_4_14, output_4_15, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_15), .y(output_3_14));
wire output_5_14, output_5_15, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_15), .y(output_4_14));
wire output_6_14, output_6_15, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_15), .y(output_5_14));
wire output_7_14, output_7_15, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_15), .y(output_6_14));
wire output_8_14, output_8_15, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_15), .y(output_7_14));
wire output_9_14, output_9_15, output_8_14;
mixer gate_output_8_14(.a(output_9_14), .b(output_9_15), .y(output_8_14));
wire output_10_14, output_10_15, output_9_14;
mixer gate_output_9_14(.a(output_10_14), .b(output_10_15), .y(output_9_14));
wire output_11_14, output_11_15, output_10_14;
mixer gate_output_10_14(.a(output_11_14), .b(output_11_15), .y(output_10_14));
wire output_12_14, output_12_15, output_11_14;
mixer gate_output_11_14(.a(output_12_14), .b(output_12_15), .y(output_11_14));
wire output_13_14, output_13_15, output_12_14;
mixer gate_output_12_14(.a(output_13_14), .b(output_13_15), .y(output_12_14));
wire output_14_14, output_14_15, output_13_14;
mixer gate_output_13_14(.a(output_14_14), .b(output_14_15), .y(output_13_14));
wire output_15_14, output_15_15, output_14_14;
mixer gate_output_14_14(.a(output_15_14), .b(output_15_15), .y(output_14_14));
wire output_16_14, output_16_15, output_15_14;
mixer gate_output_15_14(.a(output_16_14), .b(output_16_15), .y(output_15_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
wire output_9_15, output_9_0, output_8_15;
mixer gate_output_8_15(.a(output_9_15), .b(output_9_0), .y(output_8_15));
wire output_10_15, output_10_0, output_9_15;
mixer gate_output_9_15(.a(output_10_15), .b(output_10_0), .y(output_9_15));
wire output_11_15, output_11_0, output_10_15;
mixer gate_output_10_15(.a(output_11_15), .b(output_11_0), .y(output_10_15));
wire output_12_15, output_12_0, output_11_15;
mixer gate_output_11_15(.a(output_12_15), .b(output_12_0), .y(output_11_15));
wire output_13_15, output_13_0, output_12_15;
mixer gate_output_12_15(.a(output_13_15), .b(output_13_0), .y(output_12_15));
wire output_14_15, output_14_0, output_13_15;
mixer gate_output_13_15(.a(output_14_15), .b(output_14_0), .y(output_13_15));
wire output_15_15, output_15_0, output_14_15;
mixer gate_output_14_15(.a(output_15_15), .b(output_15_0), .y(output_14_15));
wire output_16_15, output_16_0, output_15_15;
mixer gate_output_15_15(.a(output_16_15), .b(output_16_0), .y(output_15_15));
assign output_0 = output_0_0;
wire output_0_16;
assign output_0_16 = input_0;
assign output_1 = output_1_0;
wire output_1_16;
assign output_1_16 = input_1;
assign output_2 = output_2_0;
wire output_2_16;
assign output_2_16 = input_2;
assign output_3 = output_3_0;
wire output_3_16;
assign output_3_16 = input_3;
assign output_4 = output_4_0;
wire output_4_16;
assign output_4_16 = input_4;
assign output_5 = output_5_0;
wire output_5_16;
assign output_5_16 = input_5;
assign output_6 = output_6_0;
wire output_6_16;
assign output_6_16 = input_6;
assign output_7 = output_7_0;
wire output_7_16;
assign output_7_16 = input_7;
assign output_8 = output_8_0;
wire output_8_16;
assign output_8_16 = input_8;
assign output_9 = output_9_0;
wire output_9_16;
assign output_9_16 = input_9;
assign output_10 = output_10_0;
wire output_10_16;
assign output_10_16 = input_10;
assign output_11 = output_11_0;
wire output_11_16;
assign output_11_16 = input_11;
assign output_12 = output_12_0;
wire output_12_16;
assign output_12_16 = input_12;
assign output_13 = output_13_0;
wire output_13_16;
assign output_13_16 = input_13;
assign output_14 = output_14_0;
wire output_14_16;
assign output_14_16 = input_14;
assign output_15 = output_15_0;
wire output_15_16;
assign output_15_16 = input_15;
endmodule
