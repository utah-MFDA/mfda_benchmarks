module Planar_Synthetic_4(
input Source1,
output Out1
);
wire flow_switch3_0_Out1;
wire flow_switch3_0_flow_switch4_10;
wire flow_switch4_9_flow_switch4_7;
wire flow_switch4_9_Filter1;
wire flow_switch4_9_Filter2;
wire flow_switch4_10_flow_switch4_8;
wire flow_switch4_10_Filter3;
wire flow_switch4_10_Filter4;
wire flow_switch4_7_flow_switch4_5;
wire flow_switch4_7_Heater1;
wire flow_switch4_7_Heater2;
wire flow_switch4_8_flow_switch4_6;
wire flow_switch4_8_Heater3;
wire flow_switch4_8_Heater4;
wire flow_switch4_5_flow_switch4_3;
wire flow_switch4_5_Mixer9;
wire flow_switch4_5_Mixer10;
wire flow_switch4_6_flow_switch4_4;
wire flow_switch4_6_Mixer11;
wire flow_switch4_6_Mixer12;
wire flow_switch4_3_flow_switch4_1;
wire flow_switch4_3_Mixer5;
wire flow_switch4_3_Mixer6;
wire flow_switch4_4_flow_switch4_2;
wire flow_switch4_4_Mixer7;
wire flow_switch4_4_Mixer8;
wire flow_switch4_1_Mixer1;
wire flow_switch4_1_Mixer2;
wire flow_switch4_2_Mixer3;
wire flow_switch4_2_Mixer4;
wire flow_switch3_1_Source1;
wire flow_switch3_1_flow_switch4_1;
wire flow_switch3_1_flow_switch4_2;
assign flow_switch3_1_Source1 = Source1;
assign Out1 = flow_switch3_0_Out1;
chamber Mixer1(.port1(flow_switch4_1_Mixer1));
chamber Mixer2(.port1(flow_switch4_1_Mixer2));
chamber Mixer3(.port0(flow_switch4_2_Mixer3));
chamber Mixer4(.port0(flow_switch4_2_Mixer4));
chamber Mixer5(.port1(flow_switch4_3_Mixer5));
chamber Mixer6(.port1(flow_switch4_3_Mixer6));
chamber Mixer7(.port0(flow_switch4_4_Mixer7));
chamber Mixer8(.port1(flow_switch4_4_Mixer8));
chamber Mixer9(.port1(flow_switch4_5_Mixer9));
chamber Mixer10(.port1(flow_switch4_5_Mixer10));
chamber Mixer11(.port0(flow_switch4_6_Mixer11));
chamber Mixer12(.port1(flow_switch4_6_Mixer12));
heater Heater1(.port0(flow_switch4_7_Heater1));
heater Heater2(.port0(flow_switch4_7_Heater2));
heater Heater3(.port1(flow_switch4_8_Heater3));
heater Heater4(.port0(flow_switch4_8_Heater4));
filter Filter1(.port0(flow_switch4_9_Filter1));
filter Filter2(.port0(flow_switch4_9_Filter2));
filter Filter3(.port0(flow_switch4_10_Filter3));
filter Filter4(.port0(flow_switch4_10_Filter4));
junction4 flow_switch3_0(.port1(flow_switch3_0_flow_switch4_10),.port3(flow_switch3_0_Out1));
junction4 flow_switch3_1(.port0(flow_switch3_1_flow_switch4_2),.port2(flow_switch3_1_Source1),.port3(flow_switch3_1_flow_switch4_1));
junction4 flow_switch4_1(.port0(flow_switch4_1_Mixer2),.port1(flow_switch4_3_flow_switch4_1),.port2(flow_switch3_1_flow_switch4_1),.port3(flow_switch4_1_Mixer1));
junction4 flow_switch4_2(.port0(flow_switch4_4_flow_switch4_2),.port1(flow_switch4_2_Mixer4),.port2(flow_switch4_2_Mixer3),.port3(flow_switch3_1_flow_switch4_2));
junction4 flow_switch4_3(.port0(flow_switch4_3_Mixer6),.port1(flow_switch4_5_flow_switch4_3),.port2(flow_switch4_3_flow_switch4_1),.port3(flow_switch4_3_Mixer5));
junction4 flow_switch4_4(.port0(flow_switch4_6_flow_switch4_4),.port1(flow_switch4_4_flow_switch4_2),.port2(flow_switch4_4_Mixer7),.port3(flow_switch4_4_Mixer8));
junction4 flow_switch4_5(.port0(flow_switch4_7_flow_switch4_5),.port1(flow_switch4_5_Mixer9),.port2(flow_switch4_5_flow_switch4_3),.port3(flow_switch4_5_Mixer10));
junction4 flow_switch4_6(.port0(flow_switch4_8_flow_switch4_6),.port1(flow_switch4_6_flow_switch4_4),.port2(flow_switch4_6_Mixer11),.port3(flow_switch4_6_Mixer12));
junction4 flow_switch4_7(.port0(flow_switch4_7_Heater2),.port1(flow_switch4_9_flow_switch4_7),.port2(flow_switch4_7_flow_switch4_5),.port3(flow_switch4_7_Heater1));
junction4 flow_switch4_8(.port0(flow_switch4_10_flow_switch4_8),.port1(flow_switch4_8_flow_switch4_6),.port2(flow_switch4_8_Heater3),.port3(flow_switch4_8_Heater4));
junction4 flow_switch4_9(.port0(flow_switch4_9_Filter2),.port2(flow_switch4_9_Filter1),.port3(flow_switch4_9_flow_switch4_7));
junction4 flow_switch4_10(.port0(flow_switch3_0_flow_switch4_10),.port1(flow_switch4_10_flow_switch4_8),.port2(flow_switch4_10_Filter3),.port3(flow_switch4_10_Filter4));
endmodule
