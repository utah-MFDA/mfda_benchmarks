module binary_tree_8_2 (
output out_0,output out_1,output out_2,output out_3,output out_4,output out_5,output out_6,output out_7,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t1_0 (.a(t1_00), .b(t1_01), .y(t1_0));
wire t1_00, t1_01;
mixer mix_t1_00 (.a(t1_000), .b(t1_001), .y(t1_00));
wire t1_000, t1_001;
mixer mix_t1_01 (.a(t1_010), .b(t1_011), .y(t1_01));
wire t1_010, t1_011;
mixer mix_t2_0 (.a(t2_00), .b(t2_01), .y(t2_0));
wire t2_00, t2_01;
mixer mix_t2_00 (.a(t2_000), .b(t2_001), .y(t2_00));
wire t2_000, t2_001;
mixer mix_t2_01 (.a(t2_010), .b(t2_011), .y(t2_01));
wire t2_010, t2_011;
mixer mix_t3_0 (.a(t3_00), .b(t3_01), .y(t3_0));
wire t3_00, t3_01;
mixer mix_t3_00 (.a(t3_000), .b(t3_001), .y(t3_00));
wire t3_000, t3_001;
mixer mix_t3_01 (.a(t3_010), .b(t3_011), .y(t3_01));
wire t3_010, t3_011;
mixer mix_t4_0 (.a(t4_00), .b(t4_01), .y(t4_0));
wire t4_00, t4_01;
mixer mix_t4_00 (.a(t4_000), .b(t4_001), .y(t4_00));
wire t4_000, t4_001;
mixer mix_t4_01 (.a(t4_010), .b(t4_011), .y(t4_01));
wire t4_010, t4_011;
mixer mix_t5_0 (.a(t5_00), .b(t5_01), .y(t5_0));
wire t5_00, t5_01;
mixer mix_t5_00 (.a(t5_000), .b(t5_001), .y(t5_00));
wire t5_000, t5_001;
mixer mix_t5_01 (.a(t5_010), .b(t5_011), .y(t5_01));
wire t5_010, t5_011;
mixer mix_t6_0 (.a(t6_00), .b(t6_01), .y(t6_0));
wire t6_00, t6_01;
mixer mix_t6_00 (.a(t6_000), .b(t6_001), .y(t6_00));
wire t6_000, t6_001;
mixer mix_t6_01 (.a(t6_010), .b(t6_011), .y(t6_01));
wire t6_010, t6_011;
mixer mix_t7_0 (.a(t7_00), .b(t7_01), .y(t7_0));
wire t7_00, t7_01;
mixer mix_t7_00 (.a(t7_000), .b(t7_001), .y(t7_00));
wire t7_000, t7_001;
mixer mix_t7_01 (.a(t7_010), .b(t7_011), .y(t7_01));
wire t7_010, t7_011;
wire t0_0;
assign out_0 = t0_0;
wire t1_0;
assign out_1 = t1_0;
wire t2_0;
assign out_2 = t2_0;
wire t3_0;
assign out_3 = t3_0;
wire t4_0;
assign out_4 = t4_0;
wire t5_0;
assign out_5 = t5_0;
wire t6_0;
assign out_6 = t6_0;
wire t7_0;
assign out_7 = t7_0;
assign input_0 = t0_000;
assign input_1 = t0_001;
assign input_2 = t0_010;
assign input_3 = t0_011;
assign input_4 = t1_000;
assign input_5 = t1_001;
assign input_6 = t1_010;
assign input_7 = t1_011;
assign input_8 = t2_000;
assign input_9 = t2_001;
assign input_10 = t2_010;
assign input_11 = t2_011;
assign input_12 = t3_000;
assign input_13 = t3_001;
assign input_14 = t3_010;
assign input_15 = t3_011;
assign input_16 = t4_000;
assign input_17 = t4_001;
assign input_18 = t4_010;
assign input_19 = t4_011;
assign input_20 = t5_000;
assign input_21 = t5_001;
assign input_22 = t5_010;
assign input_23 = t5_011;
assign input_24 = t6_000;
assign input_25 = t6_001;
assign input_26 = t6_010;
assign input_27 = t6_011;
assign input_28 = t7_000;
assign input_29 = t7_001;
assign input_30 = t7_010;
assign input_31 = t7_011;
endmodule
