module binary_tree_4_8 (
output out_0,output out_1,output out_2,output out_3,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63,input input_64,input input_65,input input_66,input input_67,input input_68,input input_69,input input_70,input input_71,input input_72,input input_73,input input_74,input input_75,input input_76,input input_77,input input_78,input input_79,input input_80,input input_81,input input_82,input input_83,input input_84,input input_85,input input_86,input input_87,input input_88,input input_89,input input_90,input input_91,input input_92,input input_93,input input_94,input input_95,input input_96,input input_97,input input_98,input input_99,input input_100,input input_101,input input_102,input input_103,input input_104,input input_105,input input_106,input input_107,input input_108,input input_109,input input_110,input input_111,input input_112,input input_113,input input_114,input input_115,input input_116,input input_117,input input_118,input input_119,input input_120,input input_121,input input_122,input input_123,input input_124,input input_125,input input_126,input input_127,input input_128,input input_129,input input_130,input input_131,input input_132,input input_133,input input_134,input input_135,input input_136,input input_137,input input_138,input input_139,input input_140,input input_141,input input_142,input input_143,input input_144,input input_145,input input_146,input input_147,input input_148,input input_149,input input_150,input input_151,input input_152,input input_153,input input_154,input input_155,input input_156,input input_157,input input_158,input input_159,input input_160,input input_161,input input_162,input input_163,input input_164,input input_165,input input_166,input input_167,input input_168,input input_169,input input_170,input input_171,input input_172,input input_173,input input_174,input input_175,input input_176,input input_177,input input_178,input input_179,input input_180,input input_181,input input_182,input input_183,input input_184,input input_185,input input_186,input input_187,input input_188,input input_189,input input_190,input input_191,input input_192,input input_193,input input_194,input input_195,input input_196,input input_197,input input_198,input input_199,input input_200,input input_201,input input_202,input input_203,input input_204,input input_205,input input_206,input input_207,input input_208,input input_209,input input_210,input input_211,input input_212,input input_213,input input_214,input input_215,input input_216,input input_217,input input_218,input input_219,input input_220,input input_221,input input_222,input input_223,input input_224,input input_225,input input_226,input input_227,input input_228,input input_229,input input_230,input input_231,input input_232,input input_233,input input_234,input input_235,input input_236,input input_237,input input_238,input input_239,input input_240,input input_241,input input_242,input input_243,input input_244,input input_245,input input_246,input input_247,input input_248,input input_249,input input_250,input input_251,input input_252,input input_253,input input_254,input input_255,input input_256,input input_257,input input_258,input input_259,input input_260,input input_261,input input_262,input input_263,input input_264,input input_265,input input_266,input input_267,input input_268,input input_269,input input_270,input input_271,input input_272,input input_273,input input_274,input input_275,input input_276,input input_277,input input_278,input input_279,input input_280,input input_281,input input_282,input input_283,input input_284,input input_285,input input_286,input input_287,input input_288,input input_289,input input_290,input input_291,input input_292,input input_293,input input_294,input input_295,input input_296,input input_297,input input_298,input input_299,input input_300,input input_301,input input_302,input input_303,input input_304,input input_305,input input_306,input input_307,input input_308,input input_309,input input_310,input input_311,input input_312,input input_313,input input_314,input input_315,input input_316,input input_317,input input_318,input input_319,input input_320,input input_321,input input_322,input input_323,input input_324,input input_325,input input_326,input input_327,input input_328,input input_329,input input_330,input input_331,input input_332,input input_333,input input_334,input input_335,input input_336,input input_337,input input_338,input input_339,input input_340,input input_341,input input_342,input input_343,input input_344,input input_345,input input_346,input input_347,input input_348,input input_349,input input_350,input input_351,input input_352,input input_353,input input_354,input input_355,input input_356,input input_357,input input_358,input input_359,input input_360,input input_361,input input_362,input input_363,input input_364,input input_365,input input_366,input input_367,input input_368,input input_369,input input_370,input input_371,input input_372,input input_373,input input_374,input input_375,input input_376,input input_377,input input_378,input input_379,input input_380,input input_381,input input_382,input input_383,input input_384,input input_385,input input_386,input input_387,input input_388,input input_389,input input_390,input input_391,input input_392,input input_393,input input_394,input input_395,input input_396,input input_397,input input_398,input input_399,input input_400,input input_401,input input_402,input input_403,input input_404,input input_405,input input_406,input input_407,input input_408,input input_409,input input_410,input input_411,input input_412,input input_413,input input_414,input input_415,input input_416,input input_417,input input_418,input input_419,input input_420,input input_421,input input_422,input input_423,input input_424,input input_425,input input_426,input input_427,input input_428,input input_429,input input_430,input input_431,input input_432,input input_433,input input_434,input input_435,input input_436,input input_437,input input_438,input input_439,input input_440,input input_441,input input_442,input input_443,input input_444,input input_445,input input_446,input input_447,input input_448,input input_449,input input_450,input input_451,input input_452,input input_453,input input_454,input input_455,input input_456,input input_457,input input_458,input input_459,input input_460,input input_461,input input_462,input input_463,input input_464,input input_465,input input_466,input input_467,input input_468,input input_469,input input_470,input input_471,input input_472,input input_473,input input_474,input input_475,input input_476,input input_477,input input_478,input input_479,input input_480,input input_481,input input_482,input input_483,input input_484,input input_485,input input_486,input input_487,input input_488,input input_489,input input_490,input input_491,input input_492,input input_493,input input_494,input input_495,input input_496,input input_497,input input_498,input input_499,input input_500,input input_501,input input_502,input input_503,input input_504,input input_505,input input_506,input input_507,input input_508,input input_509,input input_510,input input_511,input input_512,input input_513,input input_514,input input_515,input input_516,input input_517,input input_518,input input_519,input input_520,input input_521,input input_522,input input_523,input input_524,input input_525,input input_526,input input_527,input input_528,input input_529,input input_530,input input_531,input input_532,input input_533,input input_534,input input_535,input input_536,input input_537,input input_538,input input_539,input input_540,input input_541,input input_542,input input_543,input input_544,input input_545,input input_546,input input_547,input input_548,input input_549,input input_550,input input_551,input input_552,input input_553,input input_554,input input_555,input input_556,input input_557,input input_558,input input_559,input input_560,input input_561,input input_562,input input_563,input input_564,input input_565,input input_566,input input_567,input input_568,input input_569,input input_570,input input_571,input input_572,input input_573,input input_574,input input_575,input input_576,input input_577,input input_578,input input_579,input input_580,input input_581,input input_582,input input_583,input input_584,input input_585,input input_586,input input_587,input input_588,input input_589,input input_590,input input_591,input input_592,input input_593,input input_594,input input_595,input input_596,input input_597,input input_598,input input_599,input input_600,input input_601,input input_602,input input_603,input input_604,input input_605,input input_606,input input_607,input input_608,input input_609,input input_610,input input_611,input input_612,input input_613,input input_614,input input_615,input input_616,input input_617,input input_618,input input_619,input input_620,input input_621,input input_622,input input_623,input input_624,input input_625,input input_626,input input_627,input input_628,input input_629,input input_630,input input_631,input input_632,input input_633,input input_634,input input_635,input input_636,input input_637,input input_638,input input_639,input input_640,input input_641,input input_642,input input_643,input input_644,input input_645,input input_646,input input_647,input input_648,input input_649,input input_650,input input_651,input input_652,input input_653,input input_654,input input_655,input input_656,input input_657,input input_658,input input_659,input input_660,input input_661,input input_662,input input_663,input input_664,input input_665,input input_666,input input_667,input input_668,input input_669,input input_670,input input_671,input input_672,input input_673,input input_674,input input_675,input input_676,input input_677,input input_678,input input_679,input input_680,input input_681,input input_682,input input_683,input input_684,input input_685,input input_686,input input_687,input input_688,input input_689,input input_690,input input_691,input input_692,input input_693,input input_694,input input_695,input input_696,input input_697,input input_698,input input_699,input input_700,input input_701,input input_702,input input_703,input input_704,input input_705,input input_706,input input_707,input input_708,input input_709,input input_710,input input_711,input input_712,input input_713,input input_714,input input_715,input input_716,input input_717,input input_718,input input_719,input input_720,input input_721,input input_722,input input_723,input input_724,input input_725,input input_726,input input_727,input input_728,input input_729,input input_730,input input_731,input input_732,input input_733,input input_734,input input_735,input input_736,input input_737,input input_738,input input_739,input input_740,input input_741,input input_742,input input_743,input input_744,input input_745,input input_746,input input_747,input input_748,input input_749,input input_750,input input_751,input input_752,input input_753,input input_754,input input_755,input input_756,input input_757,input input_758,input input_759,input input_760,input input_761,input input_762,input input_763,input input_764,input input_765,input input_766,input input_767,input input_768,input input_769,input input_770,input input_771,input input_772,input input_773,input input_774,input input_775,input input_776,input input_777,input input_778,input input_779,input input_780,input input_781,input input_782,input input_783,input input_784,input input_785,input input_786,input input_787,input input_788,input input_789,input input_790,input input_791,input input_792,input input_793,input input_794,input input_795,input input_796,input input_797,input input_798,input input_799,input input_800,input input_801,input input_802,input input_803,input input_804,input input_805,input input_806,input input_807,input input_808,input input_809,input input_810,input input_811,input input_812,input input_813,input input_814,input input_815,input input_816,input input_817,input input_818,input input_819,input input_820,input input_821,input input_822,input input_823,input input_824,input input_825,input input_826,input input_827,input input_828,input input_829,input input_830,input input_831,input input_832,input input_833,input input_834,input input_835,input input_836,input input_837,input input_838,input input_839,input input_840,input input_841,input input_842,input input_843,input input_844,input input_845,input input_846,input input_847,input input_848,input input_849,input input_850,input input_851,input input_852,input input_853,input input_854,input input_855,input input_856,input input_857,input input_858,input input_859,input input_860,input input_861,input input_862,input input_863,input input_864,input input_865,input input_866,input input_867,input input_868,input input_869,input input_870,input input_871,input input_872,input input_873,input input_874,input input_875,input input_876,input input_877,input input_878,input input_879,input input_880,input input_881,input input_882,input input_883,input input_884,input input_885,input input_886,input input_887,input input_888,input input_889,input input_890,input input_891,input input_892,input input_893,input input_894,input input_895,input input_896,input input_897,input input_898,input input_899,input input_900,input input_901,input input_902,input input_903,input input_904,input input_905,input input_906,input input_907,input input_908,input input_909,input input_910,input input_911,input input_912,input input_913,input input_914,input input_915,input input_916,input input_917,input input_918,input input_919,input input_920,input input_921,input input_922,input input_923,input input_924,input input_925,input input_926,input input_927,input input_928,input input_929,input input_930,input input_931,input input_932,input input_933,input input_934,input input_935,input input_936,input input_937,input input_938,input input_939,input input_940,input input_941,input input_942,input input_943,input input_944,input input_945,input input_946,input input_947,input input_948,input input_949,input input_950,input input_951,input input_952,input input_953,input input_954,input input_955,input input_956,input input_957,input input_958,input input_959,input input_960,input input_961,input input_962,input input_963,input input_964,input input_965,input input_966,input input_967,input input_968,input input_969,input input_970,input input_971,input input_972,input input_973,input input_974,input input_975,input input_976,input input_977,input input_978,input input_979,input input_980,input input_981,input input_982,input input_983,input input_984,input input_985,input input_986,input input_987,input input_988,input input_989,input input_990,input input_991,input input_992,input input_993,input input_994,input input_995,input input_996,input input_997,input input_998,input input_999,input input_1000,input input_1001,input input_1002,input input_1003,input input_1004,input input_1005,input input_1006,input input_1007,input input_1008,input input_1009,input input_1010,input input_1011,input input_1012,input input_1013,input input_1014,input input_1015,input input_1016,input input_1017,input input_1018,input input_1019,input input_1020,input input_1021,input input_1022,input input_1023
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_000000 (.a(t0_0000000), .b(t0_0000001), .y(t0_000000));
wire t0_0000000, t0_0000001;
mixer mix_t0_0000000 (.a(t0_00000000), .b(t0_00000001), .y(t0_0000000));
wire t0_00000000, t0_00000001;
mixer mix_t0_00000000 (.a(t0_000000000), .b(t0_000000001), .y(t0_00000000));
wire t0_000000000, t0_000000001;
mixer mix_t0_00000001 (.a(t0_000000010), .b(t0_000000011), .y(t0_00000001));
wire t0_000000010, t0_000000011;
mixer mix_t0_0000001 (.a(t0_00000010), .b(t0_00000011), .y(t0_0000001));
wire t0_00000010, t0_00000011;
mixer mix_t0_00000010 (.a(t0_000000100), .b(t0_000000101), .y(t0_00000010));
wire t0_000000100, t0_000000101;
mixer mix_t0_00000011 (.a(t0_000000110), .b(t0_000000111), .y(t0_00000011));
wire t0_000000110, t0_000000111;
mixer mix_t0_000001 (.a(t0_0000010), .b(t0_0000011), .y(t0_000001));
wire t0_0000010, t0_0000011;
mixer mix_t0_0000010 (.a(t0_00000100), .b(t0_00000101), .y(t0_0000010));
wire t0_00000100, t0_00000101;
mixer mix_t0_00000100 (.a(t0_000001000), .b(t0_000001001), .y(t0_00000100));
wire t0_000001000, t0_000001001;
mixer mix_t0_00000101 (.a(t0_000001010), .b(t0_000001011), .y(t0_00000101));
wire t0_000001010, t0_000001011;
mixer mix_t0_0000011 (.a(t0_00000110), .b(t0_00000111), .y(t0_0000011));
wire t0_00000110, t0_00000111;
mixer mix_t0_00000110 (.a(t0_000001100), .b(t0_000001101), .y(t0_00000110));
wire t0_000001100, t0_000001101;
mixer mix_t0_00000111 (.a(t0_000001110), .b(t0_000001111), .y(t0_00000111));
wire t0_000001110, t0_000001111;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_000010 (.a(t0_0000100), .b(t0_0000101), .y(t0_000010));
wire t0_0000100, t0_0000101;
mixer mix_t0_0000100 (.a(t0_00001000), .b(t0_00001001), .y(t0_0000100));
wire t0_00001000, t0_00001001;
mixer mix_t0_00001000 (.a(t0_000010000), .b(t0_000010001), .y(t0_00001000));
wire t0_000010000, t0_000010001;
mixer mix_t0_00001001 (.a(t0_000010010), .b(t0_000010011), .y(t0_00001001));
wire t0_000010010, t0_000010011;
mixer mix_t0_0000101 (.a(t0_00001010), .b(t0_00001011), .y(t0_0000101));
wire t0_00001010, t0_00001011;
mixer mix_t0_00001010 (.a(t0_000010100), .b(t0_000010101), .y(t0_00001010));
wire t0_000010100, t0_000010101;
mixer mix_t0_00001011 (.a(t0_000010110), .b(t0_000010111), .y(t0_00001011));
wire t0_000010110, t0_000010111;
mixer mix_t0_000011 (.a(t0_0000110), .b(t0_0000111), .y(t0_000011));
wire t0_0000110, t0_0000111;
mixer mix_t0_0000110 (.a(t0_00001100), .b(t0_00001101), .y(t0_0000110));
wire t0_00001100, t0_00001101;
mixer mix_t0_00001100 (.a(t0_000011000), .b(t0_000011001), .y(t0_00001100));
wire t0_000011000, t0_000011001;
mixer mix_t0_00001101 (.a(t0_000011010), .b(t0_000011011), .y(t0_00001101));
wire t0_000011010, t0_000011011;
mixer mix_t0_0000111 (.a(t0_00001110), .b(t0_00001111), .y(t0_0000111));
wire t0_00001110, t0_00001111;
mixer mix_t0_00001110 (.a(t0_000011100), .b(t0_000011101), .y(t0_00001110));
wire t0_000011100, t0_000011101;
mixer mix_t0_00001111 (.a(t0_000011110), .b(t0_000011111), .y(t0_00001111));
wire t0_000011110, t0_000011111;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_000100 (.a(t0_0001000), .b(t0_0001001), .y(t0_000100));
wire t0_0001000, t0_0001001;
mixer mix_t0_0001000 (.a(t0_00010000), .b(t0_00010001), .y(t0_0001000));
wire t0_00010000, t0_00010001;
mixer mix_t0_00010000 (.a(t0_000100000), .b(t0_000100001), .y(t0_00010000));
wire t0_000100000, t0_000100001;
mixer mix_t0_00010001 (.a(t0_000100010), .b(t0_000100011), .y(t0_00010001));
wire t0_000100010, t0_000100011;
mixer mix_t0_0001001 (.a(t0_00010010), .b(t0_00010011), .y(t0_0001001));
wire t0_00010010, t0_00010011;
mixer mix_t0_00010010 (.a(t0_000100100), .b(t0_000100101), .y(t0_00010010));
wire t0_000100100, t0_000100101;
mixer mix_t0_00010011 (.a(t0_000100110), .b(t0_000100111), .y(t0_00010011));
wire t0_000100110, t0_000100111;
mixer mix_t0_000101 (.a(t0_0001010), .b(t0_0001011), .y(t0_000101));
wire t0_0001010, t0_0001011;
mixer mix_t0_0001010 (.a(t0_00010100), .b(t0_00010101), .y(t0_0001010));
wire t0_00010100, t0_00010101;
mixer mix_t0_00010100 (.a(t0_000101000), .b(t0_000101001), .y(t0_00010100));
wire t0_000101000, t0_000101001;
mixer mix_t0_00010101 (.a(t0_000101010), .b(t0_000101011), .y(t0_00010101));
wire t0_000101010, t0_000101011;
mixer mix_t0_0001011 (.a(t0_00010110), .b(t0_00010111), .y(t0_0001011));
wire t0_00010110, t0_00010111;
mixer mix_t0_00010110 (.a(t0_000101100), .b(t0_000101101), .y(t0_00010110));
wire t0_000101100, t0_000101101;
mixer mix_t0_00010111 (.a(t0_000101110), .b(t0_000101111), .y(t0_00010111));
wire t0_000101110, t0_000101111;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_000110 (.a(t0_0001100), .b(t0_0001101), .y(t0_000110));
wire t0_0001100, t0_0001101;
mixer mix_t0_0001100 (.a(t0_00011000), .b(t0_00011001), .y(t0_0001100));
wire t0_00011000, t0_00011001;
mixer mix_t0_00011000 (.a(t0_000110000), .b(t0_000110001), .y(t0_00011000));
wire t0_000110000, t0_000110001;
mixer mix_t0_00011001 (.a(t0_000110010), .b(t0_000110011), .y(t0_00011001));
wire t0_000110010, t0_000110011;
mixer mix_t0_0001101 (.a(t0_00011010), .b(t0_00011011), .y(t0_0001101));
wire t0_00011010, t0_00011011;
mixer mix_t0_00011010 (.a(t0_000110100), .b(t0_000110101), .y(t0_00011010));
wire t0_000110100, t0_000110101;
mixer mix_t0_00011011 (.a(t0_000110110), .b(t0_000110111), .y(t0_00011011));
wire t0_000110110, t0_000110111;
mixer mix_t0_000111 (.a(t0_0001110), .b(t0_0001111), .y(t0_000111));
wire t0_0001110, t0_0001111;
mixer mix_t0_0001110 (.a(t0_00011100), .b(t0_00011101), .y(t0_0001110));
wire t0_00011100, t0_00011101;
mixer mix_t0_00011100 (.a(t0_000111000), .b(t0_000111001), .y(t0_00011100));
wire t0_000111000, t0_000111001;
mixer mix_t0_00011101 (.a(t0_000111010), .b(t0_000111011), .y(t0_00011101));
wire t0_000111010, t0_000111011;
mixer mix_t0_0001111 (.a(t0_00011110), .b(t0_00011111), .y(t0_0001111));
wire t0_00011110, t0_00011111;
mixer mix_t0_00011110 (.a(t0_000111100), .b(t0_000111101), .y(t0_00011110));
wire t0_000111100, t0_000111101;
mixer mix_t0_00011111 (.a(t0_000111110), .b(t0_000111111), .y(t0_00011111));
wire t0_000111110, t0_000111111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_001000 (.a(t0_0010000), .b(t0_0010001), .y(t0_001000));
wire t0_0010000, t0_0010001;
mixer mix_t0_0010000 (.a(t0_00100000), .b(t0_00100001), .y(t0_0010000));
wire t0_00100000, t0_00100001;
mixer mix_t0_00100000 (.a(t0_001000000), .b(t0_001000001), .y(t0_00100000));
wire t0_001000000, t0_001000001;
mixer mix_t0_00100001 (.a(t0_001000010), .b(t0_001000011), .y(t0_00100001));
wire t0_001000010, t0_001000011;
mixer mix_t0_0010001 (.a(t0_00100010), .b(t0_00100011), .y(t0_0010001));
wire t0_00100010, t0_00100011;
mixer mix_t0_00100010 (.a(t0_001000100), .b(t0_001000101), .y(t0_00100010));
wire t0_001000100, t0_001000101;
mixer mix_t0_00100011 (.a(t0_001000110), .b(t0_001000111), .y(t0_00100011));
wire t0_001000110, t0_001000111;
mixer mix_t0_001001 (.a(t0_0010010), .b(t0_0010011), .y(t0_001001));
wire t0_0010010, t0_0010011;
mixer mix_t0_0010010 (.a(t0_00100100), .b(t0_00100101), .y(t0_0010010));
wire t0_00100100, t0_00100101;
mixer mix_t0_00100100 (.a(t0_001001000), .b(t0_001001001), .y(t0_00100100));
wire t0_001001000, t0_001001001;
mixer mix_t0_00100101 (.a(t0_001001010), .b(t0_001001011), .y(t0_00100101));
wire t0_001001010, t0_001001011;
mixer mix_t0_0010011 (.a(t0_00100110), .b(t0_00100111), .y(t0_0010011));
wire t0_00100110, t0_00100111;
mixer mix_t0_00100110 (.a(t0_001001100), .b(t0_001001101), .y(t0_00100110));
wire t0_001001100, t0_001001101;
mixer mix_t0_00100111 (.a(t0_001001110), .b(t0_001001111), .y(t0_00100111));
wire t0_001001110, t0_001001111;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_001010 (.a(t0_0010100), .b(t0_0010101), .y(t0_001010));
wire t0_0010100, t0_0010101;
mixer mix_t0_0010100 (.a(t0_00101000), .b(t0_00101001), .y(t0_0010100));
wire t0_00101000, t0_00101001;
mixer mix_t0_00101000 (.a(t0_001010000), .b(t0_001010001), .y(t0_00101000));
wire t0_001010000, t0_001010001;
mixer mix_t0_00101001 (.a(t0_001010010), .b(t0_001010011), .y(t0_00101001));
wire t0_001010010, t0_001010011;
mixer mix_t0_0010101 (.a(t0_00101010), .b(t0_00101011), .y(t0_0010101));
wire t0_00101010, t0_00101011;
mixer mix_t0_00101010 (.a(t0_001010100), .b(t0_001010101), .y(t0_00101010));
wire t0_001010100, t0_001010101;
mixer mix_t0_00101011 (.a(t0_001010110), .b(t0_001010111), .y(t0_00101011));
wire t0_001010110, t0_001010111;
mixer mix_t0_001011 (.a(t0_0010110), .b(t0_0010111), .y(t0_001011));
wire t0_0010110, t0_0010111;
mixer mix_t0_0010110 (.a(t0_00101100), .b(t0_00101101), .y(t0_0010110));
wire t0_00101100, t0_00101101;
mixer mix_t0_00101100 (.a(t0_001011000), .b(t0_001011001), .y(t0_00101100));
wire t0_001011000, t0_001011001;
mixer mix_t0_00101101 (.a(t0_001011010), .b(t0_001011011), .y(t0_00101101));
wire t0_001011010, t0_001011011;
mixer mix_t0_0010111 (.a(t0_00101110), .b(t0_00101111), .y(t0_0010111));
wire t0_00101110, t0_00101111;
mixer mix_t0_00101110 (.a(t0_001011100), .b(t0_001011101), .y(t0_00101110));
wire t0_001011100, t0_001011101;
mixer mix_t0_00101111 (.a(t0_001011110), .b(t0_001011111), .y(t0_00101111));
wire t0_001011110, t0_001011111;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_001100 (.a(t0_0011000), .b(t0_0011001), .y(t0_001100));
wire t0_0011000, t0_0011001;
mixer mix_t0_0011000 (.a(t0_00110000), .b(t0_00110001), .y(t0_0011000));
wire t0_00110000, t0_00110001;
mixer mix_t0_00110000 (.a(t0_001100000), .b(t0_001100001), .y(t0_00110000));
wire t0_001100000, t0_001100001;
mixer mix_t0_00110001 (.a(t0_001100010), .b(t0_001100011), .y(t0_00110001));
wire t0_001100010, t0_001100011;
mixer mix_t0_0011001 (.a(t0_00110010), .b(t0_00110011), .y(t0_0011001));
wire t0_00110010, t0_00110011;
mixer mix_t0_00110010 (.a(t0_001100100), .b(t0_001100101), .y(t0_00110010));
wire t0_001100100, t0_001100101;
mixer mix_t0_00110011 (.a(t0_001100110), .b(t0_001100111), .y(t0_00110011));
wire t0_001100110, t0_001100111;
mixer mix_t0_001101 (.a(t0_0011010), .b(t0_0011011), .y(t0_001101));
wire t0_0011010, t0_0011011;
mixer mix_t0_0011010 (.a(t0_00110100), .b(t0_00110101), .y(t0_0011010));
wire t0_00110100, t0_00110101;
mixer mix_t0_00110100 (.a(t0_001101000), .b(t0_001101001), .y(t0_00110100));
wire t0_001101000, t0_001101001;
mixer mix_t0_00110101 (.a(t0_001101010), .b(t0_001101011), .y(t0_00110101));
wire t0_001101010, t0_001101011;
mixer mix_t0_0011011 (.a(t0_00110110), .b(t0_00110111), .y(t0_0011011));
wire t0_00110110, t0_00110111;
mixer mix_t0_00110110 (.a(t0_001101100), .b(t0_001101101), .y(t0_00110110));
wire t0_001101100, t0_001101101;
mixer mix_t0_00110111 (.a(t0_001101110), .b(t0_001101111), .y(t0_00110111));
wire t0_001101110, t0_001101111;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_001110 (.a(t0_0011100), .b(t0_0011101), .y(t0_001110));
wire t0_0011100, t0_0011101;
mixer mix_t0_0011100 (.a(t0_00111000), .b(t0_00111001), .y(t0_0011100));
wire t0_00111000, t0_00111001;
mixer mix_t0_00111000 (.a(t0_001110000), .b(t0_001110001), .y(t0_00111000));
wire t0_001110000, t0_001110001;
mixer mix_t0_00111001 (.a(t0_001110010), .b(t0_001110011), .y(t0_00111001));
wire t0_001110010, t0_001110011;
mixer mix_t0_0011101 (.a(t0_00111010), .b(t0_00111011), .y(t0_0011101));
wire t0_00111010, t0_00111011;
mixer mix_t0_00111010 (.a(t0_001110100), .b(t0_001110101), .y(t0_00111010));
wire t0_001110100, t0_001110101;
mixer mix_t0_00111011 (.a(t0_001110110), .b(t0_001110111), .y(t0_00111011));
wire t0_001110110, t0_001110111;
mixer mix_t0_001111 (.a(t0_0011110), .b(t0_0011111), .y(t0_001111));
wire t0_0011110, t0_0011111;
mixer mix_t0_0011110 (.a(t0_00111100), .b(t0_00111101), .y(t0_0011110));
wire t0_00111100, t0_00111101;
mixer mix_t0_00111100 (.a(t0_001111000), .b(t0_001111001), .y(t0_00111100));
wire t0_001111000, t0_001111001;
mixer mix_t0_00111101 (.a(t0_001111010), .b(t0_001111011), .y(t0_00111101));
wire t0_001111010, t0_001111011;
mixer mix_t0_0011111 (.a(t0_00111110), .b(t0_00111111), .y(t0_0011111));
wire t0_00111110, t0_00111111;
mixer mix_t0_00111110 (.a(t0_001111100), .b(t0_001111101), .y(t0_00111110));
wire t0_001111100, t0_001111101;
mixer mix_t0_00111111 (.a(t0_001111110), .b(t0_001111111), .y(t0_00111111));
wire t0_001111110, t0_001111111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_010000 (.a(t0_0100000), .b(t0_0100001), .y(t0_010000));
wire t0_0100000, t0_0100001;
mixer mix_t0_0100000 (.a(t0_01000000), .b(t0_01000001), .y(t0_0100000));
wire t0_01000000, t0_01000001;
mixer mix_t0_01000000 (.a(t0_010000000), .b(t0_010000001), .y(t0_01000000));
wire t0_010000000, t0_010000001;
mixer mix_t0_01000001 (.a(t0_010000010), .b(t0_010000011), .y(t0_01000001));
wire t0_010000010, t0_010000011;
mixer mix_t0_0100001 (.a(t0_01000010), .b(t0_01000011), .y(t0_0100001));
wire t0_01000010, t0_01000011;
mixer mix_t0_01000010 (.a(t0_010000100), .b(t0_010000101), .y(t0_01000010));
wire t0_010000100, t0_010000101;
mixer mix_t0_01000011 (.a(t0_010000110), .b(t0_010000111), .y(t0_01000011));
wire t0_010000110, t0_010000111;
mixer mix_t0_010001 (.a(t0_0100010), .b(t0_0100011), .y(t0_010001));
wire t0_0100010, t0_0100011;
mixer mix_t0_0100010 (.a(t0_01000100), .b(t0_01000101), .y(t0_0100010));
wire t0_01000100, t0_01000101;
mixer mix_t0_01000100 (.a(t0_010001000), .b(t0_010001001), .y(t0_01000100));
wire t0_010001000, t0_010001001;
mixer mix_t0_01000101 (.a(t0_010001010), .b(t0_010001011), .y(t0_01000101));
wire t0_010001010, t0_010001011;
mixer mix_t0_0100011 (.a(t0_01000110), .b(t0_01000111), .y(t0_0100011));
wire t0_01000110, t0_01000111;
mixer mix_t0_01000110 (.a(t0_010001100), .b(t0_010001101), .y(t0_01000110));
wire t0_010001100, t0_010001101;
mixer mix_t0_01000111 (.a(t0_010001110), .b(t0_010001111), .y(t0_01000111));
wire t0_010001110, t0_010001111;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_010010 (.a(t0_0100100), .b(t0_0100101), .y(t0_010010));
wire t0_0100100, t0_0100101;
mixer mix_t0_0100100 (.a(t0_01001000), .b(t0_01001001), .y(t0_0100100));
wire t0_01001000, t0_01001001;
mixer mix_t0_01001000 (.a(t0_010010000), .b(t0_010010001), .y(t0_01001000));
wire t0_010010000, t0_010010001;
mixer mix_t0_01001001 (.a(t0_010010010), .b(t0_010010011), .y(t0_01001001));
wire t0_010010010, t0_010010011;
mixer mix_t0_0100101 (.a(t0_01001010), .b(t0_01001011), .y(t0_0100101));
wire t0_01001010, t0_01001011;
mixer mix_t0_01001010 (.a(t0_010010100), .b(t0_010010101), .y(t0_01001010));
wire t0_010010100, t0_010010101;
mixer mix_t0_01001011 (.a(t0_010010110), .b(t0_010010111), .y(t0_01001011));
wire t0_010010110, t0_010010111;
mixer mix_t0_010011 (.a(t0_0100110), .b(t0_0100111), .y(t0_010011));
wire t0_0100110, t0_0100111;
mixer mix_t0_0100110 (.a(t0_01001100), .b(t0_01001101), .y(t0_0100110));
wire t0_01001100, t0_01001101;
mixer mix_t0_01001100 (.a(t0_010011000), .b(t0_010011001), .y(t0_01001100));
wire t0_010011000, t0_010011001;
mixer mix_t0_01001101 (.a(t0_010011010), .b(t0_010011011), .y(t0_01001101));
wire t0_010011010, t0_010011011;
mixer mix_t0_0100111 (.a(t0_01001110), .b(t0_01001111), .y(t0_0100111));
wire t0_01001110, t0_01001111;
mixer mix_t0_01001110 (.a(t0_010011100), .b(t0_010011101), .y(t0_01001110));
wire t0_010011100, t0_010011101;
mixer mix_t0_01001111 (.a(t0_010011110), .b(t0_010011111), .y(t0_01001111));
wire t0_010011110, t0_010011111;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_010100 (.a(t0_0101000), .b(t0_0101001), .y(t0_010100));
wire t0_0101000, t0_0101001;
mixer mix_t0_0101000 (.a(t0_01010000), .b(t0_01010001), .y(t0_0101000));
wire t0_01010000, t0_01010001;
mixer mix_t0_01010000 (.a(t0_010100000), .b(t0_010100001), .y(t0_01010000));
wire t0_010100000, t0_010100001;
mixer mix_t0_01010001 (.a(t0_010100010), .b(t0_010100011), .y(t0_01010001));
wire t0_010100010, t0_010100011;
mixer mix_t0_0101001 (.a(t0_01010010), .b(t0_01010011), .y(t0_0101001));
wire t0_01010010, t0_01010011;
mixer mix_t0_01010010 (.a(t0_010100100), .b(t0_010100101), .y(t0_01010010));
wire t0_010100100, t0_010100101;
mixer mix_t0_01010011 (.a(t0_010100110), .b(t0_010100111), .y(t0_01010011));
wire t0_010100110, t0_010100111;
mixer mix_t0_010101 (.a(t0_0101010), .b(t0_0101011), .y(t0_010101));
wire t0_0101010, t0_0101011;
mixer mix_t0_0101010 (.a(t0_01010100), .b(t0_01010101), .y(t0_0101010));
wire t0_01010100, t0_01010101;
mixer mix_t0_01010100 (.a(t0_010101000), .b(t0_010101001), .y(t0_01010100));
wire t0_010101000, t0_010101001;
mixer mix_t0_01010101 (.a(t0_010101010), .b(t0_010101011), .y(t0_01010101));
wire t0_010101010, t0_010101011;
mixer mix_t0_0101011 (.a(t0_01010110), .b(t0_01010111), .y(t0_0101011));
wire t0_01010110, t0_01010111;
mixer mix_t0_01010110 (.a(t0_010101100), .b(t0_010101101), .y(t0_01010110));
wire t0_010101100, t0_010101101;
mixer mix_t0_01010111 (.a(t0_010101110), .b(t0_010101111), .y(t0_01010111));
wire t0_010101110, t0_010101111;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_010110 (.a(t0_0101100), .b(t0_0101101), .y(t0_010110));
wire t0_0101100, t0_0101101;
mixer mix_t0_0101100 (.a(t0_01011000), .b(t0_01011001), .y(t0_0101100));
wire t0_01011000, t0_01011001;
mixer mix_t0_01011000 (.a(t0_010110000), .b(t0_010110001), .y(t0_01011000));
wire t0_010110000, t0_010110001;
mixer mix_t0_01011001 (.a(t0_010110010), .b(t0_010110011), .y(t0_01011001));
wire t0_010110010, t0_010110011;
mixer mix_t0_0101101 (.a(t0_01011010), .b(t0_01011011), .y(t0_0101101));
wire t0_01011010, t0_01011011;
mixer mix_t0_01011010 (.a(t0_010110100), .b(t0_010110101), .y(t0_01011010));
wire t0_010110100, t0_010110101;
mixer mix_t0_01011011 (.a(t0_010110110), .b(t0_010110111), .y(t0_01011011));
wire t0_010110110, t0_010110111;
mixer mix_t0_010111 (.a(t0_0101110), .b(t0_0101111), .y(t0_010111));
wire t0_0101110, t0_0101111;
mixer mix_t0_0101110 (.a(t0_01011100), .b(t0_01011101), .y(t0_0101110));
wire t0_01011100, t0_01011101;
mixer mix_t0_01011100 (.a(t0_010111000), .b(t0_010111001), .y(t0_01011100));
wire t0_010111000, t0_010111001;
mixer mix_t0_01011101 (.a(t0_010111010), .b(t0_010111011), .y(t0_01011101));
wire t0_010111010, t0_010111011;
mixer mix_t0_0101111 (.a(t0_01011110), .b(t0_01011111), .y(t0_0101111));
wire t0_01011110, t0_01011111;
mixer mix_t0_01011110 (.a(t0_010111100), .b(t0_010111101), .y(t0_01011110));
wire t0_010111100, t0_010111101;
mixer mix_t0_01011111 (.a(t0_010111110), .b(t0_010111111), .y(t0_01011111));
wire t0_010111110, t0_010111111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_011000 (.a(t0_0110000), .b(t0_0110001), .y(t0_011000));
wire t0_0110000, t0_0110001;
mixer mix_t0_0110000 (.a(t0_01100000), .b(t0_01100001), .y(t0_0110000));
wire t0_01100000, t0_01100001;
mixer mix_t0_01100000 (.a(t0_011000000), .b(t0_011000001), .y(t0_01100000));
wire t0_011000000, t0_011000001;
mixer mix_t0_01100001 (.a(t0_011000010), .b(t0_011000011), .y(t0_01100001));
wire t0_011000010, t0_011000011;
mixer mix_t0_0110001 (.a(t0_01100010), .b(t0_01100011), .y(t0_0110001));
wire t0_01100010, t0_01100011;
mixer mix_t0_01100010 (.a(t0_011000100), .b(t0_011000101), .y(t0_01100010));
wire t0_011000100, t0_011000101;
mixer mix_t0_01100011 (.a(t0_011000110), .b(t0_011000111), .y(t0_01100011));
wire t0_011000110, t0_011000111;
mixer mix_t0_011001 (.a(t0_0110010), .b(t0_0110011), .y(t0_011001));
wire t0_0110010, t0_0110011;
mixer mix_t0_0110010 (.a(t0_01100100), .b(t0_01100101), .y(t0_0110010));
wire t0_01100100, t0_01100101;
mixer mix_t0_01100100 (.a(t0_011001000), .b(t0_011001001), .y(t0_01100100));
wire t0_011001000, t0_011001001;
mixer mix_t0_01100101 (.a(t0_011001010), .b(t0_011001011), .y(t0_01100101));
wire t0_011001010, t0_011001011;
mixer mix_t0_0110011 (.a(t0_01100110), .b(t0_01100111), .y(t0_0110011));
wire t0_01100110, t0_01100111;
mixer mix_t0_01100110 (.a(t0_011001100), .b(t0_011001101), .y(t0_01100110));
wire t0_011001100, t0_011001101;
mixer mix_t0_01100111 (.a(t0_011001110), .b(t0_011001111), .y(t0_01100111));
wire t0_011001110, t0_011001111;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_011010 (.a(t0_0110100), .b(t0_0110101), .y(t0_011010));
wire t0_0110100, t0_0110101;
mixer mix_t0_0110100 (.a(t0_01101000), .b(t0_01101001), .y(t0_0110100));
wire t0_01101000, t0_01101001;
mixer mix_t0_01101000 (.a(t0_011010000), .b(t0_011010001), .y(t0_01101000));
wire t0_011010000, t0_011010001;
mixer mix_t0_01101001 (.a(t0_011010010), .b(t0_011010011), .y(t0_01101001));
wire t0_011010010, t0_011010011;
mixer mix_t0_0110101 (.a(t0_01101010), .b(t0_01101011), .y(t0_0110101));
wire t0_01101010, t0_01101011;
mixer mix_t0_01101010 (.a(t0_011010100), .b(t0_011010101), .y(t0_01101010));
wire t0_011010100, t0_011010101;
mixer mix_t0_01101011 (.a(t0_011010110), .b(t0_011010111), .y(t0_01101011));
wire t0_011010110, t0_011010111;
mixer mix_t0_011011 (.a(t0_0110110), .b(t0_0110111), .y(t0_011011));
wire t0_0110110, t0_0110111;
mixer mix_t0_0110110 (.a(t0_01101100), .b(t0_01101101), .y(t0_0110110));
wire t0_01101100, t0_01101101;
mixer mix_t0_01101100 (.a(t0_011011000), .b(t0_011011001), .y(t0_01101100));
wire t0_011011000, t0_011011001;
mixer mix_t0_01101101 (.a(t0_011011010), .b(t0_011011011), .y(t0_01101101));
wire t0_011011010, t0_011011011;
mixer mix_t0_0110111 (.a(t0_01101110), .b(t0_01101111), .y(t0_0110111));
wire t0_01101110, t0_01101111;
mixer mix_t0_01101110 (.a(t0_011011100), .b(t0_011011101), .y(t0_01101110));
wire t0_011011100, t0_011011101;
mixer mix_t0_01101111 (.a(t0_011011110), .b(t0_011011111), .y(t0_01101111));
wire t0_011011110, t0_011011111;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_011100 (.a(t0_0111000), .b(t0_0111001), .y(t0_011100));
wire t0_0111000, t0_0111001;
mixer mix_t0_0111000 (.a(t0_01110000), .b(t0_01110001), .y(t0_0111000));
wire t0_01110000, t0_01110001;
mixer mix_t0_01110000 (.a(t0_011100000), .b(t0_011100001), .y(t0_01110000));
wire t0_011100000, t0_011100001;
mixer mix_t0_01110001 (.a(t0_011100010), .b(t0_011100011), .y(t0_01110001));
wire t0_011100010, t0_011100011;
mixer mix_t0_0111001 (.a(t0_01110010), .b(t0_01110011), .y(t0_0111001));
wire t0_01110010, t0_01110011;
mixer mix_t0_01110010 (.a(t0_011100100), .b(t0_011100101), .y(t0_01110010));
wire t0_011100100, t0_011100101;
mixer mix_t0_01110011 (.a(t0_011100110), .b(t0_011100111), .y(t0_01110011));
wire t0_011100110, t0_011100111;
mixer mix_t0_011101 (.a(t0_0111010), .b(t0_0111011), .y(t0_011101));
wire t0_0111010, t0_0111011;
mixer mix_t0_0111010 (.a(t0_01110100), .b(t0_01110101), .y(t0_0111010));
wire t0_01110100, t0_01110101;
mixer mix_t0_01110100 (.a(t0_011101000), .b(t0_011101001), .y(t0_01110100));
wire t0_011101000, t0_011101001;
mixer mix_t0_01110101 (.a(t0_011101010), .b(t0_011101011), .y(t0_01110101));
wire t0_011101010, t0_011101011;
mixer mix_t0_0111011 (.a(t0_01110110), .b(t0_01110111), .y(t0_0111011));
wire t0_01110110, t0_01110111;
mixer mix_t0_01110110 (.a(t0_011101100), .b(t0_011101101), .y(t0_01110110));
wire t0_011101100, t0_011101101;
mixer mix_t0_01110111 (.a(t0_011101110), .b(t0_011101111), .y(t0_01110111));
wire t0_011101110, t0_011101111;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
mixer mix_t0_011110 (.a(t0_0111100), .b(t0_0111101), .y(t0_011110));
wire t0_0111100, t0_0111101;
mixer mix_t0_0111100 (.a(t0_01111000), .b(t0_01111001), .y(t0_0111100));
wire t0_01111000, t0_01111001;
mixer mix_t0_01111000 (.a(t0_011110000), .b(t0_011110001), .y(t0_01111000));
wire t0_011110000, t0_011110001;
mixer mix_t0_01111001 (.a(t0_011110010), .b(t0_011110011), .y(t0_01111001));
wire t0_011110010, t0_011110011;
mixer mix_t0_0111101 (.a(t0_01111010), .b(t0_01111011), .y(t0_0111101));
wire t0_01111010, t0_01111011;
mixer mix_t0_01111010 (.a(t0_011110100), .b(t0_011110101), .y(t0_01111010));
wire t0_011110100, t0_011110101;
mixer mix_t0_01111011 (.a(t0_011110110), .b(t0_011110111), .y(t0_01111011));
wire t0_011110110, t0_011110111;
mixer mix_t0_011111 (.a(t0_0111110), .b(t0_0111111), .y(t0_011111));
wire t0_0111110, t0_0111111;
mixer mix_t0_0111110 (.a(t0_01111100), .b(t0_01111101), .y(t0_0111110));
wire t0_01111100, t0_01111101;
mixer mix_t0_01111100 (.a(t0_011111000), .b(t0_011111001), .y(t0_01111100));
wire t0_011111000, t0_011111001;
mixer mix_t0_01111101 (.a(t0_011111010), .b(t0_011111011), .y(t0_01111101));
wire t0_011111010, t0_011111011;
mixer mix_t0_0111111 (.a(t0_01111110), .b(t0_01111111), .y(t0_0111111));
wire t0_01111110, t0_01111111;
mixer mix_t0_01111110 (.a(t0_011111100), .b(t0_011111101), .y(t0_01111110));
wire t0_011111100, t0_011111101;
mixer mix_t0_01111111 (.a(t0_011111110), .b(t0_011111111), .y(t0_01111111));
wire t0_011111110, t0_011111111;
mixer mix_t1_0 (.a(t1_00), .b(t1_01), .y(t1_0));
wire t1_00, t1_01;
mixer mix_t1_00 (.a(t1_000), .b(t1_001), .y(t1_00));
wire t1_000, t1_001;
mixer mix_t1_000 (.a(t1_0000), .b(t1_0001), .y(t1_000));
wire t1_0000, t1_0001;
mixer mix_t1_0000 (.a(t1_00000), .b(t1_00001), .y(t1_0000));
wire t1_00000, t1_00001;
mixer mix_t1_00000 (.a(t1_000000), .b(t1_000001), .y(t1_00000));
wire t1_000000, t1_000001;
mixer mix_t1_000000 (.a(t1_0000000), .b(t1_0000001), .y(t1_000000));
wire t1_0000000, t1_0000001;
mixer mix_t1_0000000 (.a(t1_00000000), .b(t1_00000001), .y(t1_0000000));
wire t1_00000000, t1_00000001;
mixer mix_t1_00000000 (.a(t1_000000000), .b(t1_000000001), .y(t1_00000000));
wire t1_000000000, t1_000000001;
mixer mix_t1_00000001 (.a(t1_000000010), .b(t1_000000011), .y(t1_00000001));
wire t1_000000010, t1_000000011;
mixer mix_t1_0000001 (.a(t1_00000010), .b(t1_00000011), .y(t1_0000001));
wire t1_00000010, t1_00000011;
mixer mix_t1_00000010 (.a(t1_000000100), .b(t1_000000101), .y(t1_00000010));
wire t1_000000100, t1_000000101;
mixer mix_t1_00000011 (.a(t1_000000110), .b(t1_000000111), .y(t1_00000011));
wire t1_000000110, t1_000000111;
mixer mix_t1_000001 (.a(t1_0000010), .b(t1_0000011), .y(t1_000001));
wire t1_0000010, t1_0000011;
mixer mix_t1_0000010 (.a(t1_00000100), .b(t1_00000101), .y(t1_0000010));
wire t1_00000100, t1_00000101;
mixer mix_t1_00000100 (.a(t1_000001000), .b(t1_000001001), .y(t1_00000100));
wire t1_000001000, t1_000001001;
mixer mix_t1_00000101 (.a(t1_000001010), .b(t1_000001011), .y(t1_00000101));
wire t1_000001010, t1_000001011;
mixer mix_t1_0000011 (.a(t1_00000110), .b(t1_00000111), .y(t1_0000011));
wire t1_00000110, t1_00000111;
mixer mix_t1_00000110 (.a(t1_000001100), .b(t1_000001101), .y(t1_00000110));
wire t1_000001100, t1_000001101;
mixer mix_t1_00000111 (.a(t1_000001110), .b(t1_000001111), .y(t1_00000111));
wire t1_000001110, t1_000001111;
mixer mix_t1_00001 (.a(t1_000010), .b(t1_000011), .y(t1_00001));
wire t1_000010, t1_000011;
mixer mix_t1_000010 (.a(t1_0000100), .b(t1_0000101), .y(t1_000010));
wire t1_0000100, t1_0000101;
mixer mix_t1_0000100 (.a(t1_00001000), .b(t1_00001001), .y(t1_0000100));
wire t1_00001000, t1_00001001;
mixer mix_t1_00001000 (.a(t1_000010000), .b(t1_000010001), .y(t1_00001000));
wire t1_000010000, t1_000010001;
mixer mix_t1_00001001 (.a(t1_000010010), .b(t1_000010011), .y(t1_00001001));
wire t1_000010010, t1_000010011;
mixer mix_t1_0000101 (.a(t1_00001010), .b(t1_00001011), .y(t1_0000101));
wire t1_00001010, t1_00001011;
mixer mix_t1_00001010 (.a(t1_000010100), .b(t1_000010101), .y(t1_00001010));
wire t1_000010100, t1_000010101;
mixer mix_t1_00001011 (.a(t1_000010110), .b(t1_000010111), .y(t1_00001011));
wire t1_000010110, t1_000010111;
mixer mix_t1_000011 (.a(t1_0000110), .b(t1_0000111), .y(t1_000011));
wire t1_0000110, t1_0000111;
mixer mix_t1_0000110 (.a(t1_00001100), .b(t1_00001101), .y(t1_0000110));
wire t1_00001100, t1_00001101;
mixer mix_t1_00001100 (.a(t1_000011000), .b(t1_000011001), .y(t1_00001100));
wire t1_000011000, t1_000011001;
mixer mix_t1_00001101 (.a(t1_000011010), .b(t1_000011011), .y(t1_00001101));
wire t1_000011010, t1_000011011;
mixer mix_t1_0000111 (.a(t1_00001110), .b(t1_00001111), .y(t1_0000111));
wire t1_00001110, t1_00001111;
mixer mix_t1_00001110 (.a(t1_000011100), .b(t1_000011101), .y(t1_00001110));
wire t1_000011100, t1_000011101;
mixer mix_t1_00001111 (.a(t1_000011110), .b(t1_000011111), .y(t1_00001111));
wire t1_000011110, t1_000011111;
mixer mix_t1_0001 (.a(t1_00010), .b(t1_00011), .y(t1_0001));
wire t1_00010, t1_00011;
mixer mix_t1_00010 (.a(t1_000100), .b(t1_000101), .y(t1_00010));
wire t1_000100, t1_000101;
mixer mix_t1_000100 (.a(t1_0001000), .b(t1_0001001), .y(t1_000100));
wire t1_0001000, t1_0001001;
mixer mix_t1_0001000 (.a(t1_00010000), .b(t1_00010001), .y(t1_0001000));
wire t1_00010000, t1_00010001;
mixer mix_t1_00010000 (.a(t1_000100000), .b(t1_000100001), .y(t1_00010000));
wire t1_000100000, t1_000100001;
mixer mix_t1_00010001 (.a(t1_000100010), .b(t1_000100011), .y(t1_00010001));
wire t1_000100010, t1_000100011;
mixer mix_t1_0001001 (.a(t1_00010010), .b(t1_00010011), .y(t1_0001001));
wire t1_00010010, t1_00010011;
mixer mix_t1_00010010 (.a(t1_000100100), .b(t1_000100101), .y(t1_00010010));
wire t1_000100100, t1_000100101;
mixer mix_t1_00010011 (.a(t1_000100110), .b(t1_000100111), .y(t1_00010011));
wire t1_000100110, t1_000100111;
mixer mix_t1_000101 (.a(t1_0001010), .b(t1_0001011), .y(t1_000101));
wire t1_0001010, t1_0001011;
mixer mix_t1_0001010 (.a(t1_00010100), .b(t1_00010101), .y(t1_0001010));
wire t1_00010100, t1_00010101;
mixer mix_t1_00010100 (.a(t1_000101000), .b(t1_000101001), .y(t1_00010100));
wire t1_000101000, t1_000101001;
mixer mix_t1_00010101 (.a(t1_000101010), .b(t1_000101011), .y(t1_00010101));
wire t1_000101010, t1_000101011;
mixer mix_t1_0001011 (.a(t1_00010110), .b(t1_00010111), .y(t1_0001011));
wire t1_00010110, t1_00010111;
mixer mix_t1_00010110 (.a(t1_000101100), .b(t1_000101101), .y(t1_00010110));
wire t1_000101100, t1_000101101;
mixer mix_t1_00010111 (.a(t1_000101110), .b(t1_000101111), .y(t1_00010111));
wire t1_000101110, t1_000101111;
mixer mix_t1_00011 (.a(t1_000110), .b(t1_000111), .y(t1_00011));
wire t1_000110, t1_000111;
mixer mix_t1_000110 (.a(t1_0001100), .b(t1_0001101), .y(t1_000110));
wire t1_0001100, t1_0001101;
mixer mix_t1_0001100 (.a(t1_00011000), .b(t1_00011001), .y(t1_0001100));
wire t1_00011000, t1_00011001;
mixer mix_t1_00011000 (.a(t1_000110000), .b(t1_000110001), .y(t1_00011000));
wire t1_000110000, t1_000110001;
mixer mix_t1_00011001 (.a(t1_000110010), .b(t1_000110011), .y(t1_00011001));
wire t1_000110010, t1_000110011;
mixer mix_t1_0001101 (.a(t1_00011010), .b(t1_00011011), .y(t1_0001101));
wire t1_00011010, t1_00011011;
mixer mix_t1_00011010 (.a(t1_000110100), .b(t1_000110101), .y(t1_00011010));
wire t1_000110100, t1_000110101;
mixer mix_t1_00011011 (.a(t1_000110110), .b(t1_000110111), .y(t1_00011011));
wire t1_000110110, t1_000110111;
mixer mix_t1_000111 (.a(t1_0001110), .b(t1_0001111), .y(t1_000111));
wire t1_0001110, t1_0001111;
mixer mix_t1_0001110 (.a(t1_00011100), .b(t1_00011101), .y(t1_0001110));
wire t1_00011100, t1_00011101;
mixer mix_t1_00011100 (.a(t1_000111000), .b(t1_000111001), .y(t1_00011100));
wire t1_000111000, t1_000111001;
mixer mix_t1_00011101 (.a(t1_000111010), .b(t1_000111011), .y(t1_00011101));
wire t1_000111010, t1_000111011;
mixer mix_t1_0001111 (.a(t1_00011110), .b(t1_00011111), .y(t1_0001111));
wire t1_00011110, t1_00011111;
mixer mix_t1_00011110 (.a(t1_000111100), .b(t1_000111101), .y(t1_00011110));
wire t1_000111100, t1_000111101;
mixer mix_t1_00011111 (.a(t1_000111110), .b(t1_000111111), .y(t1_00011111));
wire t1_000111110, t1_000111111;
mixer mix_t1_001 (.a(t1_0010), .b(t1_0011), .y(t1_001));
wire t1_0010, t1_0011;
mixer mix_t1_0010 (.a(t1_00100), .b(t1_00101), .y(t1_0010));
wire t1_00100, t1_00101;
mixer mix_t1_00100 (.a(t1_001000), .b(t1_001001), .y(t1_00100));
wire t1_001000, t1_001001;
mixer mix_t1_001000 (.a(t1_0010000), .b(t1_0010001), .y(t1_001000));
wire t1_0010000, t1_0010001;
mixer mix_t1_0010000 (.a(t1_00100000), .b(t1_00100001), .y(t1_0010000));
wire t1_00100000, t1_00100001;
mixer mix_t1_00100000 (.a(t1_001000000), .b(t1_001000001), .y(t1_00100000));
wire t1_001000000, t1_001000001;
mixer mix_t1_00100001 (.a(t1_001000010), .b(t1_001000011), .y(t1_00100001));
wire t1_001000010, t1_001000011;
mixer mix_t1_0010001 (.a(t1_00100010), .b(t1_00100011), .y(t1_0010001));
wire t1_00100010, t1_00100011;
mixer mix_t1_00100010 (.a(t1_001000100), .b(t1_001000101), .y(t1_00100010));
wire t1_001000100, t1_001000101;
mixer mix_t1_00100011 (.a(t1_001000110), .b(t1_001000111), .y(t1_00100011));
wire t1_001000110, t1_001000111;
mixer mix_t1_001001 (.a(t1_0010010), .b(t1_0010011), .y(t1_001001));
wire t1_0010010, t1_0010011;
mixer mix_t1_0010010 (.a(t1_00100100), .b(t1_00100101), .y(t1_0010010));
wire t1_00100100, t1_00100101;
mixer mix_t1_00100100 (.a(t1_001001000), .b(t1_001001001), .y(t1_00100100));
wire t1_001001000, t1_001001001;
mixer mix_t1_00100101 (.a(t1_001001010), .b(t1_001001011), .y(t1_00100101));
wire t1_001001010, t1_001001011;
mixer mix_t1_0010011 (.a(t1_00100110), .b(t1_00100111), .y(t1_0010011));
wire t1_00100110, t1_00100111;
mixer mix_t1_00100110 (.a(t1_001001100), .b(t1_001001101), .y(t1_00100110));
wire t1_001001100, t1_001001101;
mixer mix_t1_00100111 (.a(t1_001001110), .b(t1_001001111), .y(t1_00100111));
wire t1_001001110, t1_001001111;
mixer mix_t1_00101 (.a(t1_001010), .b(t1_001011), .y(t1_00101));
wire t1_001010, t1_001011;
mixer mix_t1_001010 (.a(t1_0010100), .b(t1_0010101), .y(t1_001010));
wire t1_0010100, t1_0010101;
mixer mix_t1_0010100 (.a(t1_00101000), .b(t1_00101001), .y(t1_0010100));
wire t1_00101000, t1_00101001;
mixer mix_t1_00101000 (.a(t1_001010000), .b(t1_001010001), .y(t1_00101000));
wire t1_001010000, t1_001010001;
mixer mix_t1_00101001 (.a(t1_001010010), .b(t1_001010011), .y(t1_00101001));
wire t1_001010010, t1_001010011;
mixer mix_t1_0010101 (.a(t1_00101010), .b(t1_00101011), .y(t1_0010101));
wire t1_00101010, t1_00101011;
mixer mix_t1_00101010 (.a(t1_001010100), .b(t1_001010101), .y(t1_00101010));
wire t1_001010100, t1_001010101;
mixer mix_t1_00101011 (.a(t1_001010110), .b(t1_001010111), .y(t1_00101011));
wire t1_001010110, t1_001010111;
mixer mix_t1_001011 (.a(t1_0010110), .b(t1_0010111), .y(t1_001011));
wire t1_0010110, t1_0010111;
mixer mix_t1_0010110 (.a(t1_00101100), .b(t1_00101101), .y(t1_0010110));
wire t1_00101100, t1_00101101;
mixer mix_t1_00101100 (.a(t1_001011000), .b(t1_001011001), .y(t1_00101100));
wire t1_001011000, t1_001011001;
mixer mix_t1_00101101 (.a(t1_001011010), .b(t1_001011011), .y(t1_00101101));
wire t1_001011010, t1_001011011;
mixer mix_t1_0010111 (.a(t1_00101110), .b(t1_00101111), .y(t1_0010111));
wire t1_00101110, t1_00101111;
mixer mix_t1_00101110 (.a(t1_001011100), .b(t1_001011101), .y(t1_00101110));
wire t1_001011100, t1_001011101;
mixer mix_t1_00101111 (.a(t1_001011110), .b(t1_001011111), .y(t1_00101111));
wire t1_001011110, t1_001011111;
mixer mix_t1_0011 (.a(t1_00110), .b(t1_00111), .y(t1_0011));
wire t1_00110, t1_00111;
mixer mix_t1_00110 (.a(t1_001100), .b(t1_001101), .y(t1_00110));
wire t1_001100, t1_001101;
mixer mix_t1_001100 (.a(t1_0011000), .b(t1_0011001), .y(t1_001100));
wire t1_0011000, t1_0011001;
mixer mix_t1_0011000 (.a(t1_00110000), .b(t1_00110001), .y(t1_0011000));
wire t1_00110000, t1_00110001;
mixer mix_t1_00110000 (.a(t1_001100000), .b(t1_001100001), .y(t1_00110000));
wire t1_001100000, t1_001100001;
mixer mix_t1_00110001 (.a(t1_001100010), .b(t1_001100011), .y(t1_00110001));
wire t1_001100010, t1_001100011;
mixer mix_t1_0011001 (.a(t1_00110010), .b(t1_00110011), .y(t1_0011001));
wire t1_00110010, t1_00110011;
mixer mix_t1_00110010 (.a(t1_001100100), .b(t1_001100101), .y(t1_00110010));
wire t1_001100100, t1_001100101;
mixer mix_t1_00110011 (.a(t1_001100110), .b(t1_001100111), .y(t1_00110011));
wire t1_001100110, t1_001100111;
mixer mix_t1_001101 (.a(t1_0011010), .b(t1_0011011), .y(t1_001101));
wire t1_0011010, t1_0011011;
mixer mix_t1_0011010 (.a(t1_00110100), .b(t1_00110101), .y(t1_0011010));
wire t1_00110100, t1_00110101;
mixer mix_t1_00110100 (.a(t1_001101000), .b(t1_001101001), .y(t1_00110100));
wire t1_001101000, t1_001101001;
mixer mix_t1_00110101 (.a(t1_001101010), .b(t1_001101011), .y(t1_00110101));
wire t1_001101010, t1_001101011;
mixer mix_t1_0011011 (.a(t1_00110110), .b(t1_00110111), .y(t1_0011011));
wire t1_00110110, t1_00110111;
mixer mix_t1_00110110 (.a(t1_001101100), .b(t1_001101101), .y(t1_00110110));
wire t1_001101100, t1_001101101;
mixer mix_t1_00110111 (.a(t1_001101110), .b(t1_001101111), .y(t1_00110111));
wire t1_001101110, t1_001101111;
mixer mix_t1_00111 (.a(t1_001110), .b(t1_001111), .y(t1_00111));
wire t1_001110, t1_001111;
mixer mix_t1_001110 (.a(t1_0011100), .b(t1_0011101), .y(t1_001110));
wire t1_0011100, t1_0011101;
mixer mix_t1_0011100 (.a(t1_00111000), .b(t1_00111001), .y(t1_0011100));
wire t1_00111000, t1_00111001;
mixer mix_t1_00111000 (.a(t1_001110000), .b(t1_001110001), .y(t1_00111000));
wire t1_001110000, t1_001110001;
mixer mix_t1_00111001 (.a(t1_001110010), .b(t1_001110011), .y(t1_00111001));
wire t1_001110010, t1_001110011;
mixer mix_t1_0011101 (.a(t1_00111010), .b(t1_00111011), .y(t1_0011101));
wire t1_00111010, t1_00111011;
mixer mix_t1_00111010 (.a(t1_001110100), .b(t1_001110101), .y(t1_00111010));
wire t1_001110100, t1_001110101;
mixer mix_t1_00111011 (.a(t1_001110110), .b(t1_001110111), .y(t1_00111011));
wire t1_001110110, t1_001110111;
mixer mix_t1_001111 (.a(t1_0011110), .b(t1_0011111), .y(t1_001111));
wire t1_0011110, t1_0011111;
mixer mix_t1_0011110 (.a(t1_00111100), .b(t1_00111101), .y(t1_0011110));
wire t1_00111100, t1_00111101;
mixer mix_t1_00111100 (.a(t1_001111000), .b(t1_001111001), .y(t1_00111100));
wire t1_001111000, t1_001111001;
mixer mix_t1_00111101 (.a(t1_001111010), .b(t1_001111011), .y(t1_00111101));
wire t1_001111010, t1_001111011;
mixer mix_t1_0011111 (.a(t1_00111110), .b(t1_00111111), .y(t1_0011111));
wire t1_00111110, t1_00111111;
mixer mix_t1_00111110 (.a(t1_001111100), .b(t1_001111101), .y(t1_00111110));
wire t1_001111100, t1_001111101;
mixer mix_t1_00111111 (.a(t1_001111110), .b(t1_001111111), .y(t1_00111111));
wire t1_001111110, t1_001111111;
mixer mix_t1_01 (.a(t1_010), .b(t1_011), .y(t1_01));
wire t1_010, t1_011;
mixer mix_t1_010 (.a(t1_0100), .b(t1_0101), .y(t1_010));
wire t1_0100, t1_0101;
mixer mix_t1_0100 (.a(t1_01000), .b(t1_01001), .y(t1_0100));
wire t1_01000, t1_01001;
mixer mix_t1_01000 (.a(t1_010000), .b(t1_010001), .y(t1_01000));
wire t1_010000, t1_010001;
mixer mix_t1_010000 (.a(t1_0100000), .b(t1_0100001), .y(t1_010000));
wire t1_0100000, t1_0100001;
mixer mix_t1_0100000 (.a(t1_01000000), .b(t1_01000001), .y(t1_0100000));
wire t1_01000000, t1_01000001;
mixer mix_t1_01000000 (.a(t1_010000000), .b(t1_010000001), .y(t1_01000000));
wire t1_010000000, t1_010000001;
mixer mix_t1_01000001 (.a(t1_010000010), .b(t1_010000011), .y(t1_01000001));
wire t1_010000010, t1_010000011;
mixer mix_t1_0100001 (.a(t1_01000010), .b(t1_01000011), .y(t1_0100001));
wire t1_01000010, t1_01000011;
mixer mix_t1_01000010 (.a(t1_010000100), .b(t1_010000101), .y(t1_01000010));
wire t1_010000100, t1_010000101;
mixer mix_t1_01000011 (.a(t1_010000110), .b(t1_010000111), .y(t1_01000011));
wire t1_010000110, t1_010000111;
mixer mix_t1_010001 (.a(t1_0100010), .b(t1_0100011), .y(t1_010001));
wire t1_0100010, t1_0100011;
mixer mix_t1_0100010 (.a(t1_01000100), .b(t1_01000101), .y(t1_0100010));
wire t1_01000100, t1_01000101;
mixer mix_t1_01000100 (.a(t1_010001000), .b(t1_010001001), .y(t1_01000100));
wire t1_010001000, t1_010001001;
mixer mix_t1_01000101 (.a(t1_010001010), .b(t1_010001011), .y(t1_01000101));
wire t1_010001010, t1_010001011;
mixer mix_t1_0100011 (.a(t1_01000110), .b(t1_01000111), .y(t1_0100011));
wire t1_01000110, t1_01000111;
mixer mix_t1_01000110 (.a(t1_010001100), .b(t1_010001101), .y(t1_01000110));
wire t1_010001100, t1_010001101;
mixer mix_t1_01000111 (.a(t1_010001110), .b(t1_010001111), .y(t1_01000111));
wire t1_010001110, t1_010001111;
mixer mix_t1_01001 (.a(t1_010010), .b(t1_010011), .y(t1_01001));
wire t1_010010, t1_010011;
mixer mix_t1_010010 (.a(t1_0100100), .b(t1_0100101), .y(t1_010010));
wire t1_0100100, t1_0100101;
mixer mix_t1_0100100 (.a(t1_01001000), .b(t1_01001001), .y(t1_0100100));
wire t1_01001000, t1_01001001;
mixer mix_t1_01001000 (.a(t1_010010000), .b(t1_010010001), .y(t1_01001000));
wire t1_010010000, t1_010010001;
mixer mix_t1_01001001 (.a(t1_010010010), .b(t1_010010011), .y(t1_01001001));
wire t1_010010010, t1_010010011;
mixer mix_t1_0100101 (.a(t1_01001010), .b(t1_01001011), .y(t1_0100101));
wire t1_01001010, t1_01001011;
mixer mix_t1_01001010 (.a(t1_010010100), .b(t1_010010101), .y(t1_01001010));
wire t1_010010100, t1_010010101;
mixer mix_t1_01001011 (.a(t1_010010110), .b(t1_010010111), .y(t1_01001011));
wire t1_010010110, t1_010010111;
mixer mix_t1_010011 (.a(t1_0100110), .b(t1_0100111), .y(t1_010011));
wire t1_0100110, t1_0100111;
mixer mix_t1_0100110 (.a(t1_01001100), .b(t1_01001101), .y(t1_0100110));
wire t1_01001100, t1_01001101;
mixer mix_t1_01001100 (.a(t1_010011000), .b(t1_010011001), .y(t1_01001100));
wire t1_010011000, t1_010011001;
mixer mix_t1_01001101 (.a(t1_010011010), .b(t1_010011011), .y(t1_01001101));
wire t1_010011010, t1_010011011;
mixer mix_t1_0100111 (.a(t1_01001110), .b(t1_01001111), .y(t1_0100111));
wire t1_01001110, t1_01001111;
mixer mix_t1_01001110 (.a(t1_010011100), .b(t1_010011101), .y(t1_01001110));
wire t1_010011100, t1_010011101;
mixer mix_t1_01001111 (.a(t1_010011110), .b(t1_010011111), .y(t1_01001111));
wire t1_010011110, t1_010011111;
mixer mix_t1_0101 (.a(t1_01010), .b(t1_01011), .y(t1_0101));
wire t1_01010, t1_01011;
mixer mix_t1_01010 (.a(t1_010100), .b(t1_010101), .y(t1_01010));
wire t1_010100, t1_010101;
mixer mix_t1_010100 (.a(t1_0101000), .b(t1_0101001), .y(t1_010100));
wire t1_0101000, t1_0101001;
mixer mix_t1_0101000 (.a(t1_01010000), .b(t1_01010001), .y(t1_0101000));
wire t1_01010000, t1_01010001;
mixer mix_t1_01010000 (.a(t1_010100000), .b(t1_010100001), .y(t1_01010000));
wire t1_010100000, t1_010100001;
mixer mix_t1_01010001 (.a(t1_010100010), .b(t1_010100011), .y(t1_01010001));
wire t1_010100010, t1_010100011;
mixer mix_t1_0101001 (.a(t1_01010010), .b(t1_01010011), .y(t1_0101001));
wire t1_01010010, t1_01010011;
mixer mix_t1_01010010 (.a(t1_010100100), .b(t1_010100101), .y(t1_01010010));
wire t1_010100100, t1_010100101;
mixer mix_t1_01010011 (.a(t1_010100110), .b(t1_010100111), .y(t1_01010011));
wire t1_010100110, t1_010100111;
mixer mix_t1_010101 (.a(t1_0101010), .b(t1_0101011), .y(t1_010101));
wire t1_0101010, t1_0101011;
mixer mix_t1_0101010 (.a(t1_01010100), .b(t1_01010101), .y(t1_0101010));
wire t1_01010100, t1_01010101;
mixer mix_t1_01010100 (.a(t1_010101000), .b(t1_010101001), .y(t1_01010100));
wire t1_010101000, t1_010101001;
mixer mix_t1_01010101 (.a(t1_010101010), .b(t1_010101011), .y(t1_01010101));
wire t1_010101010, t1_010101011;
mixer mix_t1_0101011 (.a(t1_01010110), .b(t1_01010111), .y(t1_0101011));
wire t1_01010110, t1_01010111;
mixer mix_t1_01010110 (.a(t1_010101100), .b(t1_010101101), .y(t1_01010110));
wire t1_010101100, t1_010101101;
mixer mix_t1_01010111 (.a(t1_010101110), .b(t1_010101111), .y(t1_01010111));
wire t1_010101110, t1_010101111;
mixer mix_t1_01011 (.a(t1_010110), .b(t1_010111), .y(t1_01011));
wire t1_010110, t1_010111;
mixer mix_t1_010110 (.a(t1_0101100), .b(t1_0101101), .y(t1_010110));
wire t1_0101100, t1_0101101;
mixer mix_t1_0101100 (.a(t1_01011000), .b(t1_01011001), .y(t1_0101100));
wire t1_01011000, t1_01011001;
mixer mix_t1_01011000 (.a(t1_010110000), .b(t1_010110001), .y(t1_01011000));
wire t1_010110000, t1_010110001;
mixer mix_t1_01011001 (.a(t1_010110010), .b(t1_010110011), .y(t1_01011001));
wire t1_010110010, t1_010110011;
mixer mix_t1_0101101 (.a(t1_01011010), .b(t1_01011011), .y(t1_0101101));
wire t1_01011010, t1_01011011;
mixer mix_t1_01011010 (.a(t1_010110100), .b(t1_010110101), .y(t1_01011010));
wire t1_010110100, t1_010110101;
mixer mix_t1_01011011 (.a(t1_010110110), .b(t1_010110111), .y(t1_01011011));
wire t1_010110110, t1_010110111;
mixer mix_t1_010111 (.a(t1_0101110), .b(t1_0101111), .y(t1_010111));
wire t1_0101110, t1_0101111;
mixer mix_t1_0101110 (.a(t1_01011100), .b(t1_01011101), .y(t1_0101110));
wire t1_01011100, t1_01011101;
mixer mix_t1_01011100 (.a(t1_010111000), .b(t1_010111001), .y(t1_01011100));
wire t1_010111000, t1_010111001;
mixer mix_t1_01011101 (.a(t1_010111010), .b(t1_010111011), .y(t1_01011101));
wire t1_010111010, t1_010111011;
mixer mix_t1_0101111 (.a(t1_01011110), .b(t1_01011111), .y(t1_0101111));
wire t1_01011110, t1_01011111;
mixer mix_t1_01011110 (.a(t1_010111100), .b(t1_010111101), .y(t1_01011110));
wire t1_010111100, t1_010111101;
mixer mix_t1_01011111 (.a(t1_010111110), .b(t1_010111111), .y(t1_01011111));
wire t1_010111110, t1_010111111;
mixer mix_t1_011 (.a(t1_0110), .b(t1_0111), .y(t1_011));
wire t1_0110, t1_0111;
mixer mix_t1_0110 (.a(t1_01100), .b(t1_01101), .y(t1_0110));
wire t1_01100, t1_01101;
mixer mix_t1_01100 (.a(t1_011000), .b(t1_011001), .y(t1_01100));
wire t1_011000, t1_011001;
mixer mix_t1_011000 (.a(t1_0110000), .b(t1_0110001), .y(t1_011000));
wire t1_0110000, t1_0110001;
mixer mix_t1_0110000 (.a(t1_01100000), .b(t1_01100001), .y(t1_0110000));
wire t1_01100000, t1_01100001;
mixer mix_t1_01100000 (.a(t1_011000000), .b(t1_011000001), .y(t1_01100000));
wire t1_011000000, t1_011000001;
mixer mix_t1_01100001 (.a(t1_011000010), .b(t1_011000011), .y(t1_01100001));
wire t1_011000010, t1_011000011;
mixer mix_t1_0110001 (.a(t1_01100010), .b(t1_01100011), .y(t1_0110001));
wire t1_01100010, t1_01100011;
mixer mix_t1_01100010 (.a(t1_011000100), .b(t1_011000101), .y(t1_01100010));
wire t1_011000100, t1_011000101;
mixer mix_t1_01100011 (.a(t1_011000110), .b(t1_011000111), .y(t1_01100011));
wire t1_011000110, t1_011000111;
mixer mix_t1_011001 (.a(t1_0110010), .b(t1_0110011), .y(t1_011001));
wire t1_0110010, t1_0110011;
mixer mix_t1_0110010 (.a(t1_01100100), .b(t1_01100101), .y(t1_0110010));
wire t1_01100100, t1_01100101;
mixer mix_t1_01100100 (.a(t1_011001000), .b(t1_011001001), .y(t1_01100100));
wire t1_011001000, t1_011001001;
mixer mix_t1_01100101 (.a(t1_011001010), .b(t1_011001011), .y(t1_01100101));
wire t1_011001010, t1_011001011;
mixer mix_t1_0110011 (.a(t1_01100110), .b(t1_01100111), .y(t1_0110011));
wire t1_01100110, t1_01100111;
mixer mix_t1_01100110 (.a(t1_011001100), .b(t1_011001101), .y(t1_01100110));
wire t1_011001100, t1_011001101;
mixer mix_t1_01100111 (.a(t1_011001110), .b(t1_011001111), .y(t1_01100111));
wire t1_011001110, t1_011001111;
mixer mix_t1_01101 (.a(t1_011010), .b(t1_011011), .y(t1_01101));
wire t1_011010, t1_011011;
mixer mix_t1_011010 (.a(t1_0110100), .b(t1_0110101), .y(t1_011010));
wire t1_0110100, t1_0110101;
mixer mix_t1_0110100 (.a(t1_01101000), .b(t1_01101001), .y(t1_0110100));
wire t1_01101000, t1_01101001;
mixer mix_t1_01101000 (.a(t1_011010000), .b(t1_011010001), .y(t1_01101000));
wire t1_011010000, t1_011010001;
mixer mix_t1_01101001 (.a(t1_011010010), .b(t1_011010011), .y(t1_01101001));
wire t1_011010010, t1_011010011;
mixer mix_t1_0110101 (.a(t1_01101010), .b(t1_01101011), .y(t1_0110101));
wire t1_01101010, t1_01101011;
mixer mix_t1_01101010 (.a(t1_011010100), .b(t1_011010101), .y(t1_01101010));
wire t1_011010100, t1_011010101;
mixer mix_t1_01101011 (.a(t1_011010110), .b(t1_011010111), .y(t1_01101011));
wire t1_011010110, t1_011010111;
mixer mix_t1_011011 (.a(t1_0110110), .b(t1_0110111), .y(t1_011011));
wire t1_0110110, t1_0110111;
mixer mix_t1_0110110 (.a(t1_01101100), .b(t1_01101101), .y(t1_0110110));
wire t1_01101100, t1_01101101;
mixer mix_t1_01101100 (.a(t1_011011000), .b(t1_011011001), .y(t1_01101100));
wire t1_011011000, t1_011011001;
mixer mix_t1_01101101 (.a(t1_011011010), .b(t1_011011011), .y(t1_01101101));
wire t1_011011010, t1_011011011;
mixer mix_t1_0110111 (.a(t1_01101110), .b(t1_01101111), .y(t1_0110111));
wire t1_01101110, t1_01101111;
mixer mix_t1_01101110 (.a(t1_011011100), .b(t1_011011101), .y(t1_01101110));
wire t1_011011100, t1_011011101;
mixer mix_t1_01101111 (.a(t1_011011110), .b(t1_011011111), .y(t1_01101111));
wire t1_011011110, t1_011011111;
mixer mix_t1_0111 (.a(t1_01110), .b(t1_01111), .y(t1_0111));
wire t1_01110, t1_01111;
mixer mix_t1_01110 (.a(t1_011100), .b(t1_011101), .y(t1_01110));
wire t1_011100, t1_011101;
mixer mix_t1_011100 (.a(t1_0111000), .b(t1_0111001), .y(t1_011100));
wire t1_0111000, t1_0111001;
mixer mix_t1_0111000 (.a(t1_01110000), .b(t1_01110001), .y(t1_0111000));
wire t1_01110000, t1_01110001;
mixer mix_t1_01110000 (.a(t1_011100000), .b(t1_011100001), .y(t1_01110000));
wire t1_011100000, t1_011100001;
mixer mix_t1_01110001 (.a(t1_011100010), .b(t1_011100011), .y(t1_01110001));
wire t1_011100010, t1_011100011;
mixer mix_t1_0111001 (.a(t1_01110010), .b(t1_01110011), .y(t1_0111001));
wire t1_01110010, t1_01110011;
mixer mix_t1_01110010 (.a(t1_011100100), .b(t1_011100101), .y(t1_01110010));
wire t1_011100100, t1_011100101;
mixer mix_t1_01110011 (.a(t1_011100110), .b(t1_011100111), .y(t1_01110011));
wire t1_011100110, t1_011100111;
mixer mix_t1_011101 (.a(t1_0111010), .b(t1_0111011), .y(t1_011101));
wire t1_0111010, t1_0111011;
mixer mix_t1_0111010 (.a(t1_01110100), .b(t1_01110101), .y(t1_0111010));
wire t1_01110100, t1_01110101;
mixer mix_t1_01110100 (.a(t1_011101000), .b(t1_011101001), .y(t1_01110100));
wire t1_011101000, t1_011101001;
mixer mix_t1_01110101 (.a(t1_011101010), .b(t1_011101011), .y(t1_01110101));
wire t1_011101010, t1_011101011;
mixer mix_t1_0111011 (.a(t1_01110110), .b(t1_01110111), .y(t1_0111011));
wire t1_01110110, t1_01110111;
mixer mix_t1_01110110 (.a(t1_011101100), .b(t1_011101101), .y(t1_01110110));
wire t1_011101100, t1_011101101;
mixer mix_t1_01110111 (.a(t1_011101110), .b(t1_011101111), .y(t1_01110111));
wire t1_011101110, t1_011101111;
mixer mix_t1_01111 (.a(t1_011110), .b(t1_011111), .y(t1_01111));
wire t1_011110, t1_011111;
mixer mix_t1_011110 (.a(t1_0111100), .b(t1_0111101), .y(t1_011110));
wire t1_0111100, t1_0111101;
mixer mix_t1_0111100 (.a(t1_01111000), .b(t1_01111001), .y(t1_0111100));
wire t1_01111000, t1_01111001;
mixer mix_t1_01111000 (.a(t1_011110000), .b(t1_011110001), .y(t1_01111000));
wire t1_011110000, t1_011110001;
mixer mix_t1_01111001 (.a(t1_011110010), .b(t1_011110011), .y(t1_01111001));
wire t1_011110010, t1_011110011;
mixer mix_t1_0111101 (.a(t1_01111010), .b(t1_01111011), .y(t1_0111101));
wire t1_01111010, t1_01111011;
mixer mix_t1_01111010 (.a(t1_011110100), .b(t1_011110101), .y(t1_01111010));
wire t1_011110100, t1_011110101;
mixer mix_t1_01111011 (.a(t1_011110110), .b(t1_011110111), .y(t1_01111011));
wire t1_011110110, t1_011110111;
mixer mix_t1_011111 (.a(t1_0111110), .b(t1_0111111), .y(t1_011111));
wire t1_0111110, t1_0111111;
mixer mix_t1_0111110 (.a(t1_01111100), .b(t1_01111101), .y(t1_0111110));
wire t1_01111100, t1_01111101;
mixer mix_t1_01111100 (.a(t1_011111000), .b(t1_011111001), .y(t1_01111100));
wire t1_011111000, t1_011111001;
mixer mix_t1_01111101 (.a(t1_011111010), .b(t1_011111011), .y(t1_01111101));
wire t1_011111010, t1_011111011;
mixer mix_t1_0111111 (.a(t1_01111110), .b(t1_01111111), .y(t1_0111111));
wire t1_01111110, t1_01111111;
mixer mix_t1_01111110 (.a(t1_011111100), .b(t1_011111101), .y(t1_01111110));
wire t1_011111100, t1_011111101;
mixer mix_t1_01111111 (.a(t1_011111110), .b(t1_011111111), .y(t1_01111111));
wire t1_011111110, t1_011111111;
mixer mix_t2_0 (.a(t2_00), .b(t2_01), .y(t2_0));
wire t2_00, t2_01;
mixer mix_t2_00 (.a(t2_000), .b(t2_001), .y(t2_00));
wire t2_000, t2_001;
mixer mix_t2_000 (.a(t2_0000), .b(t2_0001), .y(t2_000));
wire t2_0000, t2_0001;
mixer mix_t2_0000 (.a(t2_00000), .b(t2_00001), .y(t2_0000));
wire t2_00000, t2_00001;
mixer mix_t2_00000 (.a(t2_000000), .b(t2_000001), .y(t2_00000));
wire t2_000000, t2_000001;
mixer mix_t2_000000 (.a(t2_0000000), .b(t2_0000001), .y(t2_000000));
wire t2_0000000, t2_0000001;
mixer mix_t2_0000000 (.a(t2_00000000), .b(t2_00000001), .y(t2_0000000));
wire t2_00000000, t2_00000001;
mixer mix_t2_00000000 (.a(t2_000000000), .b(t2_000000001), .y(t2_00000000));
wire t2_000000000, t2_000000001;
mixer mix_t2_00000001 (.a(t2_000000010), .b(t2_000000011), .y(t2_00000001));
wire t2_000000010, t2_000000011;
mixer mix_t2_0000001 (.a(t2_00000010), .b(t2_00000011), .y(t2_0000001));
wire t2_00000010, t2_00000011;
mixer mix_t2_00000010 (.a(t2_000000100), .b(t2_000000101), .y(t2_00000010));
wire t2_000000100, t2_000000101;
mixer mix_t2_00000011 (.a(t2_000000110), .b(t2_000000111), .y(t2_00000011));
wire t2_000000110, t2_000000111;
mixer mix_t2_000001 (.a(t2_0000010), .b(t2_0000011), .y(t2_000001));
wire t2_0000010, t2_0000011;
mixer mix_t2_0000010 (.a(t2_00000100), .b(t2_00000101), .y(t2_0000010));
wire t2_00000100, t2_00000101;
mixer mix_t2_00000100 (.a(t2_000001000), .b(t2_000001001), .y(t2_00000100));
wire t2_000001000, t2_000001001;
mixer mix_t2_00000101 (.a(t2_000001010), .b(t2_000001011), .y(t2_00000101));
wire t2_000001010, t2_000001011;
mixer mix_t2_0000011 (.a(t2_00000110), .b(t2_00000111), .y(t2_0000011));
wire t2_00000110, t2_00000111;
mixer mix_t2_00000110 (.a(t2_000001100), .b(t2_000001101), .y(t2_00000110));
wire t2_000001100, t2_000001101;
mixer mix_t2_00000111 (.a(t2_000001110), .b(t2_000001111), .y(t2_00000111));
wire t2_000001110, t2_000001111;
mixer mix_t2_00001 (.a(t2_000010), .b(t2_000011), .y(t2_00001));
wire t2_000010, t2_000011;
mixer mix_t2_000010 (.a(t2_0000100), .b(t2_0000101), .y(t2_000010));
wire t2_0000100, t2_0000101;
mixer mix_t2_0000100 (.a(t2_00001000), .b(t2_00001001), .y(t2_0000100));
wire t2_00001000, t2_00001001;
mixer mix_t2_00001000 (.a(t2_000010000), .b(t2_000010001), .y(t2_00001000));
wire t2_000010000, t2_000010001;
mixer mix_t2_00001001 (.a(t2_000010010), .b(t2_000010011), .y(t2_00001001));
wire t2_000010010, t2_000010011;
mixer mix_t2_0000101 (.a(t2_00001010), .b(t2_00001011), .y(t2_0000101));
wire t2_00001010, t2_00001011;
mixer mix_t2_00001010 (.a(t2_000010100), .b(t2_000010101), .y(t2_00001010));
wire t2_000010100, t2_000010101;
mixer mix_t2_00001011 (.a(t2_000010110), .b(t2_000010111), .y(t2_00001011));
wire t2_000010110, t2_000010111;
mixer mix_t2_000011 (.a(t2_0000110), .b(t2_0000111), .y(t2_000011));
wire t2_0000110, t2_0000111;
mixer mix_t2_0000110 (.a(t2_00001100), .b(t2_00001101), .y(t2_0000110));
wire t2_00001100, t2_00001101;
mixer mix_t2_00001100 (.a(t2_000011000), .b(t2_000011001), .y(t2_00001100));
wire t2_000011000, t2_000011001;
mixer mix_t2_00001101 (.a(t2_000011010), .b(t2_000011011), .y(t2_00001101));
wire t2_000011010, t2_000011011;
mixer mix_t2_0000111 (.a(t2_00001110), .b(t2_00001111), .y(t2_0000111));
wire t2_00001110, t2_00001111;
mixer mix_t2_00001110 (.a(t2_000011100), .b(t2_000011101), .y(t2_00001110));
wire t2_000011100, t2_000011101;
mixer mix_t2_00001111 (.a(t2_000011110), .b(t2_000011111), .y(t2_00001111));
wire t2_000011110, t2_000011111;
mixer mix_t2_0001 (.a(t2_00010), .b(t2_00011), .y(t2_0001));
wire t2_00010, t2_00011;
mixer mix_t2_00010 (.a(t2_000100), .b(t2_000101), .y(t2_00010));
wire t2_000100, t2_000101;
mixer mix_t2_000100 (.a(t2_0001000), .b(t2_0001001), .y(t2_000100));
wire t2_0001000, t2_0001001;
mixer mix_t2_0001000 (.a(t2_00010000), .b(t2_00010001), .y(t2_0001000));
wire t2_00010000, t2_00010001;
mixer mix_t2_00010000 (.a(t2_000100000), .b(t2_000100001), .y(t2_00010000));
wire t2_000100000, t2_000100001;
mixer mix_t2_00010001 (.a(t2_000100010), .b(t2_000100011), .y(t2_00010001));
wire t2_000100010, t2_000100011;
mixer mix_t2_0001001 (.a(t2_00010010), .b(t2_00010011), .y(t2_0001001));
wire t2_00010010, t2_00010011;
mixer mix_t2_00010010 (.a(t2_000100100), .b(t2_000100101), .y(t2_00010010));
wire t2_000100100, t2_000100101;
mixer mix_t2_00010011 (.a(t2_000100110), .b(t2_000100111), .y(t2_00010011));
wire t2_000100110, t2_000100111;
mixer mix_t2_000101 (.a(t2_0001010), .b(t2_0001011), .y(t2_000101));
wire t2_0001010, t2_0001011;
mixer mix_t2_0001010 (.a(t2_00010100), .b(t2_00010101), .y(t2_0001010));
wire t2_00010100, t2_00010101;
mixer mix_t2_00010100 (.a(t2_000101000), .b(t2_000101001), .y(t2_00010100));
wire t2_000101000, t2_000101001;
mixer mix_t2_00010101 (.a(t2_000101010), .b(t2_000101011), .y(t2_00010101));
wire t2_000101010, t2_000101011;
mixer mix_t2_0001011 (.a(t2_00010110), .b(t2_00010111), .y(t2_0001011));
wire t2_00010110, t2_00010111;
mixer mix_t2_00010110 (.a(t2_000101100), .b(t2_000101101), .y(t2_00010110));
wire t2_000101100, t2_000101101;
mixer mix_t2_00010111 (.a(t2_000101110), .b(t2_000101111), .y(t2_00010111));
wire t2_000101110, t2_000101111;
mixer mix_t2_00011 (.a(t2_000110), .b(t2_000111), .y(t2_00011));
wire t2_000110, t2_000111;
mixer mix_t2_000110 (.a(t2_0001100), .b(t2_0001101), .y(t2_000110));
wire t2_0001100, t2_0001101;
mixer mix_t2_0001100 (.a(t2_00011000), .b(t2_00011001), .y(t2_0001100));
wire t2_00011000, t2_00011001;
mixer mix_t2_00011000 (.a(t2_000110000), .b(t2_000110001), .y(t2_00011000));
wire t2_000110000, t2_000110001;
mixer mix_t2_00011001 (.a(t2_000110010), .b(t2_000110011), .y(t2_00011001));
wire t2_000110010, t2_000110011;
mixer mix_t2_0001101 (.a(t2_00011010), .b(t2_00011011), .y(t2_0001101));
wire t2_00011010, t2_00011011;
mixer mix_t2_00011010 (.a(t2_000110100), .b(t2_000110101), .y(t2_00011010));
wire t2_000110100, t2_000110101;
mixer mix_t2_00011011 (.a(t2_000110110), .b(t2_000110111), .y(t2_00011011));
wire t2_000110110, t2_000110111;
mixer mix_t2_000111 (.a(t2_0001110), .b(t2_0001111), .y(t2_000111));
wire t2_0001110, t2_0001111;
mixer mix_t2_0001110 (.a(t2_00011100), .b(t2_00011101), .y(t2_0001110));
wire t2_00011100, t2_00011101;
mixer mix_t2_00011100 (.a(t2_000111000), .b(t2_000111001), .y(t2_00011100));
wire t2_000111000, t2_000111001;
mixer mix_t2_00011101 (.a(t2_000111010), .b(t2_000111011), .y(t2_00011101));
wire t2_000111010, t2_000111011;
mixer mix_t2_0001111 (.a(t2_00011110), .b(t2_00011111), .y(t2_0001111));
wire t2_00011110, t2_00011111;
mixer mix_t2_00011110 (.a(t2_000111100), .b(t2_000111101), .y(t2_00011110));
wire t2_000111100, t2_000111101;
mixer mix_t2_00011111 (.a(t2_000111110), .b(t2_000111111), .y(t2_00011111));
wire t2_000111110, t2_000111111;
mixer mix_t2_001 (.a(t2_0010), .b(t2_0011), .y(t2_001));
wire t2_0010, t2_0011;
mixer mix_t2_0010 (.a(t2_00100), .b(t2_00101), .y(t2_0010));
wire t2_00100, t2_00101;
mixer mix_t2_00100 (.a(t2_001000), .b(t2_001001), .y(t2_00100));
wire t2_001000, t2_001001;
mixer mix_t2_001000 (.a(t2_0010000), .b(t2_0010001), .y(t2_001000));
wire t2_0010000, t2_0010001;
mixer mix_t2_0010000 (.a(t2_00100000), .b(t2_00100001), .y(t2_0010000));
wire t2_00100000, t2_00100001;
mixer mix_t2_00100000 (.a(t2_001000000), .b(t2_001000001), .y(t2_00100000));
wire t2_001000000, t2_001000001;
mixer mix_t2_00100001 (.a(t2_001000010), .b(t2_001000011), .y(t2_00100001));
wire t2_001000010, t2_001000011;
mixer mix_t2_0010001 (.a(t2_00100010), .b(t2_00100011), .y(t2_0010001));
wire t2_00100010, t2_00100011;
mixer mix_t2_00100010 (.a(t2_001000100), .b(t2_001000101), .y(t2_00100010));
wire t2_001000100, t2_001000101;
mixer mix_t2_00100011 (.a(t2_001000110), .b(t2_001000111), .y(t2_00100011));
wire t2_001000110, t2_001000111;
mixer mix_t2_001001 (.a(t2_0010010), .b(t2_0010011), .y(t2_001001));
wire t2_0010010, t2_0010011;
mixer mix_t2_0010010 (.a(t2_00100100), .b(t2_00100101), .y(t2_0010010));
wire t2_00100100, t2_00100101;
mixer mix_t2_00100100 (.a(t2_001001000), .b(t2_001001001), .y(t2_00100100));
wire t2_001001000, t2_001001001;
mixer mix_t2_00100101 (.a(t2_001001010), .b(t2_001001011), .y(t2_00100101));
wire t2_001001010, t2_001001011;
mixer mix_t2_0010011 (.a(t2_00100110), .b(t2_00100111), .y(t2_0010011));
wire t2_00100110, t2_00100111;
mixer mix_t2_00100110 (.a(t2_001001100), .b(t2_001001101), .y(t2_00100110));
wire t2_001001100, t2_001001101;
mixer mix_t2_00100111 (.a(t2_001001110), .b(t2_001001111), .y(t2_00100111));
wire t2_001001110, t2_001001111;
mixer mix_t2_00101 (.a(t2_001010), .b(t2_001011), .y(t2_00101));
wire t2_001010, t2_001011;
mixer mix_t2_001010 (.a(t2_0010100), .b(t2_0010101), .y(t2_001010));
wire t2_0010100, t2_0010101;
mixer mix_t2_0010100 (.a(t2_00101000), .b(t2_00101001), .y(t2_0010100));
wire t2_00101000, t2_00101001;
mixer mix_t2_00101000 (.a(t2_001010000), .b(t2_001010001), .y(t2_00101000));
wire t2_001010000, t2_001010001;
mixer mix_t2_00101001 (.a(t2_001010010), .b(t2_001010011), .y(t2_00101001));
wire t2_001010010, t2_001010011;
mixer mix_t2_0010101 (.a(t2_00101010), .b(t2_00101011), .y(t2_0010101));
wire t2_00101010, t2_00101011;
mixer mix_t2_00101010 (.a(t2_001010100), .b(t2_001010101), .y(t2_00101010));
wire t2_001010100, t2_001010101;
mixer mix_t2_00101011 (.a(t2_001010110), .b(t2_001010111), .y(t2_00101011));
wire t2_001010110, t2_001010111;
mixer mix_t2_001011 (.a(t2_0010110), .b(t2_0010111), .y(t2_001011));
wire t2_0010110, t2_0010111;
mixer mix_t2_0010110 (.a(t2_00101100), .b(t2_00101101), .y(t2_0010110));
wire t2_00101100, t2_00101101;
mixer mix_t2_00101100 (.a(t2_001011000), .b(t2_001011001), .y(t2_00101100));
wire t2_001011000, t2_001011001;
mixer mix_t2_00101101 (.a(t2_001011010), .b(t2_001011011), .y(t2_00101101));
wire t2_001011010, t2_001011011;
mixer mix_t2_0010111 (.a(t2_00101110), .b(t2_00101111), .y(t2_0010111));
wire t2_00101110, t2_00101111;
mixer mix_t2_00101110 (.a(t2_001011100), .b(t2_001011101), .y(t2_00101110));
wire t2_001011100, t2_001011101;
mixer mix_t2_00101111 (.a(t2_001011110), .b(t2_001011111), .y(t2_00101111));
wire t2_001011110, t2_001011111;
mixer mix_t2_0011 (.a(t2_00110), .b(t2_00111), .y(t2_0011));
wire t2_00110, t2_00111;
mixer mix_t2_00110 (.a(t2_001100), .b(t2_001101), .y(t2_00110));
wire t2_001100, t2_001101;
mixer mix_t2_001100 (.a(t2_0011000), .b(t2_0011001), .y(t2_001100));
wire t2_0011000, t2_0011001;
mixer mix_t2_0011000 (.a(t2_00110000), .b(t2_00110001), .y(t2_0011000));
wire t2_00110000, t2_00110001;
mixer mix_t2_00110000 (.a(t2_001100000), .b(t2_001100001), .y(t2_00110000));
wire t2_001100000, t2_001100001;
mixer mix_t2_00110001 (.a(t2_001100010), .b(t2_001100011), .y(t2_00110001));
wire t2_001100010, t2_001100011;
mixer mix_t2_0011001 (.a(t2_00110010), .b(t2_00110011), .y(t2_0011001));
wire t2_00110010, t2_00110011;
mixer mix_t2_00110010 (.a(t2_001100100), .b(t2_001100101), .y(t2_00110010));
wire t2_001100100, t2_001100101;
mixer mix_t2_00110011 (.a(t2_001100110), .b(t2_001100111), .y(t2_00110011));
wire t2_001100110, t2_001100111;
mixer mix_t2_001101 (.a(t2_0011010), .b(t2_0011011), .y(t2_001101));
wire t2_0011010, t2_0011011;
mixer mix_t2_0011010 (.a(t2_00110100), .b(t2_00110101), .y(t2_0011010));
wire t2_00110100, t2_00110101;
mixer mix_t2_00110100 (.a(t2_001101000), .b(t2_001101001), .y(t2_00110100));
wire t2_001101000, t2_001101001;
mixer mix_t2_00110101 (.a(t2_001101010), .b(t2_001101011), .y(t2_00110101));
wire t2_001101010, t2_001101011;
mixer mix_t2_0011011 (.a(t2_00110110), .b(t2_00110111), .y(t2_0011011));
wire t2_00110110, t2_00110111;
mixer mix_t2_00110110 (.a(t2_001101100), .b(t2_001101101), .y(t2_00110110));
wire t2_001101100, t2_001101101;
mixer mix_t2_00110111 (.a(t2_001101110), .b(t2_001101111), .y(t2_00110111));
wire t2_001101110, t2_001101111;
mixer mix_t2_00111 (.a(t2_001110), .b(t2_001111), .y(t2_00111));
wire t2_001110, t2_001111;
mixer mix_t2_001110 (.a(t2_0011100), .b(t2_0011101), .y(t2_001110));
wire t2_0011100, t2_0011101;
mixer mix_t2_0011100 (.a(t2_00111000), .b(t2_00111001), .y(t2_0011100));
wire t2_00111000, t2_00111001;
mixer mix_t2_00111000 (.a(t2_001110000), .b(t2_001110001), .y(t2_00111000));
wire t2_001110000, t2_001110001;
mixer mix_t2_00111001 (.a(t2_001110010), .b(t2_001110011), .y(t2_00111001));
wire t2_001110010, t2_001110011;
mixer mix_t2_0011101 (.a(t2_00111010), .b(t2_00111011), .y(t2_0011101));
wire t2_00111010, t2_00111011;
mixer mix_t2_00111010 (.a(t2_001110100), .b(t2_001110101), .y(t2_00111010));
wire t2_001110100, t2_001110101;
mixer mix_t2_00111011 (.a(t2_001110110), .b(t2_001110111), .y(t2_00111011));
wire t2_001110110, t2_001110111;
mixer mix_t2_001111 (.a(t2_0011110), .b(t2_0011111), .y(t2_001111));
wire t2_0011110, t2_0011111;
mixer mix_t2_0011110 (.a(t2_00111100), .b(t2_00111101), .y(t2_0011110));
wire t2_00111100, t2_00111101;
mixer mix_t2_00111100 (.a(t2_001111000), .b(t2_001111001), .y(t2_00111100));
wire t2_001111000, t2_001111001;
mixer mix_t2_00111101 (.a(t2_001111010), .b(t2_001111011), .y(t2_00111101));
wire t2_001111010, t2_001111011;
mixer mix_t2_0011111 (.a(t2_00111110), .b(t2_00111111), .y(t2_0011111));
wire t2_00111110, t2_00111111;
mixer mix_t2_00111110 (.a(t2_001111100), .b(t2_001111101), .y(t2_00111110));
wire t2_001111100, t2_001111101;
mixer mix_t2_00111111 (.a(t2_001111110), .b(t2_001111111), .y(t2_00111111));
wire t2_001111110, t2_001111111;
mixer mix_t2_01 (.a(t2_010), .b(t2_011), .y(t2_01));
wire t2_010, t2_011;
mixer mix_t2_010 (.a(t2_0100), .b(t2_0101), .y(t2_010));
wire t2_0100, t2_0101;
mixer mix_t2_0100 (.a(t2_01000), .b(t2_01001), .y(t2_0100));
wire t2_01000, t2_01001;
mixer mix_t2_01000 (.a(t2_010000), .b(t2_010001), .y(t2_01000));
wire t2_010000, t2_010001;
mixer mix_t2_010000 (.a(t2_0100000), .b(t2_0100001), .y(t2_010000));
wire t2_0100000, t2_0100001;
mixer mix_t2_0100000 (.a(t2_01000000), .b(t2_01000001), .y(t2_0100000));
wire t2_01000000, t2_01000001;
mixer mix_t2_01000000 (.a(t2_010000000), .b(t2_010000001), .y(t2_01000000));
wire t2_010000000, t2_010000001;
mixer mix_t2_01000001 (.a(t2_010000010), .b(t2_010000011), .y(t2_01000001));
wire t2_010000010, t2_010000011;
mixer mix_t2_0100001 (.a(t2_01000010), .b(t2_01000011), .y(t2_0100001));
wire t2_01000010, t2_01000011;
mixer mix_t2_01000010 (.a(t2_010000100), .b(t2_010000101), .y(t2_01000010));
wire t2_010000100, t2_010000101;
mixer mix_t2_01000011 (.a(t2_010000110), .b(t2_010000111), .y(t2_01000011));
wire t2_010000110, t2_010000111;
mixer mix_t2_010001 (.a(t2_0100010), .b(t2_0100011), .y(t2_010001));
wire t2_0100010, t2_0100011;
mixer mix_t2_0100010 (.a(t2_01000100), .b(t2_01000101), .y(t2_0100010));
wire t2_01000100, t2_01000101;
mixer mix_t2_01000100 (.a(t2_010001000), .b(t2_010001001), .y(t2_01000100));
wire t2_010001000, t2_010001001;
mixer mix_t2_01000101 (.a(t2_010001010), .b(t2_010001011), .y(t2_01000101));
wire t2_010001010, t2_010001011;
mixer mix_t2_0100011 (.a(t2_01000110), .b(t2_01000111), .y(t2_0100011));
wire t2_01000110, t2_01000111;
mixer mix_t2_01000110 (.a(t2_010001100), .b(t2_010001101), .y(t2_01000110));
wire t2_010001100, t2_010001101;
mixer mix_t2_01000111 (.a(t2_010001110), .b(t2_010001111), .y(t2_01000111));
wire t2_010001110, t2_010001111;
mixer mix_t2_01001 (.a(t2_010010), .b(t2_010011), .y(t2_01001));
wire t2_010010, t2_010011;
mixer mix_t2_010010 (.a(t2_0100100), .b(t2_0100101), .y(t2_010010));
wire t2_0100100, t2_0100101;
mixer mix_t2_0100100 (.a(t2_01001000), .b(t2_01001001), .y(t2_0100100));
wire t2_01001000, t2_01001001;
mixer mix_t2_01001000 (.a(t2_010010000), .b(t2_010010001), .y(t2_01001000));
wire t2_010010000, t2_010010001;
mixer mix_t2_01001001 (.a(t2_010010010), .b(t2_010010011), .y(t2_01001001));
wire t2_010010010, t2_010010011;
mixer mix_t2_0100101 (.a(t2_01001010), .b(t2_01001011), .y(t2_0100101));
wire t2_01001010, t2_01001011;
mixer mix_t2_01001010 (.a(t2_010010100), .b(t2_010010101), .y(t2_01001010));
wire t2_010010100, t2_010010101;
mixer mix_t2_01001011 (.a(t2_010010110), .b(t2_010010111), .y(t2_01001011));
wire t2_010010110, t2_010010111;
mixer mix_t2_010011 (.a(t2_0100110), .b(t2_0100111), .y(t2_010011));
wire t2_0100110, t2_0100111;
mixer mix_t2_0100110 (.a(t2_01001100), .b(t2_01001101), .y(t2_0100110));
wire t2_01001100, t2_01001101;
mixer mix_t2_01001100 (.a(t2_010011000), .b(t2_010011001), .y(t2_01001100));
wire t2_010011000, t2_010011001;
mixer mix_t2_01001101 (.a(t2_010011010), .b(t2_010011011), .y(t2_01001101));
wire t2_010011010, t2_010011011;
mixer mix_t2_0100111 (.a(t2_01001110), .b(t2_01001111), .y(t2_0100111));
wire t2_01001110, t2_01001111;
mixer mix_t2_01001110 (.a(t2_010011100), .b(t2_010011101), .y(t2_01001110));
wire t2_010011100, t2_010011101;
mixer mix_t2_01001111 (.a(t2_010011110), .b(t2_010011111), .y(t2_01001111));
wire t2_010011110, t2_010011111;
mixer mix_t2_0101 (.a(t2_01010), .b(t2_01011), .y(t2_0101));
wire t2_01010, t2_01011;
mixer mix_t2_01010 (.a(t2_010100), .b(t2_010101), .y(t2_01010));
wire t2_010100, t2_010101;
mixer mix_t2_010100 (.a(t2_0101000), .b(t2_0101001), .y(t2_010100));
wire t2_0101000, t2_0101001;
mixer mix_t2_0101000 (.a(t2_01010000), .b(t2_01010001), .y(t2_0101000));
wire t2_01010000, t2_01010001;
mixer mix_t2_01010000 (.a(t2_010100000), .b(t2_010100001), .y(t2_01010000));
wire t2_010100000, t2_010100001;
mixer mix_t2_01010001 (.a(t2_010100010), .b(t2_010100011), .y(t2_01010001));
wire t2_010100010, t2_010100011;
mixer mix_t2_0101001 (.a(t2_01010010), .b(t2_01010011), .y(t2_0101001));
wire t2_01010010, t2_01010011;
mixer mix_t2_01010010 (.a(t2_010100100), .b(t2_010100101), .y(t2_01010010));
wire t2_010100100, t2_010100101;
mixer mix_t2_01010011 (.a(t2_010100110), .b(t2_010100111), .y(t2_01010011));
wire t2_010100110, t2_010100111;
mixer mix_t2_010101 (.a(t2_0101010), .b(t2_0101011), .y(t2_010101));
wire t2_0101010, t2_0101011;
mixer mix_t2_0101010 (.a(t2_01010100), .b(t2_01010101), .y(t2_0101010));
wire t2_01010100, t2_01010101;
mixer mix_t2_01010100 (.a(t2_010101000), .b(t2_010101001), .y(t2_01010100));
wire t2_010101000, t2_010101001;
mixer mix_t2_01010101 (.a(t2_010101010), .b(t2_010101011), .y(t2_01010101));
wire t2_010101010, t2_010101011;
mixer mix_t2_0101011 (.a(t2_01010110), .b(t2_01010111), .y(t2_0101011));
wire t2_01010110, t2_01010111;
mixer mix_t2_01010110 (.a(t2_010101100), .b(t2_010101101), .y(t2_01010110));
wire t2_010101100, t2_010101101;
mixer mix_t2_01010111 (.a(t2_010101110), .b(t2_010101111), .y(t2_01010111));
wire t2_010101110, t2_010101111;
mixer mix_t2_01011 (.a(t2_010110), .b(t2_010111), .y(t2_01011));
wire t2_010110, t2_010111;
mixer mix_t2_010110 (.a(t2_0101100), .b(t2_0101101), .y(t2_010110));
wire t2_0101100, t2_0101101;
mixer mix_t2_0101100 (.a(t2_01011000), .b(t2_01011001), .y(t2_0101100));
wire t2_01011000, t2_01011001;
mixer mix_t2_01011000 (.a(t2_010110000), .b(t2_010110001), .y(t2_01011000));
wire t2_010110000, t2_010110001;
mixer mix_t2_01011001 (.a(t2_010110010), .b(t2_010110011), .y(t2_01011001));
wire t2_010110010, t2_010110011;
mixer mix_t2_0101101 (.a(t2_01011010), .b(t2_01011011), .y(t2_0101101));
wire t2_01011010, t2_01011011;
mixer mix_t2_01011010 (.a(t2_010110100), .b(t2_010110101), .y(t2_01011010));
wire t2_010110100, t2_010110101;
mixer mix_t2_01011011 (.a(t2_010110110), .b(t2_010110111), .y(t2_01011011));
wire t2_010110110, t2_010110111;
mixer mix_t2_010111 (.a(t2_0101110), .b(t2_0101111), .y(t2_010111));
wire t2_0101110, t2_0101111;
mixer mix_t2_0101110 (.a(t2_01011100), .b(t2_01011101), .y(t2_0101110));
wire t2_01011100, t2_01011101;
mixer mix_t2_01011100 (.a(t2_010111000), .b(t2_010111001), .y(t2_01011100));
wire t2_010111000, t2_010111001;
mixer mix_t2_01011101 (.a(t2_010111010), .b(t2_010111011), .y(t2_01011101));
wire t2_010111010, t2_010111011;
mixer mix_t2_0101111 (.a(t2_01011110), .b(t2_01011111), .y(t2_0101111));
wire t2_01011110, t2_01011111;
mixer mix_t2_01011110 (.a(t2_010111100), .b(t2_010111101), .y(t2_01011110));
wire t2_010111100, t2_010111101;
mixer mix_t2_01011111 (.a(t2_010111110), .b(t2_010111111), .y(t2_01011111));
wire t2_010111110, t2_010111111;
mixer mix_t2_011 (.a(t2_0110), .b(t2_0111), .y(t2_011));
wire t2_0110, t2_0111;
mixer mix_t2_0110 (.a(t2_01100), .b(t2_01101), .y(t2_0110));
wire t2_01100, t2_01101;
mixer mix_t2_01100 (.a(t2_011000), .b(t2_011001), .y(t2_01100));
wire t2_011000, t2_011001;
mixer mix_t2_011000 (.a(t2_0110000), .b(t2_0110001), .y(t2_011000));
wire t2_0110000, t2_0110001;
mixer mix_t2_0110000 (.a(t2_01100000), .b(t2_01100001), .y(t2_0110000));
wire t2_01100000, t2_01100001;
mixer mix_t2_01100000 (.a(t2_011000000), .b(t2_011000001), .y(t2_01100000));
wire t2_011000000, t2_011000001;
mixer mix_t2_01100001 (.a(t2_011000010), .b(t2_011000011), .y(t2_01100001));
wire t2_011000010, t2_011000011;
mixer mix_t2_0110001 (.a(t2_01100010), .b(t2_01100011), .y(t2_0110001));
wire t2_01100010, t2_01100011;
mixer mix_t2_01100010 (.a(t2_011000100), .b(t2_011000101), .y(t2_01100010));
wire t2_011000100, t2_011000101;
mixer mix_t2_01100011 (.a(t2_011000110), .b(t2_011000111), .y(t2_01100011));
wire t2_011000110, t2_011000111;
mixer mix_t2_011001 (.a(t2_0110010), .b(t2_0110011), .y(t2_011001));
wire t2_0110010, t2_0110011;
mixer mix_t2_0110010 (.a(t2_01100100), .b(t2_01100101), .y(t2_0110010));
wire t2_01100100, t2_01100101;
mixer mix_t2_01100100 (.a(t2_011001000), .b(t2_011001001), .y(t2_01100100));
wire t2_011001000, t2_011001001;
mixer mix_t2_01100101 (.a(t2_011001010), .b(t2_011001011), .y(t2_01100101));
wire t2_011001010, t2_011001011;
mixer mix_t2_0110011 (.a(t2_01100110), .b(t2_01100111), .y(t2_0110011));
wire t2_01100110, t2_01100111;
mixer mix_t2_01100110 (.a(t2_011001100), .b(t2_011001101), .y(t2_01100110));
wire t2_011001100, t2_011001101;
mixer mix_t2_01100111 (.a(t2_011001110), .b(t2_011001111), .y(t2_01100111));
wire t2_011001110, t2_011001111;
mixer mix_t2_01101 (.a(t2_011010), .b(t2_011011), .y(t2_01101));
wire t2_011010, t2_011011;
mixer mix_t2_011010 (.a(t2_0110100), .b(t2_0110101), .y(t2_011010));
wire t2_0110100, t2_0110101;
mixer mix_t2_0110100 (.a(t2_01101000), .b(t2_01101001), .y(t2_0110100));
wire t2_01101000, t2_01101001;
mixer mix_t2_01101000 (.a(t2_011010000), .b(t2_011010001), .y(t2_01101000));
wire t2_011010000, t2_011010001;
mixer mix_t2_01101001 (.a(t2_011010010), .b(t2_011010011), .y(t2_01101001));
wire t2_011010010, t2_011010011;
mixer mix_t2_0110101 (.a(t2_01101010), .b(t2_01101011), .y(t2_0110101));
wire t2_01101010, t2_01101011;
mixer mix_t2_01101010 (.a(t2_011010100), .b(t2_011010101), .y(t2_01101010));
wire t2_011010100, t2_011010101;
mixer mix_t2_01101011 (.a(t2_011010110), .b(t2_011010111), .y(t2_01101011));
wire t2_011010110, t2_011010111;
mixer mix_t2_011011 (.a(t2_0110110), .b(t2_0110111), .y(t2_011011));
wire t2_0110110, t2_0110111;
mixer mix_t2_0110110 (.a(t2_01101100), .b(t2_01101101), .y(t2_0110110));
wire t2_01101100, t2_01101101;
mixer mix_t2_01101100 (.a(t2_011011000), .b(t2_011011001), .y(t2_01101100));
wire t2_011011000, t2_011011001;
mixer mix_t2_01101101 (.a(t2_011011010), .b(t2_011011011), .y(t2_01101101));
wire t2_011011010, t2_011011011;
mixer mix_t2_0110111 (.a(t2_01101110), .b(t2_01101111), .y(t2_0110111));
wire t2_01101110, t2_01101111;
mixer mix_t2_01101110 (.a(t2_011011100), .b(t2_011011101), .y(t2_01101110));
wire t2_011011100, t2_011011101;
mixer mix_t2_01101111 (.a(t2_011011110), .b(t2_011011111), .y(t2_01101111));
wire t2_011011110, t2_011011111;
mixer mix_t2_0111 (.a(t2_01110), .b(t2_01111), .y(t2_0111));
wire t2_01110, t2_01111;
mixer mix_t2_01110 (.a(t2_011100), .b(t2_011101), .y(t2_01110));
wire t2_011100, t2_011101;
mixer mix_t2_011100 (.a(t2_0111000), .b(t2_0111001), .y(t2_011100));
wire t2_0111000, t2_0111001;
mixer mix_t2_0111000 (.a(t2_01110000), .b(t2_01110001), .y(t2_0111000));
wire t2_01110000, t2_01110001;
mixer mix_t2_01110000 (.a(t2_011100000), .b(t2_011100001), .y(t2_01110000));
wire t2_011100000, t2_011100001;
mixer mix_t2_01110001 (.a(t2_011100010), .b(t2_011100011), .y(t2_01110001));
wire t2_011100010, t2_011100011;
mixer mix_t2_0111001 (.a(t2_01110010), .b(t2_01110011), .y(t2_0111001));
wire t2_01110010, t2_01110011;
mixer mix_t2_01110010 (.a(t2_011100100), .b(t2_011100101), .y(t2_01110010));
wire t2_011100100, t2_011100101;
mixer mix_t2_01110011 (.a(t2_011100110), .b(t2_011100111), .y(t2_01110011));
wire t2_011100110, t2_011100111;
mixer mix_t2_011101 (.a(t2_0111010), .b(t2_0111011), .y(t2_011101));
wire t2_0111010, t2_0111011;
mixer mix_t2_0111010 (.a(t2_01110100), .b(t2_01110101), .y(t2_0111010));
wire t2_01110100, t2_01110101;
mixer mix_t2_01110100 (.a(t2_011101000), .b(t2_011101001), .y(t2_01110100));
wire t2_011101000, t2_011101001;
mixer mix_t2_01110101 (.a(t2_011101010), .b(t2_011101011), .y(t2_01110101));
wire t2_011101010, t2_011101011;
mixer mix_t2_0111011 (.a(t2_01110110), .b(t2_01110111), .y(t2_0111011));
wire t2_01110110, t2_01110111;
mixer mix_t2_01110110 (.a(t2_011101100), .b(t2_011101101), .y(t2_01110110));
wire t2_011101100, t2_011101101;
mixer mix_t2_01110111 (.a(t2_011101110), .b(t2_011101111), .y(t2_01110111));
wire t2_011101110, t2_011101111;
mixer mix_t2_01111 (.a(t2_011110), .b(t2_011111), .y(t2_01111));
wire t2_011110, t2_011111;
mixer mix_t2_011110 (.a(t2_0111100), .b(t2_0111101), .y(t2_011110));
wire t2_0111100, t2_0111101;
mixer mix_t2_0111100 (.a(t2_01111000), .b(t2_01111001), .y(t2_0111100));
wire t2_01111000, t2_01111001;
mixer mix_t2_01111000 (.a(t2_011110000), .b(t2_011110001), .y(t2_01111000));
wire t2_011110000, t2_011110001;
mixer mix_t2_01111001 (.a(t2_011110010), .b(t2_011110011), .y(t2_01111001));
wire t2_011110010, t2_011110011;
mixer mix_t2_0111101 (.a(t2_01111010), .b(t2_01111011), .y(t2_0111101));
wire t2_01111010, t2_01111011;
mixer mix_t2_01111010 (.a(t2_011110100), .b(t2_011110101), .y(t2_01111010));
wire t2_011110100, t2_011110101;
mixer mix_t2_01111011 (.a(t2_011110110), .b(t2_011110111), .y(t2_01111011));
wire t2_011110110, t2_011110111;
mixer mix_t2_011111 (.a(t2_0111110), .b(t2_0111111), .y(t2_011111));
wire t2_0111110, t2_0111111;
mixer mix_t2_0111110 (.a(t2_01111100), .b(t2_01111101), .y(t2_0111110));
wire t2_01111100, t2_01111101;
mixer mix_t2_01111100 (.a(t2_011111000), .b(t2_011111001), .y(t2_01111100));
wire t2_011111000, t2_011111001;
mixer mix_t2_01111101 (.a(t2_011111010), .b(t2_011111011), .y(t2_01111101));
wire t2_011111010, t2_011111011;
mixer mix_t2_0111111 (.a(t2_01111110), .b(t2_01111111), .y(t2_0111111));
wire t2_01111110, t2_01111111;
mixer mix_t2_01111110 (.a(t2_011111100), .b(t2_011111101), .y(t2_01111110));
wire t2_011111100, t2_011111101;
mixer mix_t2_01111111 (.a(t2_011111110), .b(t2_011111111), .y(t2_01111111));
wire t2_011111110, t2_011111111;
mixer mix_t3_0 (.a(t3_00), .b(t3_01), .y(t3_0));
wire t3_00, t3_01;
mixer mix_t3_00 (.a(t3_000), .b(t3_001), .y(t3_00));
wire t3_000, t3_001;
mixer mix_t3_000 (.a(t3_0000), .b(t3_0001), .y(t3_000));
wire t3_0000, t3_0001;
mixer mix_t3_0000 (.a(t3_00000), .b(t3_00001), .y(t3_0000));
wire t3_00000, t3_00001;
mixer mix_t3_00000 (.a(t3_000000), .b(t3_000001), .y(t3_00000));
wire t3_000000, t3_000001;
mixer mix_t3_000000 (.a(t3_0000000), .b(t3_0000001), .y(t3_000000));
wire t3_0000000, t3_0000001;
mixer mix_t3_0000000 (.a(t3_00000000), .b(t3_00000001), .y(t3_0000000));
wire t3_00000000, t3_00000001;
mixer mix_t3_00000000 (.a(t3_000000000), .b(t3_000000001), .y(t3_00000000));
wire t3_000000000, t3_000000001;
mixer mix_t3_00000001 (.a(t3_000000010), .b(t3_000000011), .y(t3_00000001));
wire t3_000000010, t3_000000011;
mixer mix_t3_0000001 (.a(t3_00000010), .b(t3_00000011), .y(t3_0000001));
wire t3_00000010, t3_00000011;
mixer mix_t3_00000010 (.a(t3_000000100), .b(t3_000000101), .y(t3_00000010));
wire t3_000000100, t3_000000101;
mixer mix_t3_00000011 (.a(t3_000000110), .b(t3_000000111), .y(t3_00000011));
wire t3_000000110, t3_000000111;
mixer mix_t3_000001 (.a(t3_0000010), .b(t3_0000011), .y(t3_000001));
wire t3_0000010, t3_0000011;
mixer mix_t3_0000010 (.a(t3_00000100), .b(t3_00000101), .y(t3_0000010));
wire t3_00000100, t3_00000101;
mixer mix_t3_00000100 (.a(t3_000001000), .b(t3_000001001), .y(t3_00000100));
wire t3_000001000, t3_000001001;
mixer mix_t3_00000101 (.a(t3_000001010), .b(t3_000001011), .y(t3_00000101));
wire t3_000001010, t3_000001011;
mixer mix_t3_0000011 (.a(t3_00000110), .b(t3_00000111), .y(t3_0000011));
wire t3_00000110, t3_00000111;
mixer mix_t3_00000110 (.a(t3_000001100), .b(t3_000001101), .y(t3_00000110));
wire t3_000001100, t3_000001101;
mixer mix_t3_00000111 (.a(t3_000001110), .b(t3_000001111), .y(t3_00000111));
wire t3_000001110, t3_000001111;
mixer mix_t3_00001 (.a(t3_000010), .b(t3_000011), .y(t3_00001));
wire t3_000010, t3_000011;
mixer mix_t3_000010 (.a(t3_0000100), .b(t3_0000101), .y(t3_000010));
wire t3_0000100, t3_0000101;
mixer mix_t3_0000100 (.a(t3_00001000), .b(t3_00001001), .y(t3_0000100));
wire t3_00001000, t3_00001001;
mixer mix_t3_00001000 (.a(t3_000010000), .b(t3_000010001), .y(t3_00001000));
wire t3_000010000, t3_000010001;
mixer mix_t3_00001001 (.a(t3_000010010), .b(t3_000010011), .y(t3_00001001));
wire t3_000010010, t3_000010011;
mixer mix_t3_0000101 (.a(t3_00001010), .b(t3_00001011), .y(t3_0000101));
wire t3_00001010, t3_00001011;
mixer mix_t3_00001010 (.a(t3_000010100), .b(t3_000010101), .y(t3_00001010));
wire t3_000010100, t3_000010101;
mixer mix_t3_00001011 (.a(t3_000010110), .b(t3_000010111), .y(t3_00001011));
wire t3_000010110, t3_000010111;
mixer mix_t3_000011 (.a(t3_0000110), .b(t3_0000111), .y(t3_000011));
wire t3_0000110, t3_0000111;
mixer mix_t3_0000110 (.a(t3_00001100), .b(t3_00001101), .y(t3_0000110));
wire t3_00001100, t3_00001101;
mixer mix_t3_00001100 (.a(t3_000011000), .b(t3_000011001), .y(t3_00001100));
wire t3_000011000, t3_000011001;
mixer mix_t3_00001101 (.a(t3_000011010), .b(t3_000011011), .y(t3_00001101));
wire t3_000011010, t3_000011011;
mixer mix_t3_0000111 (.a(t3_00001110), .b(t3_00001111), .y(t3_0000111));
wire t3_00001110, t3_00001111;
mixer mix_t3_00001110 (.a(t3_000011100), .b(t3_000011101), .y(t3_00001110));
wire t3_000011100, t3_000011101;
mixer mix_t3_00001111 (.a(t3_000011110), .b(t3_000011111), .y(t3_00001111));
wire t3_000011110, t3_000011111;
mixer mix_t3_0001 (.a(t3_00010), .b(t3_00011), .y(t3_0001));
wire t3_00010, t3_00011;
mixer mix_t3_00010 (.a(t3_000100), .b(t3_000101), .y(t3_00010));
wire t3_000100, t3_000101;
mixer mix_t3_000100 (.a(t3_0001000), .b(t3_0001001), .y(t3_000100));
wire t3_0001000, t3_0001001;
mixer mix_t3_0001000 (.a(t3_00010000), .b(t3_00010001), .y(t3_0001000));
wire t3_00010000, t3_00010001;
mixer mix_t3_00010000 (.a(t3_000100000), .b(t3_000100001), .y(t3_00010000));
wire t3_000100000, t3_000100001;
mixer mix_t3_00010001 (.a(t3_000100010), .b(t3_000100011), .y(t3_00010001));
wire t3_000100010, t3_000100011;
mixer mix_t3_0001001 (.a(t3_00010010), .b(t3_00010011), .y(t3_0001001));
wire t3_00010010, t3_00010011;
mixer mix_t3_00010010 (.a(t3_000100100), .b(t3_000100101), .y(t3_00010010));
wire t3_000100100, t3_000100101;
mixer mix_t3_00010011 (.a(t3_000100110), .b(t3_000100111), .y(t3_00010011));
wire t3_000100110, t3_000100111;
mixer mix_t3_000101 (.a(t3_0001010), .b(t3_0001011), .y(t3_000101));
wire t3_0001010, t3_0001011;
mixer mix_t3_0001010 (.a(t3_00010100), .b(t3_00010101), .y(t3_0001010));
wire t3_00010100, t3_00010101;
mixer mix_t3_00010100 (.a(t3_000101000), .b(t3_000101001), .y(t3_00010100));
wire t3_000101000, t3_000101001;
mixer mix_t3_00010101 (.a(t3_000101010), .b(t3_000101011), .y(t3_00010101));
wire t3_000101010, t3_000101011;
mixer mix_t3_0001011 (.a(t3_00010110), .b(t3_00010111), .y(t3_0001011));
wire t3_00010110, t3_00010111;
mixer mix_t3_00010110 (.a(t3_000101100), .b(t3_000101101), .y(t3_00010110));
wire t3_000101100, t3_000101101;
mixer mix_t3_00010111 (.a(t3_000101110), .b(t3_000101111), .y(t3_00010111));
wire t3_000101110, t3_000101111;
mixer mix_t3_00011 (.a(t3_000110), .b(t3_000111), .y(t3_00011));
wire t3_000110, t3_000111;
mixer mix_t3_000110 (.a(t3_0001100), .b(t3_0001101), .y(t3_000110));
wire t3_0001100, t3_0001101;
mixer mix_t3_0001100 (.a(t3_00011000), .b(t3_00011001), .y(t3_0001100));
wire t3_00011000, t3_00011001;
mixer mix_t3_00011000 (.a(t3_000110000), .b(t3_000110001), .y(t3_00011000));
wire t3_000110000, t3_000110001;
mixer mix_t3_00011001 (.a(t3_000110010), .b(t3_000110011), .y(t3_00011001));
wire t3_000110010, t3_000110011;
mixer mix_t3_0001101 (.a(t3_00011010), .b(t3_00011011), .y(t3_0001101));
wire t3_00011010, t3_00011011;
mixer mix_t3_00011010 (.a(t3_000110100), .b(t3_000110101), .y(t3_00011010));
wire t3_000110100, t3_000110101;
mixer mix_t3_00011011 (.a(t3_000110110), .b(t3_000110111), .y(t3_00011011));
wire t3_000110110, t3_000110111;
mixer mix_t3_000111 (.a(t3_0001110), .b(t3_0001111), .y(t3_000111));
wire t3_0001110, t3_0001111;
mixer mix_t3_0001110 (.a(t3_00011100), .b(t3_00011101), .y(t3_0001110));
wire t3_00011100, t3_00011101;
mixer mix_t3_00011100 (.a(t3_000111000), .b(t3_000111001), .y(t3_00011100));
wire t3_000111000, t3_000111001;
mixer mix_t3_00011101 (.a(t3_000111010), .b(t3_000111011), .y(t3_00011101));
wire t3_000111010, t3_000111011;
mixer mix_t3_0001111 (.a(t3_00011110), .b(t3_00011111), .y(t3_0001111));
wire t3_00011110, t3_00011111;
mixer mix_t3_00011110 (.a(t3_000111100), .b(t3_000111101), .y(t3_00011110));
wire t3_000111100, t3_000111101;
mixer mix_t3_00011111 (.a(t3_000111110), .b(t3_000111111), .y(t3_00011111));
wire t3_000111110, t3_000111111;
mixer mix_t3_001 (.a(t3_0010), .b(t3_0011), .y(t3_001));
wire t3_0010, t3_0011;
mixer mix_t3_0010 (.a(t3_00100), .b(t3_00101), .y(t3_0010));
wire t3_00100, t3_00101;
mixer mix_t3_00100 (.a(t3_001000), .b(t3_001001), .y(t3_00100));
wire t3_001000, t3_001001;
mixer mix_t3_001000 (.a(t3_0010000), .b(t3_0010001), .y(t3_001000));
wire t3_0010000, t3_0010001;
mixer mix_t3_0010000 (.a(t3_00100000), .b(t3_00100001), .y(t3_0010000));
wire t3_00100000, t3_00100001;
mixer mix_t3_00100000 (.a(t3_001000000), .b(t3_001000001), .y(t3_00100000));
wire t3_001000000, t3_001000001;
mixer mix_t3_00100001 (.a(t3_001000010), .b(t3_001000011), .y(t3_00100001));
wire t3_001000010, t3_001000011;
mixer mix_t3_0010001 (.a(t3_00100010), .b(t3_00100011), .y(t3_0010001));
wire t3_00100010, t3_00100011;
mixer mix_t3_00100010 (.a(t3_001000100), .b(t3_001000101), .y(t3_00100010));
wire t3_001000100, t3_001000101;
mixer mix_t3_00100011 (.a(t3_001000110), .b(t3_001000111), .y(t3_00100011));
wire t3_001000110, t3_001000111;
mixer mix_t3_001001 (.a(t3_0010010), .b(t3_0010011), .y(t3_001001));
wire t3_0010010, t3_0010011;
mixer mix_t3_0010010 (.a(t3_00100100), .b(t3_00100101), .y(t3_0010010));
wire t3_00100100, t3_00100101;
mixer mix_t3_00100100 (.a(t3_001001000), .b(t3_001001001), .y(t3_00100100));
wire t3_001001000, t3_001001001;
mixer mix_t3_00100101 (.a(t3_001001010), .b(t3_001001011), .y(t3_00100101));
wire t3_001001010, t3_001001011;
mixer mix_t3_0010011 (.a(t3_00100110), .b(t3_00100111), .y(t3_0010011));
wire t3_00100110, t3_00100111;
mixer mix_t3_00100110 (.a(t3_001001100), .b(t3_001001101), .y(t3_00100110));
wire t3_001001100, t3_001001101;
mixer mix_t3_00100111 (.a(t3_001001110), .b(t3_001001111), .y(t3_00100111));
wire t3_001001110, t3_001001111;
mixer mix_t3_00101 (.a(t3_001010), .b(t3_001011), .y(t3_00101));
wire t3_001010, t3_001011;
mixer mix_t3_001010 (.a(t3_0010100), .b(t3_0010101), .y(t3_001010));
wire t3_0010100, t3_0010101;
mixer mix_t3_0010100 (.a(t3_00101000), .b(t3_00101001), .y(t3_0010100));
wire t3_00101000, t3_00101001;
mixer mix_t3_00101000 (.a(t3_001010000), .b(t3_001010001), .y(t3_00101000));
wire t3_001010000, t3_001010001;
mixer mix_t3_00101001 (.a(t3_001010010), .b(t3_001010011), .y(t3_00101001));
wire t3_001010010, t3_001010011;
mixer mix_t3_0010101 (.a(t3_00101010), .b(t3_00101011), .y(t3_0010101));
wire t3_00101010, t3_00101011;
mixer mix_t3_00101010 (.a(t3_001010100), .b(t3_001010101), .y(t3_00101010));
wire t3_001010100, t3_001010101;
mixer mix_t3_00101011 (.a(t3_001010110), .b(t3_001010111), .y(t3_00101011));
wire t3_001010110, t3_001010111;
mixer mix_t3_001011 (.a(t3_0010110), .b(t3_0010111), .y(t3_001011));
wire t3_0010110, t3_0010111;
mixer mix_t3_0010110 (.a(t3_00101100), .b(t3_00101101), .y(t3_0010110));
wire t3_00101100, t3_00101101;
mixer mix_t3_00101100 (.a(t3_001011000), .b(t3_001011001), .y(t3_00101100));
wire t3_001011000, t3_001011001;
mixer mix_t3_00101101 (.a(t3_001011010), .b(t3_001011011), .y(t3_00101101));
wire t3_001011010, t3_001011011;
mixer mix_t3_0010111 (.a(t3_00101110), .b(t3_00101111), .y(t3_0010111));
wire t3_00101110, t3_00101111;
mixer mix_t3_00101110 (.a(t3_001011100), .b(t3_001011101), .y(t3_00101110));
wire t3_001011100, t3_001011101;
mixer mix_t3_00101111 (.a(t3_001011110), .b(t3_001011111), .y(t3_00101111));
wire t3_001011110, t3_001011111;
mixer mix_t3_0011 (.a(t3_00110), .b(t3_00111), .y(t3_0011));
wire t3_00110, t3_00111;
mixer mix_t3_00110 (.a(t3_001100), .b(t3_001101), .y(t3_00110));
wire t3_001100, t3_001101;
mixer mix_t3_001100 (.a(t3_0011000), .b(t3_0011001), .y(t3_001100));
wire t3_0011000, t3_0011001;
mixer mix_t3_0011000 (.a(t3_00110000), .b(t3_00110001), .y(t3_0011000));
wire t3_00110000, t3_00110001;
mixer mix_t3_00110000 (.a(t3_001100000), .b(t3_001100001), .y(t3_00110000));
wire t3_001100000, t3_001100001;
mixer mix_t3_00110001 (.a(t3_001100010), .b(t3_001100011), .y(t3_00110001));
wire t3_001100010, t3_001100011;
mixer mix_t3_0011001 (.a(t3_00110010), .b(t3_00110011), .y(t3_0011001));
wire t3_00110010, t3_00110011;
mixer mix_t3_00110010 (.a(t3_001100100), .b(t3_001100101), .y(t3_00110010));
wire t3_001100100, t3_001100101;
mixer mix_t3_00110011 (.a(t3_001100110), .b(t3_001100111), .y(t3_00110011));
wire t3_001100110, t3_001100111;
mixer mix_t3_001101 (.a(t3_0011010), .b(t3_0011011), .y(t3_001101));
wire t3_0011010, t3_0011011;
mixer mix_t3_0011010 (.a(t3_00110100), .b(t3_00110101), .y(t3_0011010));
wire t3_00110100, t3_00110101;
mixer mix_t3_00110100 (.a(t3_001101000), .b(t3_001101001), .y(t3_00110100));
wire t3_001101000, t3_001101001;
mixer mix_t3_00110101 (.a(t3_001101010), .b(t3_001101011), .y(t3_00110101));
wire t3_001101010, t3_001101011;
mixer mix_t3_0011011 (.a(t3_00110110), .b(t3_00110111), .y(t3_0011011));
wire t3_00110110, t3_00110111;
mixer mix_t3_00110110 (.a(t3_001101100), .b(t3_001101101), .y(t3_00110110));
wire t3_001101100, t3_001101101;
mixer mix_t3_00110111 (.a(t3_001101110), .b(t3_001101111), .y(t3_00110111));
wire t3_001101110, t3_001101111;
mixer mix_t3_00111 (.a(t3_001110), .b(t3_001111), .y(t3_00111));
wire t3_001110, t3_001111;
mixer mix_t3_001110 (.a(t3_0011100), .b(t3_0011101), .y(t3_001110));
wire t3_0011100, t3_0011101;
mixer mix_t3_0011100 (.a(t3_00111000), .b(t3_00111001), .y(t3_0011100));
wire t3_00111000, t3_00111001;
mixer mix_t3_00111000 (.a(t3_001110000), .b(t3_001110001), .y(t3_00111000));
wire t3_001110000, t3_001110001;
mixer mix_t3_00111001 (.a(t3_001110010), .b(t3_001110011), .y(t3_00111001));
wire t3_001110010, t3_001110011;
mixer mix_t3_0011101 (.a(t3_00111010), .b(t3_00111011), .y(t3_0011101));
wire t3_00111010, t3_00111011;
mixer mix_t3_00111010 (.a(t3_001110100), .b(t3_001110101), .y(t3_00111010));
wire t3_001110100, t3_001110101;
mixer mix_t3_00111011 (.a(t3_001110110), .b(t3_001110111), .y(t3_00111011));
wire t3_001110110, t3_001110111;
mixer mix_t3_001111 (.a(t3_0011110), .b(t3_0011111), .y(t3_001111));
wire t3_0011110, t3_0011111;
mixer mix_t3_0011110 (.a(t3_00111100), .b(t3_00111101), .y(t3_0011110));
wire t3_00111100, t3_00111101;
mixer mix_t3_00111100 (.a(t3_001111000), .b(t3_001111001), .y(t3_00111100));
wire t3_001111000, t3_001111001;
mixer mix_t3_00111101 (.a(t3_001111010), .b(t3_001111011), .y(t3_00111101));
wire t3_001111010, t3_001111011;
mixer mix_t3_0011111 (.a(t3_00111110), .b(t3_00111111), .y(t3_0011111));
wire t3_00111110, t3_00111111;
mixer mix_t3_00111110 (.a(t3_001111100), .b(t3_001111101), .y(t3_00111110));
wire t3_001111100, t3_001111101;
mixer mix_t3_00111111 (.a(t3_001111110), .b(t3_001111111), .y(t3_00111111));
wire t3_001111110, t3_001111111;
mixer mix_t3_01 (.a(t3_010), .b(t3_011), .y(t3_01));
wire t3_010, t3_011;
mixer mix_t3_010 (.a(t3_0100), .b(t3_0101), .y(t3_010));
wire t3_0100, t3_0101;
mixer mix_t3_0100 (.a(t3_01000), .b(t3_01001), .y(t3_0100));
wire t3_01000, t3_01001;
mixer mix_t3_01000 (.a(t3_010000), .b(t3_010001), .y(t3_01000));
wire t3_010000, t3_010001;
mixer mix_t3_010000 (.a(t3_0100000), .b(t3_0100001), .y(t3_010000));
wire t3_0100000, t3_0100001;
mixer mix_t3_0100000 (.a(t3_01000000), .b(t3_01000001), .y(t3_0100000));
wire t3_01000000, t3_01000001;
mixer mix_t3_01000000 (.a(t3_010000000), .b(t3_010000001), .y(t3_01000000));
wire t3_010000000, t3_010000001;
mixer mix_t3_01000001 (.a(t3_010000010), .b(t3_010000011), .y(t3_01000001));
wire t3_010000010, t3_010000011;
mixer mix_t3_0100001 (.a(t3_01000010), .b(t3_01000011), .y(t3_0100001));
wire t3_01000010, t3_01000011;
mixer mix_t3_01000010 (.a(t3_010000100), .b(t3_010000101), .y(t3_01000010));
wire t3_010000100, t3_010000101;
mixer mix_t3_01000011 (.a(t3_010000110), .b(t3_010000111), .y(t3_01000011));
wire t3_010000110, t3_010000111;
mixer mix_t3_010001 (.a(t3_0100010), .b(t3_0100011), .y(t3_010001));
wire t3_0100010, t3_0100011;
mixer mix_t3_0100010 (.a(t3_01000100), .b(t3_01000101), .y(t3_0100010));
wire t3_01000100, t3_01000101;
mixer mix_t3_01000100 (.a(t3_010001000), .b(t3_010001001), .y(t3_01000100));
wire t3_010001000, t3_010001001;
mixer mix_t3_01000101 (.a(t3_010001010), .b(t3_010001011), .y(t3_01000101));
wire t3_010001010, t3_010001011;
mixer mix_t3_0100011 (.a(t3_01000110), .b(t3_01000111), .y(t3_0100011));
wire t3_01000110, t3_01000111;
mixer mix_t3_01000110 (.a(t3_010001100), .b(t3_010001101), .y(t3_01000110));
wire t3_010001100, t3_010001101;
mixer mix_t3_01000111 (.a(t3_010001110), .b(t3_010001111), .y(t3_01000111));
wire t3_010001110, t3_010001111;
mixer mix_t3_01001 (.a(t3_010010), .b(t3_010011), .y(t3_01001));
wire t3_010010, t3_010011;
mixer mix_t3_010010 (.a(t3_0100100), .b(t3_0100101), .y(t3_010010));
wire t3_0100100, t3_0100101;
mixer mix_t3_0100100 (.a(t3_01001000), .b(t3_01001001), .y(t3_0100100));
wire t3_01001000, t3_01001001;
mixer mix_t3_01001000 (.a(t3_010010000), .b(t3_010010001), .y(t3_01001000));
wire t3_010010000, t3_010010001;
mixer mix_t3_01001001 (.a(t3_010010010), .b(t3_010010011), .y(t3_01001001));
wire t3_010010010, t3_010010011;
mixer mix_t3_0100101 (.a(t3_01001010), .b(t3_01001011), .y(t3_0100101));
wire t3_01001010, t3_01001011;
mixer mix_t3_01001010 (.a(t3_010010100), .b(t3_010010101), .y(t3_01001010));
wire t3_010010100, t3_010010101;
mixer mix_t3_01001011 (.a(t3_010010110), .b(t3_010010111), .y(t3_01001011));
wire t3_010010110, t3_010010111;
mixer mix_t3_010011 (.a(t3_0100110), .b(t3_0100111), .y(t3_010011));
wire t3_0100110, t3_0100111;
mixer mix_t3_0100110 (.a(t3_01001100), .b(t3_01001101), .y(t3_0100110));
wire t3_01001100, t3_01001101;
mixer mix_t3_01001100 (.a(t3_010011000), .b(t3_010011001), .y(t3_01001100));
wire t3_010011000, t3_010011001;
mixer mix_t3_01001101 (.a(t3_010011010), .b(t3_010011011), .y(t3_01001101));
wire t3_010011010, t3_010011011;
mixer mix_t3_0100111 (.a(t3_01001110), .b(t3_01001111), .y(t3_0100111));
wire t3_01001110, t3_01001111;
mixer mix_t3_01001110 (.a(t3_010011100), .b(t3_010011101), .y(t3_01001110));
wire t3_010011100, t3_010011101;
mixer mix_t3_01001111 (.a(t3_010011110), .b(t3_010011111), .y(t3_01001111));
wire t3_010011110, t3_010011111;
mixer mix_t3_0101 (.a(t3_01010), .b(t3_01011), .y(t3_0101));
wire t3_01010, t3_01011;
mixer mix_t3_01010 (.a(t3_010100), .b(t3_010101), .y(t3_01010));
wire t3_010100, t3_010101;
mixer mix_t3_010100 (.a(t3_0101000), .b(t3_0101001), .y(t3_010100));
wire t3_0101000, t3_0101001;
mixer mix_t3_0101000 (.a(t3_01010000), .b(t3_01010001), .y(t3_0101000));
wire t3_01010000, t3_01010001;
mixer mix_t3_01010000 (.a(t3_010100000), .b(t3_010100001), .y(t3_01010000));
wire t3_010100000, t3_010100001;
mixer mix_t3_01010001 (.a(t3_010100010), .b(t3_010100011), .y(t3_01010001));
wire t3_010100010, t3_010100011;
mixer mix_t3_0101001 (.a(t3_01010010), .b(t3_01010011), .y(t3_0101001));
wire t3_01010010, t3_01010011;
mixer mix_t3_01010010 (.a(t3_010100100), .b(t3_010100101), .y(t3_01010010));
wire t3_010100100, t3_010100101;
mixer mix_t3_01010011 (.a(t3_010100110), .b(t3_010100111), .y(t3_01010011));
wire t3_010100110, t3_010100111;
mixer mix_t3_010101 (.a(t3_0101010), .b(t3_0101011), .y(t3_010101));
wire t3_0101010, t3_0101011;
mixer mix_t3_0101010 (.a(t3_01010100), .b(t3_01010101), .y(t3_0101010));
wire t3_01010100, t3_01010101;
mixer mix_t3_01010100 (.a(t3_010101000), .b(t3_010101001), .y(t3_01010100));
wire t3_010101000, t3_010101001;
mixer mix_t3_01010101 (.a(t3_010101010), .b(t3_010101011), .y(t3_01010101));
wire t3_010101010, t3_010101011;
mixer mix_t3_0101011 (.a(t3_01010110), .b(t3_01010111), .y(t3_0101011));
wire t3_01010110, t3_01010111;
mixer mix_t3_01010110 (.a(t3_010101100), .b(t3_010101101), .y(t3_01010110));
wire t3_010101100, t3_010101101;
mixer mix_t3_01010111 (.a(t3_010101110), .b(t3_010101111), .y(t3_01010111));
wire t3_010101110, t3_010101111;
mixer mix_t3_01011 (.a(t3_010110), .b(t3_010111), .y(t3_01011));
wire t3_010110, t3_010111;
mixer mix_t3_010110 (.a(t3_0101100), .b(t3_0101101), .y(t3_010110));
wire t3_0101100, t3_0101101;
mixer mix_t3_0101100 (.a(t3_01011000), .b(t3_01011001), .y(t3_0101100));
wire t3_01011000, t3_01011001;
mixer mix_t3_01011000 (.a(t3_010110000), .b(t3_010110001), .y(t3_01011000));
wire t3_010110000, t3_010110001;
mixer mix_t3_01011001 (.a(t3_010110010), .b(t3_010110011), .y(t3_01011001));
wire t3_010110010, t3_010110011;
mixer mix_t3_0101101 (.a(t3_01011010), .b(t3_01011011), .y(t3_0101101));
wire t3_01011010, t3_01011011;
mixer mix_t3_01011010 (.a(t3_010110100), .b(t3_010110101), .y(t3_01011010));
wire t3_010110100, t3_010110101;
mixer mix_t3_01011011 (.a(t3_010110110), .b(t3_010110111), .y(t3_01011011));
wire t3_010110110, t3_010110111;
mixer mix_t3_010111 (.a(t3_0101110), .b(t3_0101111), .y(t3_010111));
wire t3_0101110, t3_0101111;
mixer mix_t3_0101110 (.a(t3_01011100), .b(t3_01011101), .y(t3_0101110));
wire t3_01011100, t3_01011101;
mixer mix_t3_01011100 (.a(t3_010111000), .b(t3_010111001), .y(t3_01011100));
wire t3_010111000, t3_010111001;
mixer mix_t3_01011101 (.a(t3_010111010), .b(t3_010111011), .y(t3_01011101));
wire t3_010111010, t3_010111011;
mixer mix_t3_0101111 (.a(t3_01011110), .b(t3_01011111), .y(t3_0101111));
wire t3_01011110, t3_01011111;
mixer mix_t3_01011110 (.a(t3_010111100), .b(t3_010111101), .y(t3_01011110));
wire t3_010111100, t3_010111101;
mixer mix_t3_01011111 (.a(t3_010111110), .b(t3_010111111), .y(t3_01011111));
wire t3_010111110, t3_010111111;
mixer mix_t3_011 (.a(t3_0110), .b(t3_0111), .y(t3_011));
wire t3_0110, t3_0111;
mixer mix_t3_0110 (.a(t3_01100), .b(t3_01101), .y(t3_0110));
wire t3_01100, t3_01101;
mixer mix_t3_01100 (.a(t3_011000), .b(t3_011001), .y(t3_01100));
wire t3_011000, t3_011001;
mixer mix_t3_011000 (.a(t3_0110000), .b(t3_0110001), .y(t3_011000));
wire t3_0110000, t3_0110001;
mixer mix_t3_0110000 (.a(t3_01100000), .b(t3_01100001), .y(t3_0110000));
wire t3_01100000, t3_01100001;
mixer mix_t3_01100000 (.a(t3_011000000), .b(t3_011000001), .y(t3_01100000));
wire t3_011000000, t3_011000001;
mixer mix_t3_01100001 (.a(t3_011000010), .b(t3_011000011), .y(t3_01100001));
wire t3_011000010, t3_011000011;
mixer mix_t3_0110001 (.a(t3_01100010), .b(t3_01100011), .y(t3_0110001));
wire t3_01100010, t3_01100011;
mixer mix_t3_01100010 (.a(t3_011000100), .b(t3_011000101), .y(t3_01100010));
wire t3_011000100, t3_011000101;
mixer mix_t3_01100011 (.a(t3_011000110), .b(t3_011000111), .y(t3_01100011));
wire t3_011000110, t3_011000111;
mixer mix_t3_011001 (.a(t3_0110010), .b(t3_0110011), .y(t3_011001));
wire t3_0110010, t3_0110011;
mixer mix_t3_0110010 (.a(t3_01100100), .b(t3_01100101), .y(t3_0110010));
wire t3_01100100, t3_01100101;
mixer mix_t3_01100100 (.a(t3_011001000), .b(t3_011001001), .y(t3_01100100));
wire t3_011001000, t3_011001001;
mixer mix_t3_01100101 (.a(t3_011001010), .b(t3_011001011), .y(t3_01100101));
wire t3_011001010, t3_011001011;
mixer mix_t3_0110011 (.a(t3_01100110), .b(t3_01100111), .y(t3_0110011));
wire t3_01100110, t3_01100111;
mixer mix_t3_01100110 (.a(t3_011001100), .b(t3_011001101), .y(t3_01100110));
wire t3_011001100, t3_011001101;
mixer mix_t3_01100111 (.a(t3_011001110), .b(t3_011001111), .y(t3_01100111));
wire t3_011001110, t3_011001111;
mixer mix_t3_01101 (.a(t3_011010), .b(t3_011011), .y(t3_01101));
wire t3_011010, t3_011011;
mixer mix_t3_011010 (.a(t3_0110100), .b(t3_0110101), .y(t3_011010));
wire t3_0110100, t3_0110101;
mixer mix_t3_0110100 (.a(t3_01101000), .b(t3_01101001), .y(t3_0110100));
wire t3_01101000, t3_01101001;
mixer mix_t3_01101000 (.a(t3_011010000), .b(t3_011010001), .y(t3_01101000));
wire t3_011010000, t3_011010001;
mixer mix_t3_01101001 (.a(t3_011010010), .b(t3_011010011), .y(t3_01101001));
wire t3_011010010, t3_011010011;
mixer mix_t3_0110101 (.a(t3_01101010), .b(t3_01101011), .y(t3_0110101));
wire t3_01101010, t3_01101011;
mixer mix_t3_01101010 (.a(t3_011010100), .b(t3_011010101), .y(t3_01101010));
wire t3_011010100, t3_011010101;
mixer mix_t3_01101011 (.a(t3_011010110), .b(t3_011010111), .y(t3_01101011));
wire t3_011010110, t3_011010111;
mixer mix_t3_011011 (.a(t3_0110110), .b(t3_0110111), .y(t3_011011));
wire t3_0110110, t3_0110111;
mixer mix_t3_0110110 (.a(t3_01101100), .b(t3_01101101), .y(t3_0110110));
wire t3_01101100, t3_01101101;
mixer mix_t3_01101100 (.a(t3_011011000), .b(t3_011011001), .y(t3_01101100));
wire t3_011011000, t3_011011001;
mixer mix_t3_01101101 (.a(t3_011011010), .b(t3_011011011), .y(t3_01101101));
wire t3_011011010, t3_011011011;
mixer mix_t3_0110111 (.a(t3_01101110), .b(t3_01101111), .y(t3_0110111));
wire t3_01101110, t3_01101111;
mixer mix_t3_01101110 (.a(t3_011011100), .b(t3_011011101), .y(t3_01101110));
wire t3_011011100, t3_011011101;
mixer mix_t3_01101111 (.a(t3_011011110), .b(t3_011011111), .y(t3_01101111));
wire t3_011011110, t3_011011111;
mixer mix_t3_0111 (.a(t3_01110), .b(t3_01111), .y(t3_0111));
wire t3_01110, t3_01111;
mixer mix_t3_01110 (.a(t3_011100), .b(t3_011101), .y(t3_01110));
wire t3_011100, t3_011101;
mixer mix_t3_011100 (.a(t3_0111000), .b(t3_0111001), .y(t3_011100));
wire t3_0111000, t3_0111001;
mixer mix_t3_0111000 (.a(t3_01110000), .b(t3_01110001), .y(t3_0111000));
wire t3_01110000, t3_01110001;
mixer mix_t3_01110000 (.a(t3_011100000), .b(t3_011100001), .y(t3_01110000));
wire t3_011100000, t3_011100001;
mixer mix_t3_01110001 (.a(t3_011100010), .b(t3_011100011), .y(t3_01110001));
wire t3_011100010, t3_011100011;
mixer mix_t3_0111001 (.a(t3_01110010), .b(t3_01110011), .y(t3_0111001));
wire t3_01110010, t3_01110011;
mixer mix_t3_01110010 (.a(t3_011100100), .b(t3_011100101), .y(t3_01110010));
wire t3_011100100, t3_011100101;
mixer mix_t3_01110011 (.a(t3_011100110), .b(t3_011100111), .y(t3_01110011));
wire t3_011100110, t3_011100111;
mixer mix_t3_011101 (.a(t3_0111010), .b(t3_0111011), .y(t3_011101));
wire t3_0111010, t3_0111011;
mixer mix_t3_0111010 (.a(t3_01110100), .b(t3_01110101), .y(t3_0111010));
wire t3_01110100, t3_01110101;
mixer mix_t3_01110100 (.a(t3_011101000), .b(t3_011101001), .y(t3_01110100));
wire t3_011101000, t3_011101001;
mixer mix_t3_01110101 (.a(t3_011101010), .b(t3_011101011), .y(t3_01110101));
wire t3_011101010, t3_011101011;
mixer mix_t3_0111011 (.a(t3_01110110), .b(t3_01110111), .y(t3_0111011));
wire t3_01110110, t3_01110111;
mixer mix_t3_01110110 (.a(t3_011101100), .b(t3_011101101), .y(t3_01110110));
wire t3_011101100, t3_011101101;
mixer mix_t3_01110111 (.a(t3_011101110), .b(t3_011101111), .y(t3_01110111));
wire t3_011101110, t3_011101111;
mixer mix_t3_01111 (.a(t3_011110), .b(t3_011111), .y(t3_01111));
wire t3_011110, t3_011111;
mixer mix_t3_011110 (.a(t3_0111100), .b(t3_0111101), .y(t3_011110));
wire t3_0111100, t3_0111101;
mixer mix_t3_0111100 (.a(t3_01111000), .b(t3_01111001), .y(t3_0111100));
wire t3_01111000, t3_01111001;
mixer mix_t3_01111000 (.a(t3_011110000), .b(t3_011110001), .y(t3_01111000));
wire t3_011110000, t3_011110001;
mixer mix_t3_01111001 (.a(t3_011110010), .b(t3_011110011), .y(t3_01111001));
wire t3_011110010, t3_011110011;
mixer mix_t3_0111101 (.a(t3_01111010), .b(t3_01111011), .y(t3_0111101));
wire t3_01111010, t3_01111011;
mixer mix_t3_01111010 (.a(t3_011110100), .b(t3_011110101), .y(t3_01111010));
wire t3_011110100, t3_011110101;
mixer mix_t3_01111011 (.a(t3_011110110), .b(t3_011110111), .y(t3_01111011));
wire t3_011110110, t3_011110111;
mixer mix_t3_011111 (.a(t3_0111110), .b(t3_0111111), .y(t3_011111));
wire t3_0111110, t3_0111111;
mixer mix_t3_0111110 (.a(t3_01111100), .b(t3_01111101), .y(t3_0111110));
wire t3_01111100, t3_01111101;
mixer mix_t3_01111100 (.a(t3_011111000), .b(t3_011111001), .y(t3_01111100));
wire t3_011111000, t3_011111001;
mixer mix_t3_01111101 (.a(t3_011111010), .b(t3_011111011), .y(t3_01111101));
wire t3_011111010, t3_011111011;
mixer mix_t3_0111111 (.a(t3_01111110), .b(t3_01111111), .y(t3_0111111));
wire t3_01111110, t3_01111111;
mixer mix_t3_01111110 (.a(t3_011111100), .b(t3_011111101), .y(t3_01111110));
wire t3_011111100, t3_011111101;
mixer mix_t3_01111111 (.a(t3_011111110), .b(t3_011111111), .y(t3_01111111));
wire t3_011111110, t3_011111111;
wire t0_0;
assign out_0 = t0_0;
wire t1_0;
assign out_1 = t1_0;
wire t2_0;
assign out_2 = t2_0;
wire t3_0;
assign out_3 = t3_0;
assign input_0 = t0_000000000;
assign input_1 = t0_000000001;
assign input_2 = t0_000000010;
assign input_3 = t0_000000011;
assign input_4 = t0_000000100;
assign input_5 = t0_000000101;
assign input_6 = t0_000000110;
assign input_7 = t0_000000111;
assign input_8 = t0_000001000;
assign input_9 = t0_000001001;
assign input_10 = t0_000001010;
assign input_11 = t0_000001011;
assign input_12 = t0_000001100;
assign input_13 = t0_000001101;
assign input_14 = t0_000001110;
assign input_15 = t0_000001111;
assign input_16 = t0_000010000;
assign input_17 = t0_000010001;
assign input_18 = t0_000010010;
assign input_19 = t0_000010011;
assign input_20 = t0_000010100;
assign input_21 = t0_000010101;
assign input_22 = t0_000010110;
assign input_23 = t0_000010111;
assign input_24 = t0_000011000;
assign input_25 = t0_000011001;
assign input_26 = t0_000011010;
assign input_27 = t0_000011011;
assign input_28 = t0_000011100;
assign input_29 = t0_000011101;
assign input_30 = t0_000011110;
assign input_31 = t0_000011111;
assign input_32 = t0_000100000;
assign input_33 = t0_000100001;
assign input_34 = t0_000100010;
assign input_35 = t0_000100011;
assign input_36 = t0_000100100;
assign input_37 = t0_000100101;
assign input_38 = t0_000100110;
assign input_39 = t0_000100111;
assign input_40 = t0_000101000;
assign input_41 = t0_000101001;
assign input_42 = t0_000101010;
assign input_43 = t0_000101011;
assign input_44 = t0_000101100;
assign input_45 = t0_000101101;
assign input_46 = t0_000101110;
assign input_47 = t0_000101111;
assign input_48 = t0_000110000;
assign input_49 = t0_000110001;
assign input_50 = t0_000110010;
assign input_51 = t0_000110011;
assign input_52 = t0_000110100;
assign input_53 = t0_000110101;
assign input_54 = t0_000110110;
assign input_55 = t0_000110111;
assign input_56 = t0_000111000;
assign input_57 = t0_000111001;
assign input_58 = t0_000111010;
assign input_59 = t0_000111011;
assign input_60 = t0_000111100;
assign input_61 = t0_000111101;
assign input_62 = t0_000111110;
assign input_63 = t0_000111111;
assign input_64 = t0_001000000;
assign input_65 = t0_001000001;
assign input_66 = t0_001000010;
assign input_67 = t0_001000011;
assign input_68 = t0_001000100;
assign input_69 = t0_001000101;
assign input_70 = t0_001000110;
assign input_71 = t0_001000111;
assign input_72 = t0_001001000;
assign input_73 = t0_001001001;
assign input_74 = t0_001001010;
assign input_75 = t0_001001011;
assign input_76 = t0_001001100;
assign input_77 = t0_001001101;
assign input_78 = t0_001001110;
assign input_79 = t0_001001111;
assign input_80 = t0_001010000;
assign input_81 = t0_001010001;
assign input_82 = t0_001010010;
assign input_83 = t0_001010011;
assign input_84 = t0_001010100;
assign input_85 = t0_001010101;
assign input_86 = t0_001010110;
assign input_87 = t0_001010111;
assign input_88 = t0_001011000;
assign input_89 = t0_001011001;
assign input_90 = t0_001011010;
assign input_91 = t0_001011011;
assign input_92 = t0_001011100;
assign input_93 = t0_001011101;
assign input_94 = t0_001011110;
assign input_95 = t0_001011111;
assign input_96 = t0_001100000;
assign input_97 = t0_001100001;
assign input_98 = t0_001100010;
assign input_99 = t0_001100011;
assign input_100 = t0_001100100;
assign input_101 = t0_001100101;
assign input_102 = t0_001100110;
assign input_103 = t0_001100111;
assign input_104 = t0_001101000;
assign input_105 = t0_001101001;
assign input_106 = t0_001101010;
assign input_107 = t0_001101011;
assign input_108 = t0_001101100;
assign input_109 = t0_001101101;
assign input_110 = t0_001101110;
assign input_111 = t0_001101111;
assign input_112 = t0_001110000;
assign input_113 = t0_001110001;
assign input_114 = t0_001110010;
assign input_115 = t0_001110011;
assign input_116 = t0_001110100;
assign input_117 = t0_001110101;
assign input_118 = t0_001110110;
assign input_119 = t0_001110111;
assign input_120 = t0_001111000;
assign input_121 = t0_001111001;
assign input_122 = t0_001111010;
assign input_123 = t0_001111011;
assign input_124 = t0_001111100;
assign input_125 = t0_001111101;
assign input_126 = t0_001111110;
assign input_127 = t0_001111111;
assign input_128 = t0_010000000;
assign input_129 = t0_010000001;
assign input_130 = t0_010000010;
assign input_131 = t0_010000011;
assign input_132 = t0_010000100;
assign input_133 = t0_010000101;
assign input_134 = t0_010000110;
assign input_135 = t0_010000111;
assign input_136 = t0_010001000;
assign input_137 = t0_010001001;
assign input_138 = t0_010001010;
assign input_139 = t0_010001011;
assign input_140 = t0_010001100;
assign input_141 = t0_010001101;
assign input_142 = t0_010001110;
assign input_143 = t0_010001111;
assign input_144 = t0_010010000;
assign input_145 = t0_010010001;
assign input_146 = t0_010010010;
assign input_147 = t0_010010011;
assign input_148 = t0_010010100;
assign input_149 = t0_010010101;
assign input_150 = t0_010010110;
assign input_151 = t0_010010111;
assign input_152 = t0_010011000;
assign input_153 = t0_010011001;
assign input_154 = t0_010011010;
assign input_155 = t0_010011011;
assign input_156 = t0_010011100;
assign input_157 = t0_010011101;
assign input_158 = t0_010011110;
assign input_159 = t0_010011111;
assign input_160 = t0_010100000;
assign input_161 = t0_010100001;
assign input_162 = t0_010100010;
assign input_163 = t0_010100011;
assign input_164 = t0_010100100;
assign input_165 = t0_010100101;
assign input_166 = t0_010100110;
assign input_167 = t0_010100111;
assign input_168 = t0_010101000;
assign input_169 = t0_010101001;
assign input_170 = t0_010101010;
assign input_171 = t0_010101011;
assign input_172 = t0_010101100;
assign input_173 = t0_010101101;
assign input_174 = t0_010101110;
assign input_175 = t0_010101111;
assign input_176 = t0_010110000;
assign input_177 = t0_010110001;
assign input_178 = t0_010110010;
assign input_179 = t0_010110011;
assign input_180 = t0_010110100;
assign input_181 = t0_010110101;
assign input_182 = t0_010110110;
assign input_183 = t0_010110111;
assign input_184 = t0_010111000;
assign input_185 = t0_010111001;
assign input_186 = t0_010111010;
assign input_187 = t0_010111011;
assign input_188 = t0_010111100;
assign input_189 = t0_010111101;
assign input_190 = t0_010111110;
assign input_191 = t0_010111111;
assign input_192 = t0_011000000;
assign input_193 = t0_011000001;
assign input_194 = t0_011000010;
assign input_195 = t0_011000011;
assign input_196 = t0_011000100;
assign input_197 = t0_011000101;
assign input_198 = t0_011000110;
assign input_199 = t0_011000111;
assign input_200 = t0_011001000;
assign input_201 = t0_011001001;
assign input_202 = t0_011001010;
assign input_203 = t0_011001011;
assign input_204 = t0_011001100;
assign input_205 = t0_011001101;
assign input_206 = t0_011001110;
assign input_207 = t0_011001111;
assign input_208 = t0_011010000;
assign input_209 = t0_011010001;
assign input_210 = t0_011010010;
assign input_211 = t0_011010011;
assign input_212 = t0_011010100;
assign input_213 = t0_011010101;
assign input_214 = t0_011010110;
assign input_215 = t0_011010111;
assign input_216 = t0_011011000;
assign input_217 = t0_011011001;
assign input_218 = t0_011011010;
assign input_219 = t0_011011011;
assign input_220 = t0_011011100;
assign input_221 = t0_011011101;
assign input_222 = t0_011011110;
assign input_223 = t0_011011111;
assign input_224 = t0_011100000;
assign input_225 = t0_011100001;
assign input_226 = t0_011100010;
assign input_227 = t0_011100011;
assign input_228 = t0_011100100;
assign input_229 = t0_011100101;
assign input_230 = t0_011100110;
assign input_231 = t0_011100111;
assign input_232 = t0_011101000;
assign input_233 = t0_011101001;
assign input_234 = t0_011101010;
assign input_235 = t0_011101011;
assign input_236 = t0_011101100;
assign input_237 = t0_011101101;
assign input_238 = t0_011101110;
assign input_239 = t0_011101111;
assign input_240 = t0_011110000;
assign input_241 = t0_011110001;
assign input_242 = t0_011110010;
assign input_243 = t0_011110011;
assign input_244 = t0_011110100;
assign input_245 = t0_011110101;
assign input_246 = t0_011110110;
assign input_247 = t0_011110111;
assign input_248 = t0_011111000;
assign input_249 = t0_011111001;
assign input_250 = t0_011111010;
assign input_251 = t0_011111011;
assign input_252 = t0_011111100;
assign input_253 = t0_011111101;
assign input_254 = t0_011111110;
assign input_255 = t0_011111111;
assign input_256 = t1_000000000;
assign input_257 = t1_000000001;
assign input_258 = t1_000000010;
assign input_259 = t1_000000011;
assign input_260 = t1_000000100;
assign input_261 = t1_000000101;
assign input_262 = t1_000000110;
assign input_263 = t1_000000111;
assign input_264 = t1_000001000;
assign input_265 = t1_000001001;
assign input_266 = t1_000001010;
assign input_267 = t1_000001011;
assign input_268 = t1_000001100;
assign input_269 = t1_000001101;
assign input_270 = t1_000001110;
assign input_271 = t1_000001111;
assign input_272 = t1_000010000;
assign input_273 = t1_000010001;
assign input_274 = t1_000010010;
assign input_275 = t1_000010011;
assign input_276 = t1_000010100;
assign input_277 = t1_000010101;
assign input_278 = t1_000010110;
assign input_279 = t1_000010111;
assign input_280 = t1_000011000;
assign input_281 = t1_000011001;
assign input_282 = t1_000011010;
assign input_283 = t1_000011011;
assign input_284 = t1_000011100;
assign input_285 = t1_000011101;
assign input_286 = t1_000011110;
assign input_287 = t1_000011111;
assign input_288 = t1_000100000;
assign input_289 = t1_000100001;
assign input_290 = t1_000100010;
assign input_291 = t1_000100011;
assign input_292 = t1_000100100;
assign input_293 = t1_000100101;
assign input_294 = t1_000100110;
assign input_295 = t1_000100111;
assign input_296 = t1_000101000;
assign input_297 = t1_000101001;
assign input_298 = t1_000101010;
assign input_299 = t1_000101011;
assign input_300 = t1_000101100;
assign input_301 = t1_000101101;
assign input_302 = t1_000101110;
assign input_303 = t1_000101111;
assign input_304 = t1_000110000;
assign input_305 = t1_000110001;
assign input_306 = t1_000110010;
assign input_307 = t1_000110011;
assign input_308 = t1_000110100;
assign input_309 = t1_000110101;
assign input_310 = t1_000110110;
assign input_311 = t1_000110111;
assign input_312 = t1_000111000;
assign input_313 = t1_000111001;
assign input_314 = t1_000111010;
assign input_315 = t1_000111011;
assign input_316 = t1_000111100;
assign input_317 = t1_000111101;
assign input_318 = t1_000111110;
assign input_319 = t1_000111111;
assign input_320 = t1_001000000;
assign input_321 = t1_001000001;
assign input_322 = t1_001000010;
assign input_323 = t1_001000011;
assign input_324 = t1_001000100;
assign input_325 = t1_001000101;
assign input_326 = t1_001000110;
assign input_327 = t1_001000111;
assign input_328 = t1_001001000;
assign input_329 = t1_001001001;
assign input_330 = t1_001001010;
assign input_331 = t1_001001011;
assign input_332 = t1_001001100;
assign input_333 = t1_001001101;
assign input_334 = t1_001001110;
assign input_335 = t1_001001111;
assign input_336 = t1_001010000;
assign input_337 = t1_001010001;
assign input_338 = t1_001010010;
assign input_339 = t1_001010011;
assign input_340 = t1_001010100;
assign input_341 = t1_001010101;
assign input_342 = t1_001010110;
assign input_343 = t1_001010111;
assign input_344 = t1_001011000;
assign input_345 = t1_001011001;
assign input_346 = t1_001011010;
assign input_347 = t1_001011011;
assign input_348 = t1_001011100;
assign input_349 = t1_001011101;
assign input_350 = t1_001011110;
assign input_351 = t1_001011111;
assign input_352 = t1_001100000;
assign input_353 = t1_001100001;
assign input_354 = t1_001100010;
assign input_355 = t1_001100011;
assign input_356 = t1_001100100;
assign input_357 = t1_001100101;
assign input_358 = t1_001100110;
assign input_359 = t1_001100111;
assign input_360 = t1_001101000;
assign input_361 = t1_001101001;
assign input_362 = t1_001101010;
assign input_363 = t1_001101011;
assign input_364 = t1_001101100;
assign input_365 = t1_001101101;
assign input_366 = t1_001101110;
assign input_367 = t1_001101111;
assign input_368 = t1_001110000;
assign input_369 = t1_001110001;
assign input_370 = t1_001110010;
assign input_371 = t1_001110011;
assign input_372 = t1_001110100;
assign input_373 = t1_001110101;
assign input_374 = t1_001110110;
assign input_375 = t1_001110111;
assign input_376 = t1_001111000;
assign input_377 = t1_001111001;
assign input_378 = t1_001111010;
assign input_379 = t1_001111011;
assign input_380 = t1_001111100;
assign input_381 = t1_001111101;
assign input_382 = t1_001111110;
assign input_383 = t1_001111111;
assign input_384 = t1_010000000;
assign input_385 = t1_010000001;
assign input_386 = t1_010000010;
assign input_387 = t1_010000011;
assign input_388 = t1_010000100;
assign input_389 = t1_010000101;
assign input_390 = t1_010000110;
assign input_391 = t1_010000111;
assign input_392 = t1_010001000;
assign input_393 = t1_010001001;
assign input_394 = t1_010001010;
assign input_395 = t1_010001011;
assign input_396 = t1_010001100;
assign input_397 = t1_010001101;
assign input_398 = t1_010001110;
assign input_399 = t1_010001111;
assign input_400 = t1_010010000;
assign input_401 = t1_010010001;
assign input_402 = t1_010010010;
assign input_403 = t1_010010011;
assign input_404 = t1_010010100;
assign input_405 = t1_010010101;
assign input_406 = t1_010010110;
assign input_407 = t1_010010111;
assign input_408 = t1_010011000;
assign input_409 = t1_010011001;
assign input_410 = t1_010011010;
assign input_411 = t1_010011011;
assign input_412 = t1_010011100;
assign input_413 = t1_010011101;
assign input_414 = t1_010011110;
assign input_415 = t1_010011111;
assign input_416 = t1_010100000;
assign input_417 = t1_010100001;
assign input_418 = t1_010100010;
assign input_419 = t1_010100011;
assign input_420 = t1_010100100;
assign input_421 = t1_010100101;
assign input_422 = t1_010100110;
assign input_423 = t1_010100111;
assign input_424 = t1_010101000;
assign input_425 = t1_010101001;
assign input_426 = t1_010101010;
assign input_427 = t1_010101011;
assign input_428 = t1_010101100;
assign input_429 = t1_010101101;
assign input_430 = t1_010101110;
assign input_431 = t1_010101111;
assign input_432 = t1_010110000;
assign input_433 = t1_010110001;
assign input_434 = t1_010110010;
assign input_435 = t1_010110011;
assign input_436 = t1_010110100;
assign input_437 = t1_010110101;
assign input_438 = t1_010110110;
assign input_439 = t1_010110111;
assign input_440 = t1_010111000;
assign input_441 = t1_010111001;
assign input_442 = t1_010111010;
assign input_443 = t1_010111011;
assign input_444 = t1_010111100;
assign input_445 = t1_010111101;
assign input_446 = t1_010111110;
assign input_447 = t1_010111111;
assign input_448 = t1_011000000;
assign input_449 = t1_011000001;
assign input_450 = t1_011000010;
assign input_451 = t1_011000011;
assign input_452 = t1_011000100;
assign input_453 = t1_011000101;
assign input_454 = t1_011000110;
assign input_455 = t1_011000111;
assign input_456 = t1_011001000;
assign input_457 = t1_011001001;
assign input_458 = t1_011001010;
assign input_459 = t1_011001011;
assign input_460 = t1_011001100;
assign input_461 = t1_011001101;
assign input_462 = t1_011001110;
assign input_463 = t1_011001111;
assign input_464 = t1_011010000;
assign input_465 = t1_011010001;
assign input_466 = t1_011010010;
assign input_467 = t1_011010011;
assign input_468 = t1_011010100;
assign input_469 = t1_011010101;
assign input_470 = t1_011010110;
assign input_471 = t1_011010111;
assign input_472 = t1_011011000;
assign input_473 = t1_011011001;
assign input_474 = t1_011011010;
assign input_475 = t1_011011011;
assign input_476 = t1_011011100;
assign input_477 = t1_011011101;
assign input_478 = t1_011011110;
assign input_479 = t1_011011111;
assign input_480 = t1_011100000;
assign input_481 = t1_011100001;
assign input_482 = t1_011100010;
assign input_483 = t1_011100011;
assign input_484 = t1_011100100;
assign input_485 = t1_011100101;
assign input_486 = t1_011100110;
assign input_487 = t1_011100111;
assign input_488 = t1_011101000;
assign input_489 = t1_011101001;
assign input_490 = t1_011101010;
assign input_491 = t1_011101011;
assign input_492 = t1_011101100;
assign input_493 = t1_011101101;
assign input_494 = t1_011101110;
assign input_495 = t1_011101111;
assign input_496 = t1_011110000;
assign input_497 = t1_011110001;
assign input_498 = t1_011110010;
assign input_499 = t1_011110011;
assign input_500 = t1_011110100;
assign input_501 = t1_011110101;
assign input_502 = t1_011110110;
assign input_503 = t1_011110111;
assign input_504 = t1_011111000;
assign input_505 = t1_011111001;
assign input_506 = t1_011111010;
assign input_507 = t1_011111011;
assign input_508 = t1_011111100;
assign input_509 = t1_011111101;
assign input_510 = t1_011111110;
assign input_511 = t1_011111111;
assign input_512 = t2_000000000;
assign input_513 = t2_000000001;
assign input_514 = t2_000000010;
assign input_515 = t2_000000011;
assign input_516 = t2_000000100;
assign input_517 = t2_000000101;
assign input_518 = t2_000000110;
assign input_519 = t2_000000111;
assign input_520 = t2_000001000;
assign input_521 = t2_000001001;
assign input_522 = t2_000001010;
assign input_523 = t2_000001011;
assign input_524 = t2_000001100;
assign input_525 = t2_000001101;
assign input_526 = t2_000001110;
assign input_527 = t2_000001111;
assign input_528 = t2_000010000;
assign input_529 = t2_000010001;
assign input_530 = t2_000010010;
assign input_531 = t2_000010011;
assign input_532 = t2_000010100;
assign input_533 = t2_000010101;
assign input_534 = t2_000010110;
assign input_535 = t2_000010111;
assign input_536 = t2_000011000;
assign input_537 = t2_000011001;
assign input_538 = t2_000011010;
assign input_539 = t2_000011011;
assign input_540 = t2_000011100;
assign input_541 = t2_000011101;
assign input_542 = t2_000011110;
assign input_543 = t2_000011111;
assign input_544 = t2_000100000;
assign input_545 = t2_000100001;
assign input_546 = t2_000100010;
assign input_547 = t2_000100011;
assign input_548 = t2_000100100;
assign input_549 = t2_000100101;
assign input_550 = t2_000100110;
assign input_551 = t2_000100111;
assign input_552 = t2_000101000;
assign input_553 = t2_000101001;
assign input_554 = t2_000101010;
assign input_555 = t2_000101011;
assign input_556 = t2_000101100;
assign input_557 = t2_000101101;
assign input_558 = t2_000101110;
assign input_559 = t2_000101111;
assign input_560 = t2_000110000;
assign input_561 = t2_000110001;
assign input_562 = t2_000110010;
assign input_563 = t2_000110011;
assign input_564 = t2_000110100;
assign input_565 = t2_000110101;
assign input_566 = t2_000110110;
assign input_567 = t2_000110111;
assign input_568 = t2_000111000;
assign input_569 = t2_000111001;
assign input_570 = t2_000111010;
assign input_571 = t2_000111011;
assign input_572 = t2_000111100;
assign input_573 = t2_000111101;
assign input_574 = t2_000111110;
assign input_575 = t2_000111111;
assign input_576 = t2_001000000;
assign input_577 = t2_001000001;
assign input_578 = t2_001000010;
assign input_579 = t2_001000011;
assign input_580 = t2_001000100;
assign input_581 = t2_001000101;
assign input_582 = t2_001000110;
assign input_583 = t2_001000111;
assign input_584 = t2_001001000;
assign input_585 = t2_001001001;
assign input_586 = t2_001001010;
assign input_587 = t2_001001011;
assign input_588 = t2_001001100;
assign input_589 = t2_001001101;
assign input_590 = t2_001001110;
assign input_591 = t2_001001111;
assign input_592 = t2_001010000;
assign input_593 = t2_001010001;
assign input_594 = t2_001010010;
assign input_595 = t2_001010011;
assign input_596 = t2_001010100;
assign input_597 = t2_001010101;
assign input_598 = t2_001010110;
assign input_599 = t2_001010111;
assign input_600 = t2_001011000;
assign input_601 = t2_001011001;
assign input_602 = t2_001011010;
assign input_603 = t2_001011011;
assign input_604 = t2_001011100;
assign input_605 = t2_001011101;
assign input_606 = t2_001011110;
assign input_607 = t2_001011111;
assign input_608 = t2_001100000;
assign input_609 = t2_001100001;
assign input_610 = t2_001100010;
assign input_611 = t2_001100011;
assign input_612 = t2_001100100;
assign input_613 = t2_001100101;
assign input_614 = t2_001100110;
assign input_615 = t2_001100111;
assign input_616 = t2_001101000;
assign input_617 = t2_001101001;
assign input_618 = t2_001101010;
assign input_619 = t2_001101011;
assign input_620 = t2_001101100;
assign input_621 = t2_001101101;
assign input_622 = t2_001101110;
assign input_623 = t2_001101111;
assign input_624 = t2_001110000;
assign input_625 = t2_001110001;
assign input_626 = t2_001110010;
assign input_627 = t2_001110011;
assign input_628 = t2_001110100;
assign input_629 = t2_001110101;
assign input_630 = t2_001110110;
assign input_631 = t2_001110111;
assign input_632 = t2_001111000;
assign input_633 = t2_001111001;
assign input_634 = t2_001111010;
assign input_635 = t2_001111011;
assign input_636 = t2_001111100;
assign input_637 = t2_001111101;
assign input_638 = t2_001111110;
assign input_639 = t2_001111111;
assign input_640 = t2_010000000;
assign input_641 = t2_010000001;
assign input_642 = t2_010000010;
assign input_643 = t2_010000011;
assign input_644 = t2_010000100;
assign input_645 = t2_010000101;
assign input_646 = t2_010000110;
assign input_647 = t2_010000111;
assign input_648 = t2_010001000;
assign input_649 = t2_010001001;
assign input_650 = t2_010001010;
assign input_651 = t2_010001011;
assign input_652 = t2_010001100;
assign input_653 = t2_010001101;
assign input_654 = t2_010001110;
assign input_655 = t2_010001111;
assign input_656 = t2_010010000;
assign input_657 = t2_010010001;
assign input_658 = t2_010010010;
assign input_659 = t2_010010011;
assign input_660 = t2_010010100;
assign input_661 = t2_010010101;
assign input_662 = t2_010010110;
assign input_663 = t2_010010111;
assign input_664 = t2_010011000;
assign input_665 = t2_010011001;
assign input_666 = t2_010011010;
assign input_667 = t2_010011011;
assign input_668 = t2_010011100;
assign input_669 = t2_010011101;
assign input_670 = t2_010011110;
assign input_671 = t2_010011111;
assign input_672 = t2_010100000;
assign input_673 = t2_010100001;
assign input_674 = t2_010100010;
assign input_675 = t2_010100011;
assign input_676 = t2_010100100;
assign input_677 = t2_010100101;
assign input_678 = t2_010100110;
assign input_679 = t2_010100111;
assign input_680 = t2_010101000;
assign input_681 = t2_010101001;
assign input_682 = t2_010101010;
assign input_683 = t2_010101011;
assign input_684 = t2_010101100;
assign input_685 = t2_010101101;
assign input_686 = t2_010101110;
assign input_687 = t2_010101111;
assign input_688 = t2_010110000;
assign input_689 = t2_010110001;
assign input_690 = t2_010110010;
assign input_691 = t2_010110011;
assign input_692 = t2_010110100;
assign input_693 = t2_010110101;
assign input_694 = t2_010110110;
assign input_695 = t2_010110111;
assign input_696 = t2_010111000;
assign input_697 = t2_010111001;
assign input_698 = t2_010111010;
assign input_699 = t2_010111011;
assign input_700 = t2_010111100;
assign input_701 = t2_010111101;
assign input_702 = t2_010111110;
assign input_703 = t2_010111111;
assign input_704 = t2_011000000;
assign input_705 = t2_011000001;
assign input_706 = t2_011000010;
assign input_707 = t2_011000011;
assign input_708 = t2_011000100;
assign input_709 = t2_011000101;
assign input_710 = t2_011000110;
assign input_711 = t2_011000111;
assign input_712 = t2_011001000;
assign input_713 = t2_011001001;
assign input_714 = t2_011001010;
assign input_715 = t2_011001011;
assign input_716 = t2_011001100;
assign input_717 = t2_011001101;
assign input_718 = t2_011001110;
assign input_719 = t2_011001111;
assign input_720 = t2_011010000;
assign input_721 = t2_011010001;
assign input_722 = t2_011010010;
assign input_723 = t2_011010011;
assign input_724 = t2_011010100;
assign input_725 = t2_011010101;
assign input_726 = t2_011010110;
assign input_727 = t2_011010111;
assign input_728 = t2_011011000;
assign input_729 = t2_011011001;
assign input_730 = t2_011011010;
assign input_731 = t2_011011011;
assign input_732 = t2_011011100;
assign input_733 = t2_011011101;
assign input_734 = t2_011011110;
assign input_735 = t2_011011111;
assign input_736 = t2_011100000;
assign input_737 = t2_011100001;
assign input_738 = t2_011100010;
assign input_739 = t2_011100011;
assign input_740 = t2_011100100;
assign input_741 = t2_011100101;
assign input_742 = t2_011100110;
assign input_743 = t2_011100111;
assign input_744 = t2_011101000;
assign input_745 = t2_011101001;
assign input_746 = t2_011101010;
assign input_747 = t2_011101011;
assign input_748 = t2_011101100;
assign input_749 = t2_011101101;
assign input_750 = t2_011101110;
assign input_751 = t2_011101111;
assign input_752 = t2_011110000;
assign input_753 = t2_011110001;
assign input_754 = t2_011110010;
assign input_755 = t2_011110011;
assign input_756 = t2_011110100;
assign input_757 = t2_011110101;
assign input_758 = t2_011110110;
assign input_759 = t2_011110111;
assign input_760 = t2_011111000;
assign input_761 = t2_011111001;
assign input_762 = t2_011111010;
assign input_763 = t2_011111011;
assign input_764 = t2_011111100;
assign input_765 = t2_011111101;
assign input_766 = t2_011111110;
assign input_767 = t2_011111111;
assign input_768 = t3_000000000;
assign input_769 = t3_000000001;
assign input_770 = t3_000000010;
assign input_771 = t3_000000011;
assign input_772 = t3_000000100;
assign input_773 = t3_000000101;
assign input_774 = t3_000000110;
assign input_775 = t3_000000111;
assign input_776 = t3_000001000;
assign input_777 = t3_000001001;
assign input_778 = t3_000001010;
assign input_779 = t3_000001011;
assign input_780 = t3_000001100;
assign input_781 = t3_000001101;
assign input_782 = t3_000001110;
assign input_783 = t3_000001111;
assign input_784 = t3_000010000;
assign input_785 = t3_000010001;
assign input_786 = t3_000010010;
assign input_787 = t3_000010011;
assign input_788 = t3_000010100;
assign input_789 = t3_000010101;
assign input_790 = t3_000010110;
assign input_791 = t3_000010111;
assign input_792 = t3_000011000;
assign input_793 = t3_000011001;
assign input_794 = t3_000011010;
assign input_795 = t3_000011011;
assign input_796 = t3_000011100;
assign input_797 = t3_000011101;
assign input_798 = t3_000011110;
assign input_799 = t3_000011111;
assign input_800 = t3_000100000;
assign input_801 = t3_000100001;
assign input_802 = t3_000100010;
assign input_803 = t3_000100011;
assign input_804 = t3_000100100;
assign input_805 = t3_000100101;
assign input_806 = t3_000100110;
assign input_807 = t3_000100111;
assign input_808 = t3_000101000;
assign input_809 = t3_000101001;
assign input_810 = t3_000101010;
assign input_811 = t3_000101011;
assign input_812 = t3_000101100;
assign input_813 = t3_000101101;
assign input_814 = t3_000101110;
assign input_815 = t3_000101111;
assign input_816 = t3_000110000;
assign input_817 = t3_000110001;
assign input_818 = t3_000110010;
assign input_819 = t3_000110011;
assign input_820 = t3_000110100;
assign input_821 = t3_000110101;
assign input_822 = t3_000110110;
assign input_823 = t3_000110111;
assign input_824 = t3_000111000;
assign input_825 = t3_000111001;
assign input_826 = t3_000111010;
assign input_827 = t3_000111011;
assign input_828 = t3_000111100;
assign input_829 = t3_000111101;
assign input_830 = t3_000111110;
assign input_831 = t3_000111111;
assign input_832 = t3_001000000;
assign input_833 = t3_001000001;
assign input_834 = t3_001000010;
assign input_835 = t3_001000011;
assign input_836 = t3_001000100;
assign input_837 = t3_001000101;
assign input_838 = t3_001000110;
assign input_839 = t3_001000111;
assign input_840 = t3_001001000;
assign input_841 = t3_001001001;
assign input_842 = t3_001001010;
assign input_843 = t3_001001011;
assign input_844 = t3_001001100;
assign input_845 = t3_001001101;
assign input_846 = t3_001001110;
assign input_847 = t3_001001111;
assign input_848 = t3_001010000;
assign input_849 = t3_001010001;
assign input_850 = t3_001010010;
assign input_851 = t3_001010011;
assign input_852 = t3_001010100;
assign input_853 = t3_001010101;
assign input_854 = t3_001010110;
assign input_855 = t3_001010111;
assign input_856 = t3_001011000;
assign input_857 = t3_001011001;
assign input_858 = t3_001011010;
assign input_859 = t3_001011011;
assign input_860 = t3_001011100;
assign input_861 = t3_001011101;
assign input_862 = t3_001011110;
assign input_863 = t3_001011111;
assign input_864 = t3_001100000;
assign input_865 = t3_001100001;
assign input_866 = t3_001100010;
assign input_867 = t3_001100011;
assign input_868 = t3_001100100;
assign input_869 = t3_001100101;
assign input_870 = t3_001100110;
assign input_871 = t3_001100111;
assign input_872 = t3_001101000;
assign input_873 = t3_001101001;
assign input_874 = t3_001101010;
assign input_875 = t3_001101011;
assign input_876 = t3_001101100;
assign input_877 = t3_001101101;
assign input_878 = t3_001101110;
assign input_879 = t3_001101111;
assign input_880 = t3_001110000;
assign input_881 = t3_001110001;
assign input_882 = t3_001110010;
assign input_883 = t3_001110011;
assign input_884 = t3_001110100;
assign input_885 = t3_001110101;
assign input_886 = t3_001110110;
assign input_887 = t3_001110111;
assign input_888 = t3_001111000;
assign input_889 = t3_001111001;
assign input_890 = t3_001111010;
assign input_891 = t3_001111011;
assign input_892 = t3_001111100;
assign input_893 = t3_001111101;
assign input_894 = t3_001111110;
assign input_895 = t3_001111111;
assign input_896 = t3_010000000;
assign input_897 = t3_010000001;
assign input_898 = t3_010000010;
assign input_899 = t3_010000011;
assign input_900 = t3_010000100;
assign input_901 = t3_010000101;
assign input_902 = t3_010000110;
assign input_903 = t3_010000111;
assign input_904 = t3_010001000;
assign input_905 = t3_010001001;
assign input_906 = t3_010001010;
assign input_907 = t3_010001011;
assign input_908 = t3_010001100;
assign input_909 = t3_010001101;
assign input_910 = t3_010001110;
assign input_911 = t3_010001111;
assign input_912 = t3_010010000;
assign input_913 = t3_010010001;
assign input_914 = t3_010010010;
assign input_915 = t3_010010011;
assign input_916 = t3_010010100;
assign input_917 = t3_010010101;
assign input_918 = t3_010010110;
assign input_919 = t3_010010111;
assign input_920 = t3_010011000;
assign input_921 = t3_010011001;
assign input_922 = t3_010011010;
assign input_923 = t3_010011011;
assign input_924 = t3_010011100;
assign input_925 = t3_010011101;
assign input_926 = t3_010011110;
assign input_927 = t3_010011111;
assign input_928 = t3_010100000;
assign input_929 = t3_010100001;
assign input_930 = t3_010100010;
assign input_931 = t3_010100011;
assign input_932 = t3_010100100;
assign input_933 = t3_010100101;
assign input_934 = t3_010100110;
assign input_935 = t3_010100111;
assign input_936 = t3_010101000;
assign input_937 = t3_010101001;
assign input_938 = t3_010101010;
assign input_939 = t3_010101011;
assign input_940 = t3_010101100;
assign input_941 = t3_010101101;
assign input_942 = t3_010101110;
assign input_943 = t3_010101111;
assign input_944 = t3_010110000;
assign input_945 = t3_010110001;
assign input_946 = t3_010110010;
assign input_947 = t3_010110011;
assign input_948 = t3_010110100;
assign input_949 = t3_010110101;
assign input_950 = t3_010110110;
assign input_951 = t3_010110111;
assign input_952 = t3_010111000;
assign input_953 = t3_010111001;
assign input_954 = t3_010111010;
assign input_955 = t3_010111011;
assign input_956 = t3_010111100;
assign input_957 = t3_010111101;
assign input_958 = t3_010111110;
assign input_959 = t3_010111111;
assign input_960 = t3_011000000;
assign input_961 = t3_011000001;
assign input_962 = t3_011000010;
assign input_963 = t3_011000011;
assign input_964 = t3_011000100;
assign input_965 = t3_011000101;
assign input_966 = t3_011000110;
assign input_967 = t3_011000111;
assign input_968 = t3_011001000;
assign input_969 = t3_011001001;
assign input_970 = t3_011001010;
assign input_971 = t3_011001011;
assign input_972 = t3_011001100;
assign input_973 = t3_011001101;
assign input_974 = t3_011001110;
assign input_975 = t3_011001111;
assign input_976 = t3_011010000;
assign input_977 = t3_011010001;
assign input_978 = t3_011010010;
assign input_979 = t3_011010011;
assign input_980 = t3_011010100;
assign input_981 = t3_011010101;
assign input_982 = t3_011010110;
assign input_983 = t3_011010111;
assign input_984 = t3_011011000;
assign input_985 = t3_011011001;
assign input_986 = t3_011011010;
assign input_987 = t3_011011011;
assign input_988 = t3_011011100;
assign input_989 = t3_011011101;
assign input_990 = t3_011011110;
assign input_991 = t3_011011111;
assign input_992 = t3_011100000;
assign input_993 = t3_011100001;
assign input_994 = t3_011100010;
assign input_995 = t3_011100011;
assign input_996 = t3_011100100;
assign input_997 = t3_011100101;
assign input_998 = t3_011100110;
assign input_999 = t3_011100111;
assign input_1000 = t3_011101000;
assign input_1001 = t3_011101001;
assign input_1002 = t3_011101010;
assign input_1003 = t3_011101011;
assign input_1004 = t3_011101100;
assign input_1005 = t3_011101101;
assign input_1006 = t3_011101110;
assign input_1007 = t3_011101111;
assign input_1008 = t3_011110000;
assign input_1009 = t3_011110001;
assign input_1010 = t3_011110010;
assign input_1011 = t3_011110011;
assign input_1012 = t3_011110100;
assign input_1013 = t3_011110101;
assign input_1014 = t3_011110110;
assign input_1015 = t3_011110111;
assign input_1016 = t3_011111000;
assign input_1017 = t3_011111001;
assign input_1018 = t3_011111010;
assign input_1019 = t3_011111011;
assign input_1020 = t3_011111100;
assign input_1021 = t3_011111101;
assign input_1022 = t3_011111110;
assign input_1023 = t3_011111111;
endmodule
