module fanout2_mesh_16_3 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,output output_8,output output_9,output output_10,output output_11,output output_12,output output_13,output output_14,output output_15,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15
);
wire output_1_0, output_1_1, output_0_0;
diffmix_25px_0 gate_output_0_0(.a_fluid(output_1_0), .b_fluid(output_1_1), .out_fluid(output_0_0));
wire output_2_0, output_2_1, output_1_0;
diffmix_25px_0 gate_output_1_0(.a_fluid(output_2_0), .b_fluid(output_2_1), .out_fluid(output_1_0));
wire output_3_0, output_3_1, output_2_0;
diffmix_25px_0 gate_output_2_0(.a_fluid(output_3_0), .b_fluid(output_3_1), .out_fluid(output_2_0));
wire output_4_0, output_4_1, output_3_0;
diffmix_25px_0 gate_output_3_0(.a_fluid(output_4_0), .b_fluid(output_4_1), .out_fluid(output_3_0));
wire output_5_0, output_5_1, output_4_0;
diffmix_25px_0 gate_output_4_0(.a_fluid(output_5_0), .b_fluid(output_5_1), .out_fluid(output_4_0));
wire output_6_0, output_6_1, output_5_0;
diffmix_25px_0 gate_output_5_0(.a_fluid(output_6_0), .b_fluid(output_6_1), .out_fluid(output_5_0));
wire output_7_0, output_7_1, output_6_0;
diffmix_25px_0 gate_output_6_0(.a_fluid(output_7_0), .b_fluid(output_7_1), .out_fluid(output_6_0));
wire output_8_0, output_8_1, output_7_0;
diffmix_25px_0 gate_output_7_0(.a_fluid(output_8_0), .b_fluid(output_8_1), .out_fluid(output_7_0));
wire output_9_0, output_9_1, output_8_0;
diffmix_25px_0 gate_output_8_0(.a_fluid(output_9_0), .b_fluid(output_9_1), .out_fluid(output_8_0));
wire output_10_0, output_10_1, output_9_0;
diffmix_25px_0 gate_output_9_0(.a_fluid(output_10_0), .b_fluid(output_10_1), .out_fluid(output_9_0));
wire output_11_0, output_11_1, output_10_0;
diffmix_25px_0 gate_output_10_0(.a_fluid(output_11_0), .b_fluid(output_11_1), .out_fluid(output_10_0));
wire output_12_0, output_12_1, output_11_0;
diffmix_25px_0 gate_output_11_0(.a_fluid(output_12_0), .b_fluid(output_12_1), .out_fluid(output_11_0));
wire output_13_0, output_13_1, output_12_0;
diffmix_25px_0 gate_output_12_0(.a_fluid(output_13_0), .b_fluid(output_13_1), .out_fluid(output_12_0));
wire output_14_0, output_14_1, output_13_0;
diffmix_25px_0 gate_output_13_0(.a_fluid(output_14_0), .b_fluid(output_14_1), .out_fluid(output_13_0));
wire output_15_0, output_15_1, output_14_0;
diffmix_25px_0 gate_output_14_0(.a_fluid(output_15_0), .b_fluid(output_15_1), .out_fluid(output_14_0));
wire output_16_0, output_16_1, output_15_0;
diffmix_25px_0 gate_output_15_0(.a_fluid(output_16_0), .b_fluid(output_16_1), .out_fluid(output_15_0));
wire output_1_1, output_1_2, output_0_1;
diffmix_25px_0 gate_output_0_1(.a_fluid(output_1_1), .b_fluid(output_1_2), .out_fluid(output_0_1));
wire output_2_1, output_2_2, output_1_1;
diffmix_25px_0 gate_output_1_1(.a_fluid(output_2_1), .b_fluid(output_2_2), .out_fluid(output_1_1));
wire output_3_1, output_3_2, output_2_1;
diffmix_25px_0 gate_output_2_1(.a_fluid(output_3_1), .b_fluid(output_3_2), .out_fluid(output_2_1));
wire output_4_1, output_4_2, output_3_1;
diffmix_25px_0 gate_output_3_1(.a_fluid(output_4_1), .b_fluid(output_4_2), .out_fluid(output_3_1));
wire output_5_1, output_5_2, output_4_1;
diffmix_25px_0 gate_output_4_1(.a_fluid(output_5_1), .b_fluid(output_5_2), .out_fluid(output_4_1));
wire output_6_1, output_6_2, output_5_1;
diffmix_25px_0 gate_output_5_1(.a_fluid(output_6_1), .b_fluid(output_6_2), .out_fluid(output_5_1));
wire output_7_1, output_7_2, output_6_1;
diffmix_25px_0 gate_output_6_1(.a_fluid(output_7_1), .b_fluid(output_7_2), .out_fluid(output_6_1));
wire output_8_1, output_8_2, output_7_1;
diffmix_25px_0 gate_output_7_1(.a_fluid(output_8_1), .b_fluid(output_8_2), .out_fluid(output_7_1));
wire output_9_1, output_9_2, output_8_1;
diffmix_25px_0 gate_output_8_1(.a_fluid(output_9_1), .b_fluid(output_9_2), .out_fluid(output_8_1));
wire output_10_1, output_10_2, output_9_1;
diffmix_25px_0 gate_output_9_1(.a_fluid(output_10_1), .b_fluid(output_10_2), .out_fluid(output_9_1));
wire output_11_1, output_11_2, output_10_1;
diffmix_25px_0 gate_output_10_1(.a_fluid(output_11_1), .b_fluid(output_11_2), .out_fluid(output_10_1));
wire output_12_1, output_12_2, output_11_1;
diffmix_25px_0 gate_output_11_1(.a_fluid(output_12_1), .b_fluid(output_12_2), .out_fluid(output_11_1));
wire output_13_1, output_13_2, output_12_1;
diffmix_25px_0 gate_output_12_1(.a_fluid(output_13_1), .b_fluid(output_13_2), .out_fluid(output_12_1));
wire output_14_1, output_14_2, output_13_1;
diffmix_25px_0 gate_output_13_1(.a_fluid(output_14_1), .b_fluid(output_14_2), .out_fluid(output_13_1));
wire output_15_1, output_15_2, output_14_1;
diffmix_25px_0 gate_output_14_1(.a_fluid(output_15_1), .b_fluid(output_15_2), .out_fluid(output_14_1));
wire output_16_1, output_16_2, output_15_1;
diffmix_25px_0 gate_output_15_1(.a_fluid(output_16_1), .b_fluid(output_16_2), .out_fluid(output_15_1));
wire output_1_2, output_1_3, output_0_2;
diffmix_25px_0 gate_output_0_2(.a_fluid(output_1_2), .b_fluid(output_1_3), .out_fluid(output_0_2));
wire output_2_2, output_2_3, output_1_2;
diffmix_25px_0 gate_output_1_2(.a_fluid(output_2_2), .b_fluid(output_2_3), .out_fluid(output_1_2));
wire output_3_2, output_3_3, output_2_2;
diffmix_25px_0 gate_output_2_2(.a_fluid(output_3_2), .b_fluid(output_3_3), .out_fluid(output_2_2));
wire output_4_2, output_4_3, output_3_2;
diffmix_25px_0 gate_output_3_2(.a_fluid(output_4_2), .b_fluid(output_4_3), .out_fluid(output_3_2));
wire output_5_2, output_5_3, output_4_2;
diffmix_25px_0 gate_output_4_2(.a_fluid(output_5_2), .b_fluid(output_5_3), .out_fluid(output_4_2));
wire output_6_2, output_6_3, output_5_2;
diffmix_25px_0 gate_output_5_2(.a_fluid(output_6_2), .b_fluid(output_6_3), .out_fluid(output_5_2));
wire output_7_2, output_7_3, output_6_2;
diffmix_25px_0 gate_output_6_2(.a_fluid(output_7_2), .b_fluid(output_7_3), .out_fluid(output_6_2));
wire output_8_2, output_8_3, output_7_2;
diffmix_25px_0 gate_output_7_2(.a_fluid(output_8_2), .b_fluid(output_8_3), .out_fluid(output_7_2));
wire output_9_2, output_9_3, output_8_2;
diffmix_25px_0 gate_output_8_2(.a_fluid(output_9_2), .b_fluid(output_9_3), .out_fluid(output_8_2));
wire output_10_2, output_10_3, output_9_2;
diffmix_25px_0 gate_output_9_2(.a_fluid(output_10_2), .b_fluid(output_10_3), .out_fluid(output_9_2));
wire output_11_2, output_11_3, output_10_2;
diffmix_25px_0 gate_output_10_2(.a_fluid(output_11_2), .b_fluid(output_11_3), .out_fluid(output_10_2));
wire output_12_2, output_12_3, output_11_2;
diffmix_25px_0 gate_output_11_2(.a_fluid(output_12_2), .b_fluid(output_12_3), .out_fluid(output_11_2));
wire output_13_2, output_13_3, output_12_2;
diffmix_25px_0 gate_output_12_2(.a_fluid(output_13_2), .b_fluid(output_13_3), .out_fluid(output_12_2));
wire output_14_2, output_14_3, output_13_2;
diffmix_25px_0 gate_output_13_2(.a_fluid(output_14_2), .b_fluid(output_14_3), .out_fluid(output_13_2));
wire output_15_2, output_15_3, output_14_2;
diffmix_25px_0 gate_output_14_2(.a_fluid(output_15_2), .b_fluid(output_15_3), .out_fluid(output_14_2));
wire output_16_2, output_16_3, output_15_2;
diffmix_25px_0 gate_output_15_2(.a_fluid(output_16_2), .b_fluid(output_16_3), .out_fluid(output_15_2));
assign output_0 = output_0_0;
wire output_0_3;
assign output_0_3 = input_0;
assign output_1 = output_1_0;
wire output_1_3;
assign output_1_3 = input_1;
assign output_2 = output_2_0;
wire output_2_3;
assign output_2_3 = input_2;
assign output_3 = output_3_0;
wire output_3_3;
assign output_3_3 = input_3;
assign output_4 = output_4_0;
wire output_4_3;
assign output_4_3 = input_4;
assign output_5 = output_5_0;
wire output_5_3;
assign output_5_3 = input_5;
assign output_6 = output_6_0;
wire output_6_3;
assign output_6_3 = input_6;
assign output_7 = output_7_0;
wire output_7_3;
assign output_7_3 = input_7;
assign output_8 = output_8_0;
wire output_8_3;
assign output_8_3 = input_8;
assign output_9 = output_9_0;
wire output_9_3;
assign output_9_3 = input_9;
assign output_10 = output_10_0;
wire output_10_3;
assign output_10_3 = input_10;
assign output_11 = output_11_0;
wire output_11_3;
assign output_11_3 = input_11;
assign output_12 = output_12_0;
wire output_12_3;
assign output_12_3 = input_12;
assign output_13 = output_13_0;
wire output_13_3;
assign output_13_3 = input_13;
assign output_14 = output_14_0;
wire output_14_3;
assign output_14_3 = input_14;
assign output_15 = output_15_0;
wire output_15_3;
assign output_15_3 = input_15;
endmodule
