module complete_128 (
inout io_0,inout io_1,inout io_2,inout io_3,inout io_4,inout io_5,inout io_6,inout io_7,inout io_8,inout io_9,inout io_10,inout io_11,inout io_12,inout io_13,inout io_14,inout io_15,inout io_16,inout io_17,inout io_18,inout io_19,inout io_20,inout io_21,inout io_22,inout io_23,inout io_24,inout io_25,inout io_26,inout io_27,inout io_28,inout io_29,inout io_30,inout io_31,inout io_32,inout io_33,inout io_34,inout io_35,inout io_36,inout io_37,inout io_38,inout io_39,inout io_40,inout io_41,inout io_42,inout io_43,inout io_44,inout io_45,inout io_46,inout io_47,inout io_48,inout io_49,inout io_50,inout io_51,inout io_52,inout io_53,inout io_54,inout io_55,inout io_56,inout io_57,inout io_58,inout io_59,inout io_60,inout io_61,inout io_62,inout io_63,inout io_64,inout io_65,inout io_66,inout io_67,inout io_68,inout io_69,inout io_70,inout io_71,inout io_72,inout io_73,inout io_74,inout io_75,inout io_76,inout io_77,inout io_78,inout io_79,inout io_80,inout io_81,inout io_82,inout io_83,inout io_84,inout io_85,inout io_86,inout io_87,inout io_88,inout io_89,inout io_90,inout io_91,inout io_92,inout io_93,inout io_94,inout io_95,inout io_96,inout io_97,inout io_98,inout io_99,inout io_100,inout io_101,inout io_102,inout io_103,inout io_104,inout io_105,inout io_106,inout io_107,inout io_108,inout io_109,inout io_110,inout io_111,inout io_112,inout io_113,inout io_114,inout io_115,inout io_116,inout io_117,inout io_118,inout io_119,inout io_120,inout io_121,inout io_122,inout io_123,inout io_124,inout io_125,inout io_126,inout io_127
);
assign io_0 = input_0;
assign io_0 = input_1;
assign io_0 = input_2;
assign io_0 = input_3;
assign io_0 = input_4;
assign io_0 = input_5;
assign io_0 = input_6;
assign io_0 = input_7;
assign io_0 = input_8;
assign io_0 = input_9;
assign io_0 = input_10;
assign io_0 = input_11;
assign io_0 = input_12;
assign io_0 = input_13;
assign io_0 = input_14;
assign io_0 = input_15;
assign io_0 = input_16;
assign io_0 = input_17;
assign io_0 = input_18;
assign io_0 = input_19;
assign io_0 = input_20;
assign io_0 = input_21;
assign io_0 = input_22;
assign io_0 = input_23;
assign io_0 = input_24;
assign io_0 = input_25;
assign io_0 = input_26;
assign io_0 = input_27;
assign io_0 = input_28;
assign io_0 = input_29;
assign io_0 = input_30;
assign io_0 = input_31;
assign io_0 = input_32;
assign io_0 = input_33;
assign io_0 = input_34;
assign io_0 = input_35;
assign io_0 = input_36;
assign io_0 = input_37;
assign io_0 = input_38;
assign io_0 = input_39;
assign io_0 = input_40;
assign io_0 = input_41;
assign io_0 = input_42;
assign io_0 = input_43;
assign io_0 = input_44;
assign io_0 = input_45;
assign io_0 = input_46;
assign io_0 = input_47;
assign io_0 = input_48;
assign io_0 = input_49;
assign io_0 = input_50;
assign io_0 = input_51;
assign io_0 = input_52;
assign io_0 = input_53;
assign io_0 = input_54;
assign io_0 = input_55;
assign io_0 = input_56;
assign io_0 = input_57;
assign io_0 = input_58;
assign io_0 = input_59;
assign io_0 = input_60;
assign io_0 = input_61;
assign io_0 = input_62;
assign io_0 = input_63;
assign io_0 = input_64;
assign io_0 = input_65;
assign io_0 = input_66;
assign io_0 = input_67;
assign io_0 = input_68;
assign io_0 = input_69;
assign io_0 = input_70;
assign io_0 = input_71;
assign io_0 = input_72;
assign io_0 = input_73;
assign io_0 = input_74;
assign io_0 = input_75;
assign io_0 = input_76;
assign io_0 = input_77;
assign io_0 = input_78;
assign io_0 = input_79;
assign io_0 = input_80;
assign io_0 = input_81;
assign io_0 = input_82;
assign io_0 = input_83;
assign io_0 = input_84;
assign io_0 = input_85;
assign io_0 = input_86;
assign io_0 = input_87;
assign io_0 = input_88;
assign io_0 = input_89;
assign io_0 = input_90;
assign io_0 = input_91;
assign io_0 = input_92;
assign io_0 = input_93;
assign io_0 = input_94;
assign io_0 = input_95;
assign io_0 = input_96;
assign io_0 = input_97;
assign io_0 = input_98;
assign io_0 = input_99;
assign io_0 = input_100;
assign io_0 = input_101;
assign io_0 = input_102;
assign io_0 = input_103;
assign io_0 = input_104;
assign io_0 = input_105;
assign io_0 = input_106;
assign io_0 = input_107;
assign io_0 = input_108;
assign io_0 = input_109;
assign io_0 = input_110;
assign io_0 = input_111;
assign io_0 = input_112;
assign io_0 = input_113;
assign io_0 = input_114;
assign io_0 = input_115;
assign io_0 = input_116;
assign io_0 = input_117;
assign io_0 = input_118;
assign io_0 = input_119;
assign io_0 = input_120;
assign io_0 = input_121;
assign io_0 = input_122;
assign io_0 = input_123;
assign io_0 = input_124;
assign io_0 = input_125;
assign io_0 = input_126;
assign io_0 = input_127;
assign io_1 = input_1;
assign io_1 = input_2;
assign io_1 = input_3;
assign io_1 = input_4;
assign io_1 = input_5;
assign io_1 = input_6;
assign io_1 = input_7;
assign io_1 = input_8;
assign io_1 = input_9;
assign io_1 = input_10;
assign io_1 = input_11;
assign io_1 = input_12;
assign io_1 = input_13;
assign io_1 = input_14;
assign io_1 = input_15;
assign io_1 = input_16;
assign io_1 = input_17;
assign io_1 = input_18;
assign io_1 = input_19;
assign io_1 = input_20;
assign io_1 = input_21;
assign io_1 = input_22;
assign io_1 = input_23;
assign io_1 = input_24;
assign io_1 = input_25;
assign io_1 = input_26;
assign io_1 = input_27;
assign io_1 = input_28;
assign io_1 = input_29;
assign io_1 = input_30;
assign io_1 = input_31;
assign io_1 = input_32;
assign io_1 = input_33;
assign io_1 = input_34;
assign io_1 = input_35;
assign io_1 = input_36;
assign io_1 = input_37;
assign io_1 = input_38;
assign io_1 = input_39;
assign io_1 = input_40;
assign io_1 = input_41;
assign io_1 = input_42;
assign io_1 = input_43;
assign io_1 = input_44;
assign io_1 = input_45;
assign io_1 = input_46;
assign io_1 = input_47;
assign io_1 = input_48;
assign io_1 = input_49;
assign io_1 = input_50;
assign io_1 = input_51;
assign io_1 = input_52;
assign io_1 = input_53;
assign io_1 = input_54;
assign io_1 = input_55;
assign io_1 = input_56;
assign io_1 = input_57;
assign io_1 = input_58;
assign io_1 = input_59;
assign io_1 = input_60;
assign io_1 = input_61;
assign io_1 = input_62;
assign io_1 = input_63;
assign io_1 = input_64;
assign io_1 = input_65;
assign io_1 = input_66;
assign io_1 = input_67;
assign io_1 = input_68;
assign io_1 = input_69;
assign io_1 = input_70;
assign io_1 = input_71;
assign io_1 = input_72;
assign io_1 = input_73;
assign io_1 = input_74;
assign io_1 = input_75;
assign io_1 = input_76;
assign io_1 = input_77;
assign io_1 = input_78;
assign io_1 = input_79;
assign io_1 = input_80;
assign io_1 = input_81;
assign io_1 = input_82;
assign io_1 = input_83;
assign io_1 = input_84;
assign io_1 = input_85;
assign io_1 = input_86;
assign io_1 = input_87;
assign io_1 = input_88;
assign io_1 = input_89;
assign io_1 = input_90;
assign io_1 = input_91;
assign io_1 = input_92;
assign io_1 = input_93;
assign io_1 = input_94;
assign io_1 = input_95;
assign io_1 = input_96;
assign io_1 = input_97;
assign io_1 = input_98;
assign io_1 = input_99;
assign io_1 = input_100;
assign io_1 = input_101;
assign io_1 = input_102;
assign io_1 = input_103;
assign io_1 = input_104;
assign io_1 = input_105;
assign io_1 = input_106;
assign io_1 = input_107;
assign io_1 = input_108;
assign io_1 = input_109;
assign io_1 = input_110;
assign io_1 = input_111;
assign io_1 = input_112;
assign io_1 = input_113;
assign io_1 = input_114;
assign io_1 = input_115;
assign io_1 = input_116;
assign io_1 = input_117;
assign io_1 = input_118;
assign io_1 = input_119;
assign io_1 = input_120;
assign io_1 = input_121;
assign io_1 = input_122;
assign io_1 = input_123;
assign io_1 = input_124;
assign io_1 = input_125;
assign io_1 = input_126;
assign io_1 = input_127;
assign io_2 = input_2;
assign io_2 = input_3;
assign io_2 = input_4;
assign io_2 = input_5;
assign io_2 = input_6;
assign io_2 = input_7;
assign io_2 = input_8;
assign io_2 = input_9;
assign io_2 = input_10;
assign io_2 = input_11;
assign io_2 = input_12;
assign io_2 = input_13;
assign io_2 = input_14;
assign io_2 = input_15;
assign io_2 = input_16;
assign io_2 = input_17;
assign io_2 = input_18;
assign io_2 = input_19;
assign io_2 = input_20;
assign io_2 = input_21;
assign io_2 = input_22;
assign io_2 = input_23;
assign io_2 = input_24;
assign io_2 = input_25;
assign io_2 = input_26;
assign io_2 = input_27;
assign io_2 = input_28;
assign io_2 = input_29;
assign io_2 = input_30;
assign io_2 = input_31;
assign io_2 = input_32;
assign io_2 = input_33;
assign io_2 = input_34;
assign io_2 = input_35;
assign io_2 = input_36;
assign io_2 = input_37;
assign io_2 = input_38;
assign io_2 = input_39;
assign io_2 = input_40;
assign io_2 = input_41;
assign io_2 = input_42;
assign io_2 = input_43;
assign io_2 = input_44;
assign io_2 = input_45;
assign io_2 = input_46;
assign io_2 = input_47;
assign io_2 = input_48;
assign io_2 = input_49;
assign io_2 = input_50;
assign io_2 = input_51;
assign io_2 = input_52;
assign io_2 = input_53;
assign io_2 = input_54;
assign io_2 = input_55;
assign io_2 = input_56;
assign io_2 = input_57;
assign io_2 = input_58;
assign io_2 = input_59;
assign io_2 = input_60;
assign io_2 = input_61;
assign io_2 = input_62;
assign io_2 = input_63;
assign io_2 = input_64;
assign io_2 = input_65;
assign io_2 = input_66;
assign io_2 = input_67;
assign io_2 = input_68;
assign io_2 = input_69;
assign io_2 = input_70;
assign io_2 = input_71;
assign io_2 = input_72;
assign io_2 = input_73;
assign io_2 = input_74;
assign io_2 = input_75;
assign io_2 = input_76;
assign io_2 = input_77;
assign io_2 = input_78;
assign io_2 = input_79;
assign io_2 = input_80;
assign io_2 = input_81;
assign io_2 = input_82;
assign io_2 = input_83;
assign io_2 = input_84;
assign io_2 = input_85;
assign io_2 = input_86;
assign io_2 = input_87;
assign io_2 = input_88;
assign io_2 = input_89;
assign io_2 = input_90;
assign io_2 = input_91;
assign io_2 = input_92;
assign io_2 = input_93;
assign io_2 = input_94;
assign io_2 = input_95;
assign io_2 = input_96;
assign io_2 = input_97;
assign io_2 = input_98;
assign io_2 = input_99;
assign io_2 = input_100;
assign io_2 = input_101;
assign io_2 = input_102;
assign io_2 = input_103;
assign io_2 = input_104;
assign io_2 = input_105;
assign io_2 = input_106;
assign io_2 = input_107;
assign io_2 = input_108;
assign io_2 = input_109;
assign io_2 = input_110;
assign io_2 = input_111;
assign io_2 = input_112;
assign io_2 = input_113;
assign io_2 = input_114;
assign io_2 = input_115;
assign io_2 = input_116;
assign io_2 = input_117;
assign io_2 = input_118;
assign io_2 = input_119;
assign io_2 = input_120;
assign io_2 = input_121;
assign io_2 = input_122;
assign io_2 = input_123;
assign io_2 = input_124;
assign io_2 = input_125;
assign io_2 = input_126;
assign io_2 = input_127;
assign io_3 = input_3;
assign io_3 = input_4;
assign io_3 = input_5;
assign io_3 = input_6;
assign io_3 = input_7;
assign io_3 = input_8;
assign io_3 = input_9;
assign io_3 = input_10;
assign io_3 = input_11;
assign io_3 = input_12;
assign io_3 = input_13;
assign io_3 = input_14;
assign io_3 = input_15;
assign io_3 = input_16;
assign io_3 = input_17;
assign io_3 = input_18;
assign io_3 = input_19;
assign io_3 = input_20;
assign io_3 = input_21;
assign io_3 = input_22;
assign io_3 = input_23;
assign io_3 = input_24;
assign io_3 = input_25;
assign io_3 = input_26;
assign io_3 = input_27;
assign io_3 = input_28;
assign io_3 = input_29;
assign io_3 = input_30;
assign io_3 = input_31;
assign io_3 = input_32;
assign io_3 = input_33;
assign io_3 = input_34;
assign io_3 = input_35;
assign io_3 = input_36;
assign io_3 = input_37;
assign io_3 = input_38;
assign io_3 = input_39;
assign io_3 = input_40;
assign io_3 = input_41;
assign io_3 = input_42;
assign io_3 = input_43;
assign io_3 = input_44;
assign io_3 = input_45;
assign io_3 = input_46;
assign io_3 = input_47;
assign io_3 = input_48;
assign io_3 = input_49;
assign io_3 = input_50;
assign io_3 = input_51;
assign io_3 = input_52;
assign io_3 = input_53;
assign io_3 = input_54;
assign io_3 = input_55;
assign io_3 = input_56;
assign io_3 = input_57;
assign io_3 = input_58;
assign io_3 = input_59;
assign io_3 = input_60;
assign io_3 = input_61;
assign io_3 = input_62;
assign io_3 = input_63;
assign io_3 = input_64;
assign io_3 = input_65;
assign io_3 = input_66;
assign io_3 = input_67;
assign io_3 = input_68;
assign io_3 = input_69;
assign io_3 = input_70;
assign io_3 = input_71;
assign io_3 = input_72;
assign io_3 = input_73;
assign io_3 = input_74;
assign io_3 = input_75;
assign io_3 = input_76;
assign io_3 = input_77;
assign io_3 = input_78;
assign io_3 = input_79;
assign io_3 = input_80;
assign io_3 = input_81;
assign io_3 = input_82;
assign io_3 = input_83;
assign io_3 = input_84;
assign io_3 = input_85;
assign io_3 = input_86;
assign io_3 = input_87;
assign io_3 = input_88;
assign io_3 = input_89;
assign io_3 = input_90;
assign io_3 = input_91;
assign io_3 = input_92;
assign io_3 = input_93;
assign io_3 = input_94;
assign io_3 = input_95;
assign io_3 = input_96;
assign io_3 = input_97;
assign io_3 = input_98;
assign io_3 = input_99;
assign io_3 = input_100;
assign io_3 = input_101;
assign io_3 = input_102;
assign io_3 = input_103;
assign io_3 = input_104;
assign io_3 = input_105;
assign io_3 = input_106;
assign io_3 = input_107;
assign io_3 = input_108;
assign io_3 = input_109;
assign io_3 = input_110;
assign io_3 = input_111;
assign io_3 = input_112;
assign io_3 = input_113;
assign io_3 = input_114;
assign io_3 = input_115;
assign io_3 = input_116;
assign io_3 = input_117;
assign io_3 = input_118;
assign io_3 = input_119;
assign io_3 = input_120;
assign io_3 = input_121;
assign io_3 = input_122;
assign io_3 = input_123;
assign io_3 = input_124;
assign io_3 = input_125;
assign io_3 = input_126;
assign io_3 = input_127;
assign io_4 = input_4;
assign io_4 = input_5;
assign io_4 = input_6;
assign io_4 = input_7;
assign io_4 = input_8;
assign io_4 = input_9;
assign io_4 = input_10;
assign io_4 = input_11;
assign io_4 = input_12;
assign io_4 = input_13;
assign io_4 = input_14;
assign io_4 = input_15;
assign io_4 = input_16;
assign io_4 = input_17;
assign io_4 = input_18;
assign io_4 = input_19;
assign io_4 = input_20;
assign io_4 = input_21;
assign io_4 = input_22;
assign io_4 = input_23;
assign io_4 = input_24;
assign io_4 = input_25;
assign io_4 = input_26;
assign io_4 = input_27;
assign io_4 = input_28;
assign io_4 = input_29;
assign io_4 = input_30;
assign io_4 = input_31;
assign io_4 = input_32;
assign io_4 = input_33;
assign io_4 = input_34;
assign io_4 = input_35;
assign io_4 = input_36;
assign io_4 = input_37;
assign io_4 = input_38;
assign io_4 = input_39;
assign io_4 = input_40;
assign io_4 = input_41;
assign io_4 = input_42;
assign io_4 = input_43;
assign io_4 = input_44;
assign io_4 = input_45;
assign io_4 = input_46;
assign io_4 = input_47;
assign io_4 = input_48;
assign io_4 = input_49;
assign io_4 = input_50;
assign io_4 = input_51;
assign io_4 = input_52;
assign io_4 = input_53;
assign io_4 = input_54;
assign io_4 = input_55;
assign io_4 = input_56;
assign io_4 = input_57;
assign io_4 = input_58;
assign io_4 = input_59;
assign io_4 = input_60;
assign io_4 = input_61;
assign io_4 = input_62;
assign io_4 = input_63;
assign io_4 = input_64;
assign io_4 = input_65;
assign io_4 = input_66;
assign io_4 = input_67;
assign io_4 = input_68;
assign io_4 = input_69;
assign io_4 = input_70;
assign io_4 = input_71;
assign io_4 = input_72;
assign io_4 = input_73;
assign io_4 = input_74;
assign io_4 = input_75;
assign io_4 = input_76;
assign io_4 = input_77;
assign io_4 = input_78;
assign io_4 = input_79;
assign io_4 = input_80;
assign io_4 = input_81;
assign io_4 = input_82;
assign io_4 = input_83;
assign io_4 = input_84;
assign io_4 = input_85;
assign io_4 = input_86;
assign io_4 = input_87;
assign io_4 = input_88;
assign io_4 = input_89;
assign io_4 = input_90;
assign io_4 = input_91;
assign io_4 = input_92;
assign io_4 = input_93;
assign io_4 = input_94;
assign io_4 = input_95;
assign io_4 = input_96;
assign io_4 = input_97;
assign io_4 = input_98;
assign io_4 = input_99;
assign io_4 = input_100;
assign io_4 = input_101;
assign io_4 = input_102;
assign io_4 = input_103;
assign io_4 = input_104;
assign io_4 = input_105;
assign io_4 = input_106;
assign io_4 = input_107;
assign io_4 = input_108;
assign io_4 = input_109;
assign io_4 = input_110;
assign io_4 = input_111;
assign io_4 = input_112;
assign io_4 = input_113;
assign io_4 = input_114;
assign io_4 = input_115;
assign io_4 = input_116;
assign io_4 = input_117;
assign io_4 = input_118;
assign io_4 = input_119;
assign io_4 = input_120;
assign io_4 = input_121;
assign io_4 = input_122;
assign io_4 = input_123;
assign io_4 = input_124;
assign io_4 = input_125;
assign io_4 = input_126;
assign io_4 = input_127;
assign io_5 = input_5;
assign io_5 = input_6;
assign io_5 = input_7;
assign io_5 = input_8;
assign io_5 = input_9;
assign io_5 = input_10;
assign io_5 = input_11;
assign io_5 = input_12;
assign io_5 = input_13;
assign io_5 = input_14;
assign io_5 = input_15;
assign io_5 = input_16;
assign io_5 = input_17;
assign io_5 = input_18;
assign io_5 = input_19;
assign io_5 = input_20;
assign io_5 = input_21;
assign io_5 = input_22;
assign io_5 = input_23;
assign io_5 = input_24;
assign io_5 = input_25;
assign io_5 = input_26;
assign io_5 = input_27;
assign io_5 = input_28;
assign io_5 = input_29;
assign io_5 = input_30;
assign io_5 = input_31;
assign io_5 = input_32;
assign io_5 = input_33;
assign io_5 = input_34;
assign io_5 = input_35;
assign io_5 = input_36;
assign io_5 = input_37;
assign io_5 = input_38;
assign io_5 = input_39;
assign io_5 = input_40;
assign io_5 = input_41;
assign io_5 = input_42;
assign io_5 = input_43;
assign io_5 = input_44;
assign io_5 = input_45;
assign io_5 = input_46;
assign io_5 = input_47;
assign io_5 = input_48;
assign io_5 = input_49;
assign io_5 = input_50;
assign io_5 = input_51;
assign io_5 = input_52;
assign io_5 = input_53;
assign io_5 = input_54;
assign io_5 = input_55;
assign io_5 = input_56;
assign io_5 = input_57;
assign io_5 = input_58;
assign io_5 = input_59;
assign io_5 = input_60;
assign io_5 = input_61;
assign io_5 = input_62;
assign io_5 = input_63;
assign io_5 = input_64;
assign io_5 = input_65;
assign io_5 = input_66;
assign io_5 = input_67;
assign io_5 = input_68;
assign io_5 = input_69;
assign io_5 = input_70;
assign io_5 = input_71;
assign io_5 = input_72;
assign io_5 = input_73;
assign io_5 = input_74;
assign io_5 = input_75;
assign io_5 = input_76;
assign io_5 = input_77;
assign io_5 = input_78;
assign io_5 = input_79;
assign io_5 = input_80;
assign io_5 = input_81;
assign io_5 = input_82;
assign io_5 = input_83;
assign io_5 = input_84;
assign io_5 = input_85;
assign io_5 = input_86;
assign io_5 = input_87;
assign io_5 = input_88;
assign io_5 = input_89;
assign io_5 = input_90;
assign io_5 = input_91;
assign io_5 = input_92;
assign io_5 = input_93;
assign io_5 = input_94;
assign io_5 = input_95;
assign io_5 = input_96;
assign io_5 = input_97;
assign io_5 = input_98;
assign io_5 = input_99;
assign io_5 = input_100;
assign io_5 = input_101;
assign io_5 = input_102;
assign io_5 = input_103;
assign io_5 = input_104;
assign io_5 = input_105;
assign io_5 = input_106;
assign io_5 = input_107;
assign io_5 = input_108;
assign io_5 = input_109;
assign io_5 = input_110;
assign io_5 = input_111;
assign io_5 = input_112;
assign io_5 = input_113;
assign io_5 = input_114;
assign io_5 = input_115;
assign io_5 = input_116;
assign io_5 = input_117;
assign io_5 = input_118;
assign io_5 = input_119;
assign io_5 = input_120;
assign io_5 = input_121;
assign io_5 = input_122;
assign io_5 = input_123;
assign io_5 = input_124;
assign io_5 = input_125;
assign io_5 = input_126;
assign io_5 = input_127;
assign io_6 = input_6;
assign io_6 = input_7;
assign io_6 = input_8;
assign io_6 = input_9;
assign io_6 = input_10;
assign io_6 = input_11;
assign io_6 = input_12;
assign io_6 = input_13;
assign io_6 = input_14;
assign io_6 = input_15;
assign io_6 = input_16;
assign io_6 = input_17;
assign io_6 = input_18;
assign io_6 = input_19;
assign io_6 = input_20;
assign io_6 = input_21;
assign io_6 = input_22;
assign io_6 = input_23;
assign io_6 = input_24;
assign io_6 = input_25;
assign io_6 = input_26;
assign io_6 = input_27;
assign io_6 = input_28;
assign io_6 = input_29;
assign io_6 = input_30;
assign io_6 = input_31;
assign io_6 = input_32;
assign io_6 = input_33;
assign io_6 = input_34;
assign io_6 = input_35;
assign io_6 = input_36;
assign io_6 = input_37;
assign io_6 = input_38;
assign io_6 = input_39;
assign io_6 = input_40;
assign io_6 = input_41;
assign io_6 = input_42;
assign io_6 = input_43;
assign io_6 = input_44;
assign io_6 = input_45;
assign io_6 = input_46;
assign io_6 = input_47;
assign io_6 = input_48;
assign io_6 = input_49;
assign io_6 = input_50;
assign io_6 = input_51;
assign io_6 = input_52;
assign io_6 = input_53;
assign io_6 = input_54;
assign io_6 = input_55;
assign io_6 = input_56;
assign io_6 = input_57;
assign io_6 = input_58;
assign io_6 = input_59;
assign io_6 = input_60;
assign io_6 = input_61;
assign io_6 = input_62;
assign io_6 = input_63;
assign io_6 = input_64;
assign io_6 = input_65;
assign io_6 = input_66;
assign io_6 = input_67;
assign io_6 = input_68;
assign io_6 = input_69;
assign io_6 = input_70;
assign io_6 = input_71;
assign io_6 = input_72;
assign io_6 = input_73;
assign io_6 = input_74;
assign io_6 = input_75;
assign io_6 = input_76;
assign io_6 = input_77;
assign io_6 = input_78;
assign io_6 = input_79;
assign io_6 = input_80;
assign io_6 = input_81;
assign io_6 = input_82;
assign io_6 = input_83;
assign io_6 = input_84;
assign io_6 = input_85;
assign io_6 = input_86;
assign io_6 = input_87;
assign io_6 = input_88;
assign io_6 = input_89;
assign io_6 = input_90;
assign io_6 = input_91;
assign io_6 = input_92;
assign io_6 = input_93;
assign io_6 = input_94;
assign io_6 = input_95;
assign io_6 = input_96;
assign io_6 = input_97;
assign io_6 = input_98;
assign io_6 = input_99;
assign io_6 = input_100;
assign io_6 = input_101;
assign io_6 = input_102;
assign io_6 = input_103;
assign io_6 = input_104;
assign io_6 = input_105;
assign io_6 = input_106;
assign io_6 = input_107;
assign io_6 = input_108;
assign io_6 = input_109;
assign io_6 = input_110;
assign io_6 = input_111;
assign io_6 = input_112;
assign io_6 = input_113;
assign io_6 = input_114;
assign io_6 = input_115;
assign io_6 = input_116;
assign io_6 = input_117;
assign io_6 = input_118;
assign io_6 = input_119;
assign io_6 = input_120;
assign io_6 = input_121;
assign io_6 = input_122;
assign io_6 = input_123;
assign io_6 = input_124;
assign io_6 = input_125;
assign io_6 = input_126;
assign io_6 = input_127;
assign io_7 = input_7;
assign io_7 = input_8;
assign io_7 = input_9;
assign io_7 = input_10;
assign io_7 = input_11;
assign io_7 = input_12;
assign io_7 = input_13;
assign io_7 = input_14;
assign io_7 = input_15;
assign io_7 = input_16;
assign io_7 = input_17;
assign io_7 = input_18;
assign io_7 = input_19;
assign io_7 = input_20;
assign io_7 = input_21;
assign io_7 = input_22;
assign io_7 = input_23;
assign io_7 = input_24;
assign io_7 = input_25;
assign io_7 = input_26;
assign io_7 = input_27;
assign io_7 = input_28;
assign io_7 = input_29;
assign io_7 = input_30;
assign io_7 = input_31;
assign io_7 = input_32;
assign io_7 = input_33;
assign io_7 = input_34;
assign io_7 = input_35;
assign io_7 = input_36;
assign io_7 = input_37;
assign io_7 = input_38;
assign io_7 = input_39;
assign io_7 = input_40;
assign io_7 = input_41;
assign io_7 = input_42;
assign io_7 = input_43;
assign io_7 = input_44;
assign io_7 = input_45;
assign io_7 = input_46;
assign io_7 = input_47;
assign io_7 = input_48;
assign io_7 = input_49;
assign io_7 = input_50;
assign io_7 = input_51;
assign io_7 = input_52;
assign io_7 = input_53;
assign io_7 = input_54;
assign io_7 = input_55;
assign io_7 = input_56;
assign io_7 = input_57;
assign io_7 = input_58;
assign io_7 = input_59;
assign io_7 = input_60;
assign io_7 = input_61;
assign io_7 = input_62;
assign io_7 = input_63;
assign io_7 = input_64;
assign io_7 = input_65;
assign io_7 = input_66;
assign io_7 = input_67;
assign io_7 = input_68;
assign io_7 = input_69;
assign io_7 = input_70;
assign io_7 = input_71;
assign io_7 = input_72;
assign io_7 = input_73;
assign io_7 = input_74;
assign io_7 = input_75;
assign io_7 = input_76;
assign io_7 = input_77;
assign io_7 = input_78;
assign io_7 = input_79;
assign io_7 = input_80;
assign io_7 = input_81;
assign io_7 = input_82;
assign io_7 = input_83;
assign io_7 = input_84;
assign io_7 = input_85;
assign io_7 = input_86;
assign io_7 = input_87;
assign io_7 = input_88;
assign io_7 = input_89;
assign io_7 = input_90;
assign io_7 = input_91;
assign io_7 = input_92;
assign io_7 = input_93;
assign io_7 = input_94;
assign io_7 = input_95;
assign io_7 = input_96;
assign io_7 = input_97;
assign io_7 = input_98;
assign io_7 = input_99;
assign io_7 = input_100;
assign io_7 = input_101;
assign io_7 = input_102;
assign io_7 = input_103;
assign io_7 = input_104;
assign io_7 = input_105;
assign io_7 = input_106;
assign io_7 = input_107;
assign io_7 = input_108;
assign io_7 = input_109;
assign io_7 = input_110;
assign io_7 = input_111;
assign io_7 = input_112;
assign io_7 = input_113;
assign io_7 = input_114;
assign io_7 = input_115;
assign io_7 = input_116;
assign io_7 = input_117;
assign io_7 = input_118;
assign io_7 = input_119;
assign io_7 = input_120;
assign io_7 = input_121;
assign io_7 = input_122;
assign io_7 = input_123;
assign io_7 = input_124;
assign io_7 = input_125;
assign io_7 = input_126;
assign io_7 = input_127;
assign io_8 = input_8;
assign io_8 = input_9;
assign io_8 = input_10;
assign io_8 = input_11;
assign io_8 = input_12;
assign io_8 = input_13;
assign io_8 = input_14;
assign io_8 = input_15;
assign io_8 = input_16;
assign io_8 = input_17;
assign io_8 = input_18;
assign io_8 = input_19;
assign io_8 = input_20;
assign io_8 = input_21;
assign io_8 = input_22;
assign io_8 = input_23;
assign io_8 = input_24;
assign io_8 = input_25;
assign io_8 = input_26;
assign io_8 = input_27;
assign io_8 = input_28;
assign io_8 = input_29;
assign io_8 = input_30;
assign io_8 = input_31;
assign io_8 = input_32;
assign io_8 = input_33;
assign io_8 = input_34;
assign io_8 = input_35;
assign io_8 = input_36;
assign io_8 = input_37;
assign io_8 = input_38;
assign io_8 = input_39;
assign io_8 = input_40;
assign io_8 = input_41;
assign io_8 = input_42;
assign io_8 = input_43;
assign io_8 = input_44;
assign io_8 = input_45;
assign io_8 = input_46;
assign io_8 = input_47;
assign io_8 = input_48;
assign io_8 = input_49;
assign io_8 = input_50;
assign io_8 = input_51;
assign io_8 = input_52;
assign io_8 = input_53;
assign io_8 = input_54;
assign io_8 = input_55;
assign io_8 = input_56;
assign io_8 = input_57;
assign io_8 = input_58;
assign io_8 = input_59;
assign io_8 = input_60;
assign io_8 = input_61;
assign io_8 = input_62;
assign io_8 = input_63;
assign io_8 = input_64;
assign io_8 = input_65;
assign io_8 = input_66;
assign io_8 = input_67;
assign io_8 = input_68;
assign io_8 = input_69;
assign io_8 = input_70;
assign io_8 = input_71;
assign io_8 = input_72;
assign io_8 = input_73;
assign io_8 = input_74;
assign io_8 = input_75;
assign io_8 = input_76;
assign io_8 = input_77;
assign io_8 = input_78;
assign io_8 = input_79;
assign io_8 = input_80;
assign io_8 = input_81;
assign io_8 = input_82;
assign io_8 = input_83;
assign io_8 = input_84;
assign io_8 = input_85;
assign io_8 = input_86;
assign io_8 = input_87;
assign io_8 = input_88;
assign io_8 = input_89;
assign io_8 = input_90;
assign io_8 = input_91;
assign io_8 = input_92;
assign io_8 = input_93;
assign io_8 = input_94;
assign io_8 = input_95;
assign io_8 = input_96;
assign io_8 = input_97;
assign io_8 = input_98;
assign io_8 = input_99;
assign io_8 = input_100;
assign io_8 = input_101;
assign io_8 = input_102;
assign io_8 = input_103;
assign io_8 = input_104;
assign io_8 = input_105;
assign io_8 = input_106;
assign io_8 = input_107;
assign io_8 = input_108;
assign io_8 = input_109;
assign io_8 = input_110;
assign io_8 = input_111;
assign io_8 = input_112;
assign io_8 = input_113;
assign io_8 = input_114;
assign io_8 = input_115;
assign io_8 = input_116;
assign io_8 = input_117;
assign io_8 = input_118;
assign io_8 = input_119;
assign io_8 = input_120;
assign io_8 = input_121;
assign io_8 = input_122;
assign io_8 = input_123;
assign io_8 = input_124;
assign io_8 = input_125;
assign io_8 = input_126;
assign io_8 = input_127;
assign io_9 = input_9;
assign io_9 = input_10;
assign io_9 = input_11;
assign io_9 = input_12;
assign io_9 = input_13;
assign io_9 = input_14;
assign io_9 = input_15;
assign io_9 = input_16;
assign io_9 = input_17;
assign io_9 = input_18;
assign io_9 = input_19;
assign io_9 = input_20;
assign io_9 = input_21;
assign io_9 = input_22;
assign io_9 = input_23;
assign io_9 = input_24;
assign io_9 = input_25;
assign io_9 = input_26;
assign io_9 = input_27;
assign io_9 = input_28;
assign io_9 = input_29;
assign io_9 = input_30;
assign io_9 = input_31;
assign io_9 = input_32;
assign io_9 = input_33;
assign io_9 = input_34;
assign io_9 = input_35;
assign io_9 = input_36;
assign io_9 = input_37;
assign io_9 = input_38;
assign io_9 = input_39;
assign io_9 = input_40;
assign io_9 = input_41;
assign io_9 = input_42;
assign io_9 = input_43;
assign io_9 = input_44;
assign io_9 = input_45;
assign io_9 = input_46;
assign io_9 = input_47;
assign io_9 = input_48;
assign io_9 = input_49;
assign io_9 = input_50;
assign io_9 = input_51;
assign io_9 = input_52;
assign io_9 = input_53;
assign io_9 = input_54;
assign io_9 = input_55;
assign io_9 = input_56;
assign io_9 = input_57;
assign io_9 = input_58;
assign io_9 = input_59;
assign io_9 = input_60;
assign io_9 = input_61;
assign io_9 = input_62;
assign io_9 = input_63;
assign io_9 = input_64;
assign io_9 = input_65;
assign io_9 = input_66;
assign io_9 = input_67;
assign io_9 = input_68;
assign io_9 = input_69;
assign io_9 = input_70;
assign io_9 = input_71;
assign io_9 = input_72;
assign io_9 = input_73;
assign io_9 = input_74;
assign io_9 = input_75;
assign io_9 = input_76;
assign io_9 = input_77;
assign io_9 = input_78;
assign io_9 = input_79;
assign io_9 = input_80;
assign io_9 = input_81;
assign io_9 = input_82;
assign io_9 = input_83;
assign io_9 = input_84;
assign io_9 = input_85;
assign io_9 = input_86;
assign io_9 = input_87;
assign io_9 = input_88;
assign io_9 = input_89;
assign io_9 = input_90;
assign io_9 = input_91;
assign io_9 = input_92;
assign io_9 = input_93;
assign io_9 = input_94;
assign io_9 = input_95;
assign io_9 = input_96;
assign io_9 = input_97;
assign io_9 = input_98;
assign io_9 = input_99;
assign io_9 = input_100;
assign io_9 = input_101;
assign io_9 = input_102;
assign io_9 = input_103;
assign io_9 = input_104;
assign io_9 = input_105;
assign io_9 = input_106;
assign io_9 = input_107;
assign io_9 = input_108;
assign io_9 = input_109;
assign io_9 = input_110;
assign io_9 = input_111;
assign io_9 = input_112;
assign io_9 = input_113;
assign io_9 = input_114;
assign io_9 = input_115;
assign io_9 = input_116;
assign io_9 = input_117;
assign io_9 = input_118;
assign io_9 = input_119;
assign io_9 = input_120;
assign io_9 = input_121;
assign io_9 = input_122;
assign io_9 = input_123;
assign io_9 = input_124;
assign io_9 = input_125;
assign io_9 = input_126;
assign io_9 = input_127;
assign io_10 = input_10;
assign io_10 = input_11;
assign io_10 = input_12;
assign io_10 = input_13;
assign io_10 = input_14;
assign io_10 = input_15;
assign io_10 = input_16;
assign io_10 = input_17;
assign io_10 = input_18;
assign io_10 = input_19;
assign io_10 = input_20;
assign io_10 = input_21;
assign io_10 = input_22;
assign io_10 = input_23;
assign io_10 = input_24;
assign io_10 = input_25;
assign io_10 = input_26;
assign io_10 = input_27;
assign io_10 = input_28;
assign io_10 = input_29;
assign io_10 = input_30;
assign io_10 = input_31;
assign io_10 = input_32;
assign io_10 = input_33;
assign io_10 = input_34;
assign io_10 = input_35;
assign io_10 = input_36;
assign io_10 = input_37;
assign io_10 = input_38;
assign io_10 = input_39;
assign io_10 = input_40;
assign io_10 = input_41;
assign io_10 = input_42;
assign io_10 = input_43;
assign io_10 = input_44;
assign io_10 = input_45;
assign io_10 = input_46;
assign io_10 = input_47;
assign io_10 = input_48;
assign io_10 = input_49;
assign io_10 = input_50;
assign io_10 = input_51;
assign io_10 = input_52;
assign io_10 = input_53;
assign io_10 = input_54;
assign io_10 = input_55;
assign io_10 = input_56;
assign io_10 = input_57;
assign io_10 = input_58;
assign io_10 = input_59;
assign io_10 = input_60;
assign io_10 = input_61;
assign io_10 = input_62;
assign io_10 = input_63;
assign io_10 = input_64;
assign io_10 = input_65;
assign io_10 = input_66;
assign io_10 = input_67;
assign io_10 = input_68;
assign io_10 = input_69;
assign io_10 = input_70;
assign io_10 = input_71;
assign io_10 = input_72;
assign io_10 = input_73;
assign io_10 = input_74;
assign io_10 = input_75;
assign io_10 = input_76;
assign io_10 = input_77;
assign io_10 = input_78;
assign io_10 = input_79;
assign io_10 = input_80;
assign io_10 = input_81;
assign io_10 = input_82;
assign io_10 = input_83;
assign io_10 = input_84;
assign io_10 = input_85;
assign io_10 = input_86;
assign io_10 = input_87;
assign io_10 = input_88;
assign io_10 = input_89;
assign io_10 = input_90;
assign io_10 = input_91;
assign io_10 = input_92;
assign io_10 = input_93;
assign io_10 = input_94;
assign io_10 = input_95;
assign io_10 = input_96;
assign io_10 = input_97;
assign io_10 = input_98;
assign io_10 = input_99;
assign io_10 = input_100;
assign io_10 = input_101;
assign io_10 = input_102;
assign io_10 = input_103;
assign io_10 = input_104;
assign io_10 = input_105;
assign io_10 = input_106;
assign io_10 = input_107;
assign io_10 = input_108;
assign io_10 = input_109;
assign io_10 = input_110;
assign io_10 = input_111;
assign io_10 = input_112;
assign io_10 = input_113;
assign io_10 = input_114;
assign io_10 = input_115;
assign io_10 = input_116;
assign io_10 = input_117;
assign io_10 = input_118;
assign io_10 = input_119;
assign io_10 = input_120;
assign io_10 = input_121;
assign io_10 = input_122;
assign io_10 = input_123;
assign io_10 = input_124;
assign io_10 = input_125;
assign io_10 = input_126;
assign io_10 = input_127;
assign io_11 = input_11;
assign io_11 = input_12;
assign io_11 = input_13;
assign io_11 = input_14;
assign io_11 = input_15;
assign io_11 = input_16;
assign io_11 = input_17;
assign io_11 = input_18;
assign io_11 = input_19;
assign io_11 = input_20;
assign io_11 = input_21;
assign io_11 = input_22;
assign io_11 = input_23;
assign io_11 = input_24;
assign io_11 = input_25;
assign io_11 = input_26;
assign io_11 = input_27;
assign io_11 = input_28;
assign io_11 = input_29;
assign io_11 = input_30;
assign io_11 = input_31;
assign io_11 = input_32;
assign io_11 = input_33;
assign io_11 = input_34;
assign io_11 = input_35;
assign io_11 = input_36;
assign io_11 = input_37;
assign io_11 = input_38;
assign io_11 = input_39;
assign io_11 = input_40;
assign io_11 = input_41;
assign io_11 = input_42;
assign io_11 = input_43;
assign io_11 = input_44;
assign io_11 = input_45;
assign io_11 = input_46;
assign io_11 = input_47;
assign io_11 = input_48;
assign io_11 = input_49;
assign io_11 = input_50;
assign io_11 = input_51;
assign io_11 = input_52;
assign io_11 = input_53;
assign io_11 = input_54;
assign io_11 = input_55;
assign io_11 = input_56;
assign io_11 = input_57;
assign io_11 = input_58;
assign io_11 = input_59;
assign io_11 = input_60;
assign io_11 = input_61;
assign io_11 = input_62;
assign io_11 = input_63;
assign io_11 = input_64;
assign io_11 = input_65;
assign io_11 = input_66;
assign io_11 = input_67;
assign io_11 = input_68;
assign io_11 = input_69;
assign io_11 = input_70;
assign io_11 = input_71;
assign io_11 = input_72;
assign io_11 = input_73;
assign io_11 = input_74;
assign io_11 = input_75;
assign io_11 = input_76;
assign io_11 = input_77;
assign io_11 = input_78;
assign io_11 = input_79;
assign io_11 = input_80;
assign io_11 = input_81;
assign io_11 = input_82;
assign io_11 = input_83;
assign io_11 = input_84;
assign io_11 = input_85;
assign io_11 = input_86;
assign io_11 = input_87;
assign io_11 = input_88;
assign io_11 = input_89;
assign io_11 = input_90;
assign io_11 = input_91;
assign io_11 = input_92;
assign io_11 = input_93;
assign io_11 = input_94;
assign io_11 = input_95;
assign io_11 = input_96;
assign io_11 = input_97;
assign io_11 = input_98;
assign io_11 = input_99;
assign io_11 = input_100;
assign io_11 = input_101;
assign io_11 = input_102;
assign io_11 = input_103;
assign io_11 = input_104;
assign io_11 = input_105;
assign io_11 = input_106;
assign io_11 = input_107;
assign io_11 = input_108;
assign io_11 = input_109;
assign io_11 = input_110;
assign io_11 = input_111;
assign io_11 = input_112;
assign io_11 = input_113;
assign io_11 = input_114;
assign io_11 = input_115;
assign io_11 = input_116;
assign io_11 = input_117;
assign io_11 = input_118;
assign io_11 = input_119;
assign io_11 = input_120;
assign io_11 = input_121;
assign io_11 = input_122;
assign io_11 = input_123;
assign io_11 = input_124;
assign io_11 = input_125;
assign io_11 = input_126;
assign io_11 = input_127;
assign io_12 = input_12;
assign io_12 = input_13;
assign io_12 = input_14;
assign io_12 = input_15;
assign io_12 = input_16;
assign io_12 = input_17;
assign io_12 = input_18;
assign io_12 = input_19;
assign io_12 = input_20;
assign io_12 = input_21;
assign io_12 = input_22;
assign io_12 = input_23;
assign io_12 = input_24;
assign io_12 = input_25;
assign io_12 = input_26;
assign io_12 = input_27;
assign io_12 = input_28;
assign io_12 = input_29;
assign io_12 = input_30;
assign io_12 = input_31;
assign io_12 = input_32;
assign io_12 = input_33;
assign io_12 = input_34;
assign io_12 = input_35;
assign io_12 = input_36;
assign io_12 = input_37;
assign io_12 = input_38;
assign io_12 = input_39;
assign io_12 = input_40;
assign io_12 = input_41;
assign io_12 = input_42;
assign io_12 = input_43;
assign io_12 = input_44;
assign io_12 = input_45;
assign io_12 = input_46;
assign io_12 = input_47;
assign io_12 = input_48;
assign io_12 = input_49;
assign io_12 = input_50;
assign io_12 = input_51;
assign io_12 = input_52;
assign io_12 = input_53;
assign io_12 = input_54;
assign io_12 = input_55;
assign io_12 = input_56;
assign io_12 = input_57;
assign io_12 = input_58;
assign io_12 = input_59;
assign io_12 = input_60;
assign io_12 = input_61;
assign io_12 = input_62;
assign io_12 = input_63;
assign io_12 = input_64;
assign io_12 = input_65;
assign io_12 = input_66;
assign io_12 = input_67;
assign io_12 = input_68;
assign io_12 = input_69;
assign io_12 = input_70;
assign io_12 = input_71;
assign io_12 = input_72;
assign io_12 = input_73;
assign io_12 = input_74;
assign io_12 = input_75;
assign io_12 = input_76;
assign io_12 = input_77;
assign io_12 = input_78;
assign io_12 = input_79;
assign io_12 = input_80;
assign io_12 = input_81;
assign io_12 = input_82;
assign io_12 = input_83;
assign io_12 = input_84;
assign io_12 = input_85;
assign io_12 = input_86;
assign io_12 = input_87;
assign io_12 = input_88;
assign io_12 = input_89;
assign io_12 = input_90;
assign io_12 = input_91;
assign io_12 = input_92;
assign io_12 = input_93;
assign io_12 = input_94;
assign io_12 = input_95;
assign io_12 = input_96;
assign io_12 = input_97;
assign io_12 = input_98;
assign io_12 = input_99;
assign io_12 = input_100;
assign io_12 = input_101;
assign io_12 = input_102;
assign io_12 = input_103;
assign io_12 = input_104;
assign io_12 = input_105;
assign io_12 = input_106;
assign io_12 = input_107;
assign io_12 = input_108;
assign io_12 = input_109;
assign io_12 = input_110;
assign io_12 = input_111;
assign io_12 = input_112;
assign io_12 = input_113;
assign io_12 = input_114;
assign io_12 = input_115;
assign io_12 = input_116;
assign io_12 = input_117;
assign io_12 = input_118;
assign io_12 = input_119;
assign io_12 = input_120;
assign io_12 = input_121;
assign io_12 = input_122;
assign io_12 = input_123;
assign io_12 = input_124;
assign io_12 = input_125;
assign io_12 = input_126;
assign io_12 = input_127;
assign io_13 = input_13;
assign io_13 = input_14;
assign io_13 = input_15;
assign io_13 = input_16;
assign io_13 = input_17;
assign io_13 = input_18;
assign io_13 = input_19;
assign io_13 = input_20;
assign io_13 = input_21;
assign io_13 = input_22;
assign io_13 = input_23;
assign io_13 = input_24;
assign io_13 = input_25;
assign io_13 = input_26;
assign io_13 = input_27;
assign io_13 = input_28;
assign io_13 = input_29;
assign io_13 = input_30;
assign io_13 = input_31;
assign io_13 = input_32;
assign io_13 = input_33;
assign io_13 = input_34;
assign io_13 = input_35;
assign io_13 = input_36;
assign io_13 = input_37;
assign io_13 = input_38;
assign io_13 = input_39;
assign io_13 = input_40;
assign io_13 = input_41;
assign io_13 = input_42;
assign io_13 = input_43;
assign io_13 = input_44;
assign io_13 = input_45;
assign io_13 = input_46;
assign io_13 = input_47;
assign io_13 = input_48;
assign io_13 = input_49;
assign io_13 = input_50;
assign io_13 = input_51;
assign io_13 = input_52;
assign io_13 = input_53;
assign io_13 = input_54;
assign io_13 = input_55;
assign io_13 = input_56;
assign io_13 = input_57;
assign io_13 = input_58;
assign io_13 = input_59;
assign io_13 = input_60;
assign io_13 = input_61;
assign io_13 = input_62;
assign io_13 = input_63;
assign io_13 = input_64;
assign io_13 = input_65;
assign io_13 = input_66;
assign io_13 = input_67;
assign io_13 = input_68;
assign io_13 = input_69;
assign io_13 = input_70;
assign io_13 = input_71;
assign io_13 = input_72;
assign io_13 = input_73;
assign io_13 = input_74;
assign io_13 = input_75;
assign io_13 = input_76;
assign io_13 = input_77;
assign io_13 = input_78;
assign io_13 = input_79;
assign io_13 = input_80;
assign io_13 = input_81;
assign io_13 = input_82;
assign io_13 = input_83;
assign io_13 = input_84;
assign io_13 = input_85;
assign io_13 = input_86;
assign io_13 = input_87;
assign io_13 = input_88;
assign io_13 = input_89;
assign io_13 = input_90;
assign io_13 = input_91;
assign io_13 = input_92;
assign io_13 = input_93;
assign io_13 = input_94;
assign io_13 = input_95;
assign io_13 = input_96;
assign io_13 = input_97;
assign io_13 = input_98;
assign io_13 = input_99;
assign io_13 = input_100;
assign io_13 = input_101;
assign io_13 = input_102;
assign io_13 = input_103;
assign io_13 = input_104;
assign io_13 = input_105;
assign io_13 = input_106;
assign io_13 = input_107;
assign io_13 = input_108;
assign io_13 = input_109;
assign io_13 = input_110;
assign io_13 = input_111;
assign io_13 = input_112;
assign io_13 = input_113;
assign io_13 = input_114;
assign io_13 = input_115;
assign io_13 = input_116;
assign io_13 = input_117;
assign io_13 = input_118;
assign io_13 = input_119;
assign io_13 = input_120;
assign io_13 = input_121;
assign io_13 = input_122;
assign io_13 = input_123;
assign io_13 = input_124;
assign io_13 = input_125;
assign io_13 = input_126;
assign io_13 = input_127;
assign io_14 = input_14;
assign io_14 = input_15;
assign io_14 = input_16;
assign io_14 = input_17;
assign io_14 = input_18;
assign io_14 = input_19;
assign io_14 = input_20;
assign io_14 = input_21;
assign io_14 = input_22;
assign io_14 = input_23;
assign io_14 = input_24;
assign io_14 = input_25;
assign io_14 = input_26;
assign io_14 = input_27;
assign io_14 = input_28;
assign io_14 = input_29;
assign io_14 = input_30;
assign io_14 = input_31;
assign io_14 = input_32;
assign io_14 = input_33;
assign io_14 = input_34;
assign io_14 = input_35;
assign io_14 = input_36;
assign io_14 = input_37;
assign io_14 = input_38;
assign io_14 = input_39;
assign io_14 = input_40;
assign io_14 = input_41;
assign io_14 = input_42;
assign io_14 = input_43;
assign io_14 = input_44;
assign io_14 = input_45;
assign io_14 = input_46;
assign io_14 = input_47;
assign io_14 = input_48;
assign io_14 = input_49;
assign io_14 = input_50;
assign io_14 = input_51;
assign io_14 = input_52;
assign io_14 = input_53;
assign io_14 = input_54;
assign io_14 = input_55;
assign io_14 = input_56;
assign io_14 = input_57;
assign io_14 = input_58;
assign io_14 = input_59;
assign io_14 = input_60;
assign io_14 = input_61;
assign io_14 = input_62;
assign io_14 = input_63;
assign io_14 = input_64;
assign io_14 = input_65;
assign io_14 = input_66;
assign io_14 = input_67;
assign io_14 = input_68;
assign io_14 = input_69;
assign io_14 = input_70;
assign io_14 = input_71;
assign io_14 = input_72;
assign io_14 = input_73;
assign io_14 = input_74;
assign io_14 = input_75;
assign io_14 = input_76;
assign io_14 = input_77;
assign io_14 = input_78;
assign io_14 = input_79;
assign io_14 = input_80;
assign io_14 = input_81;
assign io_14 = input_82;
assign io_14 = input_83;
assign io_14 = input_84;
assign io_14 = input_85;
assign io_14 = input_86;
assign io_14 = input_87;
assign io_14 = input_88;
assign io_14 = input_89;
assign io_14 = input_90;
assign io_14 = input_91;
assign io_14 = input_92;
assign io_14 = input_93;
assign io_14 = input_94;
assign io_14 = input_95;
assign io_14 = input_96;
assign io_14 = input_97;
assign io_14 = input_98;
assign io_14 = input_99;
assign io_14 = input_100;
assign io_14 = input_101;
assign io_14 = input_102;
assign io_14 = input_103;
assign io_14 = input_104;
assign io_14 = input_105;
assign io_14 = input_106;
assign io_14 = input_107;
assign io_14 = input_108;
assign io_14 = input_109;
assign io_14 = input_110;
assign io_14 = input_111;
assign io_14 = input_112;
assign io_14 = input_113;
assign io_14 = input_114;
assign io_14 = input_115;
assign io_14 = input_116;
assign io_14 = input_117;
assign io_14 = input_118;
assign io_14 = input_119;
assign io_14 = input_120;
assign io_14 = input_121;
assign io_14 = input_122;
assign io_14 = input_123;
assign io_14 = input_124;
assign io_14 = input_125;
assign io_14 = input_126;
assign io_14 = input_127;
assign io_15 = input_15;
assign io_15 = input_16;
assign io_15 = input_17;
assign io_15 = input_18;
assign io_15 = input_19;
assign io_15 = input_20;
assign io_15 = input_21;
assign io_15 = input_22;
assign io_15 = input_23;
assign io_15 = input_24;
assign io_15 = input_25;
assign io_15 = input_26;
assign io_15 = input_27;
assign io_15 = input_28;
assign io_15 = input_29;
assign io_15 = input_30;
assign io_15 = input_31;
assign io_15 = input_32;
assign io_15 = input_33;
assign io_15 = input_34;
assign io_15 = input_35;
assign io_15 = input_36;
assign io_15 = input_37;
assign io_15 = input_38;
assign io_15 = input_39;
assign io_15 = input_40;
assign io_15 = input_41;
assign io_15 = input_42;
assign io_15 = input_43;
assign io_15 = input_44;
assign io_15 = input_45;
assign io_15 = input_46;
assign io_15 = input_47;
assign io_15 = input_48;
assign io_15 = input_49;
assign io_15 = input_50;
assign io_15 = input_51;
assign io_15 = input_52;
assign io_15 = input_53;
assign io_15 = input_54;
assign io_15 = input_55;
assign io_15 = input_56;
assign io_15 = input_57;
assign io_15 = input_58;
assign io_15 = input_59;
assign io_15 = input_60;
assign io_15 = input_61;
assign io_15 = input_62;
assign io_15 = input_63;
assign io_15 = input_64;
assign io_15 = input_65;
assign io_15 = input_66;
assign io_15 = input_67;
assign io_15 = input_68;
assign io_15 = input_69;
assign io_15 = input_70;
assign io_15 = input_71;
assign io_15 = input_72;
assign io_15 = input_73;
assign io_15 = input_74;
assign io_15 = input_75;
assign io_15 = input_76;
assign io_15 = input_77;
assign io_15 = input_78;
assign io_15 = input_79;
assign io_15 = input_80;
assign io_15 = input_81;
assign io_15 = input_82;
assign io_15 = input_83;
assign io_15 = input_84;
assign io_15 = input_85;
assign io_15 = input_86;
assign io_15 = input_87;
assign io_15 = input_88;
assign io_15 = input_89;
assign io_15 = input_90;
assign io_15 = input_91;
assign io_15 = input_92;
assign io_15 = input_93;
assign io_15 = input_94;
assign io_15 = input_95;
assign io_15 = input_96;
assign io_15 = input_97;
assign io_15 = input_98;
assign io_15 = input_99;
assign io_15 = input_100;
assign io_15 = input_101;
assign io_15 = input_102;
assign io_15 = input_103;
assign io_15 = input_104;
assign io_15 = input_105;
assign io_15 = input_106;
assign io_15 = input_107;
assign io_15 = input_108;
assign io_15 = input_109;
assign io_15 = input_110;
assign io_15 = input_111;
assign io_15 = input_112;
assign io_15 = input_113;
assign io_15 = input_114;
assign io_15 = input_115;
assign io_15 = input_116;
assign io_15 = input_117;
assign io_15 = input_118;
assign io_15 = input_119;
assign io_15 = input_120;
assign io_15 = input_121;
assign io_15 = input_122;
assign io_15 = input_123;
assign io_15 = input_124;
assign io_15 = input_125;
assign io_15 = input_126;
assign io_15 = input_127;
assign io_16 = input_16;
assign io_16 = input_17;
assign io_16 = input_18;
assign io_16 = input_19;
assign io_16 = input_20;
assign io_16 = input_21;
assign io_16 = input_22;
assign io_16 = input_23;
assign io_16 = input_24;
assign io_16 = input_25;
assign io_16 = input_26;
assign io_16 = input_27;
assign io_16 = input_28;
assign io_16 = input_29;
assign io_16 = input_30;
assign io_16 = input_31;
assign io_16 = input_32;
assign io_16 = input_33;
assign io_16 = input_34;
assign io_16 = input_35;
assign io_16 = input_36;
assign io_16 = input_37;
assign io_16 = input_38;
assign io_16 = input_39;
assign io_16 = input_40;
assign io_16 = input_41;
assign io_16 = input_42;
assign io_16 = input_43;
assign io_16 = input_44;
assign io_16 = input_45;
assign io_16 = input_46;
assign io_16 = input_47;
assign io_16 = input_48;
assign io_16 = input_49;
assign io_16 = input_50;
assign io_16 = input_51;
assign io_16 = input_52;
assign io_16 = input_53;
assign io_16 = input_54;
assign io_16 = input_55;
assign io_16 = input_56;
assign io_16 = input_57;
assign io_16 = input_58;
assign io_16 = input_59;
assign io_16 = input_60;
assign io_16 = input_61;
assign io_16 = input_62;
assign io_16 = input_63;
assign io_16 = input_64;
assign io_16 = input_65;
assign io_16 = input_66;
assign io_16 = input_67;
assign io_16 = input_68;
assign io_16 = input_69;
assign io_16 = input_70;
assign io_16 = input_71;
assign io_16 = input_72;
assign io_16 = input_73;
assign io_16 = input_74;
assign io_16 = input_75;
assign io_16 = input_76;
assign io_16 = input_77;
assign io_16 = input_78;
assign io_16 = input_79;
assign io_16 = input_80;
assign io_16 = input_81;
assign io_16 = input_82;
assign io_16 = input_83;
assign io_16 = input_84;
assign io_16 = input_85;
assign io_16 = input_86;
assign io_16 = input_87;
assign io_16 = input_88;
assign io_16 = input_89;
assign io_16 = input_90;
assign io_16 = input_91;
assign io_16 = input_92;
assign io_16 = input_93;
assign io_16 = input_94;
assign io_16 = input_95;
assign io_16 = input_96;
assign io_16 = input_97;
assign io_16 = input_98;
assign io_16 = input_99;
assign io_16 = input_100;
assign io_16 = input_101;
assign io_16 = input_102;
assign io_16 = input_103;
assign io_16 = input_104;
assign io_16 = input_105;
assign io_16 = input_106;
assign io_16 = input_107;
assign io_16 = input_108;
assign io_16 = input_109;
assign io_16 = input_110;
assign io_16 = input_111;
assign io_16 = input_112;
assign io_16 = input_113;
assign io_16 = input_114;
assign io_16 = input_115;
assign io_16 = input_116;
assign io_16 = input_117;
assign io_16 = input_118;
assign io_16 = input_119;
assign io_16 = input_120;
assign io_16 = input_121;
assign io_16 = input_122;
assign io_16 = input_123;
assign io_16 = input_124;
assign io_16 = input_125;
assign io_16 = input_126;
assign io_16 = input_127;
assign io_17 = input_17;
assign io_17 = input_18;
assign io_17 = input_19;
assign io_17 = input_20;
assign io_17 = input_21;
assign io_17 = input_22;
assign io_17 = input_23;
assign io_17 = input_24;
assign io_17 = input_25;
assign io_17 = input_26;
assign io_17 = input_27;
assign io_17 = input_28;
assign io_17 = input_29;
assign io_17 = input_30;
assign io_17 = input_31;
assign io_17 = input_32;
assign io_17 = input_33;
assign io_17 = input_34;
assign io_17 = input_35;
assign io_17 = input_36;
assign io_17 = input_37;
assign io_17 = input_38;
assign io_17 = input_39;
assign io_17 = input_40;
assign io_17 = input_41;
assign io_17 = input_42;
assign io_17 = input_43;
assign io_17 = input_44;
assign io_17 = input_45;
assign io_17 = input_46;
assign io_17 = input_47;
assign io_17 = input_48;
assign io_17 = input_49;
assign io_17 = input_50;
assign io_17 = input_51;
assign io_17 = input_52;
assign io_17 = input_53;
assign io_17 = input_54;
assign io_17 = input_55;
assign io_17 = input_56;
assign io_17 = input_57;
assign io_17 = input_58;
assign io_17 = input_59;
assign io_17 = input_60;
assign io_17 = input_61;
assign io_17 = input_62;
assign io_17 = input_63;
assign io_17 = input_64;
assign io_17 = input_65;
assign io_17 = input_66;
assign io_17 = input_67;
assign io_17 = input_68;
assign io_17 = input_69;
assign io_17 = input_70;
assign io_17 = input_71;
assign io_17 = input_72;
assign io_17 = input_73;
assign io_17 = input_74;
assign io_17 = input_75;
assign io_17 = input_76;
assign io_17 = input_77;
assign io_17 = input_78;
assign io_17 = input_79;
assign io_17 = input_80;
assign io_17 = input_81;
assign io_17 = input_82;
assign io_17 = input_83;
assign io_17 = input_84;
assign io_17 = input_85;
assign io_17 = input_86;
assign io_17 = input_87;
assign io_17 = input_88;
assign io_17 = input_89;
assign io_17 = input_90;
assign io_17 = input_91;
assign io_17 = input_92;
assign io_17 = input_93;
assign io_17 = input_94;
assign io_17 = input_95;
assign io_17 = input_96;
assign io_17 = input_97;
assign io_17 = input_98;
assign io_17 = input_99;
assign io_17 = input_100;
assign io_17 = input_101;
assign io_17 = input_102;
assign io_17 = input_103;
assign io_17 = input_104;
assign io_17 = input_105;
assign io_17 = input_106;
assign io_17 = input_107;
assign io_17 = input_108;
assign io_17 = input_109;
assign io_17 = input_110;
assign io_17 = input_111;
assign io_17 = input_112;
assign io_17 = input_113;
assign io_17 = input_114;
assign io_17 = input_115;
assign io_17 = input_116;
assign io_17 = input_117;
assign io_17 = input_118;
assign io_17 = input_119;
assign io_17 = input_120;
assign io_17 = input_121;
assign io_17 = input_122;
assign io_17 = input_123;
assign io_17 = input_124;
assign io_17 = input_125;
assign io_17 = input_126;
assign io_17 = input_127;
assign io_18 = input_18;
assign io_18 = input_19;
assign io_18 = input_20;
assign io_18 = input_21;
assign io_18 = input_22;
assign io_18 = input_23;
assign io_18 = input_24;
assign io_18 = input_25;
assign io_18 = input_26;
assign io_18 = input_27;
assign io_18 = input_28;
assign io_18 = input_29;
assign io_18 = input_30;
assign io_18 = input_31;
assign io_18 = input_32;
assign io_18 = input_33;
assign io_18 = input_34;
assign io_18 = input_35;
assign io_18 = input_36;
assign io_18 = input_37;
assign io_18 = input_38;
assign io_18 = input_39;
assign io_18 = input_40;
assign io_18 = input_41;
assign io_18 = input_42;
assign io_18 = input_43;
assign io_18 = input_44;
assign io_18 = input_45;
assign io_18 = input_46;
assign io_18 = input_47;
assign io_18 = input_48;
assign io_18 = input_49;
assign io_18 = input_50;
assign io_18 = input_51;
assign io_18 = input_52;
assign io_18 = input_53;
assign io_18 = input_54;
assign io_18 = input_55;
assign io_18 = input_56;
assign io_18 = input_57;
assign io_18 = input_58;
assign io_18 = input_59;
assign io_18 = input_60;
assign io_18 = input_61;
assign io_18 = input_62;
assign io_18 = input_63;
assign io_18 = input_64;
assign io_18 = input_65;
assign io_18 = input_66;
assign io_18 = input_67;
assign io_18 = input_68;
assign io_18 = input_69;
assign io_18 = input_70;
assign io_18 = input_71;
assign io_18 = input_72;
assign io_18 = input_73;
assign io_18 = input_74;
assign io_18 = input_75;
assign io_18 = input_76;
assign io_18 = input_77;
assign io_18 = input_78;
assign io_18 = input_79;
assign io_18 = input_80;
assign io_18 = input_81;
assign io_18 = input_82;
assign io_18 = input_83;
assign io_18 = input_84;
assign io_18 = input_85;
assign io_18 = input_86;
assign io_18 = input_87;
assign io_18 = input_88;
assign io_18 = input_89;
assign io_18 = input_90;
assign io_18 = input_91;
assign io_18 = input_92;
assign io_18 = input_93;
assign io_18 = input_94;
assign io_18 = input_95;
assign io_18 = input_96;
assign io_18 = input_97;
assign io_18 = input_98;
assign io_18 = input_99;
assign io_18 = input_100;
assign io_18 = input_101;
assign io_18 = input_102;
assign io_18 = input_103;
assign io_18 = input_104;
assign io_18 = input_105;
assign io_18 = input_106;
assign io_18 = input_107;
assign io_18 = input_108;
assign io_18 = input_109;
assign io_18 = input_110;
assign io_18 = input_111;
assign io_18 = input_112;
assign io_18 = input_113;
assign io_18 = input_114;
assign io_18 = input_115;
assign io_18 = input_116;
assign io_18 = input_117;
assign io_18 = input_118;
assign io_18 = input_119;
assign io_18 = input_120;
assign io_18 = input_121;
assign io_18 = input_122;
assign io_18 = input_123;
assign io_18 = input_124;
assign io_18 = input_125;
assign io_18 = input_126;
assign io_18 = input_127;
assign io_19 = input_19;
assign io_19 = input_20;
assign io_19 = input_21;
assign io_19 = input_22;
assign io_19 = input_23;
assign io_19 = input_24;
assign io_19 = input_25;
assign io_19 = input_26;
assign io_19 = input_27;
assign io_19 = input_28;
assign io_19 = input_29;
assign io_19 = input_30;
assign io_19 = input_31;
assign io_19 = input_32;
assign io_19 = input_33;
assign io_19 = input_34;
assign io_19 = input_35;
assign io_19 = input_36;
assign io_19 = input_37;
assign io_19 = input_38;
assign io_19 = input_39;
assign io_19 = input_40;
assign io_19 = input_41;
assign io_19 = input_42;
assign io_19 = input_43;
assign io_19 = input_44;
assign io_19 = input_45;
assign io_19 = input_46;
assign io_19 = input_47;
assign io_19 = input_48;
assign io_19 = input_49;
assign io_19 = input_50;
assign io_19 = input_51;
assign io_19 = input_52;
assign io_19 = input_53;
assign io_19 = input_54;
assign io_19 = input_55;
assign io_19 = input_56;
assign io_19 = input_57;
assign io_19 = input_58;
assign io_19 = input_59;
assign io_19 = input_60;
assign io_19 = input_61;
assign io_19 = input_62;
assign io_19 = input_63;
assign io_19 = input_64;
assign io_19 = input_65;
assign io_19 = input_66;
assign io_19 = input_67;
assign io_19 = input_68;
assign io_19 = input_69;
assign io_19 = input_70;
assign io_19 = input_71;
assign io_19 = input_72;
assign io_19 = input_73;
assign io_19 = input_74;
assign io_19 = input_75;
assign io_19 = input_76;
assign io_19 = input_77;
assign io_19 = input_78;
assign io_19 = input_79;
assign io_19 = input_80;
assign io_19 = input_81;
assign io_19 = input_82;
assign io_19 = input_83;
assign io_19 = input_84;
assign io_19 = input_85;
assign io_19 = input_86;
assign io_19 = input_87;
assign io_19 = input_88;
assign io_19 = input_89;
assign io_19 = input_90;
assign io_19 = input_91;
assign io_19 = input_92;
assign io_19 = input_93;
assign io_19 = input_94;
assign io_19 = input_95;
assign io_19 = input_96;
assign io_19 = input_97;
assign io_19 = input_98;
assign io_19 = input_99;
assign io_19 = input_100;
assign io_19 = input_101;
assign io_19 = input_102;
assign io_19 = input_103;
assign io_19 = input_104;
assign io_19 = input_105;
assign io_19 = input_106;
assign io_19 = input_107;
assign io_19 = input_108;
assign io_19 = input_109;
assign io_19 = input_110;
assign io_19 = input_111;
assign io_19 = input_112;
assign io_19 = input_113;
assign io_19 = input_114;
assign io_19 = input_115;
assign io_19 = input_116;
assign io_19 = input_117;
assign io_19 = input_118;
assign io_19 = input_119;
assign io_19 = input_120;
assign io_19 = input_121;
assign io_19 = input_122;
assign io_19 = input_123;
assign io_19 = input_124;
assign io_19 = input_125;
assign io_19 = input_126;
assign io_19 = input_127;
assign io_20 = input_20;
assign io_20 = input_21;
assign io_20 = input_22;
assign io_20 = input_23;
assign io_20 = input_24;
assign io_20 = input_25;
assign io_20 = input_26;
assign io_20 = input_27;
assign io_20 = input_28;
assign io_20 = input_29;
assign io_20 = input_30;
assign io_20 = input_31;
assign io_20 = input_32;
assign io_20 = input_33;
assign io_20 = input_34;
assign io_20 = input_35;
assign io_20 = input_36;
assign io_20 = input_37;
assign io_20 = input_38;
assign io_20 = input_39;
assign io_20 = input_40;
assign io_20 = input_41;
assign io_20 = input_42;
assign io_20 = input_43;
assign io_20 = input_44;
assign io_20 = input_45;
assign io_20 = input_46;
assign io_20 = input_47;
assign io_20 = input_48;
assign io_20 = input_49;
assign io_20 = input_50;
assign io_20 = input_51;
assign io_20 = input_52;
assign io_20 = input_53;
assign io_20 = input_54;
assign io_20 = input_55;
assign io_20 = input_56;
assign io_20 = input_57;
assign io_20 = input_58;
assign io_20 = input_59;
assign io_20 = input_60;
assign io_20 = input_61;
assign io_20 = input_62;
assign io_20 = input_63;
assign io_20 = input_64;
assign io_20 = input_65;
assign io_20 = input_66;
assign io_20 = input_67;
assign io_20 = input_68;
assign io_20 = input_69;
assign io_20 = input_70;
assign io_20 = input_71;
assign io_20 = input_72;
assign io_20 = input_73;
assign io_20 = input_74;
assign io_20 = input_75;
assign io_20 = input_76;
assign io_20 = input_77;
assign io_20 = input_78;
assign io_20 = input_79;
assign io_20 = input_80;
assign io_20 = input_81;
assign io_20 = input_82;
assign io_20 = input_83;
assign io_20 = input_84;
assign io_20 = input_85;
assign io_20 = input_86;
assign io_20 = input_87;
assign io_20 = input_88;
assign io_20 = input_89;
assign io_20 = input_90;
assign io_20 = input_91;
assign io_20 = input_92;
assign io_20 = input_93;
assign io_20 = input_94;
assign io_20 = input_95;
assign io_20 = input_96;
assign io_20 = input_97;
assign io_20 = input_98;
assign io_20 = input_99;
assign io_20 = input_100;
assign io_20 = input_101;
assign io_20 = input_102;
assign io_20 = input_103;
assign io_20 = input_104;
assign io_20 = input_105;
assign io_20 = input_106;
assign io_20 = input_107;
assign io_20 = input_108;
assign io_20 = input_109;
assign io_20 = input_110;
assign io_20 = input_111;
assign io_20 = input_112;
assign io_20 = input_113;
assign io_20 = input_114;
assign io_20 = input_115;
assign io_20 = input_116;
assign io_20 = input_117;
assign io_20 = input_118;
assign io_20 = input_119;
assign io_20 = input_120;
assign io_20 = input_121;
assign io_20 = input_122;
assign io_20 = input_123;
assign io_20 = input_124;
assign io_20 = input_125;
assign io_20 = input_126;
assign io_20 = input_127;
assign io_21 = input_21;
assign io_21 = input_22;
assign io_21 = input_23;
assign io_21 = input_24;
assign io_21 = input_25;
assign io_21 = input_26;
assign io_21 = input_27;
assign io_21 = input_28;
assign io_21 = input_29;
assign io_21 = input_30;
assign io_21 = input_31;
assign io_21 = input_32;
assign io_21 = input_33;
assign io_21 = input_34;
assign io_21 = input_35;
assign io_21 = input_36;
assign io_21 = input_37;
assign io_21 = input_38;
assign io_21 = input_39;
assign io_21 = input_40;
assign io_21 = input_41;
assign io_21 = input_42;
assign io_21 = input_43;
assign io_21 = input_44;
assign io_21 = input_45;
assign io_21 = input_46;
assign io_21 = input_47;
assign io_21 = input_48;
assign io_21 = input_49;
assign io_21 = input_50;
assign io_21 = input_51;
assign io_21 = input_52;
assign io_21 = input_53;
assign io_21 = input_54;
assign io_21 = input_55;
assign io_21 = input_56;
assign io_21 = input_57;
assign io_21 = input_58;
assign io_21 = input_59;
assign io_21 = input_60;
assign io_21 = input_61;
assign io_21 = input_62;
assign io_21 = input_63;
assign io_21 = input_64;
assign io_21 = input_65;
assign io_21 = input_66;
assign io_21 = input_67;
assign io_21 = input_68;
assign io_21 = input_69;
assign io_21 = input_70;
assign io_21 = input_71;
assign io_21 = input_72;
assign io_21 = input_73;
assign io_21 = input_74;
assign io_21 = input_75;
assign io_21 = input_76;
assign io_21 = input_77;
assign io_21 = input_78;
assign io_21 = input_79;
assign io_21 = input_80;
assign io_21 = input_81;
assign io_21 = input_82;
assign io_21 = input_83;
assign io_21 = input_84;
assign io_21 = input_85;
assign io_21 = input_86;
assign io_21 = input_87;
assign io_21 = input_88;
assign io_21 = input_89;
assign io_21 = input_90;
assign io_21 = input_91;
assign io_21 = input_92;
assign io_21 = input_93;
assign io_21 = input_94;
assign io_21 = input_95;
assign io_21 = input_96;
assign io_21 = input_97;
assign io_21 = input_98;
assign io_21 = input_99;
assign io_21 = input_100;
assign io_21 = input_101;
assign io_21 = input_102;
assign io_21 = input_103;
assign io_21 = input_104;
assign io_21 = input_105;
assign io_21 = input_106;
assign io_21 = input_107;
assign io_21 = input_108;
assign io_21 = input_109;
assign io_21 = input_110;
assign io_21 = input_111;
assign io_21 = input_112;
assign io_21 = input_113;
assign io_21 = input_114;
assign io_21 = input_115;
assign io_21 = input_116;
assign io_21 = input_117;
assign io_21 = input_118;
assign io_21 = input_119;
assign io_21 = input_120;
assign io_21 = input_121;
assign io_21 = input_122;
assign io_21 = input_123;
assign io_21 = input_124;
assign io_21 = input_125;
assign io_21 = input_126;
assign io_21 = input_127;
assign io_22 = input_22;
assign io_22 = input_23;
assign io_22 = input_24;
assign io_22 = input_25;
assign io_22 = input_26;
assign io_22 = input_27;
assign io_22 = input_28;
assign io_22 = input_29;
assign io_22 = input_30;
assign io_22 = input_31;
assign io_22 = input_32;
assign io_22 = input_33;
assign io_22 = input_34;
assign io_22 = input_35;
assign io_22 = input_36;
assign io_22 = input_37;
assign io_22 = input_38;
assign io_22 = input_39;
assign io_22 = input_40;
assign io_22 = input_41;
assign io_22 = input_42;
assign io_22 = input_43;
assign io_22 = input_44;
assign io_22 = input_45;
assign io_22 = input_46;
assign io_22 = input_47;
assign io_22 = input_48;
assign io_22 = input_49;
assign io_22 = input_50;
assign io_22 = input_51;
assign io_22 = input_52;
assign io_22 = input_53;
assign io_22 = input_54;
assign io_22 = input_55;
assign io_22 = input_56;
assign io_22 = input_57;
assign io_22 = input_58;
assign io_22 = input_59;
assign io_22 = input_60;
assign io_22 = input_61;
assign io_22 = input_62;
assign io_22 = input_63;
assign io_22 = input_64;
assign io_22 = input_65;
assign io_22 = input_66;
assign io_22 = input_67;
assign io_22 = input_68;
assign io_22 = input_69;
assign io_22 = input_70;
assign io_22 = input_71;
assign io_22 = input_72;
assign io_22 = input_73;
assign io_22 = input_74;
assign io_22 = input_75;
assign io_22 = input_76;
assign io_22 = input_77;
assign io_22 = input_78;
assign io_22 = input_79;
assign io_22 = input_80;
assign io_22 = input_81;
assign io_22 = input_82;
assign io_22 = input_83;
assign io_22 = input_84;
assign io_22 = input_85;
assign io_22 = input_86;
assign io_22 = input_87;
assign io_22 = input_88;
assign io_22 = input_89;
assign io_22 = input_90;
assign io_22 = input_91;
assign io_22 = input_92;
assign io_22 = input_93;
assign io_22 = input_94;
assign io_22 = input_95;
assign io_22 = input_96;
assign io_22 = input_97;
assign io_22 = input_98;
assign io_22 = input_99;
assign io_22 = input_100;
assign io_22 = input_101;
assign io_22 = input_102;
assign io_22 = input_103;
assign io_22 = input_104;
assign io_22 = input_105;
assign io_22 = input_106;
assign io_22 = input_107;
assign io_22 = input_108;
assign io_22 = input_109;
assign io_22 = input_110;
assign io_22 = input_111;
assign io_22 = input_112;
assign io_22 = input_113;
assign io_22 = input_114;
assign io_22 = input_115;
assign io_22 = input_116;
assign io_22 = input_117;
assign io_22 = input_118;
assign io_22 = input_119;
assign io_22 = input_120;
assign io_22 = input_121;
assign io_22 = input_122;
assign io_22 = input_123;
assign io_22 = input_124;
assign io_22 = input_125;
assign io_22 = input_126;
assign io_22 = input_127;
assign io_23 = input_23;
assign io_23 = input_24;
assign io_23 = input_25;
assign io_23 = input_26;
assign io_23 = input_27;
assign io_23 = input_28;
assign io_23 = input_29;
assign io_23 = input_30;
assign io_23 = input_31;
assign io_23 = input_32;
assign io_23 = input_33;
assign io_23 = input_34;
assign io_23 = input_35;
assign io_23 = input_36;
assign io_23 = input_37;
assign io_23 = input_38;
assign io_23 = input_39;
assign io_23 = input_40;
assign io_23 = input_41;
assign io_23 = input_42;
assign io_23 = input_43;
assign io_23 = input_44;
assign io_23 = input_45;
assign io_23 = input_46;
assign io_23 = input_47;
assign io_23 = input_48;
assign io_23 = input_49;
assign io_23 = input_50;
assign io_23 = input_51;
assign io_23 = input_52;
assign io_23 = input_53;
assign io_23 = input_54;
assign io_23 = input_55;
assign io_23 = input_56;
assign io_23 = input_57;
assign io_23 = input_58;
assign io_23 = input_59;
assign io_23 = input_60;
assign io_23 = input_61;
assign io_23 = input_62;
assign io_23 = input_63;
assign io_23 = input_64;
assign io_23 = input_65;
assign io_23 = input_66;
assign io_23 = input_67;
assign io_23 = input_68;
assign io_23 = input_69;
assign io_23 = input_70;
assign io_23 = input_71;
assign io_23 = input_72;
assign io_23 = input_73;
assign io_23 = input_74;
assign io_23 = input_75;
assign io_23 = input_76;
assign io_23 = input_77;
assign io_23 = input_78;
assign io_23 = input_79;
assign io_23 = input_80;
assign io_23 = input_81;
assign io_23 = input_82;
assign io_23 = input_83;
assign io_23 = input_84;
assign io_23 = input_85;
assign io_23 = input_86;
assign io_23 = input_87;
assign io_23 = input_88;
assign io_23 = input_89;
assign io_23 = input_90;
assign io_23 = input_91;
assign io_23 = input_92;
assign io_23 = input_93;
assign io_23 = input_94;
assign io_23 = input_95;
assign io_23 = input_96;
assign io_23 = input_97;
assign io_23 = input_98;
assign io_23 = input_99;
assign io_23 = input_100;
assign io_23 = input_101;
assign io_23 = input_102;
assign io_23 = input_103;
assign io_23 = input_104;
assign io_23 = input_105;
assign io_23 = input_106;
assign io_23 = input_107;
assign io_23 = input_108;
assign io_23 = input_109;
assign io_23 = input_110;
assign io_23 = input_111;
assign io_23 = input_112;
assign io_23 = input_113;
assign io_23 = input_114;
assign io_23 = input_115;
assign io_23 = input_116;
assign io_23 = input_117;
assign io_23 = input_118;
assign io_23 = input_119;
assign io_23 = input_120;
assign io_23 = input_121;
assign io_23 = input_122;
assign io_23 = input_123;
assign io_23 = input_124;
assign io_23 = input_125;
assign io_23 = input_126;
assign io_23 = input_127;
assign io_24 = input_24;
assign io_24 = input_25;
assign io_24 = input_26;
assign io_24 = input_27;
assign io_24 = input_28;
assign io_24 = input_29;
assign io_24 = input_30;
assign io_24 = input_31;
assign io_24 = input_32;
assign io_24 = input_33;
assign io_24 = input_34;
assign io_24 = input_35;
assign io_24 = input_36;
assign io_24 = input_37;
assign io_24 = input_38;
assign io_24 = input_39;
assign io_24 = input_40;
assign io_24 = input_41;
assign io_24 = input_42;
assign io_24 = input_43;
assign io_24 = input_44;
assign io_24 = input_45;
assign io_24 = input_46;
assign io_24 = input_47;
assign io_24 = input_48;
assign io_24 = input_49;
assign io_24 = input_50;
assign io_24 = input_51;
assign io_24 = input_52;
assign io_24 = input_53;
assign io_24 = input_54;
assign io_24 = input_55;
assign io_24 = input_56;
assign io_24 = input_57;
assign io_24 = input_58;
assign io_24 = input_59;
assign io_24 = input_60;
assign io_24 = input_61;
assign io_24 = input_62;
assign io_24 = input_63;
assign io_24 = input_64;
assign io_24 = input_65;
assign io_24 = input_66;
assign io_24 = input_67;
assign io_24 = input_68;
assign io_24 = input_69;
assign io_24 = input_70;
assign io_24 = input_71;
assign io_24 = input_72;
assign io_24 = input_73;
assign io_24 = input_74;
assign io_24 = input_75;
assign io_24 = input_76;
assign io_24 = input_77;
assign io_24 = input_78;
assign io_24 = input_79;
assign io_24 = input_80;
assign io_24 = input_81;
assign io_24 = input_82;
assign io_24 = input_83;
assign io_24 = input_84;
assign io_24 = input_85;
assign io_24 = input_86;
assign io_24 = input_87;
assign io_24 = input_88;
assign io_24 = input_89;
assign io_24 = input_90;
assign io_24 = input_91;
assign io_24 = input_92;
assign io_24 = input_93;
assign io_24 = input_94;
assign io_24 = input_95;
assign io_24 = input_96;
assign io_24 = input_97;
assign io_24 = input_98;
assign io_24 = input_99;
assign io_24 = input_100;
assign io_24 = input_101;
assign io_24 = input_102;
assign io_24 = input_103;
assign io_24 = input_104;
assign io_24 = input_105;
assign io_24 = input_106;
assign io_24 = input_107;
assign io_24 = input_108;
assign io_24 = input_109;
assign io_24 = input_110;
assign io_24 = input_111;
assign io_24 = input_112;
assign io_24 = input_113;
assign io_24 = input_114;
assign io_24 = input_115;
assign io_24 = input_116;
assign io_24 = input_117;
assign io_24 = input_118;
assign io_24 = input_119;
assign io_24 = input_120;
assign io_24 = input_121;
assign io_24 = input_122;
assign io_24 = input_123;
assign io_24 = input_124;
assign io_24 = input_125;
assign io_24 = input_126;
assign io_24 = input_127;
assign io_25 = input_25;
assign io_25 = input_26;
assign io_25 = input_27;
assign io_25 = input_28;
assign io_25 = input_29;
assign io_25 = input_30;
assign io_25 = input_31;
assign io_25 = input_32;
assign io_25 = input_33;
assign io_25 = input_34;
assign io_25 = input_35;
assign io_25 = input_36;
assign io_25 = input_37;
assign io_25 = input_38;
assign io_25 = input_39;
assign io_25 = input_40;
assign io_25 = input_41;
assign io_25 = input_42;
assign io_25 = input_43;
assign io_25 = input_44;
assign io_25 = input_45;
assign io_25 = input_46;
assign io_25 = input_47;
assign io_25 = input_48;
assign io_25 = input_49;
assign io_25 = input_50;
assign io_25 = input_51;
assign io_25 = input_52;
assign io_25 = input_53;
assign io_25 = input_54;
assign io_25 = input_55;
assign io_25 = input_56;
assign io_25 = input_57;
assign io_25 = input_58;
assign io_25 = input_59;
assign io_25 = input_60;
assign io_25 = input_61;
assign io_25 = input_62;
assign io_25 = input_63;
assign io_25 = input_64;
assign io_25 = input_65;
assign io_25 = input_66;
assign io_25 = input_67;
assign io_25 = input_68;
assign io_25 = input_69;
assign io_25 = input_70;
assign io_25 = input_71;
assign io_25 = input_72;
assign io_25 = input_73;
assign io_25 = input_74;
assign io_25 = input_75;
assign io_25 = input_76;
assign io_25 = input_77;
assign io_25 = input_78;
assign io_25 = input_79;
assign io_25 = input_80;
assign io_25 = input_81;
assign io_25 = input_82;
assign io_25 = input_83;
assign io_25 = input_84;
assign io_25 = input_85;
assign io_25 = input_86;
assign io_25 = input_87;
assign io_25 = input_88;
assign io_25 = input_89;
assign io_25 = input_90;
assign io_25 = input_91;
assign io_25 = input_92;
assign io_25 = input_93;
assign io_25 = input_94;
assign io_25 = input_95;
assign io_25 = input_96;
assign io_25 = input_97;
assign io_25 = input_98;
assign io_25 = input_99;
assign io_25 = input_100;
assign io_25 = input_101;
assign io_25 = input_102;
assign io_25 = input_103;
assign io_25 = input_104;
assign io_25 = input_105;
assign io_25 = input_106;
assign io_25 = input_107;
assign io_25 = input_108;
assign io_25 = input_109;
assign io_25 = input_110;
assign io_25 = input_111;
assign io_25 = input_112;
assign io_25 = input_113;
assign io_25 = input_114;
assign io_25 = input_115;
assign io_25 = input_116;
assign io_25 = input_117;
assign io_25 = input_118;
assign io_25 = input_119;
assign io_25 = input_120;
assign io_25 = input_121;
assign io_25 = input_122;
assign io_25 = input_123;
assign io_25 = input_124;
assign io_25 = input_125;
assign io_25 = input_126;
assign io_25 = input_127;
assign io_26 = input_26;
assign io_26 = input_27;
assign io_26 = input_28;
assign io_26 = input_29;
assign io_26 = input_30;
assign io_26 = input_31;
assign io_26 = input_32;
assign io_26 = input_33;
assign io_26 = input_34;
assign io_26 = input_35;
assign io_26 = input_36;
assign io_26 = input_37;
assign io_26 = input_38;
assign io_26 = input_39;
assign io_26 = input_40;
assign io_26 = input_41;
assign io_26 = input_42;
assign io_26 = input_43;
assign io_26 = input_44;
assign io_26 = input_45;
assign io_26 = input_46;
assign io_26 = input_47;
assign io_26 = input_48;
assign io_26 = input_49;
assign io_26 = input_50;
assign io_26 = input_51;
assign io_26 = input_52;
assign io_26 = input_53;
assign io_26 = input_54;
assign io_26 = input_55;
assign io_26 = input_56;
assign io_26 = input_57;
assign io_26 = input_58;
assign io_26 = input_59;
assign io_26 = input_60;
assign io_26 = input_61;
assign io_26 = input_62;
assign io_26 = input_63;
assign io_26 = input_64;
assign io_26 = input_65;
assign io_26 = input_66;
assign io_26 = input_67;
assign io_26 = input_68;
assign io_26 = input_69;
assign io_26 = input_70;
assign io_26 = input_71;
assign io_26 = input_72;
assign io_26 = input_73;
assign io_26 = input_74;
assign io_26 = input_75;
assign io_26 = input_76;
assign io_26 = input_77;
assign io_26 = input_78;
assign io_26 = input_79;
assign io_26 = input_80;
assign io_26 = input_81;
assign io_26 = input_82;
assign io_26 = input_83;
assign io_26 = input_84;
assign io_26 = input_85;
assign io_26 = input_86;
assign io_26 = input_87;
assign io_26 = input_88;
assign io_26 = input_89;
assign io_26 = input_90;
assign io_26 = input_91;
assign io_26 = input_92;
assign io_26 = input_93;
assign io_26 = input_94;
assign io_26 = input_95;
assign io_26 = input_96;
assign io_26 = input_97;
assign io_26 = input_98;
assign io_26 = input_99;
assign io_26 = input_100;
assign io_26 = input_101;
assign io_26 = input_102;
assign io_26 = input_103;
assign io_26 = input_104;
assign io_26 = input_105;
assign io_26 = input_106;
assign io_26 = input_107;
assign io_26 = input_108;
assign io_26 = input_109;
assign io_26 = input_110;
assign io_26 = input_111;
assign io_26 = input_112;
assign io_26 = input_113;
assign io_26 = input_114;
assign io_26 = input_115;
assign io_26 = input_116;
assign io_26 = input_117;
assign io_26 = input_118;
assign io_26 = input_119;
assign io_26 = input_120;
assign io_26 = input_121;
assign io_26 = input_122;
assign io_26 = input_123;
assign io_26 = input_124;
assign io_26 = input_125;
assign io_26 = input_126;
assign io_26 = input_127;
assign io_27 = input_27;
assign io_27 = input_28;
assign io_27 = input_29;
assign io_27 = input_30;
assign io_27 = input_31;
assign io_27 = input_32;
assign io_27 = input_33;
assign io_27 = input_34;
assign io_27 = input_35;
assign io_27 = input_36;
assign io_27 = input_37;
assign io_27 = input_38;
assign io_27 = input_39;
assign io_27 = input_40;
assign io_27 = input_41;
assign io_27 = input_42;
assign io_27 = input_43;
assign io_27 = input_44;
assign io_27 = input_45;
assign io_27 = input_46;
assign io_27 = input_47;
assign io_27 = input_48;
assign io_27 = input_49;
assign io_27 = input_50;
assign io_27 = input_51;
assign io_27 = input_52;
assign io_27 = input_53;
assign io_27 = input_54;
assign io_27 = input_55;
assign io_27 = input_56;
assign io_27 = input_57;
assign io_27 = input_58;
assign io_27 = input_59;
assign io_27 = input_60;
assign io_27 = input_61;
assign io_27 = input_62;
assign io_27 = input_63;
assign io_27 = input_64;
assign io_27 = input_65;
assign io_27 = input_66;
assign io_27 = input_67;
assign io_27 = input_68;
assign io_27 = input_69;
assign io_27 = input_70;
assign io_27 = input_71;
assign io_27 = input_72;
assign io_27 = input_73;
assign io_27 = input_74;
assign io_27 = input_75;
assign io_27 = input_76;
assign io_27 = input_77;
assign io_27 = input_78;
assign io_27 = input_79;
assign io_27 = input_80;
assign io_27 = input_81;
assign io_27 = input_82;
assign io_27 = input_83;
assign io_27 = input_84;
assign io_27 = input_85;
assign io_27 = input_86;
assign io_27 = input_87;
assign io_27 = input_88;
assign io_27 = input_89;
assign io_27 = input_90;
assign io_27 = input_91;
assign io_27 = input_92;
assign io_27 = input_93;
assign io_27 = input_94;
assign io_27 = input_95;
assign io_27 = input_96;
assign io_27 = input_97;
assign io_27 = input_98;
assign io_27 = input_99;
assign io_27 = input_100;
assign io_27 = input_101;
assign io_27 = input_102;
assign io_27 = input_103;
assign io_27 = input_104;
assign io_27 = input_105;
assign io_27 = input_106;
assign io_27 = input_107;
assign io_27 = input_108;
assign io_27 = input_109;
assign io_27 = input_110;
assign io_27 = input_111;
assign io_27 = input_112;
assign io_27 = input_113;
assign io_27 = input_114;
assign io_27 = input_115;
assign io_27 = input_116;
assign io_27 = input_117;
assign io_27 = input_118;
assign io_27 = input_119;
assign io_27 = input_120;
assign io_27 = input_121;
assign io_27 = input_122;
assign io_27 = input_123;
assign io_27 = input_124;
assign io_27 = input_125;
assign io_27 = input_126;
assign io_27 = input_127;
assign io_28 = input_28;
assign io_28 = input_29;
assign io_28 = input_30;
assign io_28 = input_31;
assign io_28 = input_32;
assign io_28 = input_33;
assign io_28 = input_34;
assign io_28 = input_35;
assign io_28 = input_36;
assign io_28 = input_37;
assign io_28 = input_38;
assign io_28 = input_39;
assign io_28 = input_40;
assign io_28 = input_41;
assign io_28 = input_42;
assign io_28 = input_43;
assign io_28 = input_44;
assign io_28 = input_45;
assign io_28 = input_46;
assign io_28 = input_47;
assign io_28 = input_48;
assign io_28 = input_49;
assign io_28 = input_50;
assign io_28 = input_51;
assign io_28 = input_52;
assign io_28 = input_53;
assign io_28 = input_54;
assign io_28 = input_55;
assign io_28 = input_56;
assign io_28 = input_57;
assign io_28 = input_58;
assign io_28 = input_59;
assign io_28 = input_60;
assign io_28 = input_61;
assign io_28 = input_62;
assign io_28 = input_63;
assign io_28 = input_64;
assign io_28 = input_65;
assign io_28 = input_66;
assign io_28 = input_67;
assign io_28 = input_68;
assign io_28 = input_69;
assign io_28 = input_70;
assign io_28 = input_71;
assign io_28 = input_72;
assign io_28 = input_73;
assign io_28 = input_74;
assign io_28 = input_75;
assign io_28 = input_76;
assign io_28 = input_77;
assign io_28 = input_78;
assign io_28 = input_79;
assign io_28 = input_80;
assign io_28 = input_81;
assign io_28 = input_82;
assign io_28 = input_83;
assign io_28 = input_84;
assign io_28 = input_85;
assign io_28 = input_86;
assign io_28 = input_87;
assign io_28 = input_88;
assign io_28 = input_89;
assign io_28 = input_90;
assign io_28 = input_91;
assign io_28 = input_92;
assign io_28 = input_93;
assign io_28 = input_94;
assign io_28 = input_95;
assign io_28 = input_96;
assign io_28 = input_97;
assign io_28 = input_98;
assign io_28 = input_99;
assign io_28 = input_100;
assign io_28 = input_101;
assign io_28 = input_102;
assign io_28 = input_103;
assign io_28 = input_104;
assign io_28 = input_105;
assign io_28 = input_106;
assign io_28 = input_107;
assign io_28 = input_108;
assign io_28 = input_109;
assign io_28 = input_110;
assign io_28 = input_111;
assign io_28 = input_112;
assign io_28 = input_113;
assign io_28 = input_114;
assign io_28 = input_115;
assign io_28 = input_116;
assign io_28 = input_117;
assign io_28 = input_118;
assign io_28 = input_119;
assign io_28 = input_120;
assign io_28 = input_121;
assign io_28 = input_122;
assign io_28 = input_123;
assign io_28 = input_124;
assign io_28 = input_125;
assign io_28 = input_126;
assign io_28 = input_127;
assign io_29 = input_29;
assign io_29 = input_30;
assign io_29 = input_31;
assign io_29 = input_32;
assign io_29 = input_33;
assign io_29 = input_34;
assign io_29 = input_35;
assign io_29 = input_36;
assign io_29 = input_37;
assign io_29 = input_38;
assign io_29 = input_39;
assign io_29 = input_40;
assign io_29 = input_41;
assign io_29 = input_42;
assign io_29 = input_43;
assign io_29 = input_44;
assign io_29 = input_45;
assign io_29 = input_46;
assign io_29 = input_47;
assign io_29 = input_48;
assign io_29 = input_49;
assign io_29 = input_50;
assign io_29 = input_51;
assign io_29 = input_52;
assign io_29 = input_53;
assign io_29 = input_54;
assign io_29 = input_55;
assign io_29 = input_56;
assign io_29 = input_57;
assign io_29 = input_58;
assign io_29 = input_59;
assign io_29 = input_60;
assign io_29 = input_61;
assign io_29 = input_62;
assign io_29 = input_63;
assign io_29 = input_64;
assign io_29 = input_65;
assign io_29 = input_66;
assign io_29 = input_67;
assign io_29 = input_68;
assign io_29 = input_69;
assign io_29 = input_70;
assign io_29 = input_71;
assign io_29 = input_72;
assign io_29 = input_73;
assign io_29 = input_74;
assign io_29 = input_75;
assign io_29 = input_76;
assign io_29 = input_77;
assign io_29 = input_78;
assign io_29 = input_79;
assign io_29 = input_80;
assign io_29 = input_81;
assign io_29 = input_82;
assign io_29 = input_83;
assign io_29 = input_84;
assign io_29 = input_85;
assign io_29 = input_86;
assign io_29 = input_87;
assign io_29 = input_88;
assign io_29 = input_89;
assign io_29 = input_90;
assign io_29 = input_91;
assign io_29 = input_92;
assign io_29 = input_93;
assign io_29 = input_94;
assign io_29 = input_95;
assign io_29 = input_96;
assign io_29 = input_97;
assign io_29 = input_98;
assign io_29 = input_99;
assign io_29 = input_100;
assign io_29 = input_101;
assign io_29 = input_102;
assign io_29 = input_103;
assign io_29 = input_104;
assign io_29 = input_105;
assign io_29 = input_106;
assign io_29 = input_107;
assign io_29 = input_108;
assign io_29 = input_109;
assign io_29 = input_110;
assign io_29 = input_111;
assign io_29 = input_112;
assign io_29 = input_113;
assign io_29 = input_114;
assign io_29 = input_115;
assign io_29 = input_116;
assign io_29 = input_117;
assign io_29 = input_118;
assign io_29 = input_119;
assign io_29 = input_120;
assign io_29 = input_121;
assign io_29 = input_122;
assign io_29 = input_123;
assign io_29 = input_124;
assign io_29 = input_125;
assign io_29 = input_126;
assign io_29 = input_127;
assign io_30 = input_30;
assign io_30 = input_31;
assign io_30 = input_32;
assign io_30 = input_33;
assign io_30 = input_34;
assign io_30 = input_35;
assign io_30 = input_36;
assign io_30 = input_37;
assign io_30 = input_38;
assign io_30 = input_39;
assign io_30 = input_40;
assign io_30 = input_41;
assign io_30 = input_42;
assign io_30 = input_43;
assign io_30 = input_44;
assign io_30 = input_45;
assign io_30 = input_46;
assign io_30 = input_47;
assign io_30 = input_48;
assign io_30 = input_49;
assign io_30 = input_50;
assign io_30 = input_51;
assign io_30 = input_52;
assign io_30 = input_53;
assign io_30 = input_54;
assign io_30 = input_55;
assign io_30 = input_56;
assign io_30 = input_57;
assign io_30 = input_58;
assign io_30 = input_59;
assign io_30 = input_60;
assign io_30 = input_61;
assign io_30 = input_62;
assign io_30 = input_63;
assign io_30 = input_64;
assign io_30 = input_65;
assign io_30 = input_66;
assign io_30 = input_67;
assign io_30 = input_68;
assign io_30 = input_69;
assign io_30 = input_70;
assign io_30 = input_71;
assign io_30 = input_72;
assign io_30 = input_73;
assign io_30 = input_74;
assign io_30 = input_75;
assign io_30 = input_76;
assign io_30 = input_77;
assign io_30 = input_78;
assign io_30 = input_79;
assign io_30 = input_80;
assign io_30 = input_81;
assign io_30 = input_82;
assign io_30 = input_83;
assign io_30 = input_84;
assign io_30 = input_85;
assign io_30 = input_86;
assign io_30 = input_87;
assign io_30 = input_88;
assign io_30 = input_89;
assign io_30 = input_90;
assign io_30 = input_91;
assign io_30 = input_92;
assign io_30 = input_93;
assign io_30 = input_94;
assign io_30 = input_95;
assign io_30 = input_96;
assign io_30 = input_97;
assign io_30 = input_98;
assign io_30 = input_99;
assign io_30 = input_100;
assign io_30 = input_101;
assign io_30 = input_102;
assign io_30 = input_103;
assign io_30 = input_104;
assign io_30 = input_105;
assign io_30 = input_106;
assign io_30 = input_107;
assign io_30 = input_108;
assign io_30 = input_109;
assign io_30 = input_110;
assign io_30 = input_111;
assign io_30 = input_112;
assign io_30 = input_113;
assign io_30 = input_114;
assign io_30 = input_115;
assign io_30 = input_116;
assign io_30 = input_117;
assign io_30 = input_118;
assign io_30 = input_119;
assign io_30 = input_120;
assign io_30 = input_121;
assign io_30 = input_122;
assign io_30 = input_123;
assign io_30 = input_124;
assign io_30 = input_125;
assign io_30 = input_126;
assign io_30 = input_127;
assign io_31 = input_31;
assign io_31 = input_32;
assign io_31 = input_33;
assign io_31 = input_34;
assign io_31 = input_35;
assign io_31 = input_36;
assign io_31 = input_37;
assign io_31 = input_38;
assign io_31 = input_39;
assign io_31 = input_40;
assign io_31 = input_41;
assign io_31 = input_42;
assign io_31 = input_43;
assign io_31 = input_44;
assign io_31 = input_45;
assign io_31 = input_46;
assign io_31 = input_47;
assign io_31 = input_48;
assign io_31 = input_49;
assign io_31 = input_50;
assign io_31 = input_51;
assign io_31 = input_52;
assign io_31 = input_53;
assign io_31 = input_54;
assign io_31 = input_55;
assign io_31 = input_56;
assign io_31 = input_57;
assign io_31 = input_58;
assign io_31 = input_59;
assign io_31 = input_60;
assign io_31 = input_61;
assign io_31 = input_62;
assign io_31 = input_63;
assign io_31 = input_64;
assign io_31 = input_65;
assign io_31 = input_66;
assign io_31 = input_67;
assign io_31 = input_68;
assign io_31 = input_69;
assign io_31 = input_70;
assign io_31 = input_71;
assign io_31 = input_72;
assign io_31 = input_73;
assign io_31 = input_74;
assign io_31 = input_75;
assign io_31 = input_76;
assign io_31 = input_77;
assign io_31 = input_78;
assign io_31 = input_79;
assign io_31 = input_80;
assign io_31 = input_81;
assign io_31 = input_82;
assign io_31 = input_83;
assign io_31 = input_84;
assign io_31 = input_85;
assign io_31 = input_86;
assign io_31 = input_87;
assign io_31 = input_88;
assign io_31 = input_89;
assign io_31 = input_90;
assign io_31 = input_91;
assign io_31 = input_92;
assign io_31 = input_93;
assign io_31 = input_94;
assign io_31 = input_95;
assign io_31 = input_96;
assign io_31 = input_97;
assign io_31 = input_98;
assign io_31 = input_99;
assign io_31 = input_100;
assign io_31 = input_101;
assign io_31 = input_102;
assign io_31 = input_103;
assign io_31 = input_104;
assign io_31 = input_105;
assign io_31 = input_106;
assign io_31 = input_107;
assign io_31 = input_108;
assign io_31 = input_109;
assign io_31 = input_110;
assign io_31 = input_111;
assign io_31 = input_112;
assign io_31 = input_113;
assign io_31 = input_114;
assign io_31 = input_115;
assign io_31 = input_116;
assign io_31 = input_117;
assign io_31 = input_118;
assign io_31 = input_119;
assign io_31 = input_120;
assign io_31 = input_121;
assign io_31 = input_122;
assign io_31 = input_123;
assign io_31 = input_124;
assign io_31 = input_125;
assign io_31 = input_126;
assign io_31 = input_127;
assign io_32 = input_32;
assign io_32 = input_33;
assign io_32 = input_34;
assign io_32 = input_35;
assign io_32 = input_36;
assign io_32 = input_37;
assign io_32 = input_38;
assign io_32 = input_39;
assign io_32 = input_40;
assign io_32 = input_41;
assign io_32 = input_42;
assign io_32 = input_43;
assign io_32 = input_44;
assign io_32 = input_45;
assign io_32 = input_46;
assign io_32 = input_47;
assign io_32 = input_48;
assign io_32 = input_49;
assign io_32 = input_50;
assign io_32 = input_51;
assign io_32 = input_52;
assign io_32 = input_53;
assign io_32 = input_54;
assign io_32 = input_55;
assign io_32 = input_56;
assign io_32 = input_57;
assign io_32 = input_58;
assign io_32 = input_59;
assign io_32 = input_60;
assign io_32 = input_61;
assign io_32 = input_62;
assign io_32 = input_63;
assign io_32 = input_64;
assign io_32 = input_65;
assign io_32 = input_66;
assign io_32 = input_67;
assign io_32 = input_68;
assign io_32 = input_69;
assign io_32 = input_70;
assign io_32 = input_71;
assign io_32 = input_72;
assign io_32 = input_73;
assign io_32 = input_74;
assign io_32 = input_75;
assign io_32 = input_76;
assign io_32 = input_77;
assign io_32 = input_78;
assign io_32 = input_79;
assign io_32 = input_80;
assign io_32 = input_81;
assign io_32 = input_82;
assign io_32 = input_83;
assign io_32 = input_84;
assign io_32 = input_85;
assign io_32 = input_86;
assign io_32 = input_87;
assign io_32 = input_88;
assign io_32 = input_89;
assign io_32 = input_90;
assign io_32 = input_91;
assign io_32 = input_92;
assign io_32 = input_93;
assign io_32 = input_94;
assign io_32 = input_95;
assign io_32 = input_96;
assign io_32 = input_97;
assign io_32 = input_98;
assign io_32 = input_99;
assign io_32 = input_100;
assign io_32 = input_101;
assign io_32 = input_102;
assign io_32 = input_103;
assign io_32 = input_104;
assign io_32 = input_105;
assign io_32 = input_106;
assign io_32 = input_107;
assign io_32 = input_108;
assign io_32 = input_109;
assign io_32 = input_110;
assign io_32 = input_111;
assign io_32 = input_112;
assign io_32 = input_113;
assign io_32 = input_114;
assign io_32 = input_115;
assign io_32 = input_116;
assign io_32 = input_117;
assign io_32 = input_118;
assign io_32 = input_119;
assign io_32 = input_120;
assign io_32 = input_121;
assign io_32 = input_122;
assign io_32 = input_123;
assign io_32 = input_124;
assign io_32 = input_125;
assign io_32 = input_126;
assign io_32 = input_127;
assign io_33 = input_33;
assign io_33 = input_34;
assign io_33 = input_35;
assign io_33 = input_36;
assign io_33 = input_37;
assign io_33 = input_38;
assign io_33 = input_39;
assign io_33 = input_40;
assign io_33 = input_41;
assign io_33 = input_42;
assign io_33 = input_43;
assign io_33 = input_44;
assign io_33 = input_45;
assign io_33 = input_46;
assign io_33 = input_47;
assign io_33 = input_48;
assign io_33 = input_49;
assign io_33 = input_50;
assign io_33 = input_51;
assign io_33 = input_52;
assign io_33 = input_53;
assign io_33 = input_54;
assign io_33 = input_55;
assign io_33 = input_56;
assign io_33 = input_57;
assign io_33 = input_58;
assign io_33 = input_59;
assign io_33 = input_60;
assign io_33 = input_61;
assign io_33 = input_62;
assign io_33 = input_63;
assign io_33 = input_64;
assign io_33 = input_65;
assign io_33 = input_66;
assign io_33 = input_67;
assign io_33 = input_68;
assign io_33 = input_69;
assign io_33 = input_70;
assign io_33 = input_71;
assign io_33 = input_72;
assign io_33 = input_73;
assign io_33 = input_74;
assign io_33 = input_75;
assign io_33 = input_76;
assign io_33 = input_77;
assign io_33 = input_78;
assign io_33 = input_79;
assign io_33 = input_80;
assign io_33 = input_81;
assign io_33 = input_82;
assign io_33 = input_83;
assign io_33 = input_84;
assign io_33 = input_85;
assign io_33 = input_86;
assign io_33 = input_87;
assign io_33 = input_88;
assign io_33 = input_89;
assign io_33 = input_90;
assign io_33 = input_91;
assign io_33 = input_92;
assign io_33 = input_93;
assign io_33 = input_94;
assign io_33 = input_95;
assign io_33 = input_96;
assign io_33 = input_97;
assign io_33 = input_98;
assign io_33 = input_99;
assign io_33 = input_100;
assign io_33 = input_101;
assign io_33 = input_102;
assign io_33 = input_103;
assign io_33 = input_104;
assign io_33 = input_105;
assign io_33 = input_106;
assign io_33 = input_107;
assign io_33 = input_108;
assign io_33 = input_109;
assign io_33 = input_110;
assign io_33 = input_111;
assign io_33 = input_112;
assign io_33 = input_113;
assign io_33 = input_114;
assign io_33 = input_115;
assign io_33 = input_116;
assign io_33 = input_117;
assign io_33 = input_118;
assign io_33 = input_119;
assign io_33 = input_120;
assign io_33 = input_121;
assign io_33 = input_122;
assign io_33 = input_123;
assign io_33 = input_124;
assign io_33 = input_125;
assign io_33 = input_126;
assign io_33 = input_127;
assign io_34 = input_34;
assign io_34 = input_35;
assign io_34 = input_36;
assign io_34 = input_37;
assign io_34 = input_38;
assign io_34 = input_39;
assign io_34 = input_40;
assign io_34 = input_41;
assign io_34 = input_42;
assign io_34 = input_43;
assign io_34 = input_44;
assign io_34 = input_45;
assign io_34 = input_46;
assign io_34 = input_47;
assign io_34 = input_48;
assign io_34 = input_49;
assign io_34 = input_50;
assign io_34 = input_51;
assign io_34 = input_52;
assign io_34 = input_53;
assign io_34 = input_54;
assign io_34 = input_55;
assign io_34 = input_56;
assign io_34 = input_57;
assign io_34 = input_58;
assign io_34 = input_59;
assign io_34 = input_60;
assign io_34 = input_61;
assign io_34 = input_62;
assign io_34 = input_63;
assign io_34 = input_64;
assign io_34 = input_65;
assign io_34 = input_66;
assign io_34 = input_67;
assign io_34 = input_68;
assign io_34 = input_69;
assign io_34 = input_70;
assign io_34 = input_71;
assign io_34 = input_72;
assign io_34 = input_73;
assign io_34 = input_74;
assign io_34 = input_75;
assign io_34 = input_76;
assign io_34 = input_77;
assign io_34 = input_78;
assign io_34 = input_79;
assign io_34 = input_80;
assign io_34 = input_81;
assign io_34 = input_82;
assign io_34 = input_83;
assign io_34 = input_84;
assign io_34 = input_85;
assign io_34 = input_86;
assign io_34 = input_87;
assign io_34 = input_88;
assign io_34 = input_89;
assign io_34 = input_90;
assign io_34 = input_91;
assign io_34 = input_92;
assign io_34 = input_93;
assign io_34 = input_94;
assign io_34 = input_95;
assign io_34 = input_96;
assign io_34 = input_97;
assign io_34 = input_98;
assign io_34 = input_99;
assign io_34 = input_100;
assign io_34 = input_101;
assign io_34 = input_102;
assign io_34 = input_103;
assign io_34 = input_104;
assign io_34 = input_105;
assign io_34 = input_106;
assign io_34 = input_107;
assign io_34 = input_108;
assign io_34 = input_109;
assign io_34 = input_110;
assign io_34 = input_111;
assign io_34 = input_112;
assign io_34 = input_113;
assign io_34 = input_114;
assign io_34 = input_115;
assign io_34 = input_116;
assign io_34 = input_117;
assign io_34 = input_118;
assign io_34 = input_119;
assign io_34 = input_120;
assign io_34 = input_121;
assign io_34 = input_122;
assign io_34 = input_123;
assign io_34 = input_124;
assign io_34 = input_125;
assign io_34 = input_126;
assign io_34 = input_127;
assign io_35 = input_35;
assign io_35 = input_36;
assign io_35 = input_37;
assign io_35 = input_38;
assign io_35 = input_39;
assign io_35 = input_40;
assign io_35 = input_41;
assign io_35 = input_42;
assign io_35 = input_43;
assign io_35 = input_44;
assign io_35 = input_45;
assign io_35 = input_46;
assign io_35 = input_47;
assign io_35 = input_48;
assign io_35 = input_49;
assign io_35 = input_50;
assign io_35 = input_51;
assign io_35 = input_52;
assign io_35 = input_53;
assign io_35 = input_54;
assign io_35 = input_55;
assign io_35 = input_56;
assign io_35 = input_57;
assign io_35 = input_58;
assign io_35 = input_59;
assign io_35 = input_60;
assign io_35 = input_61;
assign io_35 = input_62;
assign io_35 = input_63;
assign io_35 = input_64;
assign io_35 = input_65;
assign io_35 = input_66;
assign io_35 = input_67;
assign io_35 = input_68;
assign io_35 = input_69;
assign io_35 = input_70;
assign io_35 = input_71;
assign io_35 = input_72;
assign io_35 = input_73;
assign io_35 = input_74;
assign io_35 = input_75;
assign io_35 = input_76;
assign io_35 = input_77;
assign io_35 = input_78;
assign io_35 = input_79;
assign io_35 = input_80;
assign io_35 = input_81;
assign io_35 = input_82;
assign io_35 = input_83;
assign io_35 = input_84;
assign io_35 = input_85;
assign io_35 = input_86;
assign io_35 = input_87;
assign io_35 = input_88;
assign io_35 = input_89;
assign io_35 = input_90;
assign io_35 = input_91;
assign io_35 = input_92;
assign io_35 = input_93;
assign io_35 = input_94;
assign io_35 = input_95;
assign io_35 = input_96;
assign io_35 = input_97;
assign io_35 = input_98;
assign io_35 = input_99;
assign io_35 = input_100;
assign io_35 = input_101;
assign io_35 = input_102;
assign io_35 = input_103;
assign io_35 = input_104;
assign io_35 = input_105;
assign io_35 = input_106;
assign io_35 = input_107;
assign io_35 = input_108;
assign io_35 = input_109;
assign io_35 = input_110;
assign io_35 = input_111;
assign io_35 = input_112;
assign io_35 = input_113;
assign io_35 = input_114;
assign io_35 = input_115;
assign io_35 = input_116;
assign io_35 = input_117;
assign io_35 = input_118;
assign io_35 = input_119;
assign io_35 = input_120;
assign io_35 = input_121;
assign io_35 = input_122;
assign io_35 = input_123;
assign io_35 = input_124;
assign io_35 = input_125;
assign io_35 = input_126;
assign io_35 = input_127;
assign io_36 = input_36;
assign io_36 = input_37;
assign io_36 = input_38;
assign io_36 = input_39;
assign io_36 = input_40;
assign io_36 = input_41;
assign io_36 = input_42;
assign io_36 = input_43;
assign io_36 = input_44;
assign io_36 = input_45;
assign io_36 = input_46;
assign io_36 = input_47;
assign io_36 = input_48;
assign io_36 = input_49;
assign io_36 = input_50;
assign io_36 = input_51;
assign io_36 = input_52;
assign io_36 = input_53;
assign io_36 = input_54;
assign io_36 = input_55;
assign io_36 = input_56;
assign io_36 = input_57;
assign io_36 = input_58;
assign io_36 = input_59;
assign io_36 = input_60;
assign io_36 = input_61;
assign io_36 = input_62;
assign io_36 = input_63;
assign io_36 = input_64;
assign io_36 = input_65;
assign io_36 = input_66;
assign io_36 = input_67;
assign io_36 = input_68;
assign io_36 = input_69;
assign io_36 = input_70;
assign io_36 = input_71;
assign io_36 = input_72;
assign io_36 = input_73;
assign io_36 = input_74;
assign io_36 = input_75;
assign io_36 = input_76;
assign io_36 = input_77;
assign io_36 = input_78;
assign io_36 = input_79;
assign io_36 = input_80;
assign io_36 = input_81;
assign io_36 = input_82;
assign io_36 = input_83;
assign io_36 = input_84;
assign io_36 = input_85;
assign io_36 = input_86;
assign io_36 = input_87;
assign io_36 = input_88;
assign io_36 = input_89;
assign io_36 = input_90;
assign io_36 = input_91;
assign io_36 = input_92;
assign io_36 = input_93;
assign io_36 = input_94;
assign io_36 = input_95;
assign io_36 = input_96;
assign io_36 = input_97;
assign io_36 = input_98;
assign io_36 = input_99;
assign io_36 = input_100;
assign io_36 = input_101;
assign io_36 = input_102;
assign io_36 = input_103;
assign io_36 = input_104;
assign io_36 = input_105;
assign io_36 = input_106;
assign io_36 = input_107;
assign io_36 = input_108;
assign io_36 = input_109;
assign io_36 = input_110;
assign io_36 = input_111;
assign io_36 = input_112;
assign io_36 = input_113;
assign io_36 = input_114;
assign io_36 = input_115;
assign io_36 = input_116;
assign io_36 = input_117;
assign io_36 = input_118;
assign io_36 = input_119;
assign io_36 = input_120;
assign io_36 = input_121;
assign io_36 = input_122;
assign io_36 = input_123;
assign io_36 = input_124;
assign io_36 = input_125;
assign io_36 = input_126;
assign io_36 = input_127;
assign io_37 = input_37;
assign io_37 = input_38;
assign io_37 = input_39;
assign io_37 = input_40;
assign io_37 = input_41;
assign io_37 = input_42;
assign io_37 = input_43;
assign io_37 = input_44;
assign io_37 = input_45;
assign io_37 = input_46;
assign io_37 = input_47;
assign io_37 = input_48;
assign io_37 = input_49;
assign io_37 = input_50;
assign io_37 = input_51;
assign io_37 = input_52;
assign io_37 = input_53;
assign io_37 = input_54;
assign io_37 = input_55;
assign io_37 = input_56;
assign io_37 = input_57;
assign io_37 = input_58;
assign io_37 = input_59;
assign io_37 = input_60;
assign io_37 = input_61;
assign io_37 = input_62;
assign io_37 = input_63;
assign io_37 = input_64;
assign io_37 = input_65;
assign io_37 = input_66;
assign io_37 = input_67;
assign io_37 = input_68;
assign io_37 = input_69;
assign io_37 = input_70;
assign io_37 = input_71;
assign io_37 = input_72;
assign io_37 = input_73;
assign io_37 = input_74;
assign io_37 = input_75;
assign io_37 = input_76;
assign io_37 = input_77;
assign io_37 = input_78;
assign io_37 = input_79;
assign io_37 = input_80;
assign io_37 = input_81;
assign io_37 = input_82;
assign io_37 = input_83;
assign io_37 = input_84;
assign io_37 = input_85;
assign io_37 = input_86;
assign io_37 = input_87;
assign io_37 = input_88;
assign io_37 = input_89;
assign io_37 = input_90;
assign io_37 = input_91;
assign io_37 = input_92;
assign io_37 = input_93;
assign io_37 = input_94;
assign io_37 = input_95;
assign io_37 = input_96;
assign io_37 = input_97;
assign io_37 = input_98;
assign io_37 = input_99;
assign io_37 = input_100;
assign io_37 = input_101;
assign io_37 = input_102;
assign io_37 = input_103;
assign io_37 = input_104;
assign io_37 = input_105;
assign io_37 = input_106;
assign io_37 = input_107;
assign io_37 = input_108;
assign io_37 = input_109;
assign io_37 = input_110;
assign io_37 = input_111;
assign io_37 = input_112;
assign io_37 = input_113;
assign io_37 = input_114;
assign io_37 = input_115;
assign io_37 = input_116;
assign io_37 = input_117;
assign io_37 = input_118;
assign io_37 = input_119;
assign io_37 = input_120;
assign io_37 = input_121;
assign io_37 = input_122;
assign io_37 = input_123;
assign io_37 = input_124;
assign io_37 = input_125;
assign io_37 = input_126;
assign io_37 = input_127;
assign io_38 = input_38;
assign io_38 = input_39;
assign io_38 = input_40;
assign io_38 = input_41;
assign io_38 = input_42;
assign io_38 = input_43;
assign io_38 = input_44;
assign io_38 = input_45;
assign io_38 = input_46;
assign io_38 = input_47;
assign io_38 = input_48;
assign io_38 = input_49;
assign io_38 = input_50;
assign io_38 = input_51;
assign io_38 = input_52;
assign io_38 = input_53;
assign io_38 = input_54;
assign io_38 = input_55;
assign io_38 = input_56;
assign io_38 = input_57;
assign io_38 = input_58;
assign io_38 = input_59;
assign io_38 = input_60;
assign io_38 = input_61;
assign io_38 = input_62;
assign io_38 = input_63;
assign io_38 = input_64;
assign io_38 = input_65;
assign io_38 = input_66;
assign io_38 = input_67;
assign io_38 = input_68;
assign io_38 = input_69;
assign io_38 = input_70;
assign io_38 = input_71;
assign io_38 = input_72;
assign io_38 = input_73;
assign io_38 = input_74;
assign io_38 = input_75;
assign io_38 = input_76;
assign io_38 = input_77;
assign io_38 = input_78;
assign io_38 = input_79;
assign io_38 = input_80;
assign io_38 = input_81;
assign io_38 = input_82;
assign io_38 = input_83;
assign io_38 = input_84;
assign io_38 = input_85;
assign io_38 = input_86;
assign io_38 = input_87;
assign io_38 = input_88;
assign io_38 = input_89;
assign io_38 = input_90;
assign io_38 = input_91;
assign io_38 = input_92;
assign io_38 = input_93;
assign io_38 = input_94;
assign io_38 = input_95;
assign io_38 = input_96;
assign io_38 = input_97;
assign io_38 = input_98;
assign io_38 = input_99;
assign io_38 = input_100;
assign io_38 = input_101;
assign io_38 = input_102;
assign io_38 = input_103;
assign io_38 = input_104;
assign io_38 = input_105;
assign io_38 = input_106;
assign io_38 = input_107;
assign io_38 = input_108;
assign io_38 = input_109;
assign io_38 = input_110;
assign io_38 = input_111;
assign io_38 = input_112;
assign io_38 = input_113;
assign io_38 = input_114;
assign io_38 = input_115;
assign io_38 = input_116;
assign io_38 = input_117;
assign io_38 = input_118;
assign io_38 = input_119;
assign io_38 = input_120;
assign io_38 = input_121;
assign io_38 = input_122;
assign io_38 = input_123;
assign io_38 = input_124;
assign io_38 = input_125;
assign io_38 = input_126;
assign io_38 = input_127;
assign io_39 = input_39;
assign io_39 = input_40;
assign io_39 = input_41;
assign io_39 = input_42;
assign io_39 = input_43;
assign io_39 = input_44;
assign io_39 = input_45;
assign io_39 = input_46;
assign io_39 = input_47;
assign io_39 = input_48;
assign io_39 = input_49;
assign io_39 = input_50;
assign io_39 = input_51;
assign io_39 = input_52;
assign io_39 = input_53;
assign io_39 = input_54;
assign io_39 = input_55;
assign io_39 = input_56;
assign io_39 = input_57;
assign io_39 = input_58;
assign io_39 = input_59;
assign io_39 = input_60;
assign io_39 = input_61;
assign io_39 = input_62;
assign io_39 = input_63;
assign io_39 = input_64;
assign io_39 = input_65;
assign io_39 = input_66;
assign io_39 = input_67;
assign io_39 = input_68;
assign io_39 = input_69;
assign io_39 = input_70;
assign io_39 = input_71;
assign io_39 = input_72;
assign io_39 = input_73;
assign io_39 = input_74;
assign io_39 = input_75;
assign io_39 = input_76;
assign io_39 = input_77;
assign io_39 = input_78;
assign io_39 = input_79;
assign io_39 = input_80;
assign io_39 = input_81;
assign io_39 = input_82;
assign io_39 = input_83;
assign io_39 = input_84;
assign io_39 = input_85;
assign io_39 = input_86;
assign io_39 = input_87;
assign io_39 = input_88;
assign io_39 = input_89;
assign io_39 = input_90;
assign io_39 = input_91;
assign io_39 = input_92;
assign io_39 = input_93;
assign io_39 = input_94;
assign io_39 = input_95;
assign io_39 = input_96;
assign io_39 = input_97;
assign io_39 = input_98;
assign io_39 = input_99;
assign io_39 = input_100;
assign io_39 = input_101;
assign io_39 = input_102;
assign io_39 = input_103;
assign io_39 = input_104;
assign io_39 = input_105;
assign io_39 = input_106;
assign io_39 = input_107;
assign io_39 = input_108;
assign io_39 = input_109;
assign io_39 = input_110;
assign io_39 = input_111;
assign io_39 = input_112;
assign io_39 = input_113;
assign io_39 = input_114;
assign io_39 = input_115;
assign io_39 = input_116;
assign io_39 = input_117;
assign io_39 = input_118;
assign io_39 = input_119;
assign io_39 = input_120;
assign io_39 = input_121;
assign io_39 = input_122;
assign io_39 = input_123;
assign io_39 = input_124;
assign io_39 = input_125;
assign io_39 = input_126;
assign io_39 = input_127;
assign io_40 = input_40;
assign io_40 = input_41;
assign io_40 = input_42;
assign io_40 = input_43;
assign io_40 = input_44;
assign io_40 = input_45;
assign io_40 = input_46;
assign io_40 = input_47;
assign io_40 = input_48;
assign io_40 = input_49;
assign io_40 = input_50;
assign io_40 = input_51;
assign io_40 = input_52;
assign io_40 = input_53;
assign io_40 = input_54;
assign io_40 = input_55;
assign io_40 = input_56;
assign io_40 = input_57;
assign io_40 = input_58;
assign io_40 = input_59;
assign io_40 = input_60;
assign io_40 = input_61;
assign io_40 = input_62;
assign io_40 = input_63;
assign io_40 = input_64;
assign io_40 = input_65;
assign io_40 = input_66;
assign io_40 = input_67;
assign io_40 = input_68;
assign io_40 = input_69;
assign io_40 = input_70;
assign io_40 = input_71;
assign io_40 = input_72;
assign io_40 = input_73;
assign io_40 = input_74;
assign io_40 = input_75;
assign io_40 = input_76;
assign io_40 = input_77;
assign io_40 = input_78;
assign io_40 = input_79;
assign io_40 = input_80;
assign io_40 = input_81;
assign io_40 = input_82;
assign io_40 = input_83;
assign io_40 = input_84;
assign io_40 = input_85;
assign io_40 = input_86;
assign io_40 = input_87;
assign io_40 = input_88;
assign io_40 = input_89;
assign io_40 = input_90;
assign io_40 = input_91;
assign io_40 = input_92;
assign io_40 = input_93;
assign io_40 = input_94;
assign io_40 = input_95;
assign io_40 = input_96;
assign io_40 = input_97;
assign io_40 = input_98;
assign io_40 = input_99;
assign io_40 = input_100;
assign io_40 = input_101;
assign io_40 = input_102;
assign io_40 = input_103;
assign io_40 = input_104;
assign io_40 = input_105;
assign io_40 = input_106;
assign io_40 = input_107;
assign io_40 = input_108;
assign io_40 = input_109;
assign io_40 = input_110;
assign io_40 = input_111;
assign io_40 = input_112;
assign io_40 = input_113;
assign io_40 = input_114;
assign io_40 = input_115;
assign io_40 = input_116;
assign io_40 = input_117;
assign io_40 = input_118;
assign io_40 = input_119;
assign io_40 = input_120;
assign io_40 = input_121;
assign io_40 = input_122;
assign io_40 = input_123;
assign io_40 = input_124;
assign io_40 = input_125;
assign io_40 = input_126;
assign io_40 = input_127;
assign io_41 = input_41;
assign io_41 = input_42;
assign io_41 = input_43;
assign io_41 = input_44;
assign io_41 = input_45;
assign io_41 = input_46;
assign io_41 = input_47;
assign io_41 = input_48;
assign io_41 = input_49;
assign io_41 = input_50;
assign io_41 = input_51;
assign io_41 = input_52;
assign io_41 = input_53;
assign io_41 = input_54;
assign io_41 = input_55;
assign io_41 = input_56;
assign io_41 = input_57;
assign io_41 = input_58;
assign io_41 = input_59;
assign io_41 = input_60;
assign io_41 = input_61;
assign io_41 = input_62;
assign io_41 = input_63;
assign io_41 = input_64;
assign io_41 = input_65;
assign io_41 = input_66;
assign io_41 = input_67;
assign io_41 = input_68;
assign io_41 = input_69;
assign io_41 = input_70;
assign io_41 = input_71;
assign io_41 = input_72;
assign io_41 = input_73;
assign io_41 = input_74;
assign io_41 = input_75;
assign io_41 = input_76;
assign io_41 = input_77;
assign io_41 = input_78;
assign io_41 = input_79;
assign io_41 = input_80;
assign io_41 = input_81;
assign io_41 = input_82;
assign io_41 = input_83;
assign io_41 = input_84;
assign io_41 = input_85;
assign io_41 = input_86;
assign io_41 = input_87;
assign io_41 = input_88;
assign io_41 = input_89;
assign io_41 = input_90;
assign io_41 = input_91;
assign io_41 = input_92;
assign io_41 = input_93;
assign io_41 = input_94;
assign io_41 = input_95;
assign io_41 = input_96;
assign io_41 = input_97;
assign io_41 = input_98;
assign io_41 = input_99;
assign io_41 = input_100;
assign io_41 = input_101;
assign io_41 = input_102;
assign io_41 = input_103;
assign io_41 = input_104;
assign io_41 = input_105;
assign io_41 = input_106;
assign io_41 = input_107;
assign io_41 = input_108;
assign io_41 = input_109;
assign io_41 = input_110;
assign io_41 = input_111;
assign io_41 = input_112;
assign io_41 = input_113;
assign io_41 = input_114;
assign io_41 = input_115;
assign io_41 = input_116;
assign io_41 = input_117;
assign io_41 = input_118;
assign io_41 = input_119;
assign io_41 = input_120;
assign io_41 = input_121;
assign io_41 = input_122;
assign io_41 = input_123;
assign io_41 = input_124;
assign io_41 = input_125;
assign io_41 = input_126;
assign io_41 = input_127;
assign io_42 = input_42;
assign io_42 = input_43;
assign io_42 = input_44;
assign io_42 = input_45;
assign io_42 = input_46;
assign io_42 = input_47;
assign io_42 = input_48;
assign io_42 = input_49;
assign io_42 = input_50;
assign io_42 = input_51;
assign io_42 = input_52;
assign io_42 = input_53;
assign io_42 = input_54;
assign io_42 = input_55;
assign io_42 = input_56;
assign io_42 = input_57;
assign io_42 = input_58;
assign io_42 = input_59;
assign io_42 = input_60;
assign io_42 = input_61;
assign io_42 = input_62;
assign io_42 = input_63;
assign io_42 = input_64;
assign io_42 = input_65;
assign io_42 = input_66;
assign io_42 = input_67;
assign io_42 = input_68;
assign io_42 = input_69;
assign io_42 = input_70;
assign io_42 = input_71;
assign io_42 = input_72;
assign io_42 = input_73;
assign io_42 = input_74;
assign io_42 = input_75;
assign io_42 = input_76;
assign io_42 = input_77;
assign io_42 = input_78;
assign io_42 = input_79;
assign io_42 = input_80;
assign io_42 = input_81;
assign io_42 = input_82;
assign io_42 = input_83;
assign io_42 = input_84;
assign io_42 = input_85;
assign io_42 = input_86;
assign io_42 = input_87;
assign io_42 = input_88;
assign io_42 = input_89;
assign io_42 = input_90;
assign io_42 = input_91;
assign io_42 = input_92;
assign io_42 = input_93;
assign io_42 = input_94;
assign io_42 = input_95;
assign io_42 = input_96;
assign io_42 = input_97;
assign io_42 = input_98;
assign io_42 = input_99;
assign io_42 = input_100;
assign io_42 = input_101;
assign io_42 = input_102;
assign io_42 = input_103;
assign io_42 = input_104;
assign io_42 = input_105;
assign io_42 = input_106;
assign io_42 = input_107;
assign io_42 = input_108;
assign io_42 = input_109;
assign io_42 = input_110;
assign io_42 = input_111;
assign io_42 = input_112;
assign io_42 = input_113;
assign io_42 = input_114;
assign io_42 = input_115;
assign io_42 = input_116;
assign io_42 = input_117;
assign io_42 = input_118;
assign io_42 = input_119;
assign io_42 = input_120;
assign io_42 = input_121;
assign io_42 = input_122;
assign io_42 = input_123;
assign io_42 = input_124;
assign io_42 = input_125;
assign io_42 = input_126;
assign io_42 = input_127;
assign io_43 = input_43;
assign io_43 = input_44;
assign io_43 = input_45;
assign io_43 = input_46;
assign io_43 = input_47;
assign io_43 = input_48;
assign io_43 = input_49;
assign io_43 = input_50;
assign io_43 = input_51;
assign io_43 = input_52;
assign io_43 = input_53;
assign io_43 = input_54;
assign io_43 = input_55;
assign io_43 = input_56;
assign io_43 = input_57;
assign io_43 = input_58;
assign io_43 = input_59;
assign io_43 = input_60;
assign io_43 = input_61;
assign io_43 = input_62;
assign io_43 = input_63;
assign io_43 = input_64;
assign io_43 = input_65;
assign io_43 = input_66;
assign io_43 = input_67;
assign io_43 = input_68;
assign io_43 = input_69;
assign io_43 = input_70;
assign io_43 = input_71;
assign io_43 = input_72;
assign io_43 = input_73;
assign io_43 = input_74;
assign io_43 = input_75;
assign io_43 = input_76;
assign io_43 = input_77;
assign io_43 = input_78;
assign io_43 = input_79;
assign io_43 = input_80;
assign io_43 = input_81;
assign io_43 = input_82;
assign io_43 = input_83;
assign io_43 = input_84;
assign io_43 = input_85;
assign io_43 = input_86;
assign io_43 = input_87;
assign io_43 = input_88;
assign io_43 = input_89;
assign io_43 = input_90;
assign io_43 = input_91;
assign io_43 = input_92;
assign io_43 = input_93;
assign io_43 = input_94;
assign io_43 = input_95;
assign io_43 = input_96;
assign io_43 = input_97;
assign io_43 = input_98;
assign io_43 = input_99;
assign io_43 = input_100;
assign io_43 = input_101;
assign io_43 = input_102;
assign io_43 = input_103;
assign io_43 = input_104;
assign io_43 = input_105;
assign io_43 = input_106;
assign io_43 = input_107;
assign io_43 = input_108;
assign io_43 = input_109;
assign io_43 = input_110;
assign io_43 = input_111;
assign io_43 = input_112;
assign io_43 = input_113;
assign io_43 = input_114;
assign io_43 = input_115;
assign io_43 = input_116;
assign io_43 = input_117;
assign io_43 = input_118;
assign io_43 = input_119;
assign io_43 = input_120;
assign io_43 = input_121;
assign io_43 = input_122;
assign io_43 = input_123;
assign io_43 = input_124;
assign io_43 = input_125;
assign io_43 = input_126;
assign io_43 = input_127;
assign io_44 = input_44;
assign io_44 = input_45;
assign io_44 = input_46;
assign io_44 = input_47;
assign io_44 = input_48;
assign io_44 = input_49;
assign io_44 = input_50;
assign io_44 = input_51;
assign io_44 = input_52;
assign io_44 = input_53;
assign io_44 = input_54;
assign io_44 = input_55;
assign io_44 = input_56;
assign io_44 = input_57;
assign io_44 = input_58;
assign io_44 = input_59;
assign io_44 = input_60;
assign io_44 = input_61;
assign io_44 = input_62;
assign io_44 = input_63;
assign io_44 = input_64;
assign io_44 = input_65;
assign io_44 = input_66;
assign io_44 = input_67;
assign io_44 = input_68;
assign io_44 = input_69;
assign io_44 = input_70;
assign io_44 = input_71;
assign io_44 = input_72;
assign io_44 = input_73;
assign io_44 = input_74;
assign io_44 = input_75;
assign io_44 = input_76;
assign io_44 = input_77;
assign io_44 = input_78;
assign io_44 = input_79;
assign io_44 = input_80;
assign io_44 = input_81;
assign io_44 = input_82;
assign io_44 = input_83;
assign io_44 = input_84;
assign io_44 = input_85;
assign io_44 = input_86;
assign io_44 = input_87;
assign io_44 = input_88;
assign io_44 = input_89;
assign io_44 = input_90;
assign io_44 = input_91;
assign io_44 = input_92;
assign io_44 = input_93;
assign io_44 = input_94;
assign io_44 = input_95;
assign io_44 = input_96;
assign io_44 = input_97;
assign io_44 = input_98;
assign io_44 = input_99;
assign io_44 = input_100;
assign io_44 = input_101;
assign io_44 = input_102;
assign io_44 = input_103;
assign io_44 = input_104;
assign io_44 = input_105;
assign io_44 = input_106;
assign io_44 = input_107;
assign io_44 = input_108;
assign io_44 = input_109;
assign io_44 = input_110;
assign io_44 = input_111;
assign io_44 = input_112;
assign io_44 = input_113;
assign io_44 = input_114;
assign io_44 = input_115;
assign io_44 = input_116;
assign io_44 = input_117;
assign io_44 = input_118;
assign io_44 = input_119;
assign io_44 = input_120;
assign io_44 = input_121;
assign io_44 = input_122;
assign io_44 = input_123;
assign io_44 = input_124;
assign io_44 = input_125;
assign io_44 = input_126;
assign io_44 = input_127;
assign io_45 = input_45;
assign io_45 = input_46;
assign io_45 = input_47;
assign io_45 = input_48;
assign io_45 = input_49;
assign io_45 = input_50;
assign io_45 = input_51;
assign io_45 = input_52;
assign io_45 = input_53;
assign io_45 = input_54;
assign io_45 = input_55;
assign io_45 = input_56;
assign io_45 = input_57;
assign io_45 = input_58;
assign io_45 = input_59;
assign io_45 = input_60;
assign io_45 = input_61;
assign io_45 = input_62;
assign io_45 = input_63;
assign io_45 = input_64;
assign io_45 = input_65;
assign io_45 = input_66;
assign io_45 = input_67;
assign io_45 = input_68;
assign io_45 = input_69;
assign io_45 = input_70;
assign io_45 = input_71;
assign io_45 = input_72;
assign io_45 = input_73;
assign io_45 = input_74;
assign io_45 = input_75;
assign io_45 = input_76;
assign io_45 = input_77;
assign io_45 = input_78;
assign io_45 = input_79;
assign io_45 = input_80;
assign io_45 = input_81;
assign io_45 = input_82;
assign io_45 = input_83;
assign io_45 = input_84;
assign io_45 = input_85;
assign io_45 = input_86;
assign io_45 = input_87;
assign io_45 = input_88;
assign io_45 = input_89;
assign io_45 = input_90;
assign io_45 = input_91;
assign io_45 = input_92;
assign io_45 = input_93;
assign io_45 = input_94;
assign io_45 = input_95;
assign io_45 = input_96;
assign io_45 = input_97;
assign io_45 = input_98;
assign io_45 = input_99;
assign io_45 = input_100;
assign io_45 = input_101;
assign io_45 = input_102;
assign io_45 = input_103;
assign io_45 = input_104;
assign io_45 = input_105;
assign io_45 = input_106;
assign io_45 = input_107;
assign io_45 = input_108;
assign io_45 = input_109;
assign io_45 = input_110;
assign io_45 = input_111;
assign io_45 = input_112;
assign io_45 = input_113;
assign io_45 = input_114;
assign io_45 = input_115;
assign io_45 = input_116;
assign io_45 = input_117;
assign io_45 = input_118;
assign io_45 = input_119;
assign io_45 = input_120;
assign io_45 = input_121;
assign io_45 = input_122;
assign io_45 = input_123;
assign io_45 = input_124;
assign io_45 = input_125;
assign io_45 = input_126;
assign io_45 = input_127;
assign io_46 = input_46;
assign io_46 = input_47;
assign io_46 = input_48;
assign io_46 = input_49;
assign io_46 = input_50;
assign io_46 = input_51;
assign io_46 = input_52;
assign io_46 = input_53;
assign io_46 = input_54;
assign io_46 = input_55;
assign io_46 = input_56;
assign io_46 = input_57;
assign io_46 = input_58;
assign io_46 = input_59;
assign io_46 = input_60;
assign io_46 = input_61;
assign io_46 = input_62;
assign io_46 = input_63;
assign io_46 = input_64;
assign io_46 = input_65;
assign io_46 = input_66;
assign io_46 = input_67;
assign io_46 = input_68;
assign io_46 = input_69;
assign io_46 = input_70;
assign io_46 = input_71;
assign io_46 = input_72;
assign io_46 = input_73;
assign io_46 = input_74;
assign io_46 = input_75;
assign io_46 = input_76;
assign io_46 = input_77;
assign io_46 = input_78;
assign io_46 = input_79;
assign io_46 = input_80;
assign io_46 = input_81;
assign io_46 = input_82;
assign io_46 = input_83;
assign io_46 = input_84;
assign io_46 = input_85;
assign io_46 = input_86;
assign io_46 = input_87;
assign io_46 = input_88;
assign io_46 = input_89;
assign io_46 = input_90;
assign io_46 = input_91;
assign io_46 = input_92;
assign io_46 = input_93;
assign io_46 = input_94;
assign io_46 = input_95;
assign io_46 = input_96;
assign io_46 = input_97;
assign io_46 = input_98;
assign io_46 = input_99;
assign io_46 = input_100;
assign io_46 = input_101;
assign io_46 = input_102;
assign io_46 = input_103;
assign io_46 = input_104;
assign io_46 = input_105;
assign io_46 = input_106;
assign io_46 = input_107;
assign io_46 = input_108;
assign io_46 = input_109;
assign io_46 = input_110;
assign io_46 = input_111;
assign io_46 = input_112;
assign io_46 = input_113;
assign io_46 = input_114;
assign io_46 = input_115;
assign io_46 = input_116;
assign io_46 = input_117;
assign io_46 = input_118;
assign io_46 = input_119;
assign io_46 = input_120;
assign io_46 = input_121;
assign io_46 = input_122;
assign io_46 = input_123;
assign io_46 = input_124;
assign io_46 = input_125;
assign io_46 = input_126;
assign io_46 = input_127;
assign io_47 = input_47;
assign io_47 = input_48;
assign io_47 = input_49;
assign io_47 = input_50;
assign io_47 = input_51;
assign io_47 = input_52;
assign io_47 = input_53;
assign io_47 = input_54;
assign io_47 = input_55;
assign io_47 = input_56;
assign io_47 = input_57;
assign io_47 = input_58;
assign io_47 = input_59;
assign io_47 = input_60;
assign io_47 = input_61;
assign io_47 = input_62;
assign io_47 = input_63;
assign io_47 = input_64;
assign io_47 = input_65;
assign io_47 = input_66;
assign io_47 = input_67;
assign io_47 = input_68;
assign io_47 = input_69;
assign io_47 = input_70;
assign io_47 = input_71;
assign io_47 = input_72;
assign io_47 = input_73;
assign io_47 = input_74;
assign io_47 = input_75;
assign io_47 = input_76;
assign io_47 = input_77;
assign io_47 = input_78;
assign io_47 = input_79;
assign io_47 = input_80;
assign io_47 = input_81;
assign io_47 = input_82;
assign io_47 = input_83;
assign io_47 = input_84;
assign io_47 = input_85;
assign io_47 = input_86;
assign io_47 = input_87;
assign io_47 = input_88;
assign io_47 = input_89;
assign io_47 = input_90;
assign io_47 = input_91;
assign io_47 = input_92;
assign io_47 = input_93;
assign io_47 = input_94;
assign io_47 = input_95;
assign io_47 = input_96;
assign io_47 = input_97;
assign io_47 = input_98;
assign io_47 = input_99;
assign io_47 = input_100;
assign io_47 = input_101;
assign io_47 = input_102;
assign io_47 = input_103;
assign io_47 = input_104;
assign io_47 = input_105;
assign io_47 = input_106;
assign io_47 = input_107;
assign io_47 = input_108;
assign io_47 = input_109;
assign io_47 = input_110;
assign io_47 = input_111;
assign io_47 = input_112;
assign io_47 = input_113;
assign io_47 = input_114;
assign io_47 = input_115;
assign io_47 = input_116;
assign io_47 = input_117;
assign io_47 = input_118;
assign io_47 = input_119;
assign io_47 = input_120;
assign io_47 = input_121;
assign io_47 = input_122;
assign io_47 = input_123;
assign io_47 = input_124;
assign io_47 = input_125;
assign io_47 = input_126;
assign io_47 = input_127;
assign io_48 = input_48;
assign io_48 = input_49;
assign io_48 = input_50;
assign io_48 = input_51;
assign io_48 = input_52;
assign io_48 = input_53;
assign io_48 = input_54;
assign io_48 = input_55;
assign io_48 = input_56;
assign io_48 = input_57;
assign io_48 = input_58;
assign io_48 = input_59;
assign io_48 = input_60;
assign io_48 = input_61;
assign io_48 = input_62;
assign io_48 = input_63;
assign io_48 = input_64;
assign io_48 = input_65;
assign io_48 = input_66;
assign io_48 = input_67;
assign io_48 = input_68;
assign io_48 = input_69;
assign io_48 = input_70;
assign io_48 = input_71;
assign io_48 = input_72;
assign io_48 = input_73;
assign io_48 = input_74;
assign io_48 = input_75;
assign io_48 = input_76;
assign io_48 = input_77;
assign io_48 = input_78;
assign io_48 = input_79;
assign io_48 = input_80;
assign io_48 = input_81;
assign io_48 = input_82;
assign io_48 = input_83;
assign io_48 = input_84;
assign io_48 = input_85;
assign io_48 = input_86;
assign io_48 = input_87;
assign io_48 = input_88;
assign io_48 = input_89;
assign io_48 = input_90;
assign io_48 = input_91;
assign io_48 = input_92;
assign io_48 = input_93;
assign io_48 = input_94;
assign io_48 = input_95;
assign io_48 = input_96;
assign io_48 = input_97;
assign io_48 = input_98;
assign io_48 = input_99;
assign io_48 = input_100;
assign io_48 = input_101;
assign io_48 = input_102;
assign io_48 = input_103;
assign io_48 = input_104;
assign io_48 = input_105;
assign io_48 = input_106;
assign io_48 = input_107;
assign io_48 = input_108;
assign io_48 = input_109;
assign io_48 = input_110;
assign io_48 = input_111;
assign io_48 = input_112;
assign io_48 = input_113;
assign io_48 = input_114;
assign io_48 = input_115;
assign io_48 = input_116;
assign io_48 = input_117;
assign io_48 = input_118;
assign io_48 = input_119;
assign io_48 = input_120;
assign io_48 = input_121;
assign io_48 = input_122;
assign io_48 = input_123;
assign io_48 = input_124;
assign io_48 = input_125;
assign io_48 = input_126;
assign io_48 = input_127;
assign io_49 = input_49;
assign io_49 = input_50;
assign io_49 = input_51;
assign io_49 = input_52;
assign io_49 = input_53;
assign io_49 = input_54;
assign io_49 = input_55;
assign io_49 = input_56;
assign io_49 = input_57;
assign io_49 = input_58;
assign io_49 = input_59;
assign io_49 = input_60;
assign io_49 = input_61;
assign io_49 = input_62;
assign io_49 = input_63;
assign io_49 = input_64;
assign io_49 = input_65;
assign io_49 = input_66;
assign io_49 = input_67;
assign io_49 = input_68;
assign io_49 = input_69;
assign io_49 = input_70;
assign io_49 = input_71;
assign io_49 = input_72;
assign io_49 = input_73;
assign io_49 = input_74;
assign io_49 = input_75;
assign io_49 = input_76;
assign io_49 = input_77;
assign io_49 = input_78;
assign io_49 = input_79;
assign io_49 = input_80;
assign io_49 = input_81;
assign io_49 = input_82;
assign io_49 = input_83;
assign io_49 = input_84;
assign io_49 = input_85;
assign io_49 = input_86;
assign io_49 = input_87;
assign io_49 = input_88;
assign io_49 = input_89;
assign io_49 = input_90;
assign io_49 = input_91;
assign io_49 = input_92;
assign io_49 = input_93;
assign io_49 = input_94;
assign io_49 = input_95;
assign io_49 = input_96;
assign io_49 = input_97;
assign io_49 = input_98;
assign io_49 = input_99;
assign io_49 = input_100;
assign io_49 = input_101;
assign io_49 = input_102;
assign io_49 = input_103;
assign io_49 = input_104;
assign io_49 = input_105;
assign io_49 = input_106;
assign io_49 = input_107;
assign io_49 = input_108;
assign io_49 = input_109;
assign io_49 = input_110;
assign io_49 = input_111;
assign io_49 = input_112;
assign io_49 = input_113;
assign io_49 = input_114;
assign io_49 = input_115;
assign io_49 = input_116;
assign io_49 = input_117;
assign io_49 = input_118;
assign io_49 = input_119;
assign io_49 = input_120;
assign io_49 = input_121;
assign io_49 = input_122;
assign io_49 = input_123;
assign io_49 = input_124;
assign io_49 = input_125;
assign io_49 = input_126;
assign io_49 = input_127;
assign io_50 = input_50;
assign io_50 = input_51;
assign io_50 = input_52;
assign io_50 = input_53;
assign io_50 = input_54;
assign io_50 = input_55;
assign io_50 = input_56;
assign io_50 = input_57;
assign io_50 = input_58;
assign io_50 = input_59;
assign io_50 = input_60;
assign io_50 = input_61;
assign io_50 = input_62;
assign io_50 = input_63;
assign io_50 = input_64;
assign io_50 = input_65;
assign io_50 = input_66;
assign io_50 = input_67;
assign io_50 = input_68;
assign io_50 = input_69;
assign io_50 = input_70;
assign io_50 = input_71;
assign io_50 = input_72;
assign io_50 = input_73;
assign io_50 = input_74;
assign io_50 = input_75;
assign io_50 = input_76;
assign io_50 = input_77;
assign io_50 = input_78;
assign io_50 = input_79;
assign io_50 = input_80;
assign io_50 = input_81;
assign io_50 = input_82;
assign io_50 = input_83;
assign io_50 = input_84;
assign io_50 = input_85;
assign io_50 = input_86;
assign io_50 = input_87;
assign io_50 = input_88;
assign io_50 = input_89;
assign io_50 = input_90;
assign io_50 = input_91;
assign io_50 = input_92;
assign io_50 = input_93;
assign io_50 = input_94;
assign io_50 = input_95;
assign io_50 = input_96;
assign io_50 = input_97;
assign io_50 = input_98;
assign io_50 = input_99;
assign io_50 = input_100;
assign io_50 = input_101;
assign io_50 = input_102;
assign io_50 = input_103;
assign io_50 = input_104;
assign io_50 = input_105;
assign io_50 = input_106;
assign io_50 = input_107;
assign io_50 = input_108;
assign io_50 = input_109;
assign io_50 = input_110;
assign io_50 = input_111;
assign io_50 = input_112;
assign io_50 = input_113;
assign io_50 = input_114;
assign io_50 = input_115;
assign io_50 = input_116;
assign io_50 = input_117;
assign io_50 = input_118;
assign io_50 = input_119;
assign io_50 = input_120;
assign io_50 = input_121;
assign io_50 = input_122;
assign io_50 = input_123;
assign io_50 = input_124;
assign io_50 = input_125;
assign io_50 = input_126;
assign io_50 = input_127;
assign io_51 = input_51;
assign io_51 = input_52;
assign io_51 = input_53;
assign io_51 = input_54;
assign io_51 = input_55;
assign io_51 = input_56;
assign io_51 = input_57;
assign io_51 = input_58;
assign io_51 = input_59;
assign io_51 = input_60;
assign io_51 = input_61;
assign io_51 = input_62;
assign io_51 = input_63;
assign io_51 = input_64;
assign io_51 = input_65;
assign io_51 = input_66;
assign io_51 = input_67;
assign io_51 = input_68;
assign io_51 = input_69;
assign io_51 = input_70;
assign io_51 = input_71;
assign io_51 = input_72;
assign io_51 = input_73;
assign io_51 = input_74;
assign io_51 = input_75;
assign io_51 = input_76;
assign io_51 = input_77;
assign io_51 = input_78;
assign io_51 = input_79;
assign io_51 = input_80;
assign io_51 = input_81;
assign io_51 = input_82;
assign io_51 = input_83;
assign io_51 = input_84;
assign io_51 = input_85;
assign io_51 = input_86;
assign io_51 = input_87;
assign io_51 = input_88;
assign io_51 = input_89;
assign io_51 = input_90;
assign io_51 = input_91;
assign io_51 = input_92;
assign io_51 = input_93;
assign io_51 = input_94;
assign io_51 = input_95;
assign io_51 = input_96;
assign io_51 = input_97;
assign io_51 = input_98;
assign io_51 = input_99;
assign io_51 = input_100;
assign io_51 = input_101;
assign io_51 = input_102;
assign io_51 = input_103;
assign io_51 = input_104;
assign io_51 = input_105;
assign io_51 = input_106;
assign io_51 = input_107;
assign io_51 = input_108;
assign io_51 = input_109;
assign io_51 = input_110;
assign io_51 = input_111;
assign io_51 = input_112;
assign io_51 = input_113;
assign io_51 = input_114;
assign io_51 = input_115;
assign io_51 = input_116;
assign io_51 = input_117;
assign io_51 = input_118;
assign io_51 = input_119;
assign io_51 = input_120;
assign io_51 = input_121;
assign io_51 = input_122;
assign io_51 = input_123;
assign io_51 = input_124;
assign io_51 = input_125;
assign io_51 = input_126;
assign io_51 = input_127;
assign io_52 = input_52;
assign io_52 = input_53;
assign io_52 = input_54;
assign io_52 = input_55;
assign io_52 = input_56;
assign io_52 = input_57;
assign io_52 = input_58;
assign io_52 = input_59;
assign io_52 = input_60;
assign io_52 = input_61;
assign io_52 = input_62;
assign io_52 = input_63;
assign io_52 = input_64;
assign io_52 = input_65;
assign io_52 = input_66;
assign io_52 = input_67;
assign io_52 = input_68;
assign io_52 = input_69;
assign io_52 = input_70;
assign io_52 = input_71;
assign io_52 = input_72;
assign io_52 = input_73;
assign io_52 = input_74;
assign io_52 = input_75;
assign io_52 = input_76;
assign io_52 = input_77;
assign io_52 = input_78;
assign io_52 = input_79;
assign io_52 = input_80;
assign io_52 = input_81;
assign io_52 = input_82;
assign io_52 = input_83;
assign io_52 = input_84;
assign io_52 = input_85;
assign io_52 = input_86;
assign io_52 = input_87;
assign io_52 = input_88;
assign io_52 = input_89;
assign io_52 = input_90;
assign io_52 = input_91;
assign io_52 = input_92;
assign io_52 = input_93;
assign io_52 = input_94;
assign io_52 = input_95;
assign io_52 = input_96;
assign io_52 = input_97;
assign io_52 = input_98;
assign io_52 = input_99;
assign io_52 = input_100;
assign io_52 = input_101;
assign io_52 = input_102;
assign io_52 = input_103;
assign io_52 = input_104;
assign io_52 = input_105;
assign io_52 = input_106;
assign io_52 = input_107;
assign io_52 = input_108;
assign io_52 = input_109;
assign io_52 = input_110;
assign io_52 = input_111;
assign io_52 = input_112;
assign io_52 = input_113;
assign io_52 = input_114;
assign io_52 = input_115;
assign io_52 = input_116;
assign io_52 = input_117;
assign io_52 = input_118;
assign io_52 = input_119;
assign io_52 = input_120;
assign io_52 = input_121;
assign io_52 = input_122;
assign io_52 = input_123;
assign io_52 = input_124;
assign io_52 = input_125;
assign io_52 = input_126;
assign io_52 = input_127;
assign io_53 = input_53;
assign io_53 = input_54;
assign io_53 = input_55;
assign io_53 = input_56;
assign io_53 = input_57;
assign io_53 = input_58;
assign io_53 = input_59;
assign io_53 = input_60;
assign io_53 = input_61;
assign io_53 = input_62;
assign io_53 = input_63;
assign io_53 = input_64;
assign io_53 = input_65;
assign io_53 = input_66;
assign io_53 = input_67;
assign io_53 = input_68;
assign io_53 = input_69;
assign io_53 = input_70;
assign io_53 = input_71;
assign io_53 = input_72;
assign io_53 = input_73;
assign io_53 = input_74;
assign io_53 = input_75;
assign io_53 = input_76;
assign io_53 = input_77;
assign io_53 = input_78;
assign io_53 = input_79;
assign io_53 = input_80;
assign io_53 = input_81;
assign io_53 = input_82;
assign io_53 = input_83;
assign io_53 = input_84;
assign io_53 = input_85;
assign io_53 = input_86;
assign io_53 = input_87;
assign io_53 = input_88;
assign io_53 = input_89;
assign io_53 = input_90;
assign io_53 = input_91;
assign io_53 = input_92;
assign io_53 = input_93;
assign io_53 = input_94;
assign io_53 = input_95;
assign io_53 = input_96;
assign io_53 = input_97;
assign io_53 = input_98;
assign io_53 = input_99;
assign io_53 = input_100;
assign io_53 = input_101;
assign io_53 = input_102;
assign io_53 = input_103;
assign io_53 = input_104;
assign io_53 = input_105;
assign io_53 = input_106;
assign io_53 = input_107;
assign io_53 = input_108;
assign io_53 = input_109;
assign io_53 = input_110;
assign io_53 = input_111;
assign io_53 = input_112;
assign io_53 = input_113;
assign io_53 = input_114;
assign io_53 = input_115;
assign io_53 = input_116;
assign io_53 = input_117;
assign io_53 = input_118;
assign io_53 = input_119;
assign io_53 = input_120;
assign io_53 = input_121;
assign io_53 = input_122;
assign io_53 = input_123;
assign io_53 = input_124;
assign io_53 = input_125;
assign io_53 = input_126;
assign io_53 = input_127;
assign io_54 = input_54;
assign io_54 = input_55;
assign io_54 = input_56;
assign io_54 = input_57;
assign io_54 = input_58;
assign io_54 = input_59;
assign io_54 = input_60;
assign io_54 = input_61;
assign io_54 = input_62;
assign io_54 = input_63;
assign io_54 = input_64;
assign io_54 = input_65;
assign io_54 = input_66;
assign io_54 = input_67;
assign io_54 = input_68;
assign io_54 = input_69;
assign io_54 = input_70;
assign io_54 = input_71;
assign io_54 = input_72;
assign io_54 = input_73;
assign io_54 = input_74;
assign io_54 = input_75;
assign io_54 = input_76;
assign io_54 = input_77;
assign io_54 = input_78;
assign io_54 = input_79;
assign io_54 = input_80;
assign io_54 = input_81;
assign io_54 = input_82;
assign io_54 = input_83;
assign io_54 = input_84;
assign io_54 = input_85;
assign io_54 = input_86;
assign io_54 = input_87;
assign io_54 = input_88;
assign io_54 = input_89;
assign io_54 = input_90;
assign io_54 = input_91;
assign io_54 = input_92;
assign io_54 = input_93;
assign io_54 = input_94;
assign io_54 = input_95;
assign io_54 = input_96;
assign io_54 = input_97;
assign io_54 = input_98;
assign io_54 = input_99;
assign io_54 = input_100;
assign io_54 = input_101;
assign io_54 = input_102;
assign io_54 = input_103;
assign io_54 = input_104;
assign io_54 = input_105;
assign io_54 = input_106;
assign io_54 = input_107;
assign io_54 = input_108;
assign io_54 = input_109;
assign io_54 = input_110;
assign io_54 = input_111;
assign io_54 = input_112;
assign io_54 = input_113;
assign io_54 = input_114;
assign io_54 = input_115;
assign io_54 = input_116;
assign io_54 = input_117;
assign io_54 = input_118;
assign io_54 = input_119;
assign io_54 = input_120;
assign io_54 = input_121;
assign io_54 = input_122;
assign io_54 = input_123;
assign io_54 = input_124;
assign io_54 = input_125;
assign io_54 = input_126;
assign io_54 = input_127;
assign io_55 = input_55;
assign io_55 = input_56;
assign io_55 = input_57;
assign io_55 = input_58;
assign io_55 = input_59;
assign io_55 = input_60;
assign io_55 = input_61;
assign io_55 = input_62;
assign io_55 = input_63;
assign io_55 = input_64;
assign io_55 = input_65;
assign io_55 = input_66;
assign io_55 = input_67;
assign io_55 = input_68;
assign io_55 = input_69;
assign io_55 = input_70;
assign io_55 = input_71;
assign io_55 = input_72;
assign io_55 = input_73;
assign io_55 = input_74;
assign io_55 = input_75;
assign io_55 = input_76;
assign io_55 = input_77;
assign io_55 = input_78;
assign io_55 = input_79;
assign io_55 = input_80;
assign io_55 = input_81;
assign io_55 = input_82;
assign io_55 = input_83;
assign io_55 = input_84;
assign io_55 = input_85;
assign io_55 = input_86;
assign io_55 = input_87;
assign io_55 = input_88;
assign io_55 = input_89;
assign io_55 = input_90;
assign io_55 = input_91;
assign io_55 = input_92;
assign io_55 = input_93;
assign io_55 = input_94;
assign io_55 = input_95;
assign io_55 = input_96;
assign io_55 = input_97;
assign io_55 = input_98;
assign io_55 = input_99;
assign io_55 = input_100;
assign io_55 = input_101;
assign io_55 = input_102;
assign io_55 = input_103;
assign io_55 = input_104;
assign io_55 = input_105;
assign io_55 = input_106;
assign io_55 = input_107;
assign io_55 = input_108;
assign io_55 = input_109;
assign io_55 = input_110;
assign io_55 = input_111;
assign io_55 = input_112;
assign io_55 = input_113;
assign io_55 = input_114;
assign io_55 = input_115;
assign io_55 = input_116;
assign io_55 = input_117;
assign io_55 = input_118;
assign io_55 = input_119;
assign io_55 = input_120;
assign io_55 = input_121;
assign io_55 = input_122;
assign io_55 = input_123;
assign io_55 = input_124;
assign io_55 = input_125;
assign io_55 = input_126;
assign io_55 = input_127;
assign io_56 = input_56;
assign io_56 = input_57;
assign io_56 = input_58;
assign io_56 = input_59;
assign io_56 = input_60;
assign io_56 = input_61;
assign io_56 = input_62;
assign io_56 = input_63;
assign io_56 = input_64;
assign io_56 = input_65;
assign io_56 = input_66;
assign io_56 = input_67;
assign io_56 = input_68;
assign io_56 = input_69;
assign io_56 = input_70;
assign io_56 = input_71;
assign io_56 = input_72;
assign io_56 = input_73;
assign io_56 = input_74;
assign io_56 = input_75;
assign io_56 = input_76;
assign io_56 = input_77;
assign io_56 = input_78;
assign io_56 = input_79;
assign io_56 = input_80;
assign io_56 = input_81;
assign io_56 = input_82;
assign io_56 = input_83;
assign io_56 = input_84;
assign io_56 = input_85;
assign io_56 = input_86;
assign io_56 = input_87;
assign io_56 = input_88;
assign io_56 = input_89;
assign io_56 = input_90;
assign io_56 = input_91;
assign io_56 = input_92;
assign io_56 = input_93;
assign io_56 = input_94;
assign io_56 = input_95;
assign io_56 = input_96;
assign io_56 = input_97;
assign io_56 = input_98;
assign io_56 = input_99;
assign io_56 = input_100;
assign io_56 = input_101;
assign io_56 = input_102;
assign io_56 = input_103;
assign io_56 = input_104;
assign io_56 = input_105;
assign io_56 = input_106;
assign io_56 = input_107;
assign io_56 = input_108;
assign io_56 = input_109;
assign io_56 = input_110;
assign io_56 = input_111;
assign io_56 = input_112;
assign io_56 = input_113;
assign io_56 = input_114;
assign io_56 = input_115;
assign io_56 = input_116;
assign io_56 = input_117;
assign io_56 = input_118;
assign io_56 = input_119;
assign io_56 = input_120;
assign io_56 = input_121;
assign io_56 = input_122;
assign io_56 = input_123;
assign io_56 = input_124;
assign io_56 = input_125;
assign io_56 = input_126;
assign io_56 = input_127;
assign io_57 = input_57;
assign io_57 = input_58;
assign io_57 = input_59;
assign io_57 = input_60;
assign io_57 = input_61;
assign io_57 = input_62;
assign io_57 = input_63;
assign io_57 = input_64;
assign io_57 = input_65;
assign io_57 = input_66;
assign io_57 = input_67;
assign io_57 = input_68;
assign io_57 = input_69;
assign io_57 = input_70;
assign io_57 = input_71;
assign io_57 = input_72;
assign io_57 = input_73;
assign io_57 = input_74;
assign io_57 = input_75;
assign io_57 = input_76;
assign io_57 = input_77;
assign io_57 = input_78;
assign io_57 = input_79;
assign io_57 = input_80;
assign io_57 = input_81;
assign io_57 = input_82;
assign io_57 = input_83;
assign io_57 = input_84;
assign io_57 = input_85;
assign io_57 = input_86;
assign io_57 = input_87;
assign io_57 = input_88;
assign io_57 = input_89;
assign io_57 = input_90;
assign io_57 = input_91;
assign io_57 = input_92;
assign io_57 = input_93;
assign io_57 = input_94;
assign io_57 = input_95;
assign io_57 = input_96;
assign io_57 = input_97;
assign io_57 = input_98;
assign io_57 = input_99;
assign io_57 = input_100;
assign io_57 = input_101;
assign io_57 = input_102;
assign io_57 = input_103;
assign io_57 = input_104;
assign io_57 = input_105;
assign io_57 = input_106;
assign io_57 = input_107;
assign io_57 = input_108;
assign io_57 = input_109;
assign io_57 = input_110;
assign io_57 = input_111;
assign io_57 = input_112;
assign io_57 = input_113;
assign io_57 = input_114;
assign io_57 = input_115;
assign io_57 = input_116;
assign io_57 = input_117;
assign io_57 = input_118;
assign io_57 = input_119;
assign io_57 = input_120;
assign io_57 = input_121;
assign io_57 = input_122;
assign io_57 = input_123;
assign io_57 = input_124;
assign io_57 = input_125;
assign io_57 = input_126;
assign io_57 = input_127;
assign io_58 = input_58;
assign io_58 = input_59;
assign io_58 = input_60;
assign io_58 = input_61;
assign io_58 = input_62;
assign io_58 = input_63;
assign io_58 = input_64;
assign io_58 = input_65;
assign io_58 = input_66;
assign io_58 = input_67;
assign io_58 = input_68;
assign io_58 = input_69;
assign io_58 = input_70;
assign io_58 = input_71;
assign io_58 = input_72;
assign io_58 = input_73;
assign io_58 = input_74;
assign io_58 = input_75;
assign io_58 = input_76;
assign io_58 = input_77;
assign io_58 = input_78;
assign io_58 = input_79;
assign io_58 = input_80;
assign io_58 = input_81;
assign io_58 = input_82;
assign io_58 = input_83;
assign io_58 = input_84;
assign io_58 = input_85;
assign io_58 = input_86;
assign io_58 = input_87;
assign io_58 = input_88;
assign io_58 = input_89;
assign io_58 = input_90;
assign io_58 = input_91;
assign io_58 = input_92;
assign io_58 = input_93;
assign io_58 = input_94;
assign io_58 = input_95;
assign io_58 = input_96;
assign io_58 = input_97;
assign io_58 = input_98;
assign io_58 = input_99;
assign io_58 = input_100;
assign io_58 = input_101;
assign io_58 = input_102;
assign io_58 = input_103;
assign io_58 = input_104;
assign io_58 = input_105;
assign io_58 = input_106;
assign io_58 = input_107;
assign io_58 = input_108;
assign io_58 = input_109;
assign io_58 = input_110;
assign io_58 = input_111;
assign io_58 = input_112;
assign io_58 = input_113;
assign io_58 = input_114;
assign io_58 = input_115;
assign io_58 = input_116;
assign io_58 = input_117;
assign io_58 = input_118;
assign io_58 = input_119;
assign io_58 = input_120;
assign io_58 = input_121;
assign io_58 = input_122;
assign io_58 = input_123;
assign io_58 = input_124;
assign io_58 = input_125;
assign io_58 = input_126;
assign io_58 = input_127;
assign io_59 = input_59;
assign io_59 = input_60;
assign io_59 = input_61;
assign io_59 = input_62;
assign io_59 = input_63;
assign io_59 = input_64;
assign io_59 = input_65;
assign io_59 = input_66;
assign io_59 = input_67;
assign io_59 = input_68;
assign io_59 = input_69;
assign io_59 = input_70;
assign io_59 = input_71;
assign io_59 = input_72;
assign io_59 = input_73;
assign io_59 = input_74;
assign io_59 = input_75;
assign io_59 = input_76;
assign io_59 = input_77;
assign io_59 = input_78;
assign io_59 = input_79;
assign io_59 = input_80;
assign io_59 = input_81;
assign io_59 = input_82;
assign io_59 = input_83;
assign io_59 = input_84;
assign io_59 = input_85;
assign io_59 = input_86;
assign io_59 = input_87;
assign io_59 = input_88;
assign io_59 = input_89;
assign io_59 = input_90;
assign io_59 = input_91;
assign io_59 = input_92;
assign io_59 = input_93;
assign io_59 = input_94;
assign io_59 = input_95;
assign io_59 = input_96;
assign io_59 = input_97;
assign io_59 = input_98;
assign io_59 = input_99;
assign io_59 = input_100;
assign io_59 = input_101;
assign io_59 = input_102;
assign io_59 = input_103;
assign io_59 = input_104;
assign io_59 = input_105;
assign io_59 = input_106;
assign io_59 = input_107;
assign io_59 = input_108;
assign io_59 = input_109;
assign io_59 = input_110;
assign io_59 = input_111;
assign io_59 = input_112;
assign io_59 = input_113;
assign io_59 = input_114;
assign io_59 = input_115;
assign io_59 = input_116;
assign io_59 = input_117;
assign io_59 = input_118;
assign io_59 = input_119;
assign io_59 = input_120;
assign io_59 = input_121;
assign io_59 = input_122;
assign io_59 = input_123;
assign io_59 = input_124;
assign io_59 = input_125;
assign io_59 = input_126;
assign io_59 = input_127;
assign io_60 = input_60;
assign io_60 = input_61;
assign io_60 = input_62;
assign io_60 = input_63;
assign io_60 = input_64;
assign io_60 = input_65;
assign io_60 = input_66;
assign io_60 = input_67;
assign io_60 = input_68;
assign io_60 = input_69;
assign io_60 = input_70;
assign io_60 = input_71;
assign io_60 = input_72;
assign io_60 = input_73;
assign io_60 = input_74;
assign io_60 = input_75;
assign io_60 = input_76;
assign io_60 = input_77;
assign io_60 = input_78;
assign io_60 = input_79;
assign io_60 = input_80;
assign io_60 = input_81;
assign io_60 = input_82;
assign io_60 = input_83;
assign io_60 = input_84;
assign io_60 = input_85;
assign io_60 = input_86;
assign io_60 = input_87;
assign io_60 = input_88;
assign io_60 = input_89;
assign io_60 = input_90;
assign io_60 = input_91;
assign io_60 = input_92;
assign io_60 = input_93;
assign io_60 = input_94;
assign io_60 = input_95;
assign io_60 = input_96;
assign io_60 = input_97;
assign io_60 = input_98;
assign io_60 = input_99;
assign io_60 = input_100;
assign io_60 = input_101;
assign io_60 = input_102;
assign io_60 = input_103;
assign io_60 = input_104;
assign io_60 = input_105;
assign io_60 = input_106;
assign io_60 = input_107;
assign io_60 = input_108;
assign io_60 = input_109;
assign io_60 = input_110;
assign io_60 = input_111;
assign io_60 = input_112;
assign io_60 = input_113;
assign io_60 = input_114;
assign io_60 = input_115;
assign io_60 = input_116;
assign io_60 = input_117;
assign io_60 = input_118;
assign io_60 = input_119;
assign io_60 = input_120;
assign io_60 = input_121;
assign io_60 = input_122;
assign io_60 = input_123;
assign io_60 = input_124;
assign io_60 = input_125;
assign io_60 = input_126;
assign io_60 = input_127;
assign io_61 = input_61;
assign io_61 = input_62;
assign io_61 = input_63;
assign io_61 = input_64;
assign io_61 = input_65;
assign io_61 = input_66;
assign io_61 = input_67;
assign io_61 = input_68;
assign io_61 = input_69;
assign io_61 = input_70;
assign io_61 = input_71;
assign io_61 = input_72;
assign io_61 = input_73;
assign io_61 = input_74;
assign io_61 = input_75;
assign io_61 = input_76;
assign io_61 = input_77;
assign io_61 = input_78;
assign io_61 = input_79;
assign io_61 = input_80;
assign io_61 = input_81;
assign io_61 = input_82;
assign io_61 = input_83;
assign io_61 = input_84;
assign io_61 = input_85;
assign io_61 = input_86;
assign io_61 = input_87;
assign io_61 = input_88;
assign io_61 = input_89;
assign io_61 = input_90;
assign io_61 = input_91;
assign io_61 = input_92;
assign io_61 = input_93;
assign io_61 = input_94;
assign io_61 = input_95;
assign io_61 = input_96;
assign io_61 = input_97;
assign io_61 = input_98;
assign io_61 = input_99;
assign io_61 = input_100;
assign io_61 = input_101;
assign io_61 = input_102;
assign io_61 = input_103;
assign io_61 = input_104;
assign io_61 = input_105;
assign io_61 = input_106;
assign io_61 = input_107;
assign io_61 = input_108;
assign io_61 = input_109;
assign io_61 = input_110;
assign io_61 = input_111;
assign io_61 = input_112;
assign io_61 = input_113;
assign io_61 = input_114;
assign io_61 = input_115;
assign io_61 = input_116;
assign io_61 = input_117;
assign io_61 = input_118;
assign io_61 = input_119;
assign io_61 = input_120;
assign io_61 = input_121;
assign io_61 = input_122;
assign io_61 = input_123;
assign io_61 = input_124;
assign io_61 = input_125;
assign io_61 = input_126;
assign io_61 = input_127;
assign io_62 = input_62;
assign io_62 = input_63;
assign io_62 = input_64;
assign io_62 = input_65;
assign io_62 = input_66;
assign io_62 = input_67;
assign io_62 = input_68;
assign io_62 = input_69;
assign io_62 = input_70;
assign io_62 = input_71;
assign io_62 = input_72;
assign io_62 = input_73;
assign io_62 = input_74;
assign io_62 = input_75;
assign io_62 = input_76;
assign io_62 = input_77;
assign io_62 = input_78;
assign io_62 = input_79;
assign io_62 = input_80;
assign io_62 = input_81;
assign io_62 = input_82;
assign io_62 = input_83;
assign io_62 = input_84;
assign io_62 = input_85;
assign io_62 = input_86;
assign io_62 = input_87;
assign io_62 = input_88;
assign io_62 = input_89;
assign io_62 = input_90;
assign io_62 = input_91;
assign io_62 = input_92;
assign io_62 = input_93;
assign io_62 = input_94;
assign io_62 = input_95;
assign io_62 = input_96;
assign io_62 = input_97;
assign io_62 = input_98;
assign io_62 = input_99;
assign io_62 = input_100;
assign io_62 = input_101;
assign io_62 = input_102;
assign io_62 = input_103;
assign io_62 = input_104;
assign io_62 = input_105;
assign io_62 = input_106;
assign io_62 = input_107;
assign io_62 = input_108;
assign io_62 = input_109;
assign io_62 = input_110;
assign io_62 = input_111;
assign io_62 = input_112;
assign io_62 = input_113;
assign io_62 = input_114;
assign io_62 = input_115;
assign io_62 = input_116;
assign io_62 = input_117;
assign io_62 = input_118;
assign io_62 = input_119;
assign io_62 = input_120;
assign io_62 = input_121;
assign io_62 = input_122;
assign io_62 = input_123;
assign io_62 = input_124;
assign io_62 = input_125;
assign io_62 = input_126;
assign io_62 = input_127;
assign io_63 = input_63;
assign io_63 = input_64;
assign io_63 = input_65;
assign io_63 = input_66;
assign io_63 = input_67;
assign io_63 = input_68;
assign io_63 = input_69;
assign io_63 = input_70;
assign io_63 = input_71;
assign io_63 = input_72;
assign io_63 = input_73;
assign io_63 = input_74;
assign io_63 = input_75;
assign io_63 = input_76;
assign io_63 = input_77;
assign io_63 = input_78;
assign io_63 = input_79;
assign io_63 = input_80;
assign io_63 = input_81;
assign io_63 = input_82;
assign io_63 = input_83;
assign io_63 = input_84;
assign io_63 = input_85;
assign io_63 = input_86;
assign io_63 = input_87;
assign io_63 = input_88;
assign io_63 = input_89;
assign io_63 = input_90;
assign io_63 = input_91;
assign io_63 = input_92;
assign io_63 = input_93;
assign io_63 = input_94;
assign io_63 = input_95;
assign io_63 = input_96;
assign io_63 = input_97;
assign io_63 = input_98;
assign io_63 = input_99;
assign io_63 = input_100;
assign io_63 = input_101;
assign io_63 = input_102;
assign io_63 = input_103;
assign io_63 = input_104;
assign io_63 = input_105;
assign io_63 = input_106;
assign io_63 = input_107;
assign io_63 = input_108;
assign io_63 = input_109;
assign io_63 = input_110;
assign io_63 = input_111;
assign io_63 = input_112;
assign io_63 = input_113;
assign io_63 = input_114;
assign io_63 = input_115;
assign io_63 = input_116;
assign io_63 = input_117;
assign io_63 = input_118;
assign io_63 = input_119;
assign io_63 = input_120;
assign io_63 = input_121;
assign io_63 = input_122;
assign io_63 = input_123;
assign io_63 = input_124;
assign io_63 = input_125;
assign io_63 = input_126;
assign io_63 = input_127;
assign io_64 = input_64;
assign io_64 = input_65;
assign io_64 = input_66;
assign io_64 = input_67;
assign io_64 = input_68;
assign io_64 = input_69;
assign io_64 = input_70;
assign io_64 = input_71;
assign io_64 = input_72;
assign io_64 = input_73;
assign io_64 = input_74;
assign io_64 = input_75;
assign io_64 = input_76;
assign io_64 = input_77;
assign io_64 = input_78;
assign io_64 = input_79;
assign io_64 = input_80;
assign io_64 = input_81;
assign io_64 = input_82;
assign io_64 = input_83;
assign io_64 = input_84;
assign io_64 = input_85;
assign io_64 = input_86;
assign io_64 = input_87;
assign io_64 = input_88;
assign io_64 = input_89;
assign io_64 = input_90;
assign io_64 = input_91;
assign io_64 = input_92;
assign io_64 = input_93;
assign io_64 = input_94;
assign io_64 = input_95;
assign io_64 = input_96;
assign io_64 = input_97;
assign io_64 = input_98;
assign io_64 = input_99;
assign io_64 = input_100;
assign io_64 = input_101;
assign io_64 = input_102;
assign io_64 = input_103;
assign io_64 = input_104;
assign io_64 = input_105;
assign io_64 = input_106;
assign io_64 = input_107;
assign io_64 = input_108;
assign io_64 = input_109;
assign io_64 = input_110;
assign io_64 = input_111;
assign io_64 = input_112;
assign io_64 = input_113;
assign io_64 = input_114;
assign io_64 = input_115;
assign io_64 = input_116;
assign io_64 = input_117;
assign io_64 = input_118;
assign io_64 = input_119;
assign io_64 = input_120;
assign io_64 = input_121;
assign io_64 = input_122;
assign io_64 = input_123;
assign io_64 = input_124;
assign io_64 = input_125;
assign io_64 = input_126;
assign io_64 = input_127;
assign io_65 = input_65;
assign io_65 = input_66;
assign io_65 = input_67;
assign io_65 = input_68;
assign io_65 = input_69;
assign io_65 = input_70;
assign io_65 = input_71;
assign io_65 = input_72;
assign io_65 = input_73;
assign io_65 = input_74;
assign io_65 = input_75;
assign io_65 = input_76;
assign io_65 = input_77;
assign io_65 = input_78;
assign io_65 = input_79;
assign io_65 = input_80;
assign io_65 = input_81;
assign io_65 = input_82;
assign io_65 = input_83;
assign io_65 = input_84;
assign io_65 = input_85;
assign io_65 = input_86;
assign io_65 = input_87;
assign io_65 = input_88;
assign io_65 = input_89;
assign io_65 = input_90;
assign io_65 = input_91;
assign io_65 = input_92;
assign io_65 = input_93;
assign io_65 = input_94;
assign io_65 = input_95;
assign io_65 = input_96;
assign io_65 = input_97;
assign io_65 = input_98;
assign io_65 = input_99;
assign io_65 = input_100;
assign io_65 = input_101;
assign io_65 = input_102;
assign io_65 = input_103;
assign io_65 = input_104;
assign io_65 = input_105;
assign io_65 = input_106;
assign io_65 = input_107;
assign io_65 = input_108;
assign io_65 = input_109;
assign io_65 = input_110;
assign io_65 = input_111;
assign io_65 = input_112;
assign io_65 = input_113;
assign io_65 = input_114;
assign io_65 = input_115;
assign io_65 = input_116;
assign io_65 = input_117;
assign io_65 = input_118;
assign io_65 = input_119;
assign io_65 = input_120;
assign io_65 = input_121;
assign io_65 = input_122;
assign io_65 = input_123;
assign io_65 = input_124;
assign io_65 = input_125;
assign io_65 = input_126;
assign io_65 = input_127;
assign io_66 = input_66;
assign io_66 = input_67;
assign io_66 = input_68;
assign io_66 = input_69;
assign io_66 = input_70;
assign io_66 = input_71;
assign io_66 = input_72;
assign io_66 = input_73;
assign io_66 = input_74;
assign io_66 = input_75;
assign io_66 = input_76;
assign io_66 = input_77;
assign io_66 = input_78;
assign io_66 = input_79;
assign io_66 = input_80;
assign io_66 = input_81;
assign io_66 = input_82;
assign io_66 = input_83;
assign io_66 = input_84;
assign io_66 = input_85;
assign io_66 = input_86;
assign io_66 = input_87;
assign io_66 = input_88;
assign io_66 = input_89;
assign io_66 = input_90;
assign io_66 = input_91;
assign io_66 = input_92;
assign io_66 = input_93;
assign io_66 = input_94;
assign io_66 = input_95;
assign io_66 = input_96;
assign io_66 = input_97;
assign io_66 = input_98;
assign io_66 = input_99;
assign io_66 = input_100;
assign io_66 = input_101;
assign io_66 = input_102;
assign io_66 = input_103;
assign io_66 = input_104;
assign io_66 = input_105;
assign io_66 = input_106;
assign io_66 = input_107;
assign io_66 = input_108;
assign io_66 = input_109;
assign io_66 = input_110;
assign io_66 = input_111;
assign io_66 = input_112;
assign io_66 = input_113;
assign io_66 = input_114;
assign io_66 = input_115;
assign io_66 = input_116;
assign io_66 = input_117;
assign io_66 = input_118;
assign io_66 = input_119;
assign io_66 = input_120;
assign io_66 = input_121;
assign io_66 = input_122;
assign io_66 = input_123;
assign io_66 = input_124;
assign io_66 = input_125;
assign io_66 = input_126;
assign io_66 = input_127;
assign io_67 = input_67;
assign io_67 = input_68;
assign io_67 = input_69;
assign io_67 = input_70;
assign io_67 = input_71;
assign io_67 = input_72;
assign io_67 = input_73;
assign io_67 = input_74;
assign io_67 = input_75;
assign io_67 = input_76;
assign io_67 = input_77;
assign io_67 = input_78;
assign io_67 = input_79;
assign io_67 = input_80;
assign io_67 = input_81;
assign io_67 = input_82;
assign io_67 = input_83;
assign io_67 = input_84;
assign io_67 = input_85;
assign io_67 = input_86;
assign io_67 = input_87;
assign io_67 = input_88;
assign io_67 = input_89;
assign io_67 = input_90;
assign io_67 = input_91;
assign io_67 = input_92;
assign io_67 = input_93;
assign io_67 = input_94;
assign io_67 = input_95;
assign io_67 = input_96;
assign io_67 = input_97;
assign io_67 = input_98;
assign io_67 = input_99;
assign io_67 = input_100;
assign io_67 = input_101;
assign io_67 = input_102;
assign io_67 = input_103;
assign io_67 = input_104;
assign io_67 = input_105;
assign io_67 = input_106;
assign io_67 = input_107;
assign io_67 = input_108;
assign io_67 = input_109;
assign io_67 = input_110;
assign io_67 = input_111;
assign io_67 = input_112;
assign io_67 = input_113;
assign io_67 = input_114;
assign io_67 = input_115;
assign io_67 = input_116;
assign io_67 = input_117;
assign io_67 = input_118;
assign io_67 = input_119;
assign io_67 = input_120;
assign io_67 = input_121;
assign io_67 = input_122;
assign io_67 = input_123;
assign io_67 = input_124;
assign io_67 = input_125;
assign io_67 = input_126;
assign io_67 = input_127;
assign io_68 = input_68;
assign io_68 = input_69;
assign io_68 = input_70;
assign io_68 = input_71;
assign io_68 = input_72;
assign io_68 = input_73;
assign io_68 = input_74;
assign io_68 = input_75;
assign io_68 = input_76;
assign io_68 = input_77;
assign io_68 = input_78;
assign io_68 = input_79;
assign io_68 = input_80;
assign io_68 = input_81;
assign io_68 = input_82;
assign io_68 = input_83;
assign io_68 = input_84;
assign io_68 = input_85;
assign io_68 = input_86;
assign io_68 = input_87;
assign io_68 = input_88;
assign io_68 = input_89;
assign io_68 = input_90;
assign io_68 = input_91;
assign io_68 = input_92;
assign io_68 = input_93;
assign io_68 = input_94;
assign io_68 = input_95;
assign io_68 = input_96;
assign io_68 = input_97;
assign io_68 = input_98;
assign io_68 = input_99;
assign io_68 = input_100;
assign io_68 = input_101;
assign io_68 = input_102;
assign io_68 = input_103;
assign io_68 = input_104;
assign io_68 = input_105;
assign io_68 = input_106;
assign io_68 = input_107;
assign io_68 = input_108;
assign io_68 = input_109;
assign io_68 = input_110;
assign io_68 = input_111;
assign io_68 = input_112;
assign io_68 = input_113;
assign io_68 = input_114;
assign io_68 = input_115;
assign io_68 = input_116;
assign io_68 = input_117;
assign io_68 = input_118;
assign io_68 = input_119;
assign io_68 = input_120;
assign io_68 = input_121;
assign io_68 = input_122;
assign io_68 = input_123;
assign io_68 = input_124;
assign io_68 = input_125;
assign io_68 = input_126;
assign io_68 = input_127;
assign io_69 = input_69;
assign io_69 = input_70;
assign io_69 = input_71;
assign io_69 = input_72;
assign io_69 = input_73;
assign io_69 = input_74;
assign io_69 = input_75;
assign io_69 = input_76;
assign io_69 = input_77;
assign io_69 = input_78;
assign io_69 = input_79;
assign io_69 = input_80;
assign io_69 = input_81;
assign io_69 = input_82;
assign io_69 = input_83;
assign io_69 = input_84;
assign io_69 = input_85;
assign io_69 = input_86;
assign io_69 = input_87;
assign io_69 = input_88;
assign io_69 = input_89;
assign io_69 = input_90;
assign io_69 = input_91;
assign io_69 = input_92;
assign io_69 = input_93;
assign io_69 = input_94;
assign io_69 = input_95;
assign io_69 = input_96;
assign io_69 = input_97;
assign io_69 = input_98;
assign io_69 = input_99;
assign io_69 = input_100;
assign io_69 = input_101;
assign io_69 = input_102;
assign io_69 = input_103;
assign io_69 = input_104;
assign io_69 = input_105;
assign io_69 = input_106;
assign io_69 = input_107;
assign io_69 = input_108;
assign io_69 = input_109;
assign io_69 = input_110;
assign io_69 = input_111;
assign io_69 = input_112;
assign io_69 = input_113;
assign io_69 = input_114;
assign io_69 = input_115;
assign io_69 = input_116;
assign io_69 = input_117;
assign io_69 = input_118;
assign io_69 = input_119;
assign io_69 = input_120;
assign io_69 = input_121;
assign io_69 = input_122;
assign io_69 = input_123;
assign io_69 = input_124;
assign io_69 = input_125;
assign io_69 = input_126;
assign io_69 = input_127;
assign io_70 = input_70;
assign io_70 = input_71;
assign io_70 = input_72;
assign io_70 = input_73;
assign io_70 = input_74;
assign io_70 = input_75;
assign io_70 = input_76;
assign io_70 = input_77;
assign io_70 = input_78;
assign io_70 = input_79;
assign io_70 = input_80;
assign io_70 = input_81;
assign io_70 = input_82;
assign io_70 = input_83;
assign io_70 = input_84;
assign io_70 = input_85;
assign io_70 = input_86;
assign io_70 = input_87;
assign io_70 = input_88;
assign io_70 = input_89;
assign io_70 = input_90;
assign io_70 = input_91;
assign io_70 = input_92;
assign io_70 = input_93;
assign io_70 = input_94;
assign io_70 = input_95;
assign io_70 = input_96;
assign io_70 = input_97;
assign io_70 = input_98;
assign io_70 = input_99;
assign io_70 = input_100;
assign io_70 = input_101;
assign io_70 = input_102;
assign io_70 = input_103;
assign io_70 = input_104;
assign io_70 = input_105;
assign io_70 = input_106;
assign io_70 = input_107;
assign io_70 = input_108;
assign io_70 = input_109;
assign io_70 = input_110;
assign io_70 = input_111;
assign io_70 = input_112;
assign io_70 = input_113;
assign io_70 = input_114;
assign io_70 = input_115;
assign io_70 = input_116;
assign io_70 = input_117;
assign io_70 = input_118;
assign io_70 = input_119;
assign io_70 = input_120;
assign io_70 = input_121;
assign io_70 = input_122;
assign io_70 = input_123;
assign io_70 = input_124;
assign io_70 = input_125;
assign io_70 = input_126;
assign io_70 = input_127;
assign io_71 = input_71;
assign io_71 = input_72;
assign io_71 = input_73;
assign io_71 = input_74;
assign io_71 = input_75;
assign io_71 = input_76;
assign io_71 = input_77;
assign io_71 = input_78;
assign io_71 = input_79;
assign io_71 = input_80;
assign io_71 = input_81;
assign io_71 = input_82;
assign io_71 = input_83;
assign io_71 = input_84;
assign io_71 = input_85;
assign io_71 = input_86;
assign io_71 = input_87;
assign io_71 = input_88;
assign io_71 = input_89;
assign io_71 = input_90;
assign io_71 = input_91;
assign io_71 = input_92;
assign io_71 = input_93;
assign io_71 = input_94;
assign io_71 = input_95;
assign io_71 = input_96;
assign io_71 = input_97;
assign io_71 = input_98;
assign io_71 = input_99;
assign io_71 = input_100;
assign io_71 = input_101;
assign io_71 = input_102;
assign io_71 = input_103;
assign io_71 = input_104;
assign io_71 = input_105;
assign io_71 = input_106;
assign io_71 = input_107;
assign io_71 = input_108;
assign io_71 = input_109;
assign io_71 = input_110;
assign io_71 = input_111;
assign io_71 = input_112;
assign io_71 = input_113;
assign io_71 = input_114;
assign io_71 = input_115;
assign io_71 = input_116;
assign io_71 = input_117;
assign io_71 = input_118;
assign io_71 = input_119;
assign io_71 = input_120;
assign io_71 = input_121;
assign io_71 = input_122;
assign io_71 = input_123;
assign io_71 = input_124;
assign io_71 = input_125;
assign io_71 = input_126;
assign io_71 = input_127;
assign io_72 = input_72;
assign io_72 = input_73;
assign io_72 = input_74;
assign io_72 = input_75;
assign io_72 = input_76;
assign io_72 = input_77;
assign io_72 = input_78;
assign io_72 = input_79;
assign io_72 = input_80;
assign io_72 = input_81;
assign io_72 = input_82;
assign io_72 = input_83;
assign io_72 = input_84;
assign io_72 = input_85;
assign io_72 = input_86;
assign io_72 = input_87;
assign io_72 = input_88;
assign io_72 = input_89;
assign io_72 = input_90;
assign io_72 = input_91;
assign io_72 = input_92;
assign io_72 = input_93;
assign io_72 = input_94;
assign io_72 = input_95;
assign io_72 = input_96;
assign io_72 = input_97;
assign io_72 = input_98;
assign io_72 = input_99;
assign io_72 = input_100;
assign io_72 = input_101;
assign io_72 = input_102;
assign io_72 = input_103;
assign io_72 = input_104;
assign io_72 = input_105;
assign io_72 = input_106;
assign io_72 = input_107;
assign io_72 = input_108;
assign io_72 = input_109;
assign io_72 = input_110;
assign io_72 = input_111;
assign io_72 = input_112;
assign io_72 = input_113;
assign io_72 = input_114;
assign io_72 = input_115;
assign io_72 = input_116;
assign io_72 = input_117;
assign io_72 = input_118;
assign io_72 = input_119;
assign io_72 = input_120;
assign io_72 = input_121;
assign io_72 = input_122;
assign io_72 = input_123;
assign io_72 = input_124;
assign io_72 = input_125;
assign io_72 = input_126;
assign io_72 = input_127;
assign io_73 = input_73;
assign io_73 = input_74;
assign io_73 = input_75;
assign io_73 = input_76;
assign io_73 = input_77;
assign io_73 = input_78;
assign io_73 = input_79;
assign io_73 = input_80;
assign io_73 = input_81;
assign io_73 = input_82;
assign io_73 = input_83;
assign io_73 = input_84;
assign io_73 = input_85;
assign io_73 = input_86;
assign io_73 = input_87;
assign io_73 = input_88;
assign io_73 = input_89;
assign io_73 = input_90;
assign io_73 = input_91;
assign io_73 = input_92;
assign io_73 = input_93;
assign io_73 = input_94;
assign io_73 = input_95;
assign io_73 = input_96;
assign io_73 = input_97;
assign io_73 = input_98;
assign io_73 = input_99;
assign io_73 = input_100;
assign io_73 = input_101;
assign io_73 = input_102;
assign io_73 = input_103;
assign io_73 = input_104;
assign io_73 = input_105;
assign io_73 = input_106;
assign io_73 = input_107;
assign io_73 = input_108;
assign io_73 = input_109;
assign io_73 = input_110;
assign io_73 = input_111;
assign io_73 = input_112;
assign io_73 = input_113;
assign io_73 = input_114;
assign io_73 = input_115;
assign io_73 = input_116;
assign io_73 = input_117;
assign io_73 = input_118;
assign io_73 = input_119;
assign io_73 = input_120;
assign io_73 = input_121;
assign io_73 = input_122;
assign io_73 = input_123;
assign io_73 = input_124;
assign io_73 = input_125;
assign io_73 = input_126;
assign io_73 = input_127;
assign io_74 = input_74;
assign io_74 = input_75;
assign io_74 = input_76;
assign io_74 = input_77;
assign io_74 = input_78;
assign io_74 = input_79;
assign io_74 = input_80;
assign io_74 = input_81;
assign io_74 = input_82;
assign io_74 = input_83;
assign io_74 = input_84;
assign io_74 = input_85;
assign io_74 = input_86;
assign io_74 = input_87;
assign io_74 = input_88;
assign io_74 = input_89;
assign io_74 = input_90;
assign io_74 = input_91;
assign io_74 = input_92;
assign io_74 = input_93;
assign io_74 = input_94;
assign io_74 = input_95;
assign io_74 = input_96;
assign io_74 = input_97;
assign io_74 = input_98;
assign io_74 = input_99;
assign io_74 = input_100;
assign io_74 = input_101;
assign io_74 = input_102;
assign io_74 = input_103;
assign io_74 = input_104;
assign io_74 = input_105;
assign io_74 = input_106;
assign io_74 = input_107;
assign io_74 = input_108;
assign io_74 = input_109;
assign io_74 = input_110;
assign io_74 = input_111;
assign io_74 = input_112;
assign io_74 = input_113;
assign io_74 = input_114;
assign io_74 = input_115;
assign io_74 = input_116;
assign io_74 = input_117;
assign io_74 = input_118;
assign io_74 = input_119;
assign io_74 = input_120;
assign io_74 = input_121;
assign io_74 = input_122;
assign io_74 = input_123;
assign io_74 = input_124;
assign io_74 = input_125;
assign io_74 = input_126;
assign io_74 = input_127;
assign io_75 = input_75;
assign io_75 = input_76;
assign io_75 = input_77;
assign io_75 = input_78;
assign io_75 = input_79;
assign io_75 = input_80;
assign io_75 = input_81;
assign io_75 = input_82;
assign io_75 = input_83;
assign io_75 = input_84;
assign io_75 = input_85;
assign io_75 = input_86;
assign io_75 = input_87;
assign io_75 = input_88;
assign io_75 = input_89;
assign io_75 = input_90;
assign io_75 = input_91;
assign io_75 = input_92;
assign io_75 = input_93;
assign io_75 = input_94;
assign io_75 = input_95;
assign io_75 = input_96;
assign io_75 = input_97;
assign io_75 = input_98;
assign io_75 = input_99;
assign io_75 = input_100;
assign io_75 = input_101;
assign io_75 = input_102;
assign io_75 = input_103;
assign io_75 = input_104;
assign io_75 = input_105;
assign io_75 = input_106;
assign io_75 = input_107;
assign io_75 = input_108;
assign io_75 = input_109;
assign io_75 = input_110;
assign io_75 = input_111;
assign io_75 = input_112;
assign io_75 = input_113;
assign io_75 = input_114;
assign io_75 = input_115;
assign io_75 = input_116;
assign io_75 = input_117;
assign io_75 = input_118;
assign io_75 = input_119;
assign io_75 = input_120;
assign io_75 = input_121;
assign io_75 = input_122;
assign io_75 = input_123;
assign io_75 = input_124;
assign io_75 = input_125;
assign io_75 = input_126;
assign io_75 = input_127;
assign io_76 = input_76;
assign io_76 = input_77;
assign io_76 = input_78;
assign io_76 = input_79;
assign io_76 = input_80;
assign io_76 = input_81;
assign io_76 = input_82;
assign io_76 = input_83;
assign io_76 = input_84;
assign io_76 = input_85;
assign io_76 = input_86;
assign io_76 = input_87;
assign io_76 = input_88;
assign io_76 = input_89;
assign io_76 = input_90;
assign io_76 = input_91;
assign io_76 = input_92;
assign io_76 = input_93;
assign io_76 = input_94;
assign io_76 = input_95;
assign io_76 = input_96;
assign io_76 = input_97;
assign io_76 = input_98;
assign io_76 = input_99;
assign io_76 = input_100;
assign io_76 = input_101;
assign io_76 = input_102;
assign io_76 = input_103;
assign io_76 = input_104;
assign io_76 = input_105;
assign io_76 = input_106;
assign io_76 = input_107;
assign io_76 = input_108;
assign io_76 = input_109;
assign io_76 = input_110;
assign io_76 = input_111;
assign io_76 = input_112;
assign io_76 = input_113;
assign io_76 = input_114;
assign io_76 = input_115;
assign io_76 = input_116;
assign io_76 = input_117;
assign io_76 = input_118;
assign io_76 = input_119;
assign io_76 = input_120;
assign io_76 = input_121;
assign io_76 = input_122;
assign io_76 = input_123;
assign io_76 = input_124;
assign io_76 = input_125;
assign io_76 = input_126;
assign io_76 = input_127;
assign io_77 = input_77;
assign io_77 = input_78;
assign io_77 = input_79;
assign io_77 = input_80;
assign io_77 = input_81;
assign io_77 = input_82;
assign io_77 = input_83;
assign io_77 = input_84;
assign io_77 = input_85;
assign io_77 = input_86;
assign io_77 = input_87;
assign io_77 = input_88;
assign io_77 = input_89;
assign io_77 = input_90;
assign io_77 = input_91;
assign io_77 = input_92;
assign io_77 = input_93;
assign io_77 = input_94;
assign io_77 = input_95;
assign io_77 = input_96;
assign io_77 = input_97;
assign io_77 = input_98;
assign io_77 = input_99;
assign io_77 = input_100;
assign io_77 = input_101;
assign io_77 = input_102;
assign io_77 = input_103;
assign io_77 = input_104;
assign io_77 = input_105;
assign io_77 = input_106;
assign io_77 = input_107;
assign io_77 = input_108;
assign io_77 = input_109;
assign io_77 = input_110;
assign io_77 = input_111;
assign io_77 = input_112;
assign io_77 = input_113;
assign io_77 = input_114;
assign io_77 = input_115;
assign io_77 = input_116;
assign io_77 = input_117;
assign io_77 = input_118;
assign io_77 = input_119;
assign io_77 = input_120;
assign io_77 = input_121;
assign io_77 = input_122;
assign io_77 = input_123;
assign io_77 = input_124;
assign io_77 = input_125;
assign io_77 = input_126;
assign io_77 = input_127;
assign io_78 = input_78;
assign io_78 = input_79;
assign io_78 = input_80;
assign io_78 = input_81;
assign io_78 = input_82;
assign io_78 = input_83;
assign io_78 = input_84;
assign io_78 = input_85;
assign io_78 = input_86;
assign io_78 = input_87;
assign io_78 = input_88;
assign io_78 = input_89;
assign io_78 = input_90;
assign io_78 = input_91;
assign io_78 = input_92;
assign io_78 = input_93;
assign io_78 = input_94;
assign io_78 = input_95;
assign io_78 = input_96;
assign io_78 = input_97;
assign io_78 = input_98;
assign io_78 = input_99;
assign io_78 = input_100;
assign io_78 = input_101;
assign io_78 = input_102;
assign io_78 = input_103;
assign io_78 = input_104;
assign io_78 = input_105;
assign io_78 = input_106;
assign io_78 = input_107;
assign io_78 = input_108;
assign io_78 = input_109;
assign io_78 = input_110;
assign io_78 = input_111;
assign io_78 = input_112;
assign io_78 = input_113;
assign io_78 = input_114;
assign io_78 = input_115;
assign io_78 = input_116;
assign io_78 = input_117;
assign io_78 = input_118;
assign io_78 = input_119;
assign io_78 = input_120;
assign io_78 = input_121;
assign io_78 = input_122;
assign io_78 = input_123;
assign io_78 = input_124;
assign io_78 = input_125;
assign io_78 = input_126;
assign io_78 = input_127;
assign io_79 = input_79;
assign io_79 = input_80;
assign io_79 = input_81;
assign io_79 = input_82;
assign io_79 = input_83;
assign io_79 = input_84;
assign io_79 = input_85;
assign io_79 = input_86;
assign io_79 = input_87;
assign io_79 = input_88;
assign io_79 = input_89;
assign io_79 = input_90;
assign io_79 = input_91;
assign io_79 = input_92;
assign io_79 = input_93;
assign io_79 = input_94;
assign io_79 = input_95;
assign io_79 = input_96;
assign io_79 = input_97;
assign io_79 = input_98;
assign io_79 = input_99;
assign io_79 = input_100;
assign io_79 = input_101;
assign io_79 = input_102;
assign io_79 = input_103;
assign io_79 = input_104;
assign io_79 = input_105;
assign io_79 = input_106;
assign io_79 = input_107;
assign io_79 = input_108;
assign io_79 = input_109;
assign io_79 = input_110;
assign io_79 = input_111;
assign io_79 = input_112;
assign io_79 = input_113;
assign io_79 = input_114;
assign io_79 = input_115;
assign io_79 = input_116;
assign io_79 = input_117;
assign io_79 = input_118;
assign io_79 = input_119;
assign io_79 = input_120;
assign io_79 = input_121;
assign io_79 = input_122;
assign io_79 = input_123;
assign io_79 = input_124;
assign io_79 = input_125;
assign io_79 = input_126;
assign io_79 = input_127;
assign io_80 = input_80;
assign io_80 = input_81;
assign io_80 = input_82;
assign io_80 = input_83;
assign io_80 = input_84;
assign io_80 = input_85;
assign io_80 = input_86;
assign io_80 = input_87;
assign io_80 = input_88;
assign io_80 = input_89;
assign io_80 = input_90;
assign io_80 = input_91;
assign io_80 = input_92;
assign io_80 = input_93;
assign io_80 = input_94;
assign io_80 = input_95;
assign io_80 = input_96;
assign io_80 = input_97;
assign io_80 = input_98;
assign io_80 = input_99;
assign io_80 = input_100;
assign io_80 = input_101;
assign io_80 = input_102;
assign io_80 = input_103;
assign io_80 = input_104;
assign io_80 = input_105;
assign io_80 = input_106;
assign io_80 = input_107;
assign io_80 = input_108;
assign io_80 = input_109;
assign io_80 = input_110;
assign io_80 = input_111;
assign io_80 = input_112;
assign io_80 = input_113;
assign io_80 = input_114;
assign io_80 = input_115;
assign io_80 = input_116;
assign io_80 = input_117;
assign io_80 = input_118;
assign io_80 = input_119;
assign io_80 = input_120;
assign io_80 = input_121;
assign io_80 = input_122;
assign io_80 = input_123;
assign io_80 = input_124;
assign io_80 = input_125;
assign io_80 = input_126;
assign io_80 = input_127;
assign io_81 = input_81;
assign io_81 = input_82;
assign io_81 = input_83;
assign io_81 = input_84;
assign io_81 = input_85;
assign io_81 = input_86;
assign io_81 = input_87;
assign io_81 = input_88;
assign io_81 = input_89;
assign io_81 = input_90;
assign io_81 = input_91;
assign io_81 = input_92;
assign io_81 = input_93;
assign io_81 = input_94;
assign io_81 = input_95;
assign io_81 = input_96;
assign io_81 = input_97;
assign io_81 = input_98;
assign io_81 = input_99;
assign io_81 = input_100;
assign io_81 = input_101;
assign io_81 = input_102;
assign io_81 = input_103;
assign io_81 = input_104;
assign io_81 = input_105;
assign io_81 = input_106;
assign io_81 = input_107;
assign io_81 = input_108;
assign io_81 = input_109;
assign io_81 = input_110;
assign io_81 = input_111;
assign io_81 = input_112;
assign io_81 = input_113;
assign io_81 = input_114;
assign io_81 = input_115;
assign io_81 = input_116;
assign io_81 = input_117;
assign io_81 = input_118;
assign io_81 = input_119;
assign io_81 = input_120;
assign io_81 = input_121;
assign io_81 = input_122;
assign io_81 = input_123;
assign io_81 = input_124;
assign io_81 = input_125;
assign io_81 = input_126;
assign io_81 = input_127;
assign io_82 = input_82;
assign io_82 = input_83;
assign io_82 = input_84;
assign io_82 = input_85;
assign io_82 = input_86;
assign io_82 = input_87;
assign io_82 = input_88;
assign io_82 = input_89;
assign io_82 = input_90;
assign io_82 = input_91;
assign io_82 = input_92;
assign io_82 = input_93;
assign io_82 = input_94;
assign io_82 = input_95;
assign io_82 = input_96;
assign io_82 = input_97;
assign io_82 = input_98;
assign io_82 = input_99;
assign io_82 = input_100;
assign io_82 = input_101;
assign io_82 = input_102;
assign io_82 = input_103;
assign io_82 = input_104;
assign io_82 = input_105;
assign io_82 = input_106;
assign io_82 = input_107;
assign io_82 = input_108;
assign io_82 = input_109;
assign io_82 = input_110;
assign io_82 = input_111;
assign io_82 = input_112;
assign io_82 = input_113;
assign io_82 = input_114;
assign io_82 = input_115;
assign io_82 = input_116;
assign io_82 = input_117;
assign io_82 = input_118;
assign io_82 = input_119;
assign io_82 = input_120;
assign io_82 = input_121;
assign io_82 = input_122;
assign io_82 = input_123;
assign io_82 = input_124;
assign io_82 = input_125;
assign io_82 = input_126;
assign io_82 = input_127;
assign io_83 = input_83;
assign io_83 = input_84;
assign io_83 = input_85;
assign io_83 = input_86;
assign io_83 = input_87;
assign io_83 = input_88;
assign io_83 = input_89;
assign io_83 = input_90;
assign io_83 = input_91;
assign io_83 = input_92;
assign io_83 = input_93;
assign io_83 = input_94;
assign io_83 = input_95;
assign io_83 = input_96;
assign io_83 = input_97;
assign io_83 = input_98;
assign io_83 = input_99;
assign io_83 = input_100;
assign io_83 = input_101;
assign io_83 = input_102;
assign io_83 = input_103;
assign io_83 = input_104;
assign io_83 = input_105;
assign io_83 = input_106;
assign io_83 = input_107;
assign io_83 = input_108;
assign io_83 = input_109;
assign io_83 = input_110;
assign io_83 = input_111;
assign io_83 = input_112;
assign io_83 = input_113;
assign io_83 = input_114;
assign io_83 = input_115;
assign io_83 = input_116;
assign io_83 = input_117;
assign io_83 = input_118;
assign io_83 = input_119;
assign io_83 = input_120;
assign io_83 = input_121;
assign io_83 = input_122;
assign io_83 = input_123;
assign io_83 = input_124;
assign io_83 = input_125;
assign io_83 = input_126;
assign io_83 = input_127;
assign io_84 = input_84;
assign io_84 = input_85;
assign io_84 = input_86;
assign io_84 = input_87;
assign io_84 = input_88;
assign io_84 = input_89;
assign io_84 = input_90;
assign io_84 = input_91;
assign io_84 = input_92;
assign io_84 = input_93;
assign io_84 = input_94;
assign io_84 = input_95;
assign io_84 = input_96;
assign io_84 = input_97;
assign io_84 = input_98;
assign io_84 = input_99;
assign io_84 = input_100;
assign io_84 = input_101;
assign io_84 = input_102;
assign io_84 = input_103;
assign io_84 = input_104;
assign io_84 = input_105;
assign io_84 = input_106;
assign io_84 = input_107;
assign io_84 = input_108;
assign io_84 = input_109;
assign io_84 = input_110;
assign io_84 = input_111;
assign io_84 = input_112;
assign io_84 = input_113;
assign io_84 = input_114;
assign io_84 = input_115;
assign io_84 = input_116;
assign io_84 = input_117;
assign io_84 = input_118;
assign io_84 = input_119;
assign io_84 = input_120;
assign io_84 = input_121;
assign io_84 = input_122;
assign io_84 = input_123;
assign io_84 = input_124;
assign io_84 = input_125;
assign io_84 = input_126;
assign io_84 = input_127;
assign io_85 = input_85;
assign io_85 = input_86;
assign io_85 = input_87;
assign io_85 = input_88;
assign io_85 = input_89;
assign io_85 = input_90;
assign io_85 = input_91;
assign io_85 = input_92;
assign io_85 = input_93;
assign io_85 = input_94;
assign io_85 = input_95;
assign io_85 = input_96;
assign io_85 = input_97;
assign io_85 = input_98;
assign io_85 = input_99;
assign io_85 = input_100;
assign io_85 = input_101;
assign io_85 = input_102;
assign io_85 = input_103;
assign io_85 = input_104;
assign io_85 = input_105;
assign io_85 = input_106;
assign io_85 = input_107;
assign io_85 = input_108;
assign io_85 = input_109;
assign io_85 = input_110;
assign io_85 = input_111;
assign io_85 = input_112;
assign io_85 = input_113;
assign io_85 = input_114;
assign io_85 = input_115;
assign io_85 = input_116;
assign io_85 = input_117;
assign io_85 = input_118;
assign io_85 = input_119;
assign io_85 = input_120;
assign io_85 = input_121;
assign io_85 = input_122;
assign io_85 = input_123;
assign io_85 = input_124;
assign io_85 = input_125;
assign io_85 = input_126;
assign io_85 = input_127;
assign io_86 = input_86;
assign io_86 = input_87;
assign io_86 = input_88;
assign io_86 = input_89;
assign io_86 = input_90;
assign io_86 = input_91;
assign io_86 = input_92;
assign io_86 = input_93;
assign io_86 = input_94;
assign io_86 = input_95;
assign io_86 = input_96;
assign io_86 = input_97;
assign io_86 = input_98;
assign io_86 = input_99;
assign io_86 = input_100;
assign io_86 = input_101;
assign io_86 = input_102;
assign io_86 = input_103;
assign io_86 = input_104;
assign io_86 = input_105;
assign io_86 = input_106;
assign io_86 = input_107;
assign io_86 = input_108;
assign io_86 = input_109;
assign io_86 = input_110;
assign io_86 = input_111;
assign io_86 = input_112;
assign io_86 = input_113;
assign io_86 = input_114;
assign io_86 = input_115;
assign io_86 = input_116;
assign io_86 = input_117;
assign io_86 = input_118;
assign io_86 = input_119;
assign io_86 = input_120;
assign io_86 = input_121;
assign io_86 = input_122;
assign io_86 = input_123;
assign io_86 = input_124;
assign io_86 = input_125;
assign io_86 = input_126;
assign io_86 = input_127;
assign io_87 = input_87;
assign io_87 = input_88;
assign io_87 = input_89;
assign io_87 = input_90;
assign io_87 = input_91;
assign io_87 = input_92;
assign io_87 = input_93;
assign io_87 = input_94;
assign io_87 = input_95;
assign io_87 = input_96;
assign io_87 = input_97;
assign io_87 = input_98;
assign io_87 = input_99;
assign io_87 = input_100;
assign io_87 = input_101;
assign io_87 = input_102;
assign io_87 = input_103;
assign io_87 = input_104;
assign io_87 = input_105;
assign io_87 = input_106;
assign io_87 = input_107;
assign io_87 = input_108;
assign io_87 = input_109;
assign io_87 = input_110;
assign io_87 = input_111;
assign io_87 = input_112;
assign io_87 = input_113;
assign io_87 = input_114;
assign io_87 = input_115;
assign io_87 = input_116;
assign io_87 = input_117;
assign io_87 = input_118;
assign io_87 = input_119;
assign io_87 = input_120;
assign io_87 = input_121;
assign io_87 = input_122;
assign io_87 = input_123;
assign io_87 = input_124;
assign io_87 = input_125;
assign io_87 = input_126;
assign io_87 = input_127;
assign io_88 = input_88;
assign io_88 = input_89;
assign io_88 = input_90;
assign io_88 = input_91;
assign io_88 = input_92;
assign io_88 = input_93;
assign io_88 = input_94;
assign io_88 = input_95;
assign io_88 = input_96;
assign io_88 = input_97;
assign io_88 = input_98;
assign io_88 = input_99;
assign io_88 = input_100;
assign io_88 = input_101;
assign io_88 = input_102;
assign io_88 = input_103;
assign io_88 = input_104;
assign io_88 = input_105;
assign io_88 = input_106;
assign io_88 = input_107;
assign io_88 = input_108;
assign io_88 = input_109;
assign io_88 = input_110;
assign io_88 = input_111;
assign io_88 = input_112;
assign io_88 = input_113;
assign io_88 = input_114;
assign io_88 = input_115;
assign io_88 = input_116;
assign io_88 = input_117;
assign io_88 = input_118;
assign io_88 = input_119;
assign io_88 = input_120;
assign io_88 = input_121;
assign io_88 = input_122;
assign io_88 = input_123;
assign io_88 = input_124;
assign io_88 = input_125;
assign io_88 = input_126;
assign io_88 = input_127;
assign io_89 = input_89;
assign io_89 = input_90;
assign io_89 = input_91;
assign io_89 = input_92;
assign io_89 = input_93;
assign io_89 = input_94;
assign io_89 = input_95;
assign io_89 = input_96;
assign io_89 = input_97;
assign io_89 = input_98;
assign io_89 = input_99;
assign io_89 = input_100;
assign io_89 = input_101;
assign io_89 = input_102;
assign io_89 = input_103;
assign io_89 = input_104;
assign io_89 = input_105;
assign io_89 = input_106;
assign io_89 = input_107;
assign io_89 = input_108;
assign io_89 = input_109;
assign io_89 = input_110;
assign io_89 = input_111;
assign io_89 = input_112;
assign io_89 = input_113;
assign io_89 = input_114;
assign io_89 = input_115;
assign io_89 = input_116;
assign io_89 = input_117;
assign io_89 = input_118;
assign io_89 = input_119;
assign io_89 = input_120;
assign io_89 = input_121;
assign io_89 = input_122;
assign io_89 = input_123;
assign io_89 = input_124;
assign io_89 = input_125;
assign io_89 = input_126;
assign io_89 = input_127;
assign io_90 = input_90;
assign io_90 = input_91;
assign io_90 = input_92;
assign io_90 = input_93;
assign io_90 = input_94;
assign io_90 = input_95;
assign io_90 = input_96;
assign io_90 = input_97;
assign io_90 = input_98;
assign io_90 = input_99;
assign io_90 = input_100;
assign io_90 = input_101;
assign io_90 = input_102;
assign io_90 = input_103;
assign io_90 = input_104;
assign io_90 = input_105;
assign io_90 = input_106;
assign io_90 = input_107;
assign io_90 = input_108;
assign io_90 = input_109;
assign io_90 = input_110;
assign io_90 = input_111;
assign io_90 = input_112;
assign io_90 = input_113;
assign io_90 = input_114;
assign io_90 = input_115;
assign io_90 = input_116;
assign io_90 = input_117;
assign io_90 = input_118;
assign io_90 = input_119;
assign io_90 = input_120;
assign io_90 = input_121;
assign io_90 = input_122;
assign io_90 = input_123;
assign io_90 = input_124;
assign io_90 = input_125;
assign io_90 = input_126;
assign io_90 = input_127;
assign io_91 = input_91;
assign io_91 = input_92;
assign io_91 = input_93;
assign io_91 = input_94;
assign io_91 = input_95;
assign io_91 = input_96;
assign io_91 = input_97;
assign io_91 = input_98;
assign io_91 = input_99;
assign io_91 = input_100;
assign io_91 = input_101;
assign io_91 = input_102;
assign io_91 = input_103;
assign io_91 = input_104;
assign io_91 = input_105;
assign io_91 = input_106;
assign io_91 = input_107;
assign io_91 = input_108;
assign io_91 = input_109;
assign io_91 = input_110;
assign io_91 = input_111;
assign io_91 = input_112;
assign io_91 = input_113;
assign io_91 = input_114;
assign io_91 = input_115;
assign io_91 = input_116;
assign io_91 = input_117;
assign io_91 = input_118;
assign io_91 = input_119;
assign io_91 = input_120;
assign io_91 = input_121;
assign io_91 = input_122;
assign io_91 = input_123;
assign io_91 = input_124;
assign io_91 = input_125;
assign io_91 = input_126;
assign io_91 = input_127;
assign io_92 = input_92;
assign io_92 = input_93;
assign io_92 = input_94;
assign io_92 = input_95;
assign io_92 = input_96;
assign io_92 = input_97;
assign io_92 = input_98;
assign io_92 = input_99;
assign io_92 = input_100;
assign io_92 = input_101;
assign io_92 = input_102;
assign io_92 = input_103;
assign io_92 = input_104;
assign io_92 = input_105;
assign io_92 = input_106;
assign io_92 = input_107;
assign io_92 = input_108;
assign io_92 = input_109;
assign io_92 = input_110;
assign io_92 = input_111;
assign io_92 = input_112;
assign io_92 = input_113;
assign io_92 = input_114;
assign io_92 = input_115;
assign io_92 = input_116;
assign io_92 = input_117;
assign io_92 = input_118;
assign io_92 = input_119;
assign io_92 = input_120;
assign io_92 = input_121;
assign io_92 = input_122;
assign io_92 = input_123;
assign io_92 = input_124;
assign io_92 = input_125;
assign io_92 = input_126;
assign io_92 = input_127;
assign io_93 = input_93;
assign io_93 = input_94;
assign io_93 = input_95;
assign io_93 = input_96;
assign io_93 = input_97;
assign io_93 = input_98;
assign io_93 = input_99;
assign io_93 = input_100;
assign io_93 = input_101;
assign io_93 = input_102;
assign io_93 = input_103;
assign io_93 = input_104;
assign io_93 = input_105;
assign io_93 = input_106;
assign io_93 = input_107;
assign io_93 = input_108;
assign io_93 = input_109;
assign io_93 = input_110;
assign io_93 = input_111;
assign io_93 = input_112;
assign io_93 = input_113;
assign io_93 = input_114;
assign io_93 = input_115;
assign io_93 = input_116;
assign io_93 = input_117;
assign io_93 = input_118;
assign io_93 = input_119;
assign io_93 = input_120;
assign io_93 = input_121;
assign io_93 = input_122;
assign io_93 = input_123;
assign io_93 = input_124;
assign io_93 = input_125;
assign io_93 = input_126;
assign io_93 = input_127;
assign io_94 = input_94;
assign io_94 = input_95;
assign io_94 = input_96;
assign io_94 = input_97;
assign io_94 = input_98;
assign io_94 = input_99;
assign io_94 = input_100;
assign io_94 = input_101;
assign io_94 = input_102;
assign io_94 = input_103;
assign io_94 = input_104;
assign io_94 = input_105;
assign io_94 = input_106;
assign io_94 = input_107;
assign io_94 = input_108;
assign io_94 = input_109;
assign io_94 = input_110;
assign io_94 = input_111;
assign io_94 = input_112;
assign io_94 = input_113;
assign io_94 = input_114;
assign io_94 = input_115;
assign io_94 = input_116;
assign io_94 = input_117;
assign io_94 = input_118;
assign io_94 = input_119;
assign io_94 = input_120;
assign io_94 = input_121;
assign io_94 = input_122;
assign io_94 = input_123;
assign io_94 = input_124;
assign io_94 = input_125;
assign io_94 = input_126;
assign io_94 = input_127;
assign io_95 = input_95;
assign io_95 = input_96;
assign io_95 = input_97;
assign io_95 = input_98;
assign io_95 = input_99;
assign io_95 = input_100;
assign io_95 = input_101;
assign io_95 = input_102;
assign io_95 = input_103;
assign io_95 = input_104;
assign io_95 = input_105;
assign io_95 = input_106;
assign io_95 = input_107;
assign io_95 = input_108;
assign io_95 = input_109;
assign io_95 = input_110;
assign io_95 = input_111;
assign io_95 = input_112;
assign io_95 = input_113;
assign io_95 = input_114;
assign io_95 = input_115;
assign io_95 = input_116;
assign io_95 = input_117;
assign io_95 = input_118;
assign io_95 = input_119;
assign io_95 = input_120;
assign io_95 = input_121;
assign io_95 = input_122;
assign io_95 = input_123;
assign io_95 = input_124;
assign io_95 = input_125;
assign io_95 = input_126;
assign io_95 = input_127;
assign io_96 = input_96;
assign io_96 = input_97;
assign io_96 = input_98;
assign io_96 = input_99;
assign io_96 = input_100;
assign io_96 = input_101;
assign io_96 = input_102;
assign io_96 = input_103;
assign io_96 = input_104;
assign io_96 = input_105;
assign io_96 = input_106;
assign io_96 = input_107;
assign io_96 = input_108;
assign io_96 = input_109;
assign io_96 = input_110;
assign io_96 = input_111;
assign io_96 = input_112;
assign io_96 = input_113;
assign io_96 = input_114;
assign io_96 = input_115;
assign io_96 = input_116;
assign io_96 = input_117;
assign io_96 = input_118;
assign io_96 = input_119;
assign io_96 = input_120;
assign io_96 = input_121;
assign io_96 = input_122;
assign io_96 = input_123;
assign io_96 = input_124;
assign io_96 = input_125;
assign io_96 = input_126;
assign io_96 = input_127;
assign io_97 = input_97;
assign io_97 = input_98;
assign io_97 = input_99;
assign io_97 = input_100;
assign io_97 = input_101;
assign io_97 = input_102;
assign io_97 = input_103;
assign io_97 = input_104;
assign io_97 = input_105;
assign io_97 = input_106;
assign io_97 = input_107;
assign io_97 = input_108;
assign io_97 = input_109;
assign io_97 = input_110;
assign io_97 = input_111;
assign io_97 = input_112;
assign io_97 = input_113;
assign io_97 = input_114;
assign io_97 = input_115;
assign io_97 = input_116;
assign io_97 = input_117;
assign io_97 = input_118;
assign io_97 = input_119;
assign io_97 = input_120;
assign io_97 = input_121;
assign io_97 = input_122;
assign io_97 = input_123;
assign io_97 = input_124;
assign io_97 = input_125;
assign io_97 = input_126;
assign io_97 = input_127;
assign io_98 = input_98;
assign io_98 = input_99;
assign io_98 = input_100;
assign io_98 = input_101;
assign io_98 = input_102;
assign io_98 = input_103;
assign io_98 = input_104;
assign io_98 = input_105;
assign io_98 = input_106;
assign io_98 = input_107;
assign io_98 = input_108;
assign io_98 = input_109;
assign io_98 = input_110;
assign io_98 = input_111;
assign io_98 = input_112;
assign io_98 = input_113;
assign io_98 = input_114;
assign io_98 = input_115;
assign io_98 = input_116;
assign io_98 = input_117;
assign io_98 = input_118;
assign io_98 = input_119;
assign io_98 = input_120;
assign io_98 = input_121;
assign io_98 = input_122;
assign io_98 = input_123;
assign io_98 = input_124;
assign io_98 = input_125;
assign io_98 = input_126;
assign io_98 = input_127;
assign io_99 = input_99;
assign io_99 = input_100;
assign io_99 = input_101;
assign io_99 = input_102;
assign io_99 = input_103;
assign io_99 = input_104;
assign io_99 = input_105;
assign io_99 = input_106;
assign io_99 = input_107;
assign io_99 = input_108;
assign io_99 = input_109;
assign io_99 = input_110;
assign io_99 = input_111;
assign io_99 = input_112;
assign io_99 = input_113;
assign io_99 = input_114;
assign io_99 = input_115;
assign io_99 = input_116;
assign io_99 = input_117;
assign io_99 = input_118;
assign io_99 = input_119;
assign io_99 = input_120;
assign io_99 = input_121;
assign io_99 = input_122;
assign io_99 = input_123;
assign io_99 = input_124;
assign io_99 = input_125;
assign io_99 = input_126;
assign io_99 = input_127;
assign io_100 = input_100;
assign io_100 = input_101;
assign io_100 = input_102;
assign io_100 = input_103;
assign io_100 = input_104;
assign io_100 = input_105;
assign io_100 = input_106;
assign io_100 = input_107;
assign io_100 = input_108;
assign io_100 = input_109;
assign io_100 = input_110;
assign io_100 = input_111;
assign io_100 = input_112;
assign io_100 = input_113;
assign io_100 = input_114;
assign io_100 = input_115;
assign io_100 = input_116;
assign io_100 = input_117;
assign io_100 = input_118;
assign io_100 = input_119;
assign io_100 = input_120;
assign io_100 = input_121;
assign io_100 = input_122;
assign io_100 = input_123;
assign io_100 = input_124;
assign io_100 = input_125;
assign io_100 = input_126;
assign io_100 = input_127;
assign io_101 = input_101;
assign io_101 = input_102;
assign io_101 = input_103;
assign io_101 = input_104;
assign io_101 = input_105;
assign io_101 = input_106;
assign io_101 = input_107;
assign io_101 = input_108;
assign io_101 = input_109;
assign io_101 = input_110;
assign io_101 = input_111;
assign io_101 = input_112;
assign io_101 = input_113;
assign io_101 = input_114;
assign io_101 = input_115;
assign io_101 = input_116;
assign io_101 = input_117;
assign io_101 = input_118;
assign io_101 = input_119;
assign io_101 = input_120;
assign io_101 = input_121;
assign io_101 = input_122;
assign io_101 = input_123;
assign io_101 = input_124;
assign io_101 = input_125;
assign io_101 = input_126;
assign io_101 = input_127;
assign io_102 = input_102;
assign io_102 = input_103;
assign io_102 = input_104;
assign io_102 = input_105;
assign io_102 = input_106;
assign io_102 = input_107;
assign io_102 = input_108;
assign io_102 = input_109;
assign io_102 = input_110;
assign io_102 = input_111;
assign io_102 = input_112;
assign io_102 = input_113;
assign io_102 = input_114;
assign io_102 = input_115;
assign io_102 = input_116;
assign io_102 = input_117;
assign io_102 = input_118;
assign io_102 = input_119;
assign io_102 = input_120;
assign io_102 = input_121;
assign io_102 = input_122;
assign io_102 = input_123;
assign io_102 = input_124;
assign io_102 = input_125;
assign io_102 = input_126;
assign io_102 = input_127;
assign io_103 = input_103;
assign io_103 = input_104;
assign io_103 = input_105;
assign io_103 = input_106;
assign io_103 = input_107;
assign io_103 = input_108;
assign io_103 = input_109;
assign io_103 = input_110;
assign io_103 = input_111;
assign io_103 = input_112;
assign io_103 = input_113;
assign io_103 = input_114;
assign io_103 = input_115;
assign io_103 = input_116;
assign io_103 = input_117;
assign io_103 = input_118;
assign io_103 = input_119;
assign io_103 = input_120;
assign io_103 = input_121;
assign io_103 = input_122;
assign io_103 = input_123;
assign io_103 = input_124;
assign io_103 = input_125;
assign io_103 = input_126;
assign io_103 = input_127;
assign io_104 = input_104;
assign io_104 = input_105;
assign io_104 = input_106;
assign io_104 = input_107;
assign io_104 = input_108;
assign io_104 = input_109;
assign io_104 = input_110;
assign io_104 = input_111;
assign io_104 = input_112;
assign io_104 = input_113;
assign io_104 = input_114;
assign io_104 = input_115;
assign io_104 = input_116;
assign io_104 = input_117;
assign io_104 = input_118;
assign io_104 = input_119;
assign io_104 = input_120;
assign io_104 = input_121;
assign io_104 = input_122;
assign io_104 = input_123;
assign io_104 = input_124;
assign io_104 = input_125;
assign io_104 = input_126;
assign io_104 = input_127;
assign io_105 = input_105;
assign io_105 = input_106;
assign io_105 = input_107;
assign io_105 = input_108;
assign io_105 = input_109;
assign io_105 = input_110;
assign io_105 = input_111;
assign io_105 = input_112;
assign io_105 = input_113;
assign io_105 = input_114;
assign io_105 = input_115;
assign io_105 = input_116;
assign io_105 = input_117;
assign io_105 = input_118;
assign io_105 = input_119;
assign io_105 = input_120;
assign io_105 = input_121;
assign io_105 = input_122;
assign io_105 = input_123;
assign io_105 = input_124;
assign io_105 = input_125;
assign io_105 = input_126;
assign io_105 = input_127;
assign io_106 = input_106;
assign io_106 = input_107;
assign io_106 = input_108;
assign io_106 = input_109;
assign io_106 = input_110;
assign io_106 = input_111;
assign io_106 = input_112;
assign io_106 = input_113;
assign io_106 = input_114;
assign io_106 = input_115;
assign io_106 = input_116;
assign io_106 = input_117;
assign io_106 = input_118;
assign io_106 = input_119;
assign io_106 = input_120;
assign io_106 = input_121;
assign io_106 = input_122;
assign io_106 = input_123;
assign io_106 = input_124;
assign io_106 = input_125;
assign io_106 = input_126;
assign io_106 = input_127;
assign io_107 = input_107;
assign io_107 = input_108;
assign io_107 = input_109;
assign io_107 = input_110;
assign io_107 = input_111;
assign io_107 = input_112;
assign io_107 = input_113;
assign io_107 = input_114;
assign io_107 = input_115;
assign io_107 = input_116;
assign io_107 = input_117;
assign io_107 = input_118;
assign io_107 = input_119;
assign io_107 = input_120;
assign io_107 = input_121;
assign io_107 = input_122;
assign io_107 = input_123;
assign io_107 = input_124;
assign io_107 = input_125;
assign io_107 = input_126;
assign io_107 = input_127;
assign io_108 = input_108;
assign io_108 = input_109;
assign io_108 = input_110;
assign io_108 = input_111;
assign io_108 = input_112;
assign io_108 = input_113;
assign io_108 = input_114;
assign io_108 = input_115;
assign io_108 = input_116;
assign io_108 = input_117;
assign io_108 = input_118;
assign io_108 = input_119;
assign io_108 = input_120;
assign io_108 = input_121;
assign io_108 = input_122;
assign io_108 = input_123;
assign io_108 = input_124;
assign io_108 = input_125;
assign io_108 = input_126;
assign io_108 = input_127;
assign io_109 = input_109;
assign io_109 = input_110;
assign io_109 = input_111;
assign io_109 = input_112;
assign io_109 = input_113;
assign io_109 = input_114;
assign io_109 = input_115;
assign io_109 = input_116;
assign io_109 = input_117;
assign io_109 = input_118;
assign io_109 = input_119;
assign io_109 = input_120;
assign io_109 = input_121;
assign io_109 = input_122;
assign io_109 = input_123;
assign io_109 = input_124;
assign io_109 = input_125;
assign io_109 = input_126;
assign io_109 = input_127;
assign io_110 = input_110;
assign io_110 = input_111;
assign io_110 = input_112;
assign io_110 = input_113;
assign io_110 = input_114;
assign io_110 = input_115;
assign io_110 = input_116;
assign io_110 = input_117;
assign io_110 = input_118;
assign io_110 = input_119;
assign io_110 = input_120;
assign io_110 = input_121;
assign io_110 = input_122;
assign io_110 = input_123;
assign io_110 = input_124;
assign io_110 = input_125;
assign io_110 = input_126;
assign io_110 = input_127;
assign io_111 = input_111;
assign io_111 = input_112;
assign io_111 = input_113;
assign io_111 = input_114;
assign io_111 = input_115;
assign io_111 = input_116;
assign io_111 = input_117;
assign io_111 = input_118;
assign io_111 = input_119;
assign io_111 = input_120;
assign io_111 = input_121;
assign io_111 = input_122;
assign io_111 = input_123;
assign io_111 = input_124;
assign io_111 = input_125;
assign io_111 = input_126;
assign io_111 = input_127;
assign io_112 = input_112;
assign io_112 = input_113;
assign io_112 = input_114;
assign io_112 = input_115;
assign io_112 = input_116;
assign io_112 = input_117;
assign io_112 = input_118;
assign io_112 = input_119;
assign io_112 = input_120;
assign io_112 = input_121;
assign io_112 = input_122;
assign io_112 = input_123;
assign io_112 = input_124;
assign io_112 = input_125;
assign io_112 = input_126;
assign io_112 = input_127;
assign io_113 = input_113;
assign io_113 = input_114;
assign io_113 = input_115;
assign io_113 = input_116;
assign io_113 = input_117;
assign io_113 = input_118;
assign io_113 = input_119;
assign io_113 = input_120;
assign io_113 = input_121;
assign io_113 = input_122;
assign io_113 = input_123;
assign io_113 = input_124;
assign io_113 = input_125;
assign io_113 = input_126;
assign io_113 = input_127;
assign io_114 = input_114;
assign io_114 = input_115;
assign io_114 = input_116;
assign io_114 = input_117;
assign io_114 = input_118;
assign io_114 = input_119;
assign io_114 = input_120;
assign io_114 = input_121;
assign io_114 = input_122;
assign io_114 = input_123;
assign io_114 = input_124;
assign io_114 = input_125;
assign io_114 = input_126;
assign io_114 = input_127;
assign io_115 = input_115;
assign io_115 = input_116;
assign io_115 = input_117;
assign io_115 = input_118;
assign io_115 = input_119;
assign io_115 = input_120;
assign io_115 = input_121;
assign io_115 = input_122;
assign io_115 = input_123;
assign io_115 = input_124;
assign io_115 = input_125;
assign io_115 = input_126;
assign io_115 = input_127;
assign io_116 = input_116;
assign io_116 = input_117;
assign io_116 = input_118;
assign io_116 = input_119;
assign io_116 = input_120;
assign io_116 = input_121;
assign io_116 = input_122;
assign io_116 = input_123;
assign io_116 = input_124;
assign io_116 = input_125;
assign io_116 = input_126;
assign io_116 = input_127;
assign io_117 = input_117;
assign io_117 = input_118;
assign io_117 = input_119;
assign io_117 = input_120;
assign io_117 = input_121;
assign io_117 = input_122;
assign io_117 = input_123;
assign io_117 = input_124;
assign io_117 = input_125;
assign io_117 = input_126;
assign io_117 = input_127;
assign io_118 = input_118;
assign io_118 = input_119;
assign io_118 = input_120;
assign io_118 = input_121;
assign io_118 = input_122;
assign io_118 = input_123;
assign io_118 = input_124;
assign io_118 = input_125;
assign io_118 = input_126;
assign io_118 = input_127;
assign io_119 = input_119;
assign io_119 = input_120;
assign io_119 = input_121;
assign io_119 = input_122;
assign io_119 = input_123;
assign io_119 = input_124;
assign io_119 = input_125;
assign io_119 = input_126;
assign io_119 = input_127;
assign io_120 = input_120;
assign io_120 = input_121;
assign io_120 = input_122;
assign io_120 = input_123;
assign io_120 = input_124;
assign io_120 = input_125;
assign io_120 = input_126;
assign io_120 = input_127;
assign io_121 = input_121;
assign io_121 = input_122;
assign io_121 = input_123;
assign io_121 = input_124;
assign io_121 = input_125;
assign io_121 = input_126;
assign io_121 = input_127;
assign io_122 = input_122;
assign io_122 = input_123;
assign io_122 = input_124;
assign io_122 = input_125;
assign io_122 = input_126;
assign io_122 = input_127;
assign io_123 = input_123;
assign io_123 = input_124;
assign io_123 = input_125;
assign io_123 = input_126;
assign io_123 = input_127;
assign io_124 = input_124;
assign io_124 = input_125;
assign io_124 = input_126;
assign io_124 = input_127;
assign io_125 = input_125;
assign io_125 = input_126;
assign io_125 = input_127;
assign io_126 = input_126;
assign io_126 = input_127;
assign io_127 = input_127;
endmodule
