module tutte12();
	mixer m_0(.a(e_0_1), .b(e_0_2), .y(e_0_3));
	mixer m_1(.a(e_0_1), .b(e_1_120), .y(e_1_121));
	mixer m_2(.a(e_0_2), .b(e_2_122), .y(e_2_125));
	mixer m_3(.a(e_0_3), .b(e_3_123), .y(e_3_124));
	mixer m_4(.a(e_4_36), .b(e_4_80), .y(e_4_81));
	mixer m_5(.a(e_5_36), .b(e_5_82), .y(e_5_83));
	mixer m_6(.a(e_6_37), .b(e_6_76), .y(e_6_79));
	mixer m_7(.a(e_7_37), .b(e_7_77), .y(e_7_78));
	mixer m_8(.a(e_8_38), .b(e_8_43), .y(e_8_44));
	mixer m_9(.a(e_9_38), .b(e_9_45), .y(e_9_46));
	mixer m_10(.a(e_10_39), .b(e_10_43), .y(e_10_47));
	mixer m_11(.a(e_11_42), .b(e_11_44), .y(e_11_49));
	mixer m_12(.a(e_12_40), .b(e_12_45), .y(e_12_50));
	mixer m_13(.a(e_13_41), .b(e_13_46), .y(e_13_48));
	mixer m_14(.a(e_14_40), .b(e_14_52), .y(e_14_56));
	mixer m_15(.a(e_15_42), .b(e_15_53), .y(e_15_56));
	mixer m_16(.a(e_16_39), .b(e_16_54), .y(e_16_55));
	mixer m_17(.a(e_17_41), .b(e_17_51), .y(e_17_55));
	mixer m_18(.a(e_18_47), .b(e_18_52), .y(e_18_81));
	mixer m_19(.a(e_19_50), .b(e_19_54), .y(e_19_83));
	mixer m_20(.a(e_20_48), .b(e_20_53), .y(e_20_82));
	mixer m_21(.a(e_21_49), .b(e_21_51), .y(e_21_80));
	mixer m_22(.a(e_22_57), .b(e_22_58), .y(e_22_61));
	mixer m_23(.a(e_23_57), .b(e_23_59), .y(e_23_60));
	mixer m_24(.a(e_24_65), .b(e_24_67), .y(e_24_69));
	mixer m_25(.a(e_25_64), .b(e_25_67), .y(e_25_71));
	mixer m_26(.a(e_26_62), .b(e_26_66), .y(e_26_68));
	mixer m_27(.a(e_27_63), .b(e_27_66), .y(e_27_70));
	mixer m_28(.a(e_28_60), .b(e_28_65), .y(e_28_73));
	mixer m_29(.a(e_29_58), .b(e_29_62), .y(e_29_74));
	mixer m_30(.a(e_30_61), .b(e_30_64), .y(e_30_72));
	mixer m_31(.a(e_31_59), .b(e_31_63), .y(e_31_75));
	mixer m_32(.a(e_32_68), .b(e_32_73), .y(e_32_76));
	mixer m_33(.a(e_33_69), .b(e_33_74), .y(e_33_77));
	mixer m_34(.a(e_34_71), .b(e_34_75), .y(e_34_79));
	mixer m_35(.a(e_35_70), .b(e_35_72), .y(e_35_78));
	mixer m_36(.a(e_4_36), .b(e_5_36), .y(e_36_84));
	mixer m_37(.a(e_6_37), .b(e_7_37), .y(e_37_84));
	mixer m_38(.a(e_8_38), .b(e_9_38), .y(e_38_85));
	mixer m_39(.a(e_10_39), .b(e_16_39), .y(e_39_106));
	mixer m_40(.a(e_12_40), .b(e_14_40), .y(e_40_104));
	mixer m_41(.a(e_13_41), .b(e_17_41), .y(e_41_105));
	mixer m_42(.a(e_11_42), .b(e_15_42), .y(e_42_107));
	mixer m_43(.a(e_8_43), .b(e_10_43), .y(e_43_96));
	mixer m_44(.a(e_8_44), .b(e_11_44), .y(e_44_97));
	mixer m_45(.a(e_9_45), .b(e_12_45), .y(e_45_99));
	mixer m_46(.a(e_9_46), .b(e_13_46), .y(e_46_98));
	mixer m_47(.a(e_10_47), .b(e_18_47), .y(e_47_100));
	mixer m_48(.a(e_13_48), .b(e_20_48), .y(e_48_103));
	mixer m_49(.a(e_11_49), .b(e_21_49), .y(e_49_102));
	mixer m_50(.a(e_12_50), .b(e_19_50), .y(e_50_101));
	mixer m_51(.a(e_17_51), .b(e_21_51), .y(e_51_92));
	mixer m_52(.a(e_14_52), .b(e_18_52), .y(e_52_93));
	mixer m_53(.a(e_15_53), .b(e_20_53), .y(e_53_94));
	mixer m_54(.a(e_16_54), .b(e_19_54), .y(e_54_95));
	mixer m_55(.a(e_16_55), .b(e_17_55), .y(e_55_87));
	mixer m_56(.a(e_14_56), .b(e_15_56), .y(e_56_86));
	mixer m_57(.a(e_22_57), .b(e_23_57), .y(e_57_85));
	mixer m_58(.a(e_22_58), .b(e_29_58), .y(e_58_94));
	mixer m_59(.a(e_23_59), .b(e_31_59), .y(e_59_93));
	mixer m_60(.a(e_23_60), .b(e_28_60), .y(e_60_95));
	mixer m_61(.a(e_22_61), .b(e_30_61), .y(e_61_92));
	mixer m_62(.a(e_26_62), .b(e_29_62), .y(e_62_91));
	mixer m_63(.a(e_27_63), .b(e_31_63), .y(e_63_88));
	mixer m_64(.a(e_25_64), .b(e_30_64), .y(e_64_89));
	mixer m_65(.a(e_24_65), .b(e_28_65), .y(e_65_90));
	mixer m_66(.a(e_26_66), .b(e_27_66), .y(e_66_87));
	mixer m_67(.a(e_24_67), .b(e_25_67), .y(e_67_86));
	mixer m_68(.a(e_26_68), .b(e_32_68), .y(e_68_97));
	mixer m_69(.a(e_24_69), .b(e_33_69), .y(e_69_96));
	mixer m_70(.a(e_27_70), .b(e_35_70), .y(e_70_99));
	mixer m_71(.a(e_25_71), .b(e_34_71), .y(e_71_98));
	mixer m_72(.a(e_30_72), .b(e_35_72), .y(e_72_100));
	mixer m_73(.a(e_28_73), .b(e_32_73), .y(e_73_103));
	mixer m_74(.a(e_29_74), .b(e_33_74), .y(e_74_101));
	mixer m_75(.a(e_31_75), .b(e_34_75), .y(e_75_102));
	mixer m_76(.a(e_6_76), .b(e_32_76), .y(e_76_104));
	mixer m_77(.a(e_7_77), .b(e_33_77), .y(e_77_105));
	mixer m_78(.a(e_7_78), .b(e_35_78), .y(e_78_107));
	mixer m_79(.a(e_6_79), .b(e_34_79), .y(e_79_106));
	mixer m_80(.a(e_4_80), .b(e_21_80), .y(e_80_90));
	mixer m_81(.a(e_4_81), .b(e_18_81), .y(e_81_91));
	mixer m_82(.a(e_5_82), .b(e_20_82), .y(e_82_88));
	mixer m_83(.a(e_5_83), .b(e_19_83), .y(e_83_89));
	mixer m_84(.a(e_36_84), .b(e_37_84), .y(e_84_108));
	mixer m_85(.a(e_38_85), .b(e_57_85), .y(e_85_108));
	mixer m_86(.a(e_56_86), .b(e_67_86), .y(e_86_109));
	mixer m_87(.a(e_55_87), .b(e_66_87), .y(e_87_109));
	mixer m_88(.a(e_63_88), .b(e_82_88), .y(e_88_112));
	mixer m_89(.a(e_64_89), .b(e_83_89), .y(e_89_113));
	mixer m_90(.a(e_65_90), .b(e_80_90), .y(e_90_115));
	mixer m_91(.a(e_62_91), .b(e_81_91), .y(e_91_114));
	mixer m_92(.a(e_51_92), .b(e_61_92), .y(e_92_116));
	mixer m_93(.a(e_52_93), .b(e_59_93), .y(e_93_117));
	mixer m_94(.a(e_53_94), .b(e_58_94), .y(e_94_119));
	mixer m_95(.a(e_54_95), .b(e_60_95), .y(e_95_118));
	mixer m_96(.a(e_43_96), .b(e_69_96), .y(e_96_112));
	mixer m_97(.a(e_44_97), .b(e_68_97), .y(e_97_113));
	mixer m_98(.a(e_46_98), .b(e_71_98), .y(e_98_114));
	mixer m_99(.a(e_45_99), .b(e_70_99), .y(e_99_115));
	mixer m_100(.a(e_47_100), .b(e_72_100), .y(e_100_110));
	mixer m_101(.a(e_50_101), .b(e_74_101), .y(e_101_111));
	mixer m_102(.a(e_49_102), .b(e_75_102), .y(e_102_111));
	mixer m_103(.a(e_48_103), .b(e_73_103), .y(e_103_110));
	mixer m_104(.a(e_40_104), .b(e_76_104), .y(e_104_116));
	mixer m_105(.a(e_41_105), .b(e_77_105), .y(e_105_117));
	mixer m_106(.a(e_39_106), .b(e_79_106), .y(e_106_119));
	mixer m_107(.a(e_42_107), .b(e_78_107), .y(e_107_118));
	mixer m_108(.a(e_84_108), .b(e_85_108), .y(e_108_120));
	mixer m_109(.a(e_86_109), .b(e_87_109), .y(e_109_120));
	mixer m_110(.a(e_100_110), .b(e_103_110), .y(e_110_121));
	mixer m_111(.a(e_101_111), .b(e_102_111), .y(e_111_121));
	mixer m_112(.a(e_88_112), .b(e_96_112), .y(e_112_122));
	mixer m_113(.a(e_89_113), .b(e_97_113), .y(e_113_123));
	mixer m_114(.a(e_91_114), .b(e_98_114), .y(e_114_125));
	mixer m_115(.a(e_90_115), .b(e_99_115), .y(e_115_124));
	mixer m_116(.a(e_92_116), .b(e_104_116), .y(e_116_122));
	mixer m_117(.a(e_93_117), .b(e_105_117), .y(e_117_123));
	mixer m_118(.a(e_95_118), .b(e_107_118), .y(e_118_125));
	mixer m_119(.a(e_94_119), .b(e_106_119), .y(e_119_124));
	mixer m_120(.a(e_1_120), .b(e_108_120), .y(e_109_120));
	mixer m_121(.a(e_1_121), .b(e_110_121), .y(e_111_121));
	mixer m_122(.a(e_2_122), .b(e_112_122), .y(e_116_122));
	mixer m_123(.a(e_3_123), .b(e_113_123), .y(e_117_123));
	mixer m_124(.a(e_3_124), .b(e_115_124), .y(e_119_124));
	mixer m_125(.a(e_2_125), .b(e_114_125), .y(e_118_125));
wire e_0_1,
	e_0_2,
	e_0_3,
	e_1_120,
	e_1_121,
	e_2_122,
	e_2_125,
	e_3_123,
	e_3_124,
	e_4_36,
	e_4_80,
	e_4_81,
	e_5_36,
	e_5_82,
	e_5_83,
	e_6_37,
	e_6_76,
	e_6_79,
	e_7_37,
	e_7_77,
	e_7_78,
	e_8_38,
	e_8_43,
	e_8_44,
	e_9_38,
	e_9_45,
	e_9_46,
	e_10_39,
	e_10_43,
	e_10_47,
	e_11_42,
	e_11_44,
	e_11_49,
	e_12_40,
	e_12_45,
	e_12_50,
	e_13_41,
	e_13_46,
	e_13_48,
	e_14_40,
	e_14_52,
	e_14_56,
	e_15_42,
	e_15_53,
	e_15_56,
	e_16_39,
	e_16_54,
	e_16_55,
	e_17_41,
	e_17_51,
	e_17_55,
	e_18_47,
	e_18_52,
	e_18_81,
	e_19_50,
	e_19_54,
	e_19_83,
	e_20_48,
	e_20_53,
	e_20_82,
	e_21_49,
	e_21_51,
	e_21_80,
	e_22_57,
	e_22_58,
	e_22_61,
	e_23_57,
	e_23_59,
	e_23_60,
	e_24_65,
	e_24_67,
	e_24_69,
	e_25_64,
	e_25_67,
	e_25_71,
	e_26_62,
	e_26_66,
	e_26_68,
	e_27_63,
	e_27_66,
	e_27_70,
	e_28_60,
	e_28_65,
	e_28_73,
	e_29_58,
	e_29_62,
	e_29_74,
	e_30_61,
	e_30_64,
	e_30_72,
	e_31_59,
	e_31_63,
	e_31_75,
	e_32_68,
	e_32_73,
	e_32_76,
	e_33_69,
	e_33_74,
	e_33_77,
	e_34_71,
	e_34_75,
	e_34_79,
	e_35_70,
	e_35_72,
	e_35_78,
	e_36_84,
	e_37_84,
	e_38_85,
	e_39_106,
	e_40_104,
	e_41_105,
	e_42_107,
	e_43_96,
	e_44_97,
	e_45_99,
	e_46_98,
	e_47_100,
	e_48_103,
	e_49_102,
	e_50_101,
	e_51_92,
	e_52_93,
	e_53_94,
	e_54_95,
	e_55_87,
	e_56_86,
	e_57_85,
	e_58_94,
	e_59_93,
	e_60_95,
	e_61_92,
	e_62_91,
	e_63_88,
	e_64_89,
	e_65_90,
	e_66_87,
	e_67_86,
	e_68_97,
	e_69_96,
	e_70_99,
	e_71_98,
	e_72_100,
	e_73_103,
	e_74_101,
	e_75_102,
	e_76_104,
	e_77_105,
	e_78_107,
	e_79_106,
	e_80_90,
	e_81_91,
	e_82_88,
	e_83_89,
	e_84_108,
	e_85_108,
	e_86_109,
	e_87_109,
	e_88_112,
	e_89_113,
	e_90_115,
	e_91_114,
	e_92_116,
	e_93_117,
	e_94_119,
	e_95_118,
	e_96_112,
	e_97_113,
	e_98_114,
	e_99_115,
	e_100_110,
	e_101_111,
	e_102_111,
	e_103_110,
	e_104_116,
	e_105_117,
	e_106_119,
	e_107_118,
	e_108_120,
	e_109_120,
	e_110_121,
	e_111_121,
	e_112_122,
	e_113_123,
	e_114_125,
	e_115_124,
	e_116_122,
	e_117_123,
	e_118_125,
	e_119_124;
endmodule
