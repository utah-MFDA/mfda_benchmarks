module fanout2_braid_8_16 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_1_7, output_1_0, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_0), .y(output_0_7));
wire output_2_7, output_2_0, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_0), .y(output_1_7));
wire output_3_7, output_3_0, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_0), .y(output_2_7));
wire output_4_7, output_4_0, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_0), .y(output_3_7));
wire output_5_7, output_5_0, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_0), .y(output_4_7));
wire output_6_7, output_6_0, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_0), .y(output_5_7));
wire output_7_7, output_7_0, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_0), .y(output_6_7));
wire output_8_7, output_8_0, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_0), .y(output_7_7));
wire output_1_8, output_1_1, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_1), .y(output_0_8));
wire output_2_8, output_2_1, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_1), .y(output_1_8));
wire output_3_8, output_3_1, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_1), .y(output_2_8));
wire output_4_8, output_4_1, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_1), .y(output_3_8));
wire output_5_8, output_5_1, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_1), .y(output_4_8));
wire output_6_8, output_6_1, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_1), .y(output_5_8));
wire output_7_8, output_7_1, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_1), .y(output_6_8));
wire output_8_8, output_8_1, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_1), .y(output_7_8));
wire output_1_9, output_1_2, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_2), .y(output_0_9));
wire output_2_9, output_2_2, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_2), .y(output_1_9));
wire output_3_9, output_3_2, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_2), .y(output_2_9));
wire output_4_9, output_4_2, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_2), .y(output_3_9));
wire output_5_9, output_5_2, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_2), .y(output_4_9));
wire output_6_9, output_6_2, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_2), .y(output_5_9));
wire output_7_9, output_7_2, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_2), .y(output_6_9));
wire output_8_9, output_8_2, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_2), .y(output_7_9));
wire output_1_10, output_1_3, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_3), .y(output_0_10));
wire output_2_10, output_2_3, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_3), .y(output_1_10));
wire output_3_10, output_3_3, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_3), .y(output_2_10));
wire output_4_10, output_4_3, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_3), .y(output_3_10));
wire output_5_10, output_5_3, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_3), .y(output_4_10));
wire output_6_10, output_6_3, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_3), .y(output_5_10));
wire output_7_10, output_7_3, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_3), .y(output_6_10));
wire output_8_10, output_8_3, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_3), .y(output_7_10));
wire output_1_11, output_1_4, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_4), .y(output_0_11));
wire output_2_11, output_2_4, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_4), .y(output_1_11));
wire output_3_11, output_3_4, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_4), .y(output_2_11));
wire output_4_11, output_4_4, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_4), .y(output_3_11));
wire output_5_11, output_5_4, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_4), .y(output_4_11));
wire output_6_11, output_6_4, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_4), .y(output_5_11));
wire output_7_11, output_7_4, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_4), .y(output_6_11));
wire output_8_11, output_8_4, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_4), .y(output_7_11));
wire output_1_12, output_1_5, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_5), .y(output_0_12));
wire output_2_12, output_2_5, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_5), .y(output_1_12));
wire output_3_12, output_3_5, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_5), .y(output_2_12));
wire output_4_12, output_4_5, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_5), .y(output_3_12));
wire output_5_12, output_5_5, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_5), .y(output_4_12));
wire output_6_12, output_6_5, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_5), .y(output_5_12));
wire output_7_12, output_7_5, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_5), .y(output_6_12));
wire output_8_12, output_8_5, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_5), .y(output_7_12));
wire output_1_13, output_1_6, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_6), .y(output_0_13));
wire output_2_13, output_2_6, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_6), .y(output_1_13));
wire output_3_13, output_3_6, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_6), .y(output_2_13));
wire output_4_13, output_4_6, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_6), .y(output_3_13));
wire output_5_13, output_5_6, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_6), .y(output_4_13));
wire output_6_13, output_6_6, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_6), .y(output_5_13));
wire output_7_13, output_7_6, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_6), .y(output_6_13));
wire output_8_13, output_8_6, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_6), .y(output_7_13));
wire output_1_14, output_1_7, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_7), .y(output_0_14));
wire output_2_14, output_2_7, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_7), .y(output_1_14));
wire output_3_14, output_3_7, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_7), .y(output_2_14));
wire output_4_14, output_4_7, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_7), .y(output_3_14));
wire output_5_14, output_5_7, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_7), .y(output_4_14));
wire output_6_14, output_6_7, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_7), .y(output_5_14));
wire output_7_14, output_7_7, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_7), .y(output_6_14));
wire output_8_14, output_8_7, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_7), .y(output_7_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
assign output_0 = output_0_0;
wire output_0_16;
assign output_0_16 = input_0;
assign output_1 = output_1_0;
wire output_1_16;
assign output_1_16 = input_1;
assign output_2 = output_2_0;
wire output_2_16;
assign output_2_16 = input_2;
assign output_3 = output_3_0;
wire output_3_16;
assign output_3_16 = input_3;
assign output_4 = output_4_0;
wire output_4_16;
assign output_4_16 = input_4;
assign output_5 = output_5_0;
wire output_5_16;
assign output_5_16 = input_5;
assign output_6 = output_6_0;
wire output_6_16;
assign output_6_16 = input_6;
assign output_7 = output_7_0;
wire output_7_16;
assign output_7_16 = input_7;
endmodule
