module chain_4 (
inout k0, k4
);
wire {wires};
chamber ch0 (.in(k0), .out(k1)
chamber ch1 (.in(k1), .out(k2)
chamber ch2 (.in(k2), .out(k3)
chamber ch3 (.in(k3), .out(k4)
endmodule
