module complete_96 (
inout io_0,inout io_1,inout io_2,inout io_3,inout io_4,inout io_5,inout io_6,inout io_7,inout io_8,inout io_9,inout io_10,inout io_11,inout io_12,inout io_13,inout io_14,inout io_15,inout io_16,inout io_17,inout io_18,inout io_19,inout io_20,inout io_21,inout io_22,inout io_23,inout io_24,inout io_25,inout io_26,inout io_27,inout io_28,inout io_29,inout io_30,inout io_31,inout io_32,inout io_33,inout io_34,inout io_35,inout io_36,inout io_37,inout io_38,inout io_39,inout io_40,inout io_41,inout io_42,inout io_43,inout io_44,inout io_45,inout io_46,inout io_47,inout io_48,inout io_49,inout io_50,inout io_51,inout io_52,inout io_53,inout io_54,inout io_55,inout io_56,inout io_57,inout io_58,inout io_59,inout io_60,inout io_61,inout io_62,inout io_63,inout io_64,inout io_65,inout io_66,inout io_67,inout io_68,inout io_69,inout io_70,inout io_71,inout io_72,inout io_73,inout io_74,inout io_75,inout io_76,inout io_77,inout io_78,inout io_79,inout io_80,inout io_81,inout io_82,inout io_83,inout io_84,inout io_85,inout io_86,inout io_87,inout io_88,inout io_89,inout io_90,inout io_91,inout io_92,inout io_93,inout io_94,inout io_95
);
assign io_0 = input_0;
assign io_0 = input_1;
assign io_0 = input_2;
assign io_0 = input_3;
assign io_0 = input_4;
assign io_0 = input_5;
assign io_0 = input_6;
assign io_0 = input_7;
assign io_0 = input_8;
assign io_0 = input_9;
assign io_0 = input_10;
assign io_0 = input_11;
assign io_0 = input_12;
assign io_0 = input_13;
assign io_0 = input_14;
assign io_0 = input_15;
assign io_0 = input_16;
assign io_0 = input_17;
assign io_0 = input_18;
assign io_0 = input_19;
assign io_0 = input_20;
assign io_0 = input_21;
assign io_0 = input_22;
assign io_0 = input_23;
assign io_0 = input_24;
assign io_0 = input_25;
assign io_0 = input_26;
assign io_0 = input_27;
assign io_0 = input_28;
assign io_0 = input_29;
assign io_0 = input_30;
assign io_0 = input_31;
assign io_0 = input_32;
assign io_0 = input_33;
assign io_0 = input_34;
assign io_0 = input_35;
assign io_0 = input_36;
assign io_0 = input_37;
assign io_0 = input_38;
assign io_0 = input_39;
assign io_0 = input_40;
assign io_0 = input_41;
assign io_0 = input_42;
assign io_0 = input_43;
assign io_0 = input_44;
assign io_0 = input_45;
assign io_0 = input_46;
assign io_0 = input_47;
assign io_0 = input_48;
assign io_0 = input_49;
assign io_0 = input_50;
assign io_0 = input_51;
assign io_0 = input_52;
assign io_0 = input_53;
assign io_0 = input_54;
assign io_0 = input_55;
assign io_0 = input_56;
assign io_0 = input_57;
assign io_0 = input_58;
assign io_0 = input_59;
assign io_0 = input_60;
assign io_0 = input_61;
assign io_0 = input_62;
assign io_0 = input_63;
assign io_0 = input_64;
assign io_0 = input_65;
assign io_0 = input_66;
assign io_0 = input_67;
assign io_0 = input_68;
assign io_0 = input_69;
assign io_0 = input_70;
assign io_0 = input_71;
assign io_0 = input_72;
assign io_0 = input_73;
assign io_0 = input_74;
assign io_0 = input_75;
assign io_0 = input_76;
assign io_0 = input_77;
assign io_0 = input_78;
assign io_0 = input_79;
assign io_0 = input_80;
assign io_0 = input_81;
assign io_0 = input_82;
assign io_0 = input_83;
assign io_0 = input_84;
assign io_0 = input_85;
assign io_0 = input_86;
assign io_0 = input_87;
assign io_0 = input_88;
assign io_0 = input_89;
assign io_0 = input_90;
assign io_0 = input_91;
assign io_0 = input_92;
assign io_0 = input_93;
assign io_0 = input_94;
assign io_0 = input_95;
assign io_1 = input_1;
assign io_1 = input_2;
assign io_1 = input_3;
assign io_1 = input_4;
assign io_1 = input_5;
assign io_1 = input_6;
assign io_1 = input_7;
assign io_1 = input_8;
assign io_1 = input_9;
assign io_1 = input_10;
assign io_1 = input_11;
assign io_1 = input_12;
assign io_1 = input_13;
assign io_1 = input_14;
assign io_1 = input_15;
assign io_1 = input_16;
assign io_1 = input_17;
assign io_1 = input_18;
assign io_1 = input_19;
assign io_1 = input_20;
assign io_1 = input_21;
assign io_1 = input_22;
assign io_1 = input_23;
assign io_1 = input_24;
assign io_1 = input_25;
assign io_1 = input_26;
assign io_1 = input_27;
assign io_1 = input_28;
assign io_1 = input_29;
assign io_1 = input_30;
assign io_1 = input_31;
assign io_1 = input_32;
assign io_1 = input_33;
assign io_1 = input_34;
assign io_1 = input_35;
assign io_1 = input_36;
assign io_1 = input_37;
assign io_1 = input_38;
assign io_1 = input_39;
assign io_1 = input_40;
assign io_1 = input_41;
assign io_1 = input_42;
assign io_1 = input_43;
assign io_1 = input_44;
assign io_1 = input_45;
assign io_1 = input_46;
assign io_1 = input_47;
assign io_1 = input_48;
assign io_1 = input_49;
assign io_1 = input_50;
assign io_1 = input_51;
assign io_1 = input_52;
assign io_1 = input_53;
assign io_1 = input_54;
assign io_1 = input_55;
assign io_1 = input_56;
assign io_1 = input_57;
assign io_1 = input_58;
assign io_1 = input_59;
assign io_1 = input_60;
assign io_1 = input_61;
assign io_1 = input_62;
assign io_1 = input_63;
assign io_1 = input_64;
assign io_1 = input_65;
assign io_1 = input_66;
assign io_1 = input_67;
assign io_1 = input_68;
assign io_1 = input_69;
assign io_1 = input_70;
assign io_1 = input_71;
assign io_1 = input_72;
assign io_1 = input_73;
assign io_1 = input_74;
assign io_1 = input_75;
assign io_1 = input_76;
assign io_1 = input_77;
assign io_1 = input_78;
assign io_1 = input_79;
assign io_1 = input_80;
assign io_1 = input_81;
assign io_1 = input_82;
assign io_1 = input_83;
assign io_1 = input_84;
assign io_1 = input_85;
assign io_1 = input_86;
assign io_1 = input_87;
assign io_1 = input_88;
assign io_1 = input_89;
assign io_1 = input_90;
assign io_1 = input_91;
assign io_1 = input_92;
assign io_1 = input_93;
assign io_1 = input_94;
assign io_1 = input_95;
assign io_2 = input_2;
assign io_2 = input_3;
assign io_2 = input_4;
assign io_2 = input_5;
assign io_2 = input_6;
assign io_2 = input_7;
assign io_2 = input_8;
assign io_2 = input_9;
assign io_2 = input_10;
assign io_2 = input_11;
assign io_2 = input_12;
assign io_2 = input_13;
assign io_2 = input_14;
assign io_2 = input_15;
assign io_2 = input_16;
assign io_2 = input_17;
assign io_2 = input_18;
assign io_2 = input_19;
assign io_2 = input_20;
assign io_2 = input_21;
assign io_2 = input_22;
assign io_2 = input_23;
assign io_2 = input_24;
assign io_2 = input_25;
assign io_2 = input_26;
assign io_2 = input_27;
assign io_2 = input_28;
assign io_2 = input_29;
assign io_2 = input_30;
assign io_2 = input_31;
assign io_2 = input_32;
assign io_2 = input_33;
assign io_2 = input_34;
assign io_2 = input_35;
assign io_2 = input_36;
assign io_2 = input_37;
assign io_2 = input_38;
assign io_2 = input_39;
assign io_2 = input_40;
assign io_2 = input_41;
assign io_2 = input_42;
assign io_2 = input_43;
assign io_2 = input_44;
assign io_2 = input_45;
assign io_2 = input_46;
assign io_2 = input_47;
assign io_2 = input_48;
assign io_2 = input_49;
assign io_2 = input_50;
assign io_2 = input_51;
assign io_2 = input_52;
assign io_2 = input_53;
assign io_2 = input_54;
assign io_2 = input_55;
assign io_2 = input_56;
assign io_2 = input_57;
assign io_2 = input_58;
assign io_2 = input_59;
assign io_2 = input_60;
assign io_2 = input_61;
assign io_2 = input_62;
assign io_2 = input_63;
assign io_2 = input_64;
assign io_2 = input_65;
assign io_2 = input_66;
assign io_2 = input_67;
assign io_2 = input_68;
assign io_2 = input_69;
assign io_2 = input_70;
assign io_2 = input_71;
assign io_2 = input_72;
assign io_2 = input_73;
assign io_2 = input_74;
assign io_2 = input_75;
assign io_2 = input_76;
assign io_2 = input_77;
assign io_2 = input_78;
assign io_2 = input_79;
assign io_2 = input_80;
assign io_2 = input_81;
assign io_2 = input_82;
assign io_2 = input_83;
assign io_2 = input_84;
assign io_2 = input_85;
assign io_2 = input_86;
assign io_2 = input_87;
assign io_2 = input_88;
assign io_2 = input_89;
assign io_2 = input_90;
assign io_2 = input_91;
assign io_2 = input_92;
assign io_2 = input_93;
assign io_2 = input_94;
assign io_2 = input_95;
assign io_3 = input_3;
assign io_3 = input_4;
assign io_3 = input_5;
assign io_3 = input_6;
assign io_3 = input_7;
assign io_3 = input_8;
assign io_3 = input_9;
assign io_3 = input_10;
assign io_3 = input_11;
assign io_3 = input_12;
assign io_3 = input_13;
assign io_3 = input_14;
assign io_3 = input_15;
assign io_3 = input_16;
assign io_3 = input_17;
assign io_3 = input_18;
assign io_3 = input_19;
assign io_3 = input_20;
assign io_3 = input_21;
assign io_3 = input_22;
assign io_3 = input_23;
assign io_3 = input_24;
assign io_3 = input_25;
assign io_3 = input_26;
assign io_3 = input_27;
assign io_3 = input_28;
assign io_3 = input_29;
assign io_3 = input_30;
assign io_3 = input_31;
assign io_3 = input_32;
assign io_3 = input_33;
assign io_3 = input_34;
assign io_3 = input_35;
assign io_3 = input_36;
assign io_3 = input_37;
assign io_3 = input_38;
assign io_3 = input_39;
assign io_3 = input_40;
assign io_3 = input_41;
assign io_3 = input_42;
assign io_3 = input_43;
assign io_3 = input_44;
assign io_3 = input_45;
assign io_3 = input_46;
assign io_3 = input_47;
assign io_3 = input_48;
assign io_3 = input_49;
assign io_3 = input_50;
assign io_3 = input_51;
assign io_3 = input_52;
assign io_3 = input_53;
assign io_3 = input_54;
assign io_3 = input_55;
assign io_3 = input_56;
assign io_3 = input_57;
assign io_3 = input_58;
assign io_3 = input_59;
assign io_3 = input_60;
assign io_3 = input_61;
assign io_3 = input_62;
assign io_3 = input_63;
assign io_3 = input_64;
assign io_3 = input_65;
assign io_3 = input_66;
assign io_3 = input_67;
assign io_3 = input_68;
assign io_3 = input_69;
assign io_3 = input_70;
assign io_3 = input_71;
assign io_3 = input_72;
assign io_3 = input_73;
assign io_3 = input_74;
assign io_3 = input_75;
assign io_3 = input_76;
assign io_3 = input_77;
assign io_3 = input_78;
assign io_3 = input_79;
assign io_3 = input_80;
assign io_3 = input_81;
assign io_3 = input_82;
assign io_3 = input_83;
assign io_3 = input_84;
assign io_3 = input_85;
assign io_3 = input_86;
assign io_3 = input_87;
assign io_3 = input_88;
assign io_3 = input_89;
assign io_3 = input_90;
assign io_3 = input_91;
assign io_3 = input_92;
assign io_3 = input_93;
assign io_3 = input_94;
assign io_3 = input_95;
assign io_4 = input_4;
assign io_4 = input_5;
assign io_4 = input_6;
assign io_4 = input_7;
assign io_4 = input_8;
assign io_4 = input_9;
assign io_4 = input_10;
assign io_4 = input_11;
assign io_4 = input_12;
assign io_4 = input_13;
assign io_4 = input_14;
assign io_4 = input_15;
assign io_4 = input_16;
assign io_4 = input_17;
assign io_4 = input_18;
assign io_4 = input_19;
assign io_4 = input_20;
assign io_4 = input_21;
assign io_4 = input_22;
assign io_4 = input_23;
assign io_4 = input_24;
assign io_4 = input_25;
assign io_4 = input_26;
assign io_4 = input_27;
assign io_4 = input_28;
assign io_4 = input_29;
assign io_4 = input_30;
assign io_4 = input_31;
assign io_4 = input_32;
assign io_4 = input_33;
assign io_4 = input_34;
assign io_4 = input_35;
assign io_4 = input_36;
assign io_4 = input_37;
assign io_4 = input_38;
assign io_4 = input_39;
assign io_4 = input_40;
assign io_4 = input_41;
assign io_4 = input_42;
assign io_4 = input_43;
assign io_4 = input_44;
assign io_4 = input_45;
assign io_4 = input_46;
assign io_4 = input_47;
assign io_4 = input_48;
assign io_4 = input_49;
assign io_4 = input_50;
assign io_4 = input_51;
assign io_4 = input_52;
assign io_4 = input_53;
assign io_4 = input_54;
assign io_4 = input_55;
assign io_4 = input_56;
assign io_4 = input_57;
assign io_4 = input_58;
assign io_4 = input_59;
assign io_4 = input_60;
assign io_4 = input_61;
assign io_4 = input_62;
assign io_4 = input_63;
assign io_4 = input_64;
assign io_4 = input_65;
assign io_4 = input_66;
assign io_4 = input_67;
assign io_4 = input_68;
assign io_4 = input_69;
assign io_4 = input_70;
assign io_4 = input_71;
assign io_4 = input_72;
assign io_4 = input_73;
assign io_4 = input_74;
assign io_4 = input_75;
assign io_4 = input_76;
assign io_4 = input_77;
assign io_4 = input_78;
assign io_4 = input_79;
assign io_4 = input_80;
assign io_4 = input_81;
assign io_4 = input_82;
assign io_4 = input_83;
assign io_4 = input_84;
assign io_4 = input_85;
assign io_4 = input_86;
assign io_4 = input_87;
assign io_4 = input_88;
assign io_4 = input_89;
assign io_4 = input_90;
assign io_4 = input_91;
assign io_4 = input_92;
assign io_4 = input_93;
assign io_4 = input_94;
assign io_4 = input_95;
assign io_5 = input_5;
assign io_5 = input_6;
assign io_5 = input_7;
assign io_5 = input_8;
assign io_5 = input_9;
assign io_5 = input_10;
assign io_5 = input_11;
assign io_5 = input_12;
assign io_5 = input_13;
assign io_5 = input_14;
assign io_5 = input_15;
assign io_5 = input_16;
assign io_5 = input_17;
assign io_5 = input_18;
assign io_5 = input_19;
assign io_5 = input_20;
assign io_5 = input_21;
assign io_5 = input_22;
assign io_5 = input_23;
assign io_5 = input_24;
assign io_5 = input_25;
assign io_5 = input_26;
assign io_5 = input_27;
assign io_5 = input_28;
assign io_5 = input_29;
assign io_5 = input_30;
assign io_5 = input_31;
assign io_5 = input_32;
assign io_5 = input_33;
assign io_5 = input_34;
assign io_5 = input_35;
assign io_5 = input_36;
assign io_5 = input_37;
assign io_5 = input_38;
assign io_5 = input_39;
assign io_5 = input_40;
assign io_5 = input_41;
assign io_5 = input_42;
assign io_5 = input_43;
assign io_5 = input_44;
assign io_5 = input_45;
assign io_5 = input_46;
assign io_5 = input_47;
assign io_5 = input_48;
assign io_5 = input_49;
assign io_5 = input_50;
assign io_5 = input_51;
assign io_5 = input_52;
assign io_5 = input_53;
assign io_5 = input_54;
assign io_5 = input_55;
assign io_5 = input_56;
assign io_5 = input_57;
assign io_5 = input_58;
assign io_5 = input_59;
assign io_5 = input_60;
assign io_5 = input_61;
assign io_5 = input_62;
assign io_5 = input_63;
assign io_5 = input_64;
assign io_5 = input_65;
assign io_5 = input_66;
assign io_5 = input_67;
assign io_5 = input_68;
assign io_5 = input_69;
assign io_5 = input_70;
assign io_5 = input_71;
assign io_5 = input_72;
assign io_5 = input_73;
assign io_5 = input_74;
assign io_5 = input_75;
assign io_5 = input_76;
assign io_5 = input_77;
assign io_5 = input_78;
assign io_5 = input_79;
assign io_5 = input_80;
assign io_5 = input_81;
assign io_5 = input_82;
assign io_5 = input_83;
assign io_5 = input_84;
assign io_5 = input_85;
assign io_5 = input_86;
assign io_5 = input_87;
assign io_5 = input_88;
assign io_5 = input_89;
assign io_5 = input_90;
assign io_5 = input_91;
assign io_5 = input_92;
assign io_5 = input_93;
assign io_5 = input_94;
assign io_5 = input_95;
assign io_6 = input_6;
assign io_6 = input_7;
assign io_6 = input_8;
assign io_6 = input_9;
assign io_6 = input_10;
assign io_6 = input_11;
assign io_6 = input_12;
assign io_6 = input_13;
assign io_6 = input_14;
assign io_6 = input_15;
assign io_6 = input_16;
assign io_6 = input_17;
assign io_6 = input_18;
assign io_6 = input_19;
assign io_6 = input_20;
assign io_6 = input_21;
assign io_6 = input_22;
assign io_6 = input_23;
assign io_6 = input_24;
assign io_6 = input_25;
assign io_6 = input_26;
assign io_6 = input_27;
assign io_6 = input_28;
assign io_6 = input_29;
assign io_6 = input_30;
assign io_6 = input_31;
assign io_6 = input_32;
assign io_6 = input_33;
assign io_6 = input_34;
assign io_6 = input_35;
assign io_6 = input_36;
assign io_6 = input_37;
assign io_6 = input_38;
assign io_6 = input_39;
assign io_6 = input_40;
assign io_6 = input_41;
assign io_6 = input_42;
assign io_6 = input_43;
assign io_6 = input_44;
assign io_6 = input_45;
assign io_6 = input_46;
assign io_6 = input_47;
assign io_6 = input_48;
assign io_6 = input_49;
assign io_6 = input_50;
assign io_6 = input_51;
assign io_6 = input_52;
assign io_6 = input_53;
assign io_6 = input_54;
assign io_6 = input_55;
assign io_6 = input_56;
assign io_6 = input_57;
assign io_6 = input_58;
assign io_6 = input_59;
assign io_6 = input_60;
assign io_6 = input_61;
assign io_6 = input_62;
assign io_6 = input_63;
assign io_6 = input_64;
assign io_6 = input_65;
assign io_6 = input_66;
assign io_6 = input_67;
assign io_6 = input_68;
assign io_6 = input_69;
assign io_6 = input_70;
assign io_6 = input_71;
assign io_6 = input_72;
assign io_6 = input_73;
assign io_6 = input_74;
assign io_6 = input_75;
assign io_6 = input_76;
assign io_6 = input_77;
assign io_6 = input_78;
assign io_6 = input_79;
assign io_6 = input_80;
assign io_6 = input_81;
assign io_6 = input_82;
assign io_6 = input_83;
assign io_6 = input_84;
assign io_6 = input_85;
assign io_6 = input_86;
assign io_6 = input_87;
assign io_6 = input_88;
assign io_6 = input_89;
assign io_6 = input_90;
assign io_6 = input_91;
assign io_6 = input_92;
assign io_6 = input_93;
assign io_6 = input_94;
assign io_6 = input_95;
assign io_7 = input_7;
assign io_7 = input_8;
assign io_7 = input_9;
assign io_7 = input_10;
assign io_7 = input_11;
assign io_7 = input_12;
assign io_7 = input_13;
assign io_7 = input_14;
assign io_7 = input_15;
assign io_7 = input_16;
assign io_7 = input_17;
assign io_7 = input_18;
assign io_7 = input_19;
assign io_7 = input_20;
assign io_7 = input_21;
assign io_7 = input_22;
assign io_7 = input_23;
assign io_7 = input_24;
assign io_7 = input_25;
assign io_7 = input_26;
assign io_7 = input_27;
assign io_7 = input_28;
assign io_7 = input_29;
assign io_7 = input_30;
assign io_7 = input_31;
assign io_7 = input_32;
assign io_7 = input_33;
assign io_7 = input_34;
assign io_7 = input_35;
assign io_7 = input_36;
assign io_7 = input_37;
assign io_7 = input_38;
assign io_7 = input_39;
assign io_7 = input_40;
assign io_7 = input_41;
assign io_7 = input_42;
assign io_7 = input_43;
assign io_7 = input_44;
assign io_7 = input_45;
assign io_7 = input_46;
assign io_7 = input_47;
assign io_7 = input_48;
assign io_7 = input_49;
assign io_7 = input_50;
assign io_7 = input_51;
assign io_7 = input_52;
assign io_7 = input_53;
assign io_7 = input_54;
assign io_7 = input_55;
assign io_7 = input_56;
assign io_7 = input_57;
assign io_7 = input_58;
assign io_7 = input_59;
assign io_7 = input_60;
assign io_7 = input_61;
assign io_7 = input_62;
assign io_7 = input_63;
assign io_7 = input_64;
assign io_7 = input_65;
assign io_7 = input_66;
assign io_7 = input_67;
assign io_7 = input_68;
assign io_7 = input_69;
assign io_7 = input_70;
assign io_7 = input_71;
assign io_7 = input_72;
assign io_7 = input_73;
assign io_7 = input_74;
assign io_7 = input_75;
assign io_7 = input_76;
assign io_7 = input_77;
assign io_7 = input_78;
assign io_7 = input_79;
assign io_7 = input_80;
assign io_7 = input_81;
assign io_7 = input_82;
assign io_7 = input_83;
assign io_7 = input_84;
assign io_7 = input_85;
assign io_7 = input_86;
assign io_7 = input_87;
assign io_7 = input_88;
assign io_7 = input_89;
assign io_7 = input_90;
assign io_7 = input_91;
assign io_7 = input_92;
assign io_7 = input_93;
assign io_7 = input_94;
assign io_7 = input_95;
assign io_8 = input_8;
assign io_8 = input_9;
assign io_8 = input_10;
assign io_8 = input_11;
assign io_8 = input_12;
assign io_8 = input_13;
assign io_8 = input_14;
assign io_8 = input_15;
assign io_8 = input_16;
assign io_8 = input_17;
assign io_8 = input_18;
assign io_8 = input_19;
assign io_8 = input_20;
assign io_8 = input_21;
assign io_8 = input_22;
assign io_8 = input_23;
assign io_8 = input_24;
assign io_8 = input_25;
assign io_8 = input_26;
assign io_8 = input_27;
assign io_8 = input_28;
assign io_8 = input_29;
assign io_8 = input_30;
assign io_8 = input_31;
assign io_8 = input_32;
assign io_8 = input_33;
assign io_8 = input_34;
assign io_8 = input_35;
assign io_8 = input_36;
assign io_8 = input_37;
assign io_8 = input_38;
assign io_8 = input_39;
assign io_8 = input_40;
assign io_8 = input_41;
assign io_8 = input_42;
assign io_8 = input_43;
assign io_8 = input_44;
assign io_8 = input_45;
assign io_8 = input_46;
assign io_8 = input_47;
assign io_8 = input_48;
assign io_8 = input_49;
assign io_8 = input_50;
assign io_8 = input_51;
assign io_8 = input_52;
assign io_8 = input_53;
assign io_8 = input_54;
assign io_8 = input_55;
assign io_8 = input_56;
assign io_8 = input_57;
assign io_8 = input_58;
assign io_8 = input_59;
assign io_8 = input_60;
assign io_8 = input_61;
assign io_8 = input_62;
assign io_8 = input_63;
assign io_8 = input_64;
assign io_8 = input_65;
assign io_8 = input_66;
assign io_8 = input_67;
assign io_8 = input_68;
assign io_8 = input_69;
assign io_8 = input_70;
assign io_8 = input_71;
assign io_8 = input_72;
assign io_8 = input_73;
assign io_8 = input_74;
assign io_8 = input_75;
assign io_8 = input_76;
assign io_8 = input_77;
assign io_8 = input_78;
assign io_8 = input_79;
assign io_8 = input_80;
assign io_8 = input_81;
assign io_8 = input_82;
assign io_8 = input_83;
assign io_8 = input_84;
assign io_8 = input_85;
assign io_8 = input_86;
assign io_8 = input_87;
assign io_8 = input_88;
assign io_8 = input_89;
assign io_8 = input_90;
assign io_8 = input_91;
assign io_8 = input_92;
assign io_8 = input_93;
assign io_8 = input_94;
assign io_8 = input_95;
assign io_9 = input_9;
assign io_9 = input_10;
assign io_9 = input_11;
assign io_9 = input_12;
assign io_9 = input_13;
assign io_9 = input_14;
assign io_9 = input_15;
assign io_9 = input_16;
assign io_9 = input_17;
assign io_9 = input_18;
assign io_9 = input_19;
assign io_9 = input_20;
assign io_9 = input_21;
assign io_9 = input_22;
assign io_9 = input_23;
assign io_9 = input_24;
assign io_9 = input_25;
assign io_9 = input_26;
assign io_9 = input_27;
assign io_9 = input_28;
assign io_9 = input_29;
assign io_9 = input_30;
assign io_9 = input_31;
assign io_9 = input_32;
assign io_9 = input_33;
assign io_9 = input_34;
assign io_9 = input_35;
assign io_9 = input_36;
assign io_9 = input_37;
assign io_9 = input_38;
assign io_9 = input_39;
assign io_9 = input_40;
assign io_9 = input_41;
assign io_9 = input_42;
assign io_9 = input_43;
assign io_9 = input_44;
assign io_9 = input_45;
assign io_9 = input_46;
assign io_9 = input_47;
assign io_9 = input_48;
assign io_9 = input_49;
assign io_9 = input_50;
assign io_9 = input_51;
assign io_9 = input_52;
assign io_9 = input_53;
assign io_9 = input_54;
assign io_9 = input_55;
assign io_9 = input_56;
assign io_9 = input_57;
assign io_9 = input_58;
assign io_9 = input_59;
assign io_9 = input_60;
assign io_9 = input_61;
assign io_9 = input_62;
assign io_9 = input_63;
assign io_9 = input_64;
assign io_9 = input_65;
assign io_9 = input_66;
assign io_9 = input_67;
assign io_9 = input_68;
assign io_9 = input_69;
assign io_9 = input_70;
assign io_9 = input_71;
assign io_9 = input_72;
assign io_9 = input_73;
assign io_9 = input_74;
assign io_9 = input_75;
assign io_9 = input_76;
assign io_9 = input_77;
assign io_9 = input_78;
assign io_9 = input_79;
assign io_9 = input_80;
assign io_9 = input_81;
assign io_9 = input_82;
assign io_9 = input_83;
assign io_9 = input_84;
assign io_9 = input_85;
assign io_9 = input_86;
assign io_9 = input_87;
assign io_9 = input_88;
assign io_9 = input_89;
assign io_9 = input_90;
assign io_9 = input_91;
assign io_9 = input_92;
assign io_9 = input_93;
assign io_9 = input_94;
assign io_9 = input_95;
assign io_10 = input_10;
assign io_10 = input_11;
assign io_10 = input_12;
assign io_10 = input_13;
assign io_10 = input_14;
assign io_10 = input_15;
assign io_10 = input_16;
assign io_10 = input_17;
assign io_10 = input_18;
assign io_10 = input_19;
assign io_10 = input_20;
assign io_10 = input_21;
assign io_10 = input_22;
assign io_10 = input_23;
assign io_10 = input_24;
assign io_10 = input_25;
assign io_10 = input_26;
assign io_10 = input_27;
assign io_10 = input_28;
assign io_10 = input_29;
assign io_10 = input_30;
assign io_10 = input_31;
assign io_10 = input_32;
assign io_10 = input_33;
assign io_10 = input_34;
assign io_10 = input_35;
assign io_10 = input_36;
assign io_10 = input_37;
assign io_10 = input_38;
assign io_10 = input_39;
assign io_10 = input_40;
assign io_10 = input_41;
assign io_10 = input_42;
assign io_10 = input_43;
assign io_10 = input_44;
assign io_10 = input_45;
assign io_10 = input_46;
assign io_10 = input_47;
assign io_10 = input_48;
assign io_10 = input_49;
assign io_10 = input_50;
assign io_10 = input_51;
assign io_10 = input_52;
assign io_10 = input_53;
assign io_10 = input_54;
assign io_10 = input_55;
assign io_10 = input_56;
assign io_10 = input_57;
assign io_10 = input_58;
assign io_10 = input_59;
assign io_10 = input_60;
assign io_10 = input_61;
assign io_10 = input_62;
assign io_10 = input_63;
assign io_10 = input_64;
assign io_10 = input_65;
assign io_10 = input_66;
assign io_10 = input_67;
assign io_10 = input_68;
assign io_10 = input_69;
assign io_10 = input_70;
assign io_10 = input_71;
assign io_10 = input_72;
assign io_10 = input_73;
assign io_10 = input_74;
assign io_10 = input_75;
assign io_10 = input_76;
assign io_10 = input_77;
assign io_10 = input_78;
assign io_10 = input_79;
assign io_10 = input_80;
assign io_10 = input_81;
assign io_10 = input_82;
assign io_10 = input_83;
assign io_10 = input_84;
assign io_10 = input_85;
assign io_10 = input_86;
assign io_10 = input_87;
assign io_10 = input_88;
assign io_10 = input_89;
assign io_10 = input_90;
assign io_10 = input_91;
assign io_10 = input_92;
assign io_10 = input_93;
assign io_10 = input_94;
assign io_10 = input_95;
assign io_11 = input_11;
assign io_11 = input_12;
assign io_11 = input_13;
assign io_11 = input_14;
assign io_11 = input_15;
assign io_11 = input_16;
assign io_11 = input_17;
assign io_11 = input_18;
assign io_11 = input_19;
assign io_11 = input_20;
assign io_11 = input_21;
assign io_11 = input_22;
assign io_11 = input_23;
assign io_11 = input_24;
assign io_11 = input_25;
assign io_11 = input_26;
assign io_11 = input_27;
assign io_11 = input_28;
assign io_11 = input_29;
assign io_11 = input_30;
assign io_11 = input_31;
assign io_11 = input_32;
assign io_11 = input_33;
assign io_11 = input_34;
assign io_11 = input_35;
assign io_11 = input_36;
assign io_11 = input_37;
assign io_11 = input_38;
assign io_11 = input_39;
assign io_11 = input_40;
assign io_11 = input_41;
assign io_11 = input_42;
assign io_11 = input_43;
assign io_11 = input_44;
assign io_11 = input_45;
assign io_11 = input_46;
assign io_11 = input_47;
assign io_11 = input_48;
assign io_11 = input_49;
assign io_11 = input_50;
assign io_11 = input_51;
assign io_11 = input_52;
assign io_11 = input_53;
assign io_11 = input_54;
assign io_11 = input_55;
assign io_11 = input_56;
assign io_11 = input_57;
assign io_11 = input_58;
assign io_11 = input_59;
assign io_11 = input_60;
assign io_11 = input_61;
assign io_11 = input_62;
assign io_11 = input_63;
assign io_11 = input_64;
assign io_11 = input_65;
assign io_11 = input_66;
assign io_11 = input_67;
assign io_11 = input_68;
assign io_11 = input_69;
assign io_11 = input_70;
assign io_11 = input_71;
assign io_11 = input_72;
assign io_11 = input_73;
assign io_11 = input_74;
assign io_11 = input_75;
assign io_11 = input_76;
assign io_11 = input_77;
assign io_11 = input_78;
assign io_11 = input_79;
assign io_11 = input_80;
assign io_11 = input_81;
assign io_11 = input_82;
assign io_11 = input_83;
assign io_11 = input_84;
assign io_11 = input_85;
assign io_11 = input_86;
assign io_11 = input_87;
assign io_11 = input_88;
assign io_11 = input_89;
assign io_11 = input_90;
assign io_11 = input_91;
assign io_11 = input_92;
assign io_11 = input_93;
assign io_11 = input_94;
assign io_11 = input_95;
assign io_12 = input_12;
assign io_12 = input_13;
assign io_12 = input_14;
assign io_12 = input_15;
assign io_12 = input_16;
assign io_12 = input_17;
assign io_12 = input_18;
assign io_12 = input_19;
assign io_12 = input_20;
assign io_12 = input_21;
assign io_12 = input_22;
assign io_12 = input_23;
assign io_12 = input_24;
assign io_12 = input_25;
assign io_12 = input_26;
assign io_12 = input_27;
assign io_12 = input_28;
assign io_12 = input_29;
assign io_12 = input_30;
assign io_12 = input_31;
assign io_12 = input_32;
assign io_12 = input_33;
assign io_12 = input_34;
assign io_12 = input_35;
assign io_12 = input_36;
assign io_12 = input_37;
assign io_12 = input_38;
assign io_12 = input_39;
assign io_12 = input_40;
assign io_12 = input_41;
assign io_12 = input_42;
assign io_12 = input_43;
assign io_12 = input_44;
assign io_12 = input_45;
assign io_12 = input_46;
assign io_12 = input_47;
assign io_12 = input_48;
assign io_12 = input_49;
assign io_12 = input_50;
assign io_12 = input_51;
assign io_12 = input_52;
assign io_12 = input_53;
assign io_12 = input_54;
assign io_12 = input_55;
assign io_12 = input_56;
assign io_12 = input_57;
assign io_12 = input_58;
assign io_12 = input_59;
assign io_12 = input_60;
assign io_12 = input_61;
assign io_12 = input_62;
assign io_12 = input_63;
assign io_12 = input_64;
assign io_12 = input_65;
assign io_12 = input_66;
assign io_12 = input_67;
assign io_12 = input_68;
assign io_12 = input_69;
assign io_12 = input_70;
assign io_12 = input_71;
assign io_12 = input_72;
assign io_12 = input_73;
assign io_12 = input_74;
assign io_12 = input_75;
assign io_12 = input_76;
assign io_12 = input_77;
assign io_12 = input_78;
assign io_12 = input_79;
assign io_12 = input_80;
assign io_12 = input_81;
assign io_12 = input_82;
assign io_12 = input_83;
assign io_12 = input_84;
assign io_12 = input_85;
assign io_12 = input_86;
assign io_12 = input_87;
assign io_12 = input_88;
assign io_12 = input_89;
assign io_12 = input_90;
assign io_12 = input_91;
assign io_12 = input_92;
assign io_12 = input_93;
assign io_12 = input_94;
assign io_12 = input_95;
assign io_13 = input_13;
assign io_13 = input_14;
assign io_13 = input_15;
assign io_13 = input_16;
assign io_13 = input_17;
assign io_13 = input_18;
assign io_13 = input_19;
assign io_13 = input_20;
assign io_13 = input_21;
assign io_13 = input_22;
assign io_13 = input_23;
assign io_13 = input_24;
assign io_13 = input_25;
assign io_13 = input_26;
assign io_13 = input_27;
assign io_13 = input_28;
assign io_13 = input_29;
assign io_13 = input_30;
assign io_13 = input_31;
assign io_13 = input_32;
assign io_13 = input_33;
assign io_13 = input_34;
assign io_13 = input_35;
assign io_13 = input_36;
assign io_13 = input_37;
assign io_13 = input_38;
assign io_13 = input_39;
assign io_13 = input_40;
assign io_13 = input_41;
assign io_13 = input_42;
assign io_13 = input_43;
assign io_13 = input_44;
assign io_13 = input_45;
assign io_13 = input_46;
assign io_13 = input_47;
assign io_13 = input_48;
assign io_13 = input_49;
assign io_13 = input_50;
assign io_13 = input_51;
assign io_13 = input_52;
assign io_13 = input_53;
assign io_13 = input_54;
assign io_13 = input_55;
assign io_13 = input_56;
assign io_13 = input_57;
assign io_13 = input_58;
assign io_13 = input_59;
assign io_13 = input_60;
assign io_13 = input_61;
assign io_13 = input_62;
assign io_13 = input_63;
assign io_13 = input_64;
assign io_13 = input_65;
assign io_13 = input_66;
assign io_13 = input_67;
assign io_13 = input_68;
assign io_13 = input_69;
assign io_13 = input_70;
assign io_13 = input_71;
assign io_13 = input_72;
assign io_13 = input_73;
assign io_13 = input_74;
assign io_13 = input_75;
assign io_13 = input_76;
assign io_13 = input_77;
assign io_13 = input_78;
assign io_13 = input_79;
assign io_13 = input_80;
assign io_13 = input_81;
assign io_13 = input_82;
assign io_13 = input_83;
assign io_13 = input_84;
assign io_13 = input_85;
assign io_13 = input_86;
assign io_13 = input_87;
assign io_13 = input_88;
assign io_13 = input_89;
assign io_13 = input_90;
assign io_13 = input_91;
assign io_13 = input_92;
assign io_13 = input_93;
assign io_13 = input_94;
assign io_13 = input_95;
assign io_14 = input_14;
assign io_14 = input_15;
assign io_14 = input_16;
assign io_14 = input_17;
assign io_14 = input_18;
assign io_14 = input_19;
assign io_14 = input_20;
assign io_14 = input_21;
assign io_14 = input_22;
assign io_14 = input_23;
assign io_14 = input_24;
assign io_14 = input_25;
assign io_14 = input_26;
assign io_14 = input_27;
assign io_14 = input_28;
assign io_14 = input_29;
assign io_14 = input_30;
assign io_14 = input_31;
assign io_14 = input_32;
assign io_14 = input_33;
assign io_14 = input_34;
assign io_14 = input_35;
assign io_14 = input_36;
assign io_14 = input_37;
assign io_14 = input_38;
assign io_14 = input_39;
assign io_14 = input_40;
assign io_14 = input_41;
assign io_14 = input_42;
assign io_14 = input_43;
assign io_14 = input_44;
assign io_14 = input_45;
assign io_14 = input_46;
assign io_14 = input_47;
assign io_14 = input_48;
assign io_14 = input_49;
assign io_14 = input_50;
assign io_14 = input_51;
assign io_14 = input_52;
assign io_14 = input_53;
assign io_14 = input_54;
assign io_14 = input_55;
assign io_14 = input_56;
assign io_14 = input_57;
assign io_14 = input_58;
assign io_14 = input_59;
assign io_14 = input_60;
assign io_14 = input_61;
assign io_14 = input_62;
assign io_14 = input_63;
assign io_14 = input_64;
assign io_14 = input_65;
assign io_14 = input_66;
assign io_14 = input_67;
assign io_14 = input_68;
assign io_14 = input_69;
assign io_14 = input_70;
assign io_14 = input_71;
assign io_14 = input_72;
assign io_14 = input_73;
assign io_14 = input_74;
assign io_14 = input_75;
assign io_14 = input_76;
assign io_14 = input_77;
assign io_14 = input_78;
assign io_14 = input_79;
assign io_14 = input_80;
assign io_14 = input_81;
assign io_14 = input_82;
assign io_14 = input_83;
assign io_14 = input_84;
assign io_14 = input_85;
assign io_14 = input_86;
assign io_14 = input_87;
assign io_14 = input_88;
assign io_14 = input_89;
assign io_14 = input_90;
assign io_14 = input_91;
assign io_14 = input_92;
assign io_14 = input_93;
assign io_14 = input_94;
assign io_14 = input_95;
assign io_15 = input_15;
assign io_15 = input_16;
assign io_15 = input_17;
assign io_15 = input_18;
assign io_15 = input_19;
assign io_15 = input_20;
assign io_15 = input_21;
assign io_15 = input_22;
assign io_15 = input_23;
assign io_15 = input_24;
assign io_15 = input_25;
assign io_15 = input_26;
assign io_15 = input_27;
assign io_15 = input_28;
assign io_15 = input_29;
assign io_15 = input_30;
assign io_15 = input_31;
assign io_15 = input_32;
assign io_15 = input_33;
assign io_15 = input_34;
assign io_15 = input_35;
assign io_15 = input_36;
assign io_15 = input_37;
assign io_15 = input_38;
assign io_15 = input_39;
assign io_15 = input_40;
assign io_15 = input_41;
assign io_15 = input_42;
assign io_15 = input_43;
assign io_15 = input_44;
assign io_15 = input_45;
assign io_15 = input_46;
assign io_15 = input_47;
assign io_15 = input_48;
assign io_15 = input_49;
assign io_15 = input_50;
assign io_15 = input_51;
assign io_15 = input_52;
assign io_15 = input_53;
assign io_15 = input_54;
assign io_15 = input_55;
assign io_15 = input_56;
assign io_15 = input_57;
assign io_15 = input_58;
assign io_15 = input_59;
assign io_15 = input_60;
assign io_15 = input_61;
assign io_15 = input_62;
assign io_15 = input_63;
assign io_15 = input_64;
assign io_15 = input_65;
assign io_15 = input_66;
assign io_15 = input_67;
assign io_15 = input_68;
assign io_15 = input_69;
assign io_15 = input_70;
assign io_15 = input_71;
assign io_15 = input_72;
assign io_15 = input_73;
assign io_15 = input_74;
assign io_15 = input_75;
assign io_15 = input_76;
assign io_15 = input_77;
assign io_15 = input_78;
assign io_15 = input_79;
assign io_15 = input_80;
assign io_15 = input_81;
assign io_15 = input_82;
assign io_15 = input_83;
assign io_15 = input_84;
assign io_15 = input_85;
assign io_15 = input_86;
assign io_15 = input_87;
assign io_15 = input_88;
assign io_15 = input_89;
assign io_15 = input_90;
assign io_15 = input_91;
assign io_15 = input_92;
assign io_15 = input_93;
assign io_15 = input_94;
assign io_15 = input_95;
assign io_16 = input_16;
assign io_16 = input_17;
assign io_16 = input_18;
assign io_16 = input_19;
assign io_16 = input_20;
assign io_16 = input_21;
assign io_16 = input_22;
assign io_16 = input_23;
assign io_16 = input_24;
assign io_16 = input_25;
assign io_16 = input_26;
assign io_16 = input_27;
assign io_16 = input_28;
assign io_16 = input_29;
assign io_16 = input_30;
assign io_16 = input_31;
assign io_16 = input_32;
assign io_16 = input_33;
assign io_16 = input_34;
assign io_16 = input_35;
assign io_16 = input_36;
assign io_16 = input_37;
assign io_16 = input_38;
assign io_16 = input_39;
assign io_16 = input_40;
assign io_16 = input_41;
assign io_16 = input_42;
assign io_16 = input_43;
assign io_16 = input_44;
assign io_16 = input_45;
assign io_16 = input_46;
assign io_16 = input_47;
assign io_16 = input_48;
assign io_16 = input_49;
assign io_16 = input_50;
assign io_16 = input_51;
assign io_16 = input_52;
assign io_16 = input_53;
assign io_16 = input_54;
assign io_16 = input_55;
assign io_16 = input_56;
assign io_16 = input_57;
assign io_16 = input_58;
assign io_16 = input_59;
assign io_16 = input_60;
assign io_16 = input_61;
assign io_16 = input_62;
assign io_16 = input_63;
assign io_16 = input_64;
assign io_16 = input_65;
assign io_16 = input_66;
assign io_16 = input_67;
assign io_16 = input_68;
assign io_16 = input_69;
assign io_16 = input_70;
assign io_16 = input_71;
assign io_16 = input_72;
assign io_16 = input_73;
assign io_16 = input_74;
assign io_16 = input_75;
assign io_16 = input_76;
assign io_16 = input_77;
assign io_16 = input_78;
assign io_16 = input_79;
assign io_16 = input_80;
assign io_16 = input_81;
assign io_16 = input_82;
assign io_16 = input_83;
assign io_16 = input_84;
assign io_16 = input_85;
assign io_16 = input_86;
assign io_16 = input_87;
assign io_16 = input_88;
assign io_16 = input_89;
assign io_16 = input_90;
assign io_16 = input_91;
assign io_16 = input_92;
assign io_16 = input_93;
assign io_16 = input_94;
assign io_16 = input_95;
assign io_17 = input_17;
assign io_17 = input_18;
assign io_17 = input_19;
assign io_17 = input_20;
assign io_17 = input_21;
assign io_17 = input_22;
assign io_17 = input_23;
assign io_17 = input_24;
assign io_17 = input_25;
assign io_17 = input_26;
assign io_17 = input_27;
assign io_17 = input_28;
assign io_17 = input_29;
assign io_17 = input_30;
assign io_17 = input_31;
assign io_17 = input_32;
assign io_17 = input_33;
assign io_17 = input_34;
assign io_17 = input_35;
assign io_17 = input_36;
assign io_17 = input_37;
assign io_17 = input_38;
assign io_17 = input_39;
assign io_17 = input_40;
assign io_17 = input_41;
assign io_17 = input_42;
assign io_17 = input_43;
assign io_17 = input_44;
assign io_17 = input_45;
assign io_17 = input_46;
assign io_17 = input_47;
assign io_17 = input_48;
assign io_17 = input_49;
assign io_17 = input_50;
assign io_17 = input_51;
assign io_17 = input_52;
assign io_17 = input_53;
assign io_17 = input_54;
assign io_17 = input_55;
assign io_17 = input_56;
assign io_17 = input_57;
assign io_17 = input_58;
assign io_17 = input_59;
assign io_17 = input_60;
assign io_17 = input_61;
assign io_17 = input_62;
assign io_17 = input_63;
assign io_17 = input_64;
assign io_17 = input_65;
assign io_17 = input_66;
assign io_17 = input_67;
assign io_17 = input_68;
assign io_17 = input_69;
assign io_17 = input_70;
assign io_17 = input_71;
assign io_17 = input_72;
assign io_17 = input_73;
assign io_17 = input_74;
assign io_17 = input_75;
assign io_17 = input_76;
assign io_17 = input_77;
assign io_17 = input_78;
assign io_17 = input_79;
assign io_17 = input_80;
assign io_17 = input_81;
assign io_17 = input_82;
assign io_17 = input_83;
assign io_17 = input_84;
assign io_17 = input_85;
assign io_17 = input_86;
assign io_17 = input_87;
assign io_17 = input_88;
assign io_17 = input_89;
assign io_17 = input_90;
assign io_17 = input_91;
assign io_17 = input_92;
assign io_17 = input_93;
assign io_17 = input_94;
assign io_17 = input_95;
assign io_18 = input_18;
assign io_18 = input_19;
assign io_18 = input_20;
assign io_18 = input_21;
assign io_18 = input_22;
assign io_18 = input_23;
assign io_18 = input_24;
assign io_18 = input_25;
assign io_18 = input_26;
assign io_18 = input_27;
assign io_18 = input_28;
assign io_18 = input_29;
assign io_18 = input_30;
assign io_18 = input_31;
assign io_18 = input_32;
assign io_18 = input_33;
assign io_18 = input_34;
assign io_18 = input_35;
assign io_18 = input_36;
assign io_18 = input_37;
assign io_18 = input_38;
assign io_18 = input_39;
assign io_18 = input_40;
assign io_18 = input_41;
assign io_18 = input_42;
assign io_18 = input_43;
assign io_18 = input_44;
assign io_18 = input_45;
assign io_18 = input_46;
assign io_18 = input_47;
assign io_18 = input_48;
assign io_18 = input_49;
assign io_18 = input_50;
assign io_18 = input_51;
assign io_18 = input_52;
assign io_18 = input_53;
assign io_18 = input_54;
assign io_18 = input_55;
assign io_18 = input_56;
assign io_18 = input_57;
assign io_18 = input_58;
assign io_18 = input_59;
assign io_18 = input_60;
assign io_18 = input_61;
assign io_18 = input_62;
assign io_18 = input_63;
assign io_18 = input_64;
assign io_18 = input_65;
assign io_18 = input_66;
assign io_18 = input_67;
assign io_18 = input_68;
assign io_18 = input_69;
assign io_18 = input_70;
assign io_18 = input_71;
assign io_18 = input_72;
assign io_18 = input_73;
assign io_18 = input_74;
assign io_18 = input_75;
assign io_18 = input_76;
assign io_18 = input_77;
assign io_18 = input_78;
assign io_18 = input_79;
assign io_18 = input_80;
assign io_18 = input_81;
assign io_18 = input_82;
assign io_18 = input_83;
assign io_18 = input_84;
assign io_18 = input_85;
assign io_18 = input_86;
assign io_18 = input_87;
assign io_18 = input_88;
assign io_18 = input_89;
assign io_18 = input_90;
assign io_18 = input_91;
assign io_18 = input_92;
assign io_18 = input_93;
assign io_18 = input_94;
assign io_18 = input_95;
assign io_19 = input_19;
assign io_19 = input_20;
assign io_19 = input_21;
assign io_19 = input_22;
assign io_19 = input_23;
assign io_19 = input_24;
assign io_19 = input_25;
assign io_19 = input_26;
assign io_19 = input_27;
assign io_19 = input_28;
assign io_19 = input_29;
assign io_19 = input_30;
assign io_19 = input_31;
assign io_19 = input_32;
assign io_19 = input_33;
assign io_19 = input_34;
assign io_19 = input_35;
assign io_19 = input_36;
assign io_19 = input_37;
assign io_19 = input_38;
assign io_19 = input_39;
assign io_19 = input_40;
assign io_19 = input_41;
assign io_19 = input_42;
assign io_19 = input_43;
assign io_19 = input_44;
assign io_19 = input_45;
assign io_19 = input_46;
assign io_19 = input_47;
assign io_19 = input_48;
assign io_19 = input_49;
assign io_19 = input_50;
assign io_19 = input_51;
assign io_19 = input_52;
assign io_19 = input_53;
assign io_19 = input_54;
assign io_19 = input_55;
assign io_19 = input_56;
assign io_19 = input_57;
assign io_19 = input_58;
assign io_19 = input_59;
assign io_19 = input_60;
assign io_19 = input_61;
assign io_19 = input_62;
assign io_19 = input_63;
assign io_19 = input_64;
assign io_19 = input_65;
assign io_19 = input_66;
assign io_19 = input_67;
assign io_19 = input_68;
assign io_19 = input_69;
assign io_19 = input_70;
assign io_19 = input_71;
assign io_19 = input_72;
assign io_19 = input_73;
assign io_19 = input_74;
assign io_19 = input_75;
assign io_19 = input_76;
assign io_19 = input_77;
assign io_19 = input_78;
assign io_19 = input_79;
assign io_19 = input_80;
assign io_19 = input_81;
assign io_19 = input_82;
assign io_19 = input_83;
assign io_19 = input_84;
assign io_19 = input_85;
assign io_19 = input_86;
assign io_19 = input_87;
assign io_19 = input_88;
assign io_19 = input_89;
assign io_19 = input_90;
assign io_19 = input_91;
assign io_19 = input_92;
assign io_19 = input_93;
assign io_19 = input_94;
assign io_19 = input_95;
assign io_20 = input_20;
assign io_20 = input_21;
assign io_20 = input_22;
assign io_20 = input_23;
assign io_20 = input_24;
assign io_20 = input_25;
assign io_20 = input_26;
assign io_20 = input_27;
assign io_20 = input_28;
assign io_20 = input_29;
assign io_20 = input_30;
assign io_20 = input_31;
assign io_20 = input_32;
assign io_20 = input_33;
assign io_20 = input_34;
assign io_20 = input_35;
assign io_20 = input_36;
assign io_20 = input_37;
assign io_20 = input_38;
assign io_20 = input_39;
assign io_20 = input_40;
assign io_20 = input_41;
assign io_20 = input_42;
assign io_20 = input_43;
assign io_20 = input_44;
assign io_20 = input_45;
assign io_20 = input_46;
assign io_20 = input_47;
assign io_20 = input_48;
assign io_20 = input_49;
assign io_20 = input_50;
assign io_20 = input_51;
assign io_20 = input_52;
assign io_20 = input_53;
assign io_20 = input_54;
assign io_20 = input_55;
assign io_20 = input_56;
assign io_20 = input_57;
assign io_20 = input_58;
assign io_20 = input_59;
assign io_20 = input_60;
assign io_20 = input_61;
assign io_20 = input_62;
assign io_20 = input_63;
assign io_20 = input_64;
assign io_20 = input_65;
assign io_20 = input_66;
assign io_20 = input_67;
assign io_20 = input_68;
assign io_20 = input_69;
assign io_20 = input_70;
assign io_20 = input_71;
assign io_20 = input_72;
assign io_20 = input_73;
assign io_20 = input_74;
assign io_20 = input_75;
assign io_20 = input_76;
assign io_20 = input_77;
assign io_20 = input_78;
assign io_20 = input_79;
assign io_20 = input_80;
assign io_20 = input_81;
assign io_20 = input_82;
assign io_20 = input_83;
assign io_20 = input_84;
assign io_20 = input_85;
assign io_20 = input_86;
assign io_20 = input_87;
assign io_20 = input_88;
assign io_20 = input_89;
assign io_20 = input_90;
assign io_20 = input_91;
assign io_20 = input_92;
assign io_20 = input_93;
assign io_20 = input_94;
assign io_20 = input_95;
assign io_21 = input_21;
assign io_21 = input_22;
assign io_21 = input_23;
assign io_21 = input_24;
assign io_21 = input_25;
assign io_21 = input_26;
assign io_21 = input_27;
assign io_21 = input_28;
assign io_21 = input_29;
assign io_21 = input_30;
assign io_21 = input_31;
assign io_21 = input_32;
assign io_21 = input_33;
assign io_21 = input_34;
assign io_21 = input_35;
assign io_21 = input_36;
assign io_21 = input_37;
assign io_21 = input_38;
assign io_21 = input_39;
assign io_21 = input_40;
assign io_21 = input_41;
assign io_21 = input_42;
assign io_21 = input_43;
assign io_21 = input_44;
assign io_21 = input_45;
assign io_21 = input_46;
assign io_21 = input_47;
assign io_21 = input_48;
assign io_21 = input_49;
assign io_21 = input_50;
assign io_21 = input_51;
assign io_21 = input_52;
assign io_21 = input_53;
assign io_21 = input_54;
assign io_21 = input_55;
assign io_21 = input_56;
assign io_21 = input_57;
assign io_21 = input_58;
assign io_21 = input_59;
assign io_21 = input_60;
assign io_21 = input_61;
assign io_21 = input_62;
assign io_21 = input_63;
assign io_21 = input_64;
assign io_21 = input_65;
assign io_21 = input_66;
assign io_21 = input_67;
assign io_21 = input_68;
assign io_21 = input_69;
assign io_21 = input_70;
assign io_21 = input_71;
assign io_21 = input_72;
assign io_21 = input_73;
assign io_21 = input_74;
assign io_21 = input_75;
assign io_21 = input_76;
assign io_21 = input_77;
assign io_21 = input_78;
assign io_21 = input_79;
assign io_21 = input_80;
assign io_21 = input_81;
assign io_21 = input_82;
assign io_21 = input_83;
assign io_21 = input_84;
assign io_21 = input_85;
assign io_21 = input_86;
assign io_21 = input_87;
assign io_21 = input_88;
assign io_21 = input_89;
assign io_21 = input_90;
assign io_21 = input_91;
assign io_21 = input_92;
assign io_21 = input_93;
assign io_21 = input_94;
assign io_21 = input_95;
assign io_22 = input_22;
assign io_22 = input_23;
assign io_22 = input_24;
assign io_22 = input_25;
assign io_22 = input_26;
assign io_22 = input_27;
assign io_22 = input_28;
assign io_22 = input_29;
assign io_22 = input_30;
assign io_22 = input_31;
assign io_22 = input_32;
assign io_22 = input_33;
assign io_22 = input_34;
assign io_22 = input_35;
assign io_22 = input_36;
assign io_22 = input_37;
assign io_22 = input_38;
assign io_22 = input_39;
assign io_22 = input_40;
assign io_22 = input_41;
assign io_22 = input_42;
assign io_22 = input_43;
assign io_22 = input_44;
assign io_22 = input_45;
assign io_22 = input_46;
assign io_22 = input_47;
assign io_22 = input_48;
assign io_22 = input_49;
assign io_22 = input_50;
assign io_22 = input_51;
assign io_22 = input_52;
assign io_22 = input_53;
assign io_22 = input_54;
assign io_22 = input_55;
assign io_22 = input_56;
assign io_22 = input_57;
assign io_22 = input_58;
assign io_22 = input_59;
assign io_22 = input_60;
assign io_22 = input_61;
assign io_22 = input_62;
assign io_22 = input_63;
assign io_22 = input_64;
assign io_22 = input_65;
assign io_22 = input_66;
assign io_22 = input_67;
assign io_22 = input_68;
assign io_22 = input_69;
assign io_22 = input_70;
assign io_22 = input_71;
assign io_22 = input_72;
assign io_22 = input_73;
assign io_22 = input_74;
assign io_22 = input_75;
assign io_22 = input_76;
assign io_22 = input_77;
assign io_22 = input_78;
assign io_22 = input_79;
assign io_22 = input_80;
assign io_22 = input_81;
assign io_22 = input_82;
assign io_22 = input_83;
assign io_22 = input_84;
assign io_22 = input_85;
assign io_22 = input_86;
assign io_22 = input_87;
assign io_22 = input_88;
assign io_22 = input_89;
assign io_22 = input_90;
assign io_22 = input_91;
assign io_22 = input_92;
assign io_22 = input_93;
assign io_22 = input_94;
assign io_22 = input_95;
assign io_23 = input_23;
assign io_23 = input_24;
assign io_23 = input_25;
assign io_23 = input_26;
assign io_23 = input_27;
assign io_23 = input_28;
assign io_23 = input_29;
assign io_23 = input_30;
assign io_23 = input_31;
assign io_23 = input_32;
assign io_23 = input_33;
assign io_23 = input_34;
assign io_23 = input_35;
assign io_23 = input_36;
assign io_23 = input_37;
assign io_23 = input_38;
assign io_23 = input_39;
assign io_23 = input_40;
assign io_23 = input_41;
assign io_23 = input_42;
assign io_23 = input_43;
assign io_23 = input_44;
assign io_23 = input_45;
assign io_23 = input_46;
assign io_23 = input_47;
assign io_23 = input_48;
assign io_23 = input_49;
assign io_23 = input_50;
assign io_23 = input_51;
assign io_23 = input_52;
assign io_23 = input_53;
assign io_23 = input_54;
assign io_23 = input_55;
assign io_23 = input_56;
assign io_23 = input_57;
assign io_23 = input_58;
assign io_23 = input_59;
assign io_23 = input_60;
assign io_23 = input_61;
assign io_23 = input_62;
assign io_23 = input_63;
assign io_23 = input_64;
assign io_23 = input_65;
assign io_23 = input_66;
assign io_23 = input_67;
assign io_23 = input_68;
assign io_23 = input_69;
assign io_23 = input_70;
assign io_23 = input_71;
assign io_23 = input_72;
assign io_23 = input_73;
assign io_23 = input_74;
assign io_23 = input_75;
assign io_23 = input_76;
assign io_23 = input_77;
assign io_23 = input_78;
assign io_23 = input_79;
assign io_23 = input_80;
assign io_23 = input_81;
assign io_23 = input_82;
assign io_23 = input_83;
assign io_23 = input_84;
assign io_23 = input_85;
assign io_23 = input_86;
assign io_23 = input_87;
assign io_23 = input_88;
assign io_23 = input_89;
assign io_23 = input_90;
assign io_23 = input_91;
assign io_23 = input_92;
assign io_23 = input_93;
assign io_23 = input_94;
assign io_23 = input_95;
assign io_24 = input_24;
assign io_24 = input_25;
assign io_24 = input_26;
assign io_24 = input_27;
assign io_24 = input_28;
assign io_24 = input_29;
assign io_24 = input_30;
assign io_24 = input_31;
assign io_24 = input_32;
assign io_24 = input_33;
assign io_24 = input_34;
assign io_24 = input_35;
assign io_24 = input_36;
assign io_24 = input_37;
assign io_24 = input_38;
assign io_24 = input_39;
assign io_24 = input_40;
assign io_24 = input_41;
assign io_24 = input_42;
assign io_24 = input_43;
assign io_24 = input_44;
assign io_24 = input_45;
assign io_24 = input_46;
assign io_24 = input_47;
assign io_24 = input_48;
assign io_24 = input_49;
assign io_24 = input_50;
assign io_24 = input_51;
assign io_24 = input_52;
assign io_24 = input_53;
assign io_24 = input_54;
assign io_24 = input_55;
assign io_24 = input_56;
assign io_24 = input_57;
assign io_24 = input_58;
assign io_24 = input_59;
assign io_24 = input_60;
assign io_24 = input_61;
assign io_24 = input_62;
assign io_24 = input_63;
assign io_24 = input_64;
assign io_24 = input_65;
assign io_24 = input_66;
assign io_24 = input_67;
assign io_24 = input_68;
assign io_24 = input_69;
assign io_24 = input_70;
assign io_24 = input_71;
assign io_24 = input_72;
assign io_24 = input_73;
assign io_24 = input_74;
assign io_24 = input_75;
assign io_24 = input_76;
assign io_24 = input_77;
assign io_24 = input_78;
assign io_24 = input_79;
assign io_24 = input_80;
assign io_24 = input_81;
assign io_24 = input_82;
assign io_24 = input_83;
assign io_24 = input_84;
assign io_24 = input_85;
assign io_24 = input_86;
assign io_24 = input_87;
assign io_24 = input_88;
assign io_24 = input_89;
assign io_24 = input_90;
assign io_24 = input_91;
assign io_24 = input_92;
assign io_24 = input_93;
assign io_24 = input_94;
assign io_24 = input_95;
assign io_25 = input_25;
assign io_25 = input_26;
assign io_25 = input_27;
assign io_25 = input_28;
assign io_25 = input_29;
assign io_25 = input_30;
assign io_25 = input_31;
assign io_25 = input_32;
assign io_25 = input_33;
assign io_25 = input_34;
assign io_25 = input_35;
assign io_25 = input_36;
assign io_25 = input_37;
assign io_25 = input_38;
assign io_25 = input_39;
assign io_25 = input_40;
assign io_25 = input_41;
assign io_25 = input_42;
assign io_25 = input_43;
assign io_25 = input_44;
assign io_25 = input_45;
assign io_25 = input_46;
assign io_25 = input_47;
assign io_25 = input_48;
assign io_25 = input_49;
assign io_25 = input_50;
assign io_25 = input_51;
assign io_25 = input_52;
assign io_25 = input_53;
assign io_25 = input_54;
assign io_25 = input_55;
assign io_25 = input_56;
assign io_25 = input_57;
assign io_25 = input_58;
assign io_25 = input_59;
assign io_25 = input_60;
assign io_25 = input_61;
assign io_25 = input_62;
assign io_25 = input_63;
assign io_25 = input_64;
assign io_25 = input_65;
assign io_25 = input_66;
assign io_25 = input_67;
assign io_25 = input_68;
assign io_25 = input_69;
assign io_25 = input_70;
assign io_25 = input_71;
assign io_25 = input_72;
assign io_25 = input_73;
assign io_25 = input_74;
assign io_25 = input_75;
assign io_25 = input_76;
assign io_25 = input_77;
assign io_25 = input_78;
assign io_25 = input_79;
assign io_25 = input_80;
assign io_25 = input_81;
assign io_25 = input_82;
assign io_25 = input_83;
assign io_25 = input_84;
assign io_25 = input_85;
assign io_25 = input_86;
assign io_25 = input_87;
assign io_25 = input_88;
assign io_25 = input_89;
assign io_25 = input_90;
assign io_25 = input_91;
assign io_25 = input_92;
assign io_25 = input_93;
assign io_25 = input_94;
assign io_25 = input_95;
assign io_26 = input_26;
assign io_26 = input_27;
assign io_26 = input_28;
assign io_26 = input_29;
assign io_26 = input_30;
assign io_26 = input_31;
assign io_26 = input_32;
assign io_26 = input_33;
assign io_26 = input_34;
assign io_26 = input_35;
assign io_26 = input_36;
assign io_26 = input_37;
assign io_26 = input_38;
assign io_26 = input_39;
assign io_26 = input_40;
assign io_26 = input_41;
assign io_26 = input_42;
assign io_26 = input_43;
assign io_26 = input_44;
assign io_26 = input_45;
assign io_26 = input_46;
assign io_26 = input_47;
assign io_26 = input_48;
assign io_26 = input_49;
assign io_26 = input_50;
assign io_26 = input_51;
assign io_26 = input_52;
assign io_26 = input_53;
assign io_26 = input_54;
assign io_26 = input_55;
assign io_26 = input_56;
assign io_26 = input_57;
assign io_26 = input_58;
assign io_26 = input_59;
assign io_26 = input_60;
assign io_26 = input_61;
assign io_26 = input_62;
assign io_26 = input_63;
assign io_26 = input_64;
assign io_26 = input_65;
assign io_26 = input_66;
assign io_26 = input_67;
assign io_26 = input_68;
assign io_26 = input_69;
assign io_26 = input_70;
assign io_26 = input_71;
assign io_26 = input_72;
assign io_26 = input_73;
assign io_26 = input_74;
assign io_26 = input_75;
assign io_26 = input_76;
assign io_26 = input_77;
assign io_26 = input_78;
assign io_26 = input_79;
assign io_26 = input_80;
assign io_26 = input_81;
assign io_26 = input_82;
assign io_26 = input_83;
assign io_26 = input_84;
assign io_26 = input_85;
assign io_26 = input_86;
assign io_26 = input_87;
assign io_26 = input_88;
assign io_26 = input_89;
assign io_26 = input_90;
assign io_26 = input_91;
assign io_26 = input_92;
assign io_26 = input_93;
assign io_26 = input_94;
assign io_26 = input_95;
assign io_27 = input_27;
assign io_27 = input_28;
assign io_27 = input_29;
assign io_27 = input_30;
assign io_27 = input_31;
assign io_27 = input_32;
assign io_27 = input_33;
assign io_27 = input_34;
assign io_27 = input_35;
assign io_27 = input_36;
assign io_27 = input_37;
assign io_27 = input_38;
assign io_27 = input_39;
assign io_27 = input_40;
assign io_27 = input_41;
assign io_27 = input_42;
assign io_27 = input_43;
assign io_27 = input_44;
assign io_27 = input_45;
assign io_27 = input_46;
assign io_27 = input_47;
assign io_27 = input_48;
assign io_27 = input_49;
assign io_27 = input_50;
assign io_27 = input_51;
assign io_27 = input_52;
assign io_27 = input_53;
assign io_27 = input_54;
assign io_27 = input_55;
assign io_27 = input_56;
assign io_27 = input_57;
assign io_27 = input_58;
assign io_27 = input_59;
assign io_27 = input_60;
assign io_27 = input_61;
assign io_27 = input_62;
assign io_27 = input_63;
assign io_27 = input_64;
assign io_27 = input_65;
assign io_27 = input_66;
assign io_27 = input_67;
assign io_27 = input_68;
assign io_27 = input_69;
assign io_27 = input_70;
assign io_27 = input_71;
assign io_27 = input_72;
assign io_27 = input_73;
assign io_27 = input_74;
assign io_27 = input_75;
assign io_27 = input_76;
assign io_27 = input_77;
assign io_27 = input_78;
assign io_27 = input_79;
assign io_27 = input_80;
assign io_27 = input_81;
assign io_27 = input_82;
assign io_27 = input_83;
assign io_27 = input_84;
assign io_27 = input_85;
assign io_27 = input_86;
assign io_27 = input_87;
assign io_27 = input_88;
assign io_27 = input_89;
assign io_27 = input_90;
assign io_27 = input_91;
assign io_27 = input_92;
assign io_27 = input_93;
assign io_27 = input_94;
assign io_27 = input_95;
assign io_28 = input_28;
assign io_28 = input_29;
assign io_28 = input_30;
assign io_28 = input_31;
assign io_28 = input_32;
assign io_28 = input_33;
assign io_28 = input_34;
assign io_28 = input_35;
assign io_28 = input_36;
assign io_28 = input_37;
assign io_28 = input_38;
assign io_28 = input_39;
assign io_28 = input_40;
assign io_28 = input_41;
assign io_28 = input_42;
assign io_28 = input_43;
assign io_28 = input_44;
assign io_28 = input_45;
assign io_28 = input_46;
assign io_28 = input_47;
assign io_28 = input_48;
assign io_28 = input_49;
assign io_28 = input_50;
assign io_28 = input_51;
assign io_28 = input_52;
assign io_28 = input_53;
assign io_28 = input_54;
assign io_28 = input_55;
assign io_28 = input_56;
assign io_28 = input_57;
assign io_28 = input_58;
assign io_28 = input_59;
assign io_28 = input_60;
assign io_28 = input_61;
assign io_28 = input_62;
assign io_28 = input_63;
assign io_28 = input_64;
assign io_28 = input_65;
assign io_28 = input_66;
assign io_28 = input_67;
assign io_28 = input_68;
assign io_28 = input_69;
assign io_28 = input_70;
assign io_28 = input_71;
assign io_28 = input_72;
assign io_28 = input_73;
assign io_28 = input_74;
assign io_28 = input_75;
assign io_28 = input_76;
assign io_28 = input_77;
assign io_28 = input_78;
assign io_28 = input_79;
assign io_28 = input_80;
assign io_28 = input_81;
assign io_28 = input_82;
assign io_28 = input_83;
assign io_28 = input_84;
assign io_28 = input_85;
assign io_28 = input_86;
assign io_28 = input_87;
assign io_28 = input_88;
assign io_28 = input_89;
assign io_28 = input_90;
assign io_28 = input_91;
assign io_28 = input_92;
assign io_28 = input_93;
assign io_28 = input_94;
assign io_28 = input_95;
assign io_29 = input_29;
assign io_29 = input_30;
assign io_29 = input_31;
assign io_29 = input_32;
assign io_29 = input_33;
assign io_29 = input_34;
assign io_29 = input_35;
assign io_29 = input_36;
assign io_29 = input_37;
assign io_29 = input_38;
assign io_29 = input_39;
assign io_29 = input_40;
assign io_29 = input_41;
assign io_29 = input_42;
assign io_29 = input_43;
assign io_29 = input_44;
assign io_29 = input_45;
assign io_29 = input_46;
assign io_29 = input_47;
assign io_29 = input_48;
assign io_29 = input_49;
assign io_29 = input_50;
assign io_29 = input_51;
assign io_29 = input_52;
assign io_29 = input_53;
assign io_29 = input_54;
assign io_29 = input_55;
assign io_29 = input_56;
assign io_29 = input_57;
assign io_29 = input_58;
assign io_29 = input_59;
assign io_29 = input_60;
assign io_29 = input_61;
assign io_29 = input_62;
assign io_29 = input_63;
assign io_29 = input_64;
assign io_29 = input_65;
assign io_29 = input_66;
assign io_29 = input_67;
assign io_29 = input_68;
assign io_29 = input_69;
assign io_29 = input_70;
assign io_29 = input_71;
assign io_29 = input_72;
assign io_29 = input_73;
assign io_29 = input_74;
assign io_29 = input_75;
assign io_29 = input_76;
assign io_29 = input_77;
assign io_29 = input_78;
assign io_29 = input_79;
assign io_29 = input_80;
assign io_29 = input_81;
assign io_29 = input_82;
assign io_29 = input_83;
assign io_29 = input_84;
assign io_29 = input_85;
assign io_29 = input_86;
assign io_29 = input_87;
assign io_29 = input_88;
assign io_29 = input_89;
assign io_29 = input_90;
assign io_29 = input_91;
assign io_29 = input_92;
assign io_29 = input_93;
assign io_29 = input_94;
assign io_29 = input_95;
assign io_30 = input_30;
assign io_30 = input_31;
assign io_30 = input_32;
assign io_30 = input_33;
assign io_30 = input_34;
assign io_30 = input_35;
assign io_30 = input_36;
assign io_30 = input_37;
assign io_30 = input_38;
assign io_30 = input_39;
assign io_30 = input_40;
assign io_30 = input_41;
assign io_30 = input_42;
assign io_30 = input_43;
assign io_30 = input_44;
assign io_30 = input_45;
assign io_30 = input_46;
assign io_30 = input_47;
assign io_30 = input_48;
assign io_30 = input_49;
assign io_30 = input_50;
assign io_30 = input_51;
assign io_30 = input_52;
assign io_30 = input_53;
assign io_30 = input_54;
assign io_30 = input_55;
assign io_30 = input_56;
assign io_30 = input_57;
assign io_30 = input_58;
assign io_30 = input_59;
assign io_30 = input_60;
assign io_30 = input_61;
assign io_30 = input_62;
assign io_30 = input_63;
assign io_30 = input_64;
assign io_30 = input_65;
assign io_30 = input_66;
assign io_30 = input_67;
assign io_30 = input_68;
assign io_30 = input_69;
assign io_30 = input_70;
assign io_30 = input_71;
assign io_30 = input_72;
assign io_30 = input_73;
assign io_30 = input_74;
assign io_30 = input_75;
assign io_30 = input_76;
assign io_30 = input_77;
assign io_30 = input_78;
assign io_30 = input_79;
assign io_30 = input_80;
assign io_30 = input_81;
assign io_30 = input_82;
assign io_30 = input_83;
assign io_30 = input_84;
assign io_30 = input_85;
assign io_30 = input_86;
assign io_30 = input_87;
assign io_30 = input_88;
assign io_30 = input_89;
assign io_30 = input_90;
assign io_30 = input_91;
assign io_30 = input_92;
assign io_30 = input_93;
assign io_30 = input_94;
assign io_30 = input_95;
assign io_31 = input_31;
assign io_31 = input_32;
assign io_31 = input_33;
assign io_31 = input_34;
assign io_31 = input_35;
assign io_31 = input_36;
assign io_31 = input_37;
assign io_31 = input_38;
assign io_31 = input_39;
assign io_31 = input_40;
assign io_31 = input_41;
assign io_31 = input_42;
assign io_31 = input_43;
assign io_31 = input_44;
assign io_31 = input_45;
assign io_31 = input_46;
assign io_31 = input_47;
assign io_31 = input_48;
assign io_31 = input_49;
assign io_31 = input_50;
assign io_31 = input_51;
assign io_31 = input_52;
assign io_31 = input_53;
assign io_31 = input_54;
assign io_31 = input_55;
assign io_31 = input_56;
assign io_31 = input_57;
assign io_31 = input_58;
assign io_31 = input_59;
assign io_31 = input_60;
assign io_31 = input_61;
assign io_31 = input_62;
assign io_31 = input_63;
assign io_31 = input_64;
assign io_31 = input_65;
assign io_31 = input_66;
assign io_31 = input_67;
assign io_31 = input_68;
assign io_31 = input_69;
assign io_31 = input_70;
assign io_31 = input_71;
assign io_31 = input_72;
assign io_31 = input_73;
assign io_31 = input_74;
assign io_31 = input_75;
assign io_31 = input_76;
assign io_31 = input_77;
assign io_31 = input_78;
assign io_31 = input_79;
assign io_31 = input_80;
assign io_31 = input_81;
assign io_31 = input_82;
assign io_31 = input_83;
assign io_31 = input_84;
assign io_31 = input_85;
assign io_31 = input_86;
assign io_31 = input_87;
assign io_31 = input_88;
assign io_31 = input_89;
assign io_31 = input_90;
assign io_31 = input_91;
assign io_31 = input_92;
assign io_31 = input_93;
assign io_31 = input_94;
assign io_31 = input_95;
assign io_32 = input_32;
assign io_32 = input_33;
assign io_32 = input_34;
assign io_32 = input_35;
assign io_32 = input_36;
assign io_32 = input_37;
assign io_32 = input_38;
assign io_32 = input_39;
assign io_32 = input_40;
assign io_32 = input_41;
assign io_32 = input_42;
assign io_32 = input_43;
assign io_32 = input_44;
assign io_32 = input_45;
assign io_32 = input_46;
assign io_32 = input_47;
assign io_32 = input_48;
assign io_32 = input_49;
assign io_32 = input_50;
assign io_32 = input_51;
assign io_32 = input_52;
assign io_32 = input_53;
assign io_32 = input_54;
assign io_32 = input_55;
assign io_32 = input_56;
assign io_32 = input_57;
assign io_32 = input_58;
assign io_32 = input_59;
assign io_32 = input_60;
assign io_32 = input_61;
assign io_32 = input_62;
assign io_32 = input_63;
assign io_32 = input_64;
assign io_32 = input_65;
assign io_32 = input_66;
assign io_32 = input_67;
assign io_32 = input_68;
assign io_32 = input_69;
assign io_32 = input_70;
assign io_32 = input_71;
assign io_32 = input_72;
assign io_32 = input_73;
assign io_32 = input_74;
assign io_32 = input_75;
assign io_32 = input_76;
assign io_32 = input_77;
assign io_32 = input_78;
assign io_32 = input_79;
assign io_32 = input_80;
assign io_32 = input_81;
assign io_32 = input_82;
assign io_32 = input_83;
assign io_32 = input_84;
assign io_32 = input_85;
assign io_32 = input_86;
assign io_32 = input_87;
assign io_32 = input_88;
assign io_32 = input_89;
assign io_32 = input_90;
assign io_32 = input_91;
assign io_32 = input_92;
assign io_32 = input_93;
assign io_32 = input_94;
assign io_32 = input_95;
assign io_33 = input_33;
assign io_33 = input_34;
assign io_33 = input_35;
assign io_33 = input_36;
assign io_33 = input_37;
assign io_33 = input_38;
assign io_33 = input_39;
assign io_33 = input_40;
assign io_33 = input_41;
assign io_33 = input_42;
assign io_33 = input_43;
assign io_33 = input_44;
assign io_33 = input_45;
assign io_33 = input_46;
assign io_33 = input_47;
assign io_33 = input_48;
assign io_33 = input_49;
assign io_33 = input_50;
assign io_33 = input_51;
assign io_33 = input_52;
assign io_33 = input_53;
assign io_33 = input_54;
assign io_33 = input_55;
assign io_33 = input_56;
assign io_33 = input_57;
assign io_33 = input_58;
assign io_33 = input_59;
assign io_33 = input_60;
assign io_33 = input_61;
assign io_33 = input_62;
assign io_33 = input_63;
assign io_33 = input_64;
assign io_33 = input_65;
assign io_33 = input_66;
assign io_33 = input_67;
assign io_33 = input_68;
assign io_33 = input_69;
assign io_33 = input_70;
assign io_33 = input_71;
assign io_33 = input_72;
assign io_33 = input_73;
assign io_33 = input_74;
assign io_33 = input_75;
assign io_33 = input_76;
assign io_33 = input_77;
assign io_33 = input_78;
assign io_33 = input_79;
assign io_33 = input_80;
assign io_33 = input_81;
assign io_33 = input_82;
assign io_33 = input_83;
assign io_33 = input_84;
assign io_33 = input_85;
assign io_33 = input_86;
assign io_33 = input_87;
assign io_33 = input_88;
assign io_33 = input_89;
assign io_33 = input_90;
assign io_33 = input_91;
assign io_33 = input_92;
assign io_33 = input_93;
assign io_33 = input_94;
assign io_33 = input_95;
assign io_34 = input_34;
assign io_34 = input_35;
assign io_34 = input_36;
assign io_34 = input_37;
assign io_34 = input_38;
assign io_34 = input_39;
assign io_34 = input_40;
assign io_34 = input_41;
assign io_34 = input_42;
assign io_34 = input_43;
assign io_34 = input_44;
assign io_34 = input_45;
assign io_34 = input_46;
assign io_34 = input_47;
assign io_34 = input_48;
assign io_34 = input_49;
assign io_34 = input_50;
assign io_34 = input_51;
assign io_34 = input_52;
assign io_34 = input_53;
assign io_34 = input_54;
assign io_34 = input_55;
assign io_34 = input_56;
assign io_34 = input_57;
assign io_34 = input_58;
assign io_34 = input_59;
assign io_34 = input_60;
assign io_34 = input_61;
assign io_34 = input_62;
assign io_34 = input_63;
assign io_34 = input_64;
assign io_34 = input_65;
assign io_34 = input_66;
assign io_34 = input_67;
assign io_34 = input_68;
assign io_34 = input_69;
assign io_34 = input_70;
assign io_34 = input_71;
assign io_34 = input_72;
assign io_34 = input_73;
assign io_34 = input_74;
assign io_34 = input_75;
assign io_34 = input_76;
assign io_34 = input_77;
assign io_34 = input_78;
assign io_34 = input_79;
assign io_34 = input_80;
assign io_34 = input_81;
assign io_34 = input_82;
assign io_34 = input_83;
assign io_34 = input_84;
assign io_34 = input_85;
assign io_34 = input_86;
assign io_34 = input_87;
assign io_34 = input_88;
assign io_34 = input_89;
assign io_34 = input_90;
assign io_34 = input_91;
assign io_34 = input_92;
assign io_34 = input_93;
assign io_34 = input_94;
assign io_34 = input_95;
assign io_35 = input_35;
assign io_35 = input_36;
assign io_35 = input_37;
assign io_35 = input_38;
assign io_35 = input_39;
assign io_35 = input_40;
assign io_35 = input_41;
assign io_35 = input_42;
assign io_35 = input_43;
assign io_35 = input_44;
assign io_35 = input_45;
assign io_35 = input_46;
assign io_35 = input_47;
assign io_35 = input_48;
assign io_35 = input_49;
assign io_35 = input_50;
assign io_35 = input_51;
assign io_35 = input_52;
assign io_35 = input_53;
assign io_35 = input_54;
assign io_35 = input_55;
assign io_35 = input_56;
assign io_35 = input_57;
assign io_35 = input_58;
assign io_35 = input_59;
assign io_35 = input_60;
assign io_35 = input_61;
assign io_35 = input_62;
assign io_35 = input_63;
assign io_35 = input_64;
assign io_35 = input_65;
assign io_35 = input_66;
assign io_35 = input_67;
assign io_35 = input_68;
assign io_35 = input_69;
assign io_35 = input_70;
assign io_35 = input_71;
assign io_35 = input_72;
assign io_35 = input_73;
assign io_35 = input_74;
assign io_35 = input_75;
assign io_35 = input_76;
assign io_35 = input_77;
assign io_35 = input_78;
assign io_35 = input_79;
assign io_35 = input_80;
assign io_35 = input_81;
assign io_35 = input_82;
assign io_35 = input_83;
assign io_35 = input_84;
assign io_35 = input_85;
assign io_35 = input_86;
assign io_35 = input_87;
assign io_35 = input_88;
assign io_35 = input_89;
assign io_35 = input_90;
assign io_35 = input_91;
assign io_35 = input_92;
assign io_35 = input_93;
assign io_35 = input_94;
assign io_35 = input_95;
assign io_36 = input_36;
assign io_36 = input_37;
assign io_36 = input_38;
assign io_36 = input_39;
assign io_36 = input_40;
assign io_36 = input_41;
assign io_36 = input_42;
assign io_36 = input_43;
assign io_36 = input_44;
assign io_36 = input_45;
assign io_36 = input_46;
assign io_36 = input_47;
assign io_36 = input_48;
assign io_36 = input_49;
assign io_36 = input_50;
assign io_36 = input_51;
assign io_36 = input_52;
assign io_36 = input_53;
assign io_36 = input_54;
assign io_36 = input_55;
assign io_36 = input_56;
assign io_36 = input_57;
assign io_36 = input_58;
assign io_36 = input_59;
assign io_36 = input_60;
assign io_36 = input_61;
assign io_36 = input_62;
assign io_36 = input_63;
assign io_36 = input_64;
assign io_36 = input_65;
assign io_36 = input_66;
assign io_36 = input_67;
assign io_36 = input_68;
assign io_36 = input_69;
assign io_36 = input_70;
assign io_36 = input_71;
assign io_36 = input_72;
assign io_36 = input_73;
assign io_36 = input_74;
assign io_36 = input_75;
assign io_36 = input_76;
assign io_36 = input_77;
assign io_36 = input_78;
assign io_36 = input_79;
assign io_36 = input_80;
assign io_36 = input_81;
assign io_36 = input_82;
assign io_36 = input_83;
assign io_36 = input_84;
assign io_36 = input_85;
assign io_36 = input_86;
assign io_36 = input_87;
assign io_36 = input_88;
assign io_36 = input_89;
assign io_36 = input_90;
assign io_36 = input_91;
assign io_36 = input_92;
assign io_36 = input_93;
assign io_36 = input_94;
assign io_36 = input_95;
assign io_37 = input_37;
assign io_37 = input_38;
assign io_37 = input_39;
assign io_37 = input_40;
assign io_37 = input_41;
assign io_37 = input_42;
assign io_37 = input_43;
assign io_37 = input_44;
assign io_37 = input_45;
assign io_37 = input_46;
assign io_37 = input_47;
assign io_37 = input_48;
assign io_37 = input_49;
assign io_37 = input_50;
assign io_37 = input_51;
assign io_37 = input_52;
assign io_37 = input_53;
assign io_37 = input_54;
assign io_37 = input_55;
assign io_37 = input_56;
assign io_37 = input_57;
assign io_37 = input_58;
assign io_37 = input_59;
assign io_37 = input_60;
assign io_37 = input_61;
assign io_37 = input_62;
assign io_37 = input_63;
assign io_37 = input_64;
assign io_37 = input_65;
assign io_37 = input_66;
assign io_37 = input_67;
assign io_37 = input_68;
assign io_37 = input_69;
assign io_37 = input_70;
assign io_37 = input_71;
assign io_37 = input_72;
assign io_37 = input_73;
assign io_37 = input_74;
assign io_37 = input_75;
assign io_37 = input_76;
assign io_37 = input_77;
assign io_37 = input_78;
assign io_37 = input_79;
assign io_37 = input_80;
assign io_37 = input_81;
assign io_37 = input_82;
assign io_37 = input_83;
assign io_37 = input_84;
assign io_37 = input_85;
assign io_37 = input_86;
assign io_37 = input_87;
assign io_37 = input_88;
assign io_37 = input_89;
assign io_37 = input_90;
assign io_37 = input_91;
assign io_37 = input_92;
assign io_37 = input_93;
assign io_37 = input_94;
assign io_37 = input_95;
assign io_38 = input_38;
assign io_38 = input_39;
assign io_38 = input_40;
assign io_38 = input_41;
assign io_38 = input_42;
assign io_38 = input_43;
assign io_38 = input_44;
assign io_38 = input_45;
assign io_38 = input_46;
assign io_38 = input_47;
assign io_38 = input_48;
assign io_38 = input_49;
assign io_38 = input_50;
assign io_38 = input_51;
assign io_38 = input_52;
assign io_38 = input_53;
assign io_38 = input_54;
assign io_38 = input_55;
assign io_38 = input_56;
assign io_38 = input_57;
assign io_38 = input_58;
assign io_38 = input_59;
assign io_38 = input_60;
assign io_38 = input_61;
assign io_38 = input_62;
assign io_38 = input_63;
assign io_38 = input_64;
assign io_38 = input_65;
assign io_38 = input_66;
assign io_38 = input_67;
assign io_38 = input_68;
assign io_38 = input_69;
assign io_38 = input_70;
assign io_38 = input_71;
assign io_38 = input_72;
assign io_38 = input_73;
assign io_38 = input_74;
assign io_38 = input_75;
assign io_38 = input_76;
assign io_38 = input_77;
assign io_38 = input_78;
assign io_38 = input_79;
assign io_38 = input_80;
assign io_38 = input_81;
assign io_38 = input_82;
assign io_38 = input_83;
assign io_38 = input_84;
assign io_38 = input_85;
assign io_38 = input_86;
assign io_38 = input_87;
assign io_38 = input_88;
assign io_38 = input_89;
assign io_38 = input_90;
assign io_38 = input_91;
assign io_38 = input_92;
assign io_38 = input_93;
assign io_38 = input_94;
assign io_38 = input_95;
assign io_39 = input_39;
assign io_39 = input_40;
assign io_39 = input_41;
assign io_39 = input_42;
assign io_39 = input_43;
assign io_39 = input_44;
assign io_39 = input_45;
assign io_39 = input_46;
assign io_39 = input_47;
assign io_39 = input_48;
assign io_39 = input_49;
assign io_39 = input_50;
assign io_39 = input_51;
assign io_39 = input_52;
assign io_39 = input_53;
assign io_39 = input_54;
assign io_39 = input_55;
assign io_39 = input_56;
assign io_39 = input_57;
assign io_39 = input_58;
assign io_39 = input_59;
assign io_39 = input_60;
assign io_39 = input_61;
assign io_39 = input_62;
assign io_39 = input_63;
assign io_39 = input_64;
assign io_39 = input_65;
assign io_39 = input_66;
assign io_39 = input_67;
assign io_39 = input_68;
assign io_39 = input_69;
assign io_39 = input_70;
assign io_39 = input_71;
assign io_39 = input_72;
assign io_39 = input_73;
assign io_39 = input_74;
assign io_39 = input_75;
assign io_39 = input_76;
assign io_39 = input_77;
assign io_39 = input_78;
assign io_39 = input_79;
assign io_39 = input_80;
assign io_39 = input_81;
assign io_39 = input_82;
assign io_39 = input_83;
assign io_39 = input_84;
assign io_39 = input_85;
assign io_39 = input_86;
assign io_39 = input_87;
assign io_39 = input_88;
assign io_39 = input_89;
assign io_39 = input_90;
assign io_39 = input_91;
assign io_39 = input_92;
assign io_39 = input_93;
assign io_39 = input_94;
assign io_39 = input_95;
assign io_40 = input_40;
assign io_40 = input_41;
assign io_40 = input_42;
assign io_40 = input_43;
assign io_40 = input_44;
assign io_40 = input_45;
assign io_40 = input_46;
assign io_40 = input_47;
assign io_40 = input_48;
assign io_40 = input_49;
assign io_40 = input_50;
assign io_40 = input_51;
assign io_40 = input_52;
assign io_40 = input_53;
assign io_40 = input_54;
assign io_40 = input_55;
assign io_40 = input_56;
assign io_40 = input_57;
assign io_40 = input_58;
assign io_40 = input_59;
assign io_40 = input_60;
assign io_40 = input_61;
assign io_40 = input_62;
assign io_40 = input_63;
assign io_40 = input_64;
assign io_40 = input_65;
assign io_40 = input_66;
assign io_40 = input_67;
assign io_40 = input_68;
assign io_40 = input_69;
assign io_40 = input_70;
assign io_40 = input_71;
assign io_40 = input_72;
assign io_40 = input_73;
assign io_40 = input_74;
assign io_40 = input_75;
assign io_40 = input_76;
assign io_40 = input_77;
assign io_40 = input_78;
assign io_40 = input_79;
assign io_40 = input_80;
assign io_40 = input_81;
assign io_40 = input_82;
assign io_40 = input_83;
assign io_40 = input_84;
assign io_40 = input_85;
assign io_40 = input_86;
assign io_40 = input_87;
assign io_40 = input_88;
assign io_40 = input_89;
assign io_40 = input_90;
assign io_40 = input_91;
assign io_40 = input_92;
assign io_40 = input_93;
assign io_40 = input_94;
assign io_40 = input_95;
assign io_41 = input_41;
assign io_41 = input_42;
assign io_41 = input_43;
assign io_41 = input_44;
assign io_41 = input_45;
assign io_41 = input_46;
assign io_41 = input_47;
assign io_41 = input_48;
assign io_41 = input_49;
assign io_41 = input_50;
assign io_41 = input_51;
assign io_41 = input_52;
assign io_41 = input_53;
assign io_41 = input_54;
assign io_41 = input_55;
assign io_41 = input_56;
assign io_41 = input_57;
assign io_41 = input_58;
assign io_41 = input_59;
assign io_41 = input_60;
assign io_41 = input_61;
assign io_41 = input_62;
assign io_41 = input_63;
assign io_41 = input_64;
assign io_41 = input_65;
assign io_41 = input_66;
assign io_41 = input_67;
assign io_41 = input_68;
assign io_41 = input_69;
assign io_41 = input_70;
assign io_41 = input_71;
assign io_41 = input_72;
assign io_41 = input_73;
assign io_41 = input_74;
assign io_41 = input_75;
assign io_41 = input_76;
assign io_41 = input_77;
assign io_41 = input_78;
assign io_41 = input_79;
assign io_41 = input_80;
assign io_41 = input_81;
assign io_41 = input_82;
assign io_41 = input_83;
assign io_41 = input_84;
assign io_41 = input_85;
assign io_41 = input_86;
assign io_41 = input_87;
assign io_41 = input_88;
assign io_41 = input_89;
assign io_41 = input_90;
assign io_41 = input_91;
assign io_41 = input_92;
assign io_41 = input_93;
assign io_41 = input_94;
assign io_41 = input_95;
assign io_42 = input_42;
assign io_42 = input_43;
assign io_42 = input_44;
assign io_42 = input_45;
assign io_42 = input_46;
assign io_42 = input_47;
assign io_42 = input_48;
assign io_42 = input_49;
assign io_42 = input_50;
assign io_42 = input_51;
assign io_42 = input_52;
assign io_42 = input_53;
assign io_42 = input_54;
assign io_42 = input_55;
assign io_42 = input_56;
assign io_42 = input_57;
assign io_42 = input_58;
assign io_42 = input_59;
assign io_42 = input_60;
assign io_42 = input_61;
assign io_42 = input_62;
assign io_42 = input_63;
assign io_42 = input_64;
assign io_42 = input_65;
assign io_42 = input_66;
assign io_42 = input_67;
assign io_42 = input_68;
assign io_42 = input_69;
assign io_42 = input_70;
assign io_42 = input_71;
assign io_42 = input_72;
assign io_42 = input_73;
assign io_42 = input_74;
assign io_42 = input_75;
assign io_42 = input_76;
assign io_42 = input_77;
assign io_42 = input_78;
assign io_42 = input_79;
assign io_42 = input_80;
assign io_42 = input_81;
assign io_42 = input_82;
assign io_42 = input_83;
assign io_42 = input_84;
assign io_42 = input_85;
assign io_42 = input_86;
assign io_42 = input_87;
assign io_42 = input_88;
assign io_42 = input_89;
assign io_42 = input_90;
assign io_42 = input_91;
assign io_42 = input_92;
assign io_42 = input_93;
assign io_42 = input_94;
assign io_42 = input_95;
assign io_43 = input_43;
assign io_43 = input_44;
assign io_43 = input_45;
assign io_43 = input_46;
assign io_43 = input_47;
assign io_43 = input_48;
assign io_43 = input_49;
assign io_43 = input_50;
assign io_43 = input_51;
assign io_43 = input_52;
assign io_43 = input_53;
assign io_43 = input_54;
assign io_43 = input_55;
assign io_43 = input_56;
assign io_43 = input_57;
assign io_43 = input_58;
assign io_43 = input_59;
assign io_43 = input_60;
assign io_43 = input_61;
assign io_43 = input_62;
assign io_43 = input_63;
assign io_43 = input_64;
assign io_43 = input_65;
assign io_43 = input_66;
assign io_43 = input_67;
assign io_43 = input_68;
assign io_43 = input_69;
assign io_43 = input_70;
assign io_43 = input_71;
assign io_43 = input_72;
assign io_43 = input_73;
assign io_43 = input_74;
assign io_43 = input_75;
assign io_43 = input_76;
assign io_43 = input_77;
assign io_43 = input_78;
assign io_43 = input_79;
assign io_43 = input_80;
assign io_43 = input_81;
assign io_43 = input_82;
assign io_43 = input_83;
assign io_43 = input_84;
assign io_43 = input_85;
assign io_43 = input_86;
assign io_43 = input_87;
assign io_43 = input_88;
assign io_43 = input_89;
assign io_43 = input_90;
assign io_43 = input_91;
assign io_43 = input_92;
assign io_43 = input_93;
assign io_43 = input_94;
assign io_43 = input_95;
assign io_44 = input_44;
assign io_44 = input_45;
assign io_44 = input_46;
assign io_44 = input_47;
assign io_44 = input_48;
assign io_44 = input_49;
assign io_44 = input_50;
assign io_44 = input_51;
assign io_44 = input_52;
assign io_44 = input_53;
assign io_44 = input_54;
assign io_44 = input_55;
assign io_44 = input_56;
assign io_44 = input_57;
assign io_44 = input_58;
assign io_44 = input_59;
assign io_44 = input_60;
assign io_44 = input_61;
assign io_44 = input_62;
assign io_44 = input_63;
assign io_44 = input_64;
assign io_44 = input_65;
assign io_44 = input_66;
assign io_44 = input_67;
assign io_44 = input_68;
assign io_44 = input_69;
assign io_44 = input_70;
assign io_44 = input_71;
assign io_44 = input_72;
assign io_44 = input_73;
assign io_44 = input_74;
assign io_44 = input_75;
assign io_44 = input_76;
assign io_44 = input_77;
assign io_44 = input_78;
assign io_44 = input_79;
assign io_44 = input_80;
assign io_44 = input_81;
assign io_44 = input_82;
assign io_44 = input_83;
assign io_44 = input_84;
assign io_44 = input_85;
assign io_44 = input_86;
assign io_44 = input_87;
assign io_44 = input_88;
assign io_44 = input_89;
assign io_44 = input_90;
assign io_44 = input_91;
assign io_44 = input_92;
assign io_44 = input_93;
assign io_44 = input_94;
assign io_44 = input_95;
assign io_45 = input_45;
assign io_45 = input_46;
assign io_45 = input_47;
assign io_45 = input_48;
assign io_45 = input_49;
assign io_45 = input_50;
assign io_45 = input_51;
assign io_45 = input_52;
assign io_45 = input_53;
assign io_45 = input_54;
assign io_45 = input_55;
assign io_45 = input_56;
assign io_45 = input_57;
assign io_45 = input_58;
assign io_45 = input_59;
assign io_45 = input_60;
assign io_45 = input_61;
assign io_45 = input_62;
assign io_45 = input_63;
assign io_45 = input_64;
assign io_45 = input_65;
assign io_45 = input_66;
assign io_45 = input_67;
assign io_45 = input_68;
assign io_45 = input_69;
assign io_45 = input_70;
assign io_45 = input_71;
assign io_45 = input_72;
assign io_45 = input_73;
assign io_45 = input_74;
assign io_45 = input_75;
assign io_45 = input_76;
assign io_45 = input_77;
assign io_45 = input_78;
assign io_45 = input_79;
assign io_45 = input_80;
assign io_45 = input_81;
assign io_45 = input_82;
assign io_45 = input_83;
assign io_45 = input_84;
assign io_45 = input_85;
assign io_45 = input_86;
assign io_45 = input_87;
assign io_45 = input_88;
assign io_45 = input_89;
assign io_45 = input_90;
assign io_45 = input_91;
assign io_45 = input_92;
assign io_45 = input_93;
assign io_45 = input_94;
assign io_45 = input_95;
assign io_46 = input_46;
assign io_46 = input_47;
assign io_46 = input_48;
assign io_46 = input_49;
assign io_46 = input_50;
assign io_46 = input_51;
assign io_46 = input_52;
assign io_46 = input_53;
assign io_46 = input_54;
assign io_46 = input_55;
assign io_46 = input_56;
assign io_46 = input_57;
assign io_46 = input_58;
assign io_46 = input_59;
assign io_46 = input_60;
assign io_46 = input_61;
assign io_46 = input_62;
assign io_46 = input_63;
assign io_46 = input_64;
assign io_46 = input_65;
assign io_46 = input_66;
assign io_46 = input_67;
assign io_46 = input_68;
assign io_46 = input_69;
assign io_46 = input_70;
assign io_46 = input_71;
assign io_46 = input_72;
assign io_46 = input_73;
assign io_46 = input_74;
assign io_46 = input_75;
assign io_46 = input_76;
assign io_46 = input_77;
assign io_46 = input_78;
assign io_46 = input_79;
assign io_46 = input_80;
assign io_46 = input_81;
assign io_46 = input_82;
assign io_46 = input_83;
assign io_46 = input_84;
assign io_46 = input_85;
assign io_46 = input_86;
assign io_46 = input_87;
assign io_46 = input_88;
assign io_46 = input_89;
assign io_46 = input_90;
assign io_46 = input_91;
assign io_46 = input_92;
assign io_46 = input_93;
assign io_46 = input_94;
assign io_46 = input_95;
assign io_47 = input_47;
assign io_47 = input_48;
assign io_47 = input_49;
assign io_47 = input_50;
assign io_47 = input_51;
assign io_47 = input_52;
assign io_47 = input_53;
assign io_47 = input_54;
assign io_47 = input_55;
assign io_47 = input_56;
assign io_47 = input_57;
assign io_47 = input_58;
assign io_47 = input_59;
assign io_47 = input_60;
assign io_47 = input_61;
assign io_47 = input_62;
assign io_47 = input_63;
assign io_47 = input_64;
assign io_47 = input_65;
assign io_47 = input_66;
assign io_47 = input_67;
assign io_47 = input_68;
assign io_47 = input_69;
assign io_47 = input_70;
assign io_47 = input_71;
assign io_47 = input_72;
assign io_47 = input_73;
assign io_47 = input_74;
assign io_47 = input_75;
assign io_47 = input_76;
assign io_47 = input_77;
assign io_47 = input_78;
assign io_47 = input_79;
assign io_47 = input_80;
assign io_47 = input_81;
assign io_47 = input_82;
assign io_47 = input_83;
assign io_47 = input_84;
assign io_47 = input_85;
assign io_47 = input_86;
assign io_47 = input_87;
assign io_47 = input_88;
assign io_47 = input_89;
assign io_47 = input_90;
assign io_47 = input_91;
assign io_47 = input_92;
assign io_47 = input_93;
assign io_47 = input_94;
assign io_47 = input_95;
assign io_48 = input_48;
assign io_48 = input_49;
assign io_48 = input_50;
assign io_48 = input_51;
assign io_48 = input_52;
assign io_48 = input_53;
assign io_48 = input_54;
assign io_48 = input_55;
assign io_48 = input_56;
assign io_48 = input_57;
assign io_48 = input_58;
assign io_48 = input_59;
assign io_48 = input_60;
assign io_48 = input_61;
assign io_48 = input_62;
assign io_48 = input_63;
assign io_48 = input_64;
assign io_48 = input_65;
assign io_48 = input_66;
assign io_48 = input_67;
assign io_48 = input_68;
assign io_48 = input_69;
assign io_48 = input_70;
assign io_48 = input_71;
assign io_48 = input_72;
assign io_48 = input_73;
assign io_48 = input_74;
assign io_48 = input_75;
assign io_48 = input_76;
assign io_48 = input_77;
assign io_48 = input_78;
assign io_48 = input_79;
assign io_48 = input_80;
assign io_48 = input_81;
assign io_48 = input_82;
assign io_48 = input_83;
assign io_48 = input_84;
assign io_48 = input_85;
assign io_48 = input_86;
assign io_48 = input_87;
assign io_48 = input_88;
assign io_48 = input_89;
assign io_48 = input_90;
assign io_48 = input_91;
assign io_48 = input_92;
assign io_48 = input_93;
assign io_48 = input_94;
assign io_48 = input_95;
assign io_49 = input_49;
assign io_49 = input_50;
assign io_49 = input_51;
assign io_49 = input_52;
assign io_49 = input_53;
assign io_49 = input_54;
assign io_49 = input_55;
assign io_49 = input_56;
assign io_49 = input_57;
assign io_49 = input_58;
assign io_49 = input_59;
assign io_49 = input_60;
assign io_49 = input_61;
assign io_49 = input_62;
assign io_49 = input_63;
assign io_49 = input_64;
assign io_49 = input_65;
assign io_49 = input_66;
assign io_49 = input_67;
assign io_49 = input_68;
assign io_49 = input_69;
assign io_49 = input_70;
assign io_49 = input_71;
assign io_49 = input_72;
assign io_49 = input_73;
assign io_49 = input_74;
assign io_49 = input_75;
assign io_49 = input_76;
assign io_49 = input_77;
assign io_49 = input_78;
assign io_49 = input_79;
assign io_49 = input_80;
assign io_49 = input_81;
assign io_49 = input_82;
assign io_49 = input_83;
assign io_49 = input_84;
assign io_49 = input_85;
assign io_49 = input_86;
assign io_49 = input_87;
assign io_49 = input_88;
assign io_49 = input_89;
assign io_49 = input_90;
assign io_49 = input_91;
assign io_49 = input_92;
assign io_49 = input_93;
assign io_49 = input_94;
assign io_49 = input_95;
assign io_50 = input_50;
assign io_50 = input_51;
assign io_50 = input_52;
assign io_50 = input_53;
assign io_50 = input_54;
assign io_50 = input_55;
assign io_50 = input_56;
assign io_50 = input_57;
assign io_50 = input_58;
assign io_50 = input_59;
assign io_50 = input_60;
assign io_50 = input_61;
assign io_50 = input_62;
assign io_50 = input_63;
assign io_50 = input_64;
assign io_50 = input_65;
assign io_50 = input_66;
assign io_50 = input_67;
assign io_50 = input_68;
assign io_50 = input_69;
assign io_50 = input_70;
assign io_50 = input_71;
assign io_50 = input_72;
assign io_50 = input_73;
assign io_50 = input_74;
assign io_50 = input_75;
assign io_50 = input_76;
assign io_50 = input_77;
assign io_50 = input_78;
assign io_50 = input_79;
assign io_50 = input_80;
assign io_50 = input_81;
assign io_50 = input_82;
assign io_50 = input_83;
assign io_50 = input_84;
assign io_50 = input_85;
assign io_50 = input_86;
assign io_50 = input_87;
assign io_50 = input_88;
assign io_50 = input_89;
assign io_50 = input_90;
assign io_50 = input_91;
assign io_50 = input_92;
assign io_50 = input_93;
assign io_50 = input_94;
assign io_50 = input_95;
assign io_51 = input_51;
assign io_51 = input_52;
assign io_51 = input_53;
assign io_51 = input_54;
assign io_51 = input_55;
assign io_51 = input_56;
assign io_51 = input_57;
assign io_51 = input_58;
assign io_51 = input_59;
assign io_51 = input_60;
assign io_51 = input_61;
assign io_51 = input_62;
assign io_51 = input_63;
assign io_51 = input_64;
assign io_51 = input_65;
assign io_51 = input_66;
assign io_51 = input_67;
assign io_51 = input_68;
assign io_51 = input_69;
assign io_51 = input_70;
assign io_51 = input_71;
assign io_51 = input_72;
assign io_51 = input_73;
assign io_51 = input_74;
assign io_51 = input_75;
assign io_51 = input_76;
assign io_51 = input_77;
assign io_51 = input_78;
assign io_51 = input_79;
assign io_51 = input_80;
assign io_51 = input_81;
assign io_51 = input_82;
assign io_51 = input_83;
assign io_51 = input_84;
assign io_51 = input_85;
assign io_51 = input_86;
assign io_51 = input_87;
assign io_51 = input_88;
assign io_51 = input_89;
assign io_51 = input_90;
assign io_51 = input_91;
assign io_51 = input_92;
assign io_51 = input_93;
assign io_51 = input_94;
assign io_51 = input_95;
assign io_52 = input_52;
assign io_52 = input_53;
assign io_52 = input_54;
assign io_52 = input_55;
assign io_52 = input_56;
assign io_52 = input_57;
assign io_52 = input_58;
assign io_52 = input_59;
assign io_52 = input_60;
assign io_52 = input_61;
assign io_52 = input_62;
assign io_52 = input_63;
assign io_52 = input_64;
assign io_52 = input_65;
assign io_52 = input_66;
assign io_52 = input_67;
assign io_52 = input_68;
assign io_52 = input_69;
assign io_52 = input_70;
assign io_52 = input_71;
assign io_52 = input_72;
assign io_52 = input_73;
assign io_52 = input_74;
assign io_52 = input_75;
assign io_52 = input_76;
assign io_52 = input_77;
assign io_52 = input_78;
assign io_52 = input_79;
assign io_52 = input_80;
assign io_52 = input_81;
assign io_52 = input_82;
assign io_52 = input_83;
assign io_52 = input_84;
assign io_52 = input_85;
assign io_52 = input_86;
assign io_52 = input_87;
assign io_52 = input_88;
assign io_52 = input_89;
assign io_52 = input_90;
assign io_52 = input_91;
assign io_52 = input_92;
assign io_52 = input_93;
assign io_52 = input_94;
assign io_52 = input_95;
assign io_53 = input_53;
assign io_53 = input_54;
assign io_53 = input_55;
assign io_53 = input_56;
assign io_53 = input_57;
assign io_53 = input_58;
assign io_53 = input_59;
assign io_53 = input_60;
assign io_53 = input_61;
assign io_53 = input_62;
assign io_53 = input_63;
assign io_53 = input_64;
assign io_53 = input_65;
assign io_53 = input_66;
assign io_53 = input_67;
assign io_53 = input_68;
assign io_53 = input_69;
assign io_53 = input_70;
assign io_53 = input_71;
assign io_53 = input_72;
assign io_53 = input_73;
assign io_53 = input_74;
assign io_53 = input_75;
assign io_53 = input_76;
assign io_53 = input_77;
assign io_53 = input_78;
assign io_53 = input_79;
assign io_53 = input_80;
assign io_53 = input_81;
assign io_53 = input_82;
assign io_53 = input_83;
assign io_53 = input_84;
assign io_53 = input_85;
assign io_53 = input_86;
assign io_53 = input_87;
assign io_53 = input_88;
assign io_53 = input_89;
assign io_53 = input_90;
assign io_53 = input_91;
assign io_53 = input_92;
assign io_53 = input_93;
assign io_53 = input_94;
assign io_53 = input_95;
assign io_54 = input_54;
assign io_54 = input_55;
assign io_54 = input_56;
assign io_54 = input_57;
assign io_54 = input_58;
assign io_54 = input_59;
assign io_54 = input_60;
assign io_54 = input_61;
assign io_54 = input_62;
assign io_54 = input_63;
assign io_54 = input_64;
assign io_54 = input_65;
assign io_54 = input_66;
assign io_54 = input_67;
assign io_54 = input_68;
assign io_54 = input_69;
assign io_54 = input_70;
assign io_54 = input_71;
assign io_54 = input_72;
assign io_54 = input_73;
assign io_54 = input_74;
assign io_54 = input_75;
assign io_54 = input_76;
assign io_54 = input_77;
assign io_54 = input_78;
assign io_54 = input_79;
assign io_54 = input_80;
assign io_54 = input_81;
assign io_54 = input_82;
assign io_54 = input_83;
assign io_54 = input_84;
assign io_54 = input_85;
assign io_54 = input_86;
assign io_54 = input_87;
assign io_54 = input_88;
assign io_54 = input_89;
assign io_54 = input_90;
assign io_54 = input_91;
assign io_54 = input_92;
assign io_54 = input_93;
assign io_54 = input_94;
assign io_54 = input_95;
assign io_55 = input_55;
assign io_55 = input_56;
assign io_55 = input_57;
assign io_55 = input_58;
assign io_55 = input_59;
assign io_55 = input_60;
assign io_55 = input_61;
assign io_55 = input_62;
assign io_55 = input_63;
assign io_55 = input_64;
assign io_55 = input_65;
assign io_55 = input_66;
assign io_55 = input_67;
assign io_55 = input_68;
assign io_55 = input_69;
assign io_55 = input_70;
assign io_55 = input_71;
assign io_55 = input_72;
assign io_55 = input_73;
assign io_55 = input_74;
assign io_55 = input_75;
assign io_55 = input_76;
assign io_55 = input_77;
assign io_55 = input_78;
assign io_55 = input_79;
assign io_55 = input_80;
assign io_55 = input_81;
assign io_55 = input_82;
assign io_55 = input_83;
assign io_55 = input_84;
assign io_55 = input_85;
assign io_55 = input_86;
assign io_55 = input_87;
assign io_55 = input_88;
assign io_55 = input_89;
assign io_55 = input_90;
assign io_55 = input_91;
assign io_55 = input_92;
assign io_55 = input_93;
assign io_55 = input_94;
assign io_55 = input_95;
assign io_56 = input_56;
assign io_56 = input_57;
assign io_56 = input_58;
assign io_56 = input_59;
assign io_56 = input_60;
assign io_56 = input_61;
assign io_56 = input_62;
assign io_56 = input_63;
assign io_56 = input_64;
assign io_56 = input_65;
assign io_56 = input_66;
assign io_56 = input_67;
assign io_56 = input_68;
assign io_56 = input_69;
assign io_56 = input_70;
assign io_56 = input_71;
assign io_56 = input_72;
assign io_56 = input_73;
assign io_56 = input_74;
assign io_56 = input_75;
assign io_56 = input_76;
assign io_56 = input_77;
assign io_56 = input_78;
assign io_56 = input_79;
assign io_56 = input_80;
assign io_56 = input_81;
assign io_56 = input_82;
assign io_56 = input_83;
assign io_56 = input_84;
assign io_56 = input_85;
assign io_56 = input_86;
assign io_56 = input_87;
assign io_56 = input_88;
assign io_56 = input_89;
assign io_56 = input_90;
assign io_56 = input_91;
assign io_56 = input_92;
assign io_56 = input_93;
assign io_56 = input_94;
assign io_56 = input_95;
assign io_57 = input_57;
assign io_57 = input_58;
assign io_57 = input_59;
assign io_57 = input_60;
assign io_57 = input_61;
assign io_57 = input_62;
assign io_57 = input_63;
assign io_57 = input_64;
assign io_57 = input_65;
assign io_57 = input_66;
assign io_57 = input_67;
assign io_57 = input_68;
assign io_57 = input_69;
assign io_57 = input_70;
assign io_57 = input_71;
assign io_57 = input_72;
assign io_57 = input_73;
assign io_57 = input_74;
assign io_57 = input_75;
assign io_57 = input_76;
assign io_57 = input_77;
assign io_57 = input_78;
assign io_57 = input_79;
assign io_57 = input_80;
assign io_57 = input_81;
assign io_57 = input_82;
assign io_57 = input_83;
assign io_57 = input_84;
assign io_57 = input_85;
assign io_57 = input_86;
assign io_57 = input_87;
assign io_57 = input_88;
assign io_57 = input_89;
assign io_57 = input_90;
assign io_57 = input_91;
assign io_57 = input_92;
assign io_57 = input_93;
assign io_57 = input_94;
assign io_57 = input_95;
assign io_58 = input_58;
assign io_58 = input_59;
assign io_58 = input_60;
assign io_58 = input_61;
assign io_58 = input_62;
assign io_58 = input_63;
assign io_58 = input_64;
assign io_58 = input_65;
assign io_58 = input_66;
assign io_58 = input_67;
assign io_58 = input_68;
assign io_58 = input_69;
assign io_58 = input_70;
assign io_58 = input_71;
assign io_58 = input_72;
assign io_58 = input_73;
assign io_58 = input_74;
assign io_58 = input_75;
assign io_58 = input_76;
assign io_58 = input_77;
assign io_58 = input_78;
assign io_58 = input_79;
assign io_58 = input_80;
assign io_58 = input_81;
assign io_58 = input_82;
assign io_58 = input_83;
assign io_58 = input_84;
assign io_58 = input_85;
assign io_58 = input_86;
assign io_58 = input_87;
assign io_58 = input_88;
assign io_58 = input_89;
assign io_58 = input_90;
assign io_58 = input_91;
assign io_58 = input_92;
assign io_58 = input_93;
assign io_58 = input_94;
assign io_58 = input_95;
assign io_59 = input_59;
assign io_59 = input_60;
assign io_59 = input_61;
assign io_59 = input_62;
assign io_59 = input_63;
assign io_59 = input_64;
assign io_59 = input_65;
assign io_59 = input_66;
assign io_59 = input_67;
assign io_59 = input_68;
assign io_59 = input_69;
assign io_59 = input_70;
assign io_59 = input_71;
assign io_59 = input_72;
assign io_59 = input_73;
assign io_59 = input_74;
assign io_59 = input_75;
assign io_59 = input_76;
assign io_59 = input_77;
assign io_59 = input_78;
assign io_59 = input_79;
assign io_59 = input_80;
assign io_59 = input_81;
assign io_59 = input_82;
assign io_59 = input_83;
assign io_59 = input_84;
assign io_59 = input_85;
assign io_59 = input_86;
assign io_59 = input_87;
assign io_59 = input_88;
assign io_59 = input_89;
assign io_59 = input_90;
assign io_59 = input_91;
assign io_59 = input_92;
assign io_59 = input_93;
assign io_59 = input_94;
assign io_59 = input_95;
assign io_60 = input_60;
assign io_60 = input_61;
assign io_60 = input_62;
assign io_60 = input_63;
assign io_60 = input_64;
assign io_60 = input_65;
assign io_60 = input_66;
assign io_60 = input_67;
assign io_60 = input_68;
assign io_60 = input_69;
assign io_60 = input_70;
assign io_60 = input_71;
assign io_60 = input_72;
assign io_60 = input_73;
assign io_60 = input_74;
assign io_60 = input_75;
assign io_60 = input_76;
assign io_60 = input_77;
assign io_60 = input_78;
assign io_60 = input_79;
assign io_60 = input_80;
assign io_60 = input_81;
assign io_60 = input_82;
assign io_60 = input_83;
assign io_60 = input_84;
assign io_60 = input_85;
assign io_60 = input_86;
assign io_60 = input_87;
assign io_60 = input_88;
assign io_60 = input_89;
assign io_60 = input_90;
assign io_60 = input_91;
assign io_60 = input_92;
assign io_60 = input_93;
assign io_60 = input_94;
assign io_60 = input_95;
assign io_61 = input_61;
assign io_61 = input_62;
assign io_61 = input_63;
assign io_61 = input_64;
assign io_61 = input_65;
assign io_61 = input_66;
assign io_61 = input_67;
assign io_61 = input_68;
assign io_61 = input_69;
assign io_61 = input_70;
assign io_61 = input_71;
assign io_61 = input_72;
assign io_61 = input_73;
assign io_61 = input_74;
assign io_61 = input_75;
assign io_61 = input_76;
assign io_61 = input_77;
assign io_61 = input_78;
assign io_61 = input_79;
assign io_61 = input_80;
assign io_61 = input_81;
assign io_61 = input_82;
assign io_61 = input_83;
assign io_61 = input_84;
assign io_61 = input_85;
assign io_61 = input_86;
assign io_61 = input_87;
assign io_61 = input_88;
assign io_61 = input_89;
assign io_61 = input_90;
assign io_61 = input_91;
assign io_61 = input_92;
assign io_61 = input_93;
assign io_61 = input_94;
assign io_61 = input_95;
assign io_62 = input_62;
assign io_62 = input_63;
assign io_62 = input_64;
assign io_62 = input_65;
assign io_62 = input_66;
assign io_62 = input_67;
assign io_62 = input_68;
assign io_62 = input_69;
assign io_62 = input_70;
assign io_62 = input_71;
assign io_62 = input_72;
assign io_62 = input_73;
assign io_62 = input_74;
assign io_62 = input_75;
assign io_62 = input_76;
assign io_62 = input_77;
assign io_62 = input_78;
assign io_62 = input_79;
assign io_62 = input_80;
assign io_62 = input_81;
assign io_62 = input_82;
assign io_62 = input_83;
assign io_62 = input_84;
assign io_62 = input_85;
assign io_62 = input_86;
assign io_62 = input_87;
assign io_62 = input_88;
assign io_62 = input_89;
assign io_62 = input_90;
assign io_62 = input_91;
assign io_62 = input_92;
assign io_62 = input_93;
assign io_62 = input_94;
assign io_62 = input_95;
assign io_63 = input_63;
assign io_63 = input_64;
assign io_63 = input_65;
assign io_63 = input_66;
assign io_63 = input_67;
assign io_63 = input_68;
assign io_63 = input_69;
assign io_63 = input_70;
assign io_63 = input_71;
assign io_63 = input_72;
assign io_63 = input_73;
assign io_63 = input_74;
assign io_63 = input_75;
assign io_63 = input_76;
assign io_63 = input_77;
assign io_63 = input_78;
assign io_63 = input_79;
assign io_63 = input_80;
assign io_63 = input_81;
assign io_63 = input_82;
assign io_63 = input_83;
assign io_63 = input_84;
assign io_63 = input_85;
assign io_63 = input_86;
assign io_63 = input_87;
assign io_63 = input_88;
assign io_63 = input_89;
assign io_63 = input_90;
assign io_63 = input_91;
assign io_63 = input_92;
assign io_63 = input_93;
assign io_63 = input_94;
assign io_63 = input_95;
assign io_64 = input_64;
assign io_64 = input_65;
assign io_64 = input_66;
assign io_64 = input_67;
assign io_64 = input_68;
assign io_64 = input_69;
assign io_64 = input_70;
assign io_64 = input_71;
assign io_64 = input_72;
assign io_64 = input_73;
assign io_64 = input_74;
assign io_64 = input_75;
assign io_64 = input_76;
assign io_64 = input_77;
assign io_64 = input_78;
assign io_64 = input_79;
assign io_64 = input_80;
assign io_64 = input_81;
assign io_64 = input_82;
assign io_64 = input_83;
assign io_64 = input_84;
assign io_64 = input_85;
assign io_64 = input_86;
assign io_64 = input_87;
assign io_64 = input_88;
assign io_64 = input_89;
assign io_64 = input_90;
assign io_64 = input_91;
assign io_64 = input_92;
assign io_64 = input_93;
assign io_64 = input_94;
assign io_64 = input_95;
assign io_65 = input_65;
assign io_65 = input_66;
assign io_65 = input_67;
assign io_65 = input_68;
assign io_65 = input_69;
assign io_65 = input_70;
assign io_65 = input_71;
assign io_65 = input_72;
assign io_65 = input_73;
assign io_65 = input_74;
assign io_65 = input_75;
assign io_65 = input_76;
assign io_65 = input_77;
assign io_65 = input_78;
assign io_65 = input_79;
assign io_65 = input_80;
assign io_65 = input_81;
assign io_65 = input_82;
assign io_65 = input_83;
assign io_65 = input_84;
assign io_65 = input_85;
assign io_65 = input_86;
assign io_65 = input_87;
assign io_65 = input_88;
assign io_65 = input_89;
assign io_65 = input_90;
assign io_65 = input_91;
assign io_65 = input_92;
assign io_65 = input_93;
assign io_65 = input_94;
assign io_65 = input_95;
assign io_66 = input_66;
assign io_66 = input_67;
assign io_66 = input_68;
assign io_66 = input_69;
assign io_66 = input_70;
assign io_66 = input_71;
assign io_66 = input_72;
assign io_66 = input_73;
assign io_66 = input_74;
assign io_66 = input_75;
assign io_66 = input_76;
assign io_66 = input_77;
assign io_66 = input_78;
assign io_66 = input_79;
assign io_66 = input_80;
assign io_66 = input_81;
assign io_66 = input_82;
assign io_66 = input_83;
assign io_66 = input_84;
assign io_66 = input_85;
assign io_66 = input_86;
assign io_66 = input_87;
assign io_66 = input_88;
assign io_66 = input_89;
assign io_66 = input_90;
assign io_66 = input_91;
assign io_66 = input_92;
assign io_66 = input_93;
assign io_66 = input_94;
assign io_66 = input_95;
assign io_67 = input_67;
assign io_67 = input_68;
assign io_67 = input_69;
assign io_67 = input_70;
assign io_67 = input_71;
assign io_67 = input_72;
assign io_67 = input_73;
assign io_67 = input_74;
assign io_67 = input_75;
assign io_67 = input_76;
assign io_67 = input_77;
assign io_67 = input_78;
assign io_67 = input_79;
assign io_67 = input_80;
assign io_67 = input_81;
assign io_67 = input_82;
assign io_67 = input_83;
assign io_67 = input_84;
assign io_67 = input_85;
assign io_67 = input_86;
assign io_67 = input_87;
assign io_67 = input_88;
assign io_67 = input_89;
assign io_67 = input_90;
assign io_67 = input_91;
assign io_67 = input_92;
assign io_67 = input_93;
assign io_67 = input_94;
assign io_67 = input_95;
assign io_68 = input_68;
assign io_68 = input_69;
assign io_68 = input_70;
assign io_68 = input_71;
assign io_68 = input_72;
assign io_68 = input_73;
assign io_68 = input_74;
assign io_68 = input_75;
assign io_68 = input_76;
assign io_68 = input_77;
assign io_68 = input_78;
assign io_68 = input_79;
assign io_68 = input_80;
assign io_68 = input_81;
assign io_68 = input_82;
assign io_68 = input_83;
assign io_68 = input_84;
assign io_68 = input_85;
assign io_68 = input_86;
assign io_68 = input_87;
assign io_68 = input_88;
assign io_68 = input_89;
assign io_68 = input_90;
assign io_68 = input_91;
assign io_68 = input_92;
assign io_68 = input_93;
assign io_68 = input_94;
assign io_68 = input_95;
assign io_69 = input_69;
assign io_69 = input_70;
assign io_69 = input_71;
assign io_69 = input_72;
assign io_69 = input_73;
assign io_69 = input_74;
assign io_69 = input_75;
assign io_69 = input_76;
assign io_69 = input_77;
assign io_69 = input_78;
assign io_69 = input_79;
assign io_69 = input_80;
assign io_69 = input_81;
assign io_69 = input_82;
assign io_69 = input_83;
assign io_69 = input_84;
assign io_69 = input_85;
assign io_69 = input_86;
assign io_69 = input_87;
assign io_69 = input_88;
assign io_69 = input_89;
assign io_69 = input_90;
assign io_69 = input_91;
assign io_69 = input_92;
assign io_69 = input_93;
assign io_69 = input_94;
assign io_69 = input_95;
assign io_70 = input_70;
assign io_70 = input_71;
assign io_70 = input_72;
assign io_70 = input_73;
assign io_70 = input_74;
assign io_70 = input_75;
assign io_70 = input_76;
assign io_70 = input_77;
assign io_70 = input_78;
assign io_70 = input_79;
assign io_70 = input_80;
assign io_70 = input_81;
assign io_70 = input_82;
assign io_70 = input_83;
assign io_70 = input_84;
assign io_70 = input_85;
assign io_70 = input_86;
assign io_70 = input_87;
assign io_70 = input_88;
assign io_70 = input_89;
assign io_70 = input_90;
assign io_70 = input_91;
assign io_70 = input_92;
assign io_70 = input_93;
assign io_70 = input_94;
assign io_70 = input_95;
assign io_71 = input_71;
assign io_71 = input_72;
assign io_71 = input_73;
assign io_71 = input_74;
assign io_71 = input_75;
assign io_71 = input_76;
assign io_71 = input_77;
assign io_71 = input_78;
assign io_71 = input_79;
assign io_71 = input_80;
assign io_71 = input_81;
assign io_71 = input_82;
assign io_71 = input_83;
assign io_71 = input_84;
assign io_71 = input_85;
assign io_71 = input_86;
assign io_71 = input_87;
assign io_71 = input_88;
assign io_71 = input_89;
assign io_71 = input_90;
assign io_71 = input_91;
assign io_71 = input_92;
assign io_71 = input_93;
assign io_71 = input_94;
assign io_71 = input_95;
assign io_72 = input_72;
assign io_72 = input_73;
assign io_72 = input_74;
assign io_72 = input_75;
assign io_72 = input_76;
assign io_72 = input_77;
assign io_72 = input_78;
assign io_72 = input_79;
assign io_72 = input_80;
assign io_72 = input_81;
assign io_72 = input_82;
assign io_72 = input_83;
assign io_72 = input_84;
assign io_72 = input_85;
assign io_72 = input_86;
assign io_72 = input_87;
assign io_72 = input_88;
assign io_72 = input_89;
assign io_72 = input_90;
assign io_72 = input_91;
assign io_72 = input_92;
assign io_72 = input_93;
assign io_72 = input_94;
assign io_72 = input_95;
assign io_73 = input_73;
assign io_73 = input_74;
assign io_73 = input_75;
assign io_73 = input_76;
assign io_73 = input_77;
assign io_73 = input_78;
assign io_73 = input_79;
assign io_73 = input_80;
assign io_73 = input_81;
assign io_73 = input_82;
assign io_73 = input_83;
assign io_73 = input_84;
assign io_73 = input_85;
assign io_73 = input_86;
assign io_73 = input_87;
assign io_73 = input_88;
assign io_73 = input_89;
assign io_73 = input_90;
assign io_73 = input_91;
assign io_73 = input_92;
assign io_73 = input_93;
assign io_73 = input_94;
assign io_73 = input_95;
assign io_74 = input_74;
assign io_74 = input_75;
assign io_74 = input_76;
assign io_74 = input_77;
assign io_74 = input_78;
assign io_74 = input_79;
assign io_74 = input_80;
assign io_74 = input_81;
assign io_74 = input_82;
assign io_74 = input_83;
assign io_74 = input_84;
assign io_74 = input_85;
assign io_74 = input_86;
assign io_74 = input_87;
assign io_74 = input_88;
assign io_74 = input_89;
assign io_74 = input_90;
assign io_74 = input_91;
assign io_74 = input_92;
assign io_74 = input_93;
assign io_74 = input_94;
assign io_74 = input_95;
assign io_75 = input_75;
assign io_75 = input_76;
assign io_75 = input_77;
assign io_75 = input_78;
assign io_75 = input_79;
assign io_75 = input_80;
assign io_75 = input_81;
assign io_75 = input_82;
assign io_75 = input_83;
assign io_75 = input_84;
assign io_75 = input_85;
assign io_75 = input_86;
assign io_75 = input_87;
assign io_75 = input_88;
assign io_75 = input_89;
assign io_75 = input_90;
assign io_75 = input_91;
assign io_75 = input_92;
assign io_75 = input_93;
assign io_75 = input_94;
assign io_75 = input_95;
assign io_76 = input_76;
assign io_76 = input_77;
assign io_76 = input_78;
assign io_76 = input_79;
assign io_76 = input_80;
assign io_76 = input_81;
assign io_76 = input_82;
assign io_76 = input_83;
assign io_76 = input_84;
assign io_76 = input_85;
assign io_76 = input_86;
assign io_76 = input_87;
assign io_76 = input_88;
assign io_76 = input_89;
assign io_76 = input_90;
assign io_76 = input_91;
assign io_76 = input_92;
assign io_76 = input_93;
assign io_76 = input_94;
assign io_76 = input_95;
assign io_77 = input_77;
assign io_77 = input_78;
assign io_77 = input_79;
assign io_77 = input_80;
assign io_77 = input_81;
assign io_77 = input_82;
assign io_77 = input_83;
assign io_77 = input_84;
assign io_77 = input_85;
assign io_77 = input_86;
assign io_77 = input_87;
assign io_77 = input_88;
assign io_77 = input_89;
assign io_77 = input_90;
assign io_77 = input_91;
assign io_77 = input_92;
assign io_77 = input_93;
assign io_77 = input_94;
assign io_77 = input_95;
assign io_78 = input_78;
assign io_78 = input_79;
assign io_78 = input_80;
assign io_78 = input_81;
assign io_78 = input_82;
assign io_78 = input_83;
assign io_78 = input_84;
assign io_78 = input_85;
assign io_78 = input_86;
assign io_78 = input_87;
assign io_78 = input_88;
assign io_78 = input_89;
assign io_78 = input_90;
assign io_78 = input_91;
assign io_78 = input_92;
assign io_78 = input_93;
assign io_78 = input_94;
assign io_78 = input_95;
assign io_79 = input_79;
assign io_79 = input_80;
assign io_79 = input_81;
assign io_79 = input_82;
assign io_79 = input_83;
assign io_79 = input_84;
assign io_79 = input_85;
assign io_79 = input_86;
assign io_79 = input_87;
assign io_79 = input_88;
assign io_79 = input_89;
assign io_79 = input_90;
assign io_79 = input_91;
assign io_79 = input_92;
assign io_79 = input_93;
assign io_79 = input_94;
assign io_79 = input_95;
assign io_80 = input_80;
assign io_80 = input_81;
assign io_80 = input_82;
assign io_80 = input_83;
assign io_80 = input_84;
assign io_80 = input_85;
assign io_80 = input_86;
assign io_80 = input_87;
assign io_80 = input_88;
assign io_80 = input_89;
assign io_80 = input_90;
assign io_80 = input_91;
assign io_80 = input_92;
assign io_80 = input_93;
assign io_80 = input_94;
assign io_80 = input_95;
assign io_81 = input_81;
assign io_81 = input_82;
assign io_81 = input_83;
assign io_81 = input_84;
assign io_81 = input_85;
assign io_81 = input_86;
assign io_81 = input_87;
assign io_81 = input_88;
assign io_81 = input_89;
assign io_81 = input_90;
assign io_81 = input_91;
assign io_81 = input_92;
assign io_81 = input_93;
assign io_81 = input_94;
assign io_81 = input_95;
assign io_82 = input_82;
assign io_82 = input_83;
assign io_82 = input_84;
assign io_82 = input_85;
assign io_82 = input_86;
assign io_82 = input_87;
assign io_82 = input_88;
assign io_82 = input_89;
assign io_82 = input_90;
assign io_82 = input_91;
assign io_82 = input_92;
assign io_82 = input_93;
assign io_82 = input_94;
assign io_82 = input_95;
assign io_83 = input_83;
assign io_83 = input_84;
assign io_83 = input_85;
assign io_83 = input_86;
assign io_83 = input_87;
assign io_83 = input_88;
assign io_83 = input_89;
assign io_83 = input_90;
assign io_83 = input_91;
assign io_83 = input_92;
assign io_83 = input_93;
assign io_83 = input_94;
assign io_83 = input_95;
assign io_84 = input_84;
assign io_84 = input_85;
assign io_84 = input_86;
assign io_84 = input_87;
assign io_84 = input_88;
assign io_84 = input_89;
assign io_84 = input_90;
assign io_84 = input_91;
assign io_84 = input_92;
assign io_84 = input_93;
assign io_84 = input_94;
assign io_84 = input_95;
assign io_85 = input_85;
assign io_85 = input_86;
assign io_85 = input_87;
assign io_85 = input_88;
assign io_85 = input_89;
assign io_85 = input_90;
assign io_85 = input_91;
assign io_85 = input_92;
assign io_85 = input_93;
assign io_85 = input_94;
assign io_85 = input_95;
assign io_86 = input_86;
assign io_86 = input_87;
assign io_86 = input_88;
assign io_86 = input_89;
assign io_86 = input_90;
assign io_86 = input_91;
assign io_86 = input_92;
assign io_86 = input_93;
assign io_86 = input_94;
assign io_86 = input_95;
assign io_87 = input_87;
assign io_87 = input_88;
assign io_87 = input_89;
assign io_87 = input_90;
assign io_87 = input_91;
assign io_87 = input_92;
assign io_87 = input_93;
assign io_87 = input_94;
assign io_87 = input_95;
assign io_88 = input_88;
assign io_88 = input_89;
assign io_88 = input_90;
assign io_88 = input_91;
assign io_88 = input_92;
assign io_88 = input_93;
assign io_88 = input_94;
assign io_88 = input_95;
assign io_89 = input_89;
assign io_89 = input_90;
assign io_89 = input_91;
assign io_89 = input_92;
assign io_89 = input_93;
assign io_89 = input_94;
assign io_89 = input_95;
assign io_90 = input_90;
assign io_90 = input_91;
assign io_90 = input_92;
assign io_90 = input_93;
assign io_90 = input_94;
assign io_90 = input_95;
assign io_91 = input_91;
assign io_91 = input_92;
assign io_91 = input_93;
assign io_91 = input_94;
assign io_91 = input_95;
assign io_92 = input_92;
assign io_92 = input_93;
assign io_92 = input_94;
assign io_92 = input_95;
assign io_93 = input_93;
assign io_93 = input_94;
assign io_93 = input_95;
assign io_94 = input_94;
assign io_94 = input_95;
assign io_95 = input_95;
endmodule
