module fanout2_braid_3_16 (
output output_0,output output_1,output output_2,input input_0,input input_1,input input_2
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_1_2, output_1_0, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_0), .y(output_0_2));
wire output_2_2, output_2_0, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_0), .y(output_1_2));
wire output_3_2, output_3_0, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_0), .y(output_2_2));
wire output_1_3, output_1_1, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_1), .y(output_0_3));
wire output_2_3, output_2_1, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_1), .y(output_1_3));
wire output_3_3, output_3_1, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_1), .y(output_2_3));
wire output_1_4, output_1_2, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_2), .y(output_0_4));
wire output_2_4, output_2_2, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_2), .y(output_1_4));
wire output_3_4, output_3_2, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_2), .y(output_2_4));
wire output_1_5, output_1_0, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_0), .y(output_0_5));
wire output_2_5, output_2_0, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_0), .y(output_1_5));
wire output_3_5, output_3_0, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_0), .y(output_2_5));
wire output_1_6, output_1_1, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_1), .y(output_0_6));
wire output_2_6, output_2_1, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_1), .y(output_1_6));
wire output_3_6, output_3_1, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_1), .y(output_2_6));
wire output_1_7, output_1_2, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_2), .y(output_0_7));
wire output_2_7, output_2_2, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_2), .y(output_1_7));
wire output_3_7, output_3_2, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_2), .y(output_2_7));
wire output_1_8, output_1_0, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_0), .y(output_0_8));
wire output_2_8, output_2_0, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_0), .y(output_1_8));
wire output_3_8, output_3_0, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_0), .y(output_2_8));
wire output_1_9, output_1_1, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_1), .y(output_0_9));
wire output_2_9, output_2_1, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_1), .y(output_1_9));
wire output_3_9, output_3_1, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_1), .y(output_2_9));
wire output_1_10, output_1_2, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_2), .y(output_0_10));
wire output_2_10, output_2_2, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_2), .y(output_1_10));
wire output_3_10, output_3_2, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_2), .y(output_2_10));
wire output_1_11, output_1_0, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_0), .y(output_0_11));
wire output_2_11, output_2_0, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_0), .y(output_1_11));
wire output_3_11, output_3_0, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_0), .y(output_2_11));
wire output_1_12, output_1_1, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_1), .y(output_0_12));
wire output_2_12, output_2_1, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_1), .y(output_1_12));
wire output_3_12, output_3_1, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_1), .y(output_2_12));
wire output_1_13, output_1_2, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_2), .y(output_0_13));
wire output_2_13, output_2_2, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_2), .y(output_1_13));
wire output_3_13, output_3_2, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_2), .y(output_2_13));
wire output_1_14, output_1_0, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_0), .y(output_0_14));
wire output_2_14, output_2_0, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_0), .y(output_1_14));
wire output_3_14, output_3_0, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_0), .y(output_2_14));
wire output_1_15, output_1_1, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_1), .y(output_0_15));
wire output_2_15, output_2_1, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_1), .y(output_1_15));
wire output_3_15, output_3_1, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_1), .y(output_2_15));
assign output_0 = output_0_0;
wire output_0_16;
assign output_0_16 = input_0;
assign output_1 = output_1_0;
wire output_1_16;
assign output_1_16 = input_1;
assign output_2 = output_2_0;
wire output_2_16;
assign output_2_16 = input_2;
endmodule
