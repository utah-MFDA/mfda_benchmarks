// Device H
module logic04 (
inout b0_1, b0_2, b0_3, b0_3, b0_4, b0_5, b0_6, b0_7, b0_8, b4_1, b4_2, b4_3, b4_4, b4_5, b5_1, b5_2, b5_3, b5_4, b1_1, b1_2, b1_3, b1_4, b1_5, b3_1, b3_2, b3_3, b3_4, b3_5, b2_1, b2_2, b2_3, b2_4, b2_5, b2_6, b2_7, b2_8, b2_9, b2_10
);
wire c0;
wire c1;
wire c2;
wire c3;
wire c4;
wire c5;
wire c6;
wire c7;
wire c8;
wire c9;
wire c10;
wire c11;
wire cc21;
wire cc22;
wire cc23;
wire cc24;
wire cc25;
wire cc26;
wire cca;
wire ccb;
wire ccc;
wire cc10;
wire cc11;
wire cc9;
wire cc12;
wire cc8;
wire cc13;
wire cc7;
wire cc14;
wire cc6;
wire cc15;
wire cc1;
wire cc5;
wire cc2;
wire cc4;
wire cc3;
wire cc16;
wire cc17;
wire cc18;
wire cc19;
wire cc20;
LOGIC ARRAY la(.port1(c3),.port24(cca),.port25(ccb),.port26(ccc),.port13(cc10),.port14(cc11),.port12(cc9),.port15(cc12),.port11(cc8),.port16(cc13),.port10(cc7),.port17(cc14),.port9(cc6),.port18(cc15),.port3(c1),.port3(c1),.port4(cc1),.port8(cc5),.port5(cc2),.port7(cc4),.port6(cc3),.port19(cc16),.port20(cc17),.port21(cc18),.port22(cc19),.port23(cc20));
assign c4 = b0_1;
assign c5 = b0_2;
assign c6 = b0_3;
assign c6 = b0_3;
assign c7 = b0_4;
assign c8 = b0_5;
assign c9 = b0_6;
assign c10 = b0_7;
assign c11 = b0_8;
MUX m1(.port9(c0),.port10(cc21),.port11(cc22),.port12(cc23),.port13(cc24),.port14(cc25),.port15(cc26),.port1(c4),.port2(c5),.port3(c6),.port4(c7),.port5(c8),.port6(c9),.port7(c10),.port8(c11));
NODE n1(.port0(c1),.port0(c1),.port0(c0),.port0(c3));
assign cc21 = b4_1;
assign cc23 = b4_2;
assign cc25 = b4_3;
assign cca = b4_4;
assign ccb = b4_5;
assign cc22 = b5_1;
assign cc24 = b5_2;
assign cc26 = b5_3;
assign ccc = b5_4;
assign cc1 = b1_1;
assign cc2 = b1_2;
assign cc3 = b1_3;
assign cc4 = b1_4;
assign cc5 = b1_5;
assign cc16 = b3_1;
assign cc17 = b3_2;
assign cc18 = b3_3;
assign cc19 = b3_4;
assign cc20 = b3_5;
assign cc6 = b2_1;
assign cc7 = b2_2;
assign cc8 = b2_3;
assign cc9 = b2_4;
assign cc10 = b2_5;
assign cc11 = b2_6;
assign cc12 = b2_7;
assign cc13 = b2_8;
assign cc14 = b2_9;
assign cc15 = b2_10;
endmodule
