module fanout2_braid_4_256 (
output output_0,output output_1,output output_2,output output_3,input input_0,input input_1,input input_2,input input_3
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_1_3, output_1_0, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_0), .y(output_0_3));
wire output_2_3, output_2_0, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_0), .y(output_1_3));
wire output_3_3, output_3_0, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_0), .y(output_2_3));
wire output_4_3, output_4_0, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_0), .y(output_3_3));
wire output_1_4, output_1_1, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_1), .y(output_0_4));
wire output_2_4, output_2_1, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_1), .y(output_1_4));
wire output_3_4, output_3_1, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_1), .y(output_2_4));
wire output_4_4, output_4_1, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_1), .y(output_3_4));
wire output_1_5, output_1_2, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_2), .y(output_0_5));
wire output_2_5, output_2_2, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_2), .y(output_1_5));
wire output_3_5, output_3_2, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_2), .y(output_2_5));
wire output_4_5, output_4_2, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_2), .y(output_3_5));
wire output_1_6, output_1_3, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_3), .y(output_0_6));
wire output_2_6, output_2_3, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_3), .y(output_1_6));
wire output_3_6, output_3_3, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_3), .y(output_2_6));
wire output_4_6, output_4_3, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_3), .y(output_3_6));
wire output_1_7, output_1_0, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_0), .y(output_0_7));
wire output_2_7, output_2_0, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_0), .y(output_1_7));
wire output_3_7, output_3_0, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_0), .y(output_2_7));
wire output_4_7, output_4_0, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_0), .y(output_3_7));
wire output_1_8, output_1_1, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_1), .y(output_0_8));
wire output_2_8, output_2_1, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_1), .y(output_1_8));
wire output_3_8, output_3_1, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_1), .y(output_2_8));
wire output_4_8, output_4_1, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_1), .y(output_3_8));
wire output_1_9, output_1_2, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_2), .y(output_0_9));
wire output_2_9, output_2_2, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_2), .y(output_1_9));
wire output_3_9, output_3_2, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_2), .y(output_2_9));
wire output_4_9, output_4_2, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_2), .y(output_3_9));
wire output_1_10, output_1_3, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_3), .y(output_0_10));
wire output_2_10, output_2_3, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_3), .y(output_1_10));
wire output_3_10, output_3_3, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_3), .y(output_2_10));
wire output_4_10, output_4_3, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_3), .y(output_3_10));
wire output_1_11, output_1_0, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_0), .y(output_0_11));
wire output_2_11, output_2_0, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_0), .y(output_1_11));
wire output_3_11, output_3_0, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_0), .y(output_2_11));
wire output_4_11, output_4_0, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_0), .y(output_3_11));
wire output_1_12, output_1_1, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_1), .y(output_0_12));
wire output_2_12, output_2_1, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_1), .y(output_1_12));
wire output_3_12, output_3_1, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_1), .y(output_2_12));
wire output_4_12, output_4_1, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_1), .y(output_3_12));
wire output_1_13, output_1_2, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_2), .y(output_0_13));
wire output_2_13, output_2_2, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_2), .y(output_1_13));
wire output_3_13, output_3_2, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_2), .y(output_2_13));
wire output_4_13, output_4_2, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_2), .y(output_3_13));
wire output_1_14, output_1_3, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_3), .y(output_0_14));
wire output_2_14, output_2_3, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_3), .y(output_1_14));
wire output_3_14, output_3_3, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_3), .y(output_2_14));
wire output_4_14, output_4_3, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_3), .y(output_3_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_1_16, output_1_1, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_1), .y(output_0_16));
wire output_2_16, output_2_1, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_1), .y(output_1_16));
wire output_3_16, output_3_1, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_1), .y(output_2_16));
wire output_4_16, output_4_1, output_3_16;
mixer gate_output_3_16(.a(output_4_16), .b(output_4_1), .y(output_3_16));
wire output_1_17, output_1_2, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_2), .y(output_0_17));
wire output_2_17, output_2_2, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_2), .y(output_1_17));
wire output_3_17, output_3_2, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_2), .y(output_2_17));
wire output_4_17, output_4_2, output_3_17;
mixer gate_output_3_17(.a(output_4_17), .b(output_4_2), .y(output_3_17));
wire output_1_18, output_1_3, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_3), .y(output_0_18));
wire output_2_18, output_2_3, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_3), .y(output_1_18));
wire output_3_18, output_3_3, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_3), .y(output_2_18));
wire output_4_18, output_4_3, output_3_18;
mixer gate_output_3_18(.a(output_4_18), .b(output_4_3), .y(output_3_18));
wire output_1_19, output_1_0, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_0), .y(output_0_19));
wire output_2_19, output_2_0, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_0), .y(output_1_19));
wire output_3_19, output_3_0, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_0), .y(output_2_19));
wire output_4_19, output_4_0, output_3_19;
mixer gate_output_3_19(.a(output_4_19), .b(output_4_0), .y(output_3_19));
wire output_1_20, output_1_1, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_1), .y(output_0_20));
wire output_2_20, output_2_1, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_1), .y(output_1_20));
wire output_3_20, output_3_1, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_1), .y(output_2_20));
wire output_4_20, output_4_1, output_3_20;
mixer gate_output_3_20(.a(output_4_20), .b(output_4_1), .y(output_3_20));
wire output_1_21, output_1_2, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_2), .y(output_0_21));
wire output_2_21, output_2_2, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_2), .y(output_1_21));
wire output_3_21, output_3_2, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_2), .y(output_2_21));
wire output_4_21, output_4_2, output_3_21;
mixer gate_output_3_21(.a(output_4_21), .b(output_4_2), .y(output_3_21));
wire output_1_22, output_1_3, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_3), .y(output_0_22));
wire output_2_22, output_2_3, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_3), .y(output_1_22));
wire output_3_22, output_3_3, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_3), .y(output_2_22));
wire output_4_22, output_4_3, output_3_22;
mixer gate_output_3_22(.a(output_4_22), .b(output_4_3), .y(output_3_22));
wire output_1_23, output_1_0, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_0), .y(output_0_23));
wire output_2_23, output_2_0, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_0), .y(output_1_23));
wire output_3_23, output_3_0, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_0), .y(output_2_23));
wire output_4_23, output_4_0, output_3_23;
mixer gate_output_3_23(.a(output_4_23), .b(output_4_0), .y(output_3_23));
wire output_1_24, output_1_1, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_1), .y(output_0_24));
wire output_2_24, output_2_1, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_1), .y(output_1_24));
wire output_3_24, output_3_1, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_1), .y(output_2_24));
wire output_4_24, output_4_1, output_3_24;
mixer gate_output_3_24(.a(output_4_24), .b(output_4_1), .y(output_3_24));
wire output_1_25, output_1_2, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_2), .y(output_0_25));
wire output_2_25, output_2_2, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_2), .y(output_1_25));
wire output_3_25, output_3_2, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_2), .y(output_2_25));
wire output_4_25, output_4_2, output_3_25;
mixer gate_output_3_25(.a(output_4_25), .b(output_4_2), .y(output_3_25));
wire output_1_26, output_1_3, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_3), .y(output_0_26));
wire output_2_26, output_2_3, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_3), .y(output_1_26));
wire output_3_26, output_3_3, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_3), .y(output_2_26));
wire output_4_26, output_4_3, output_3_26;
mixer gate_output_3_26(.a(output_4_26), .b(output_4_3), .y(output_3_26));
wire output_1_27, output_1_0, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_0), .y(output_0_27));
wire output_2_27, output_2_0, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_0), .y(output_1_27));
wire output_3_27, output_3_0, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_0), .y(output_2_27));
wire output_4_27, output_4_0, output_3_27;
mixer gate_output_3_27(.a(output_4_27), .b(output_4_0), .y(output_3_27));
wire output_1_28, output_1_1, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_1), .y(output_0_28));
wire output_2_28, output_2_1, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_1), .y(output_1_28));
wire output_3_28, output_3_1, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_1), .y(output_2_28));
wire output_4_28, output_4_1, output_3_28;
mixer gate_output_3_28(.a(output_4_28), .b(output_4_1), .y(output_3_28));
wire output_1_29, output_1_2, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_2), .y(output_0_29));
wire output_2_29, output_2_2, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_2), .y(output_1_29));
wire output_3_29, output_3_2, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_2), .y(output_2_29));
wire output_4_29, output_4_2, output_3_29;
mixer gate_output_3_29(.a(output_4_29), .b(output_4_2), .y(output_3_29));
wire output_1_30, output_1_3, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_3), .y(output_0_30));
wire output_2_30, output_2_3, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_3), .y(output_1_30));
wire output_3_30, output_3_3, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_3), .y(output_2_30));
wire output_4_30, output_4_3, output_3_30;
mixer gate_output_3_30(.a(output_4_30), .b(output_4_3), .y(output_3_30));
wire output_1_31, output_1_0, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_0), .y(output_0_31));
wire output_2_31, output_2_0, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_0), .y(output_1_31));
wire output_3_31, output_3_0, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_0), .y(output_2_31));
wire output_4_31, output_4_0, output_3_31;
mixer gate_output_3_31(.a(output_4_31), .b(output_4_0), .y(output_3_31));
wire output_1_32, output_1_1, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_1), .y(output_0_32));
wire output_2_32, output_2_1, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_1), .y(output_1_32));
wire output_3_32, output_3_1, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_1), .y(output_2_32));
wire output_4_32, output_4_1, output_3_32;
mixer gate_output_3_32(.a(output_4_32), .b(output_4_1), .y(output_3_32));
wire output_1_33, output_1_2, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_2), .y(output_0_33));
wire output_2_33, output_2_2, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_2), .y(output_1_33));
wire output_3_33, output_3_2, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_2), .y(output_2_33));
wire output_4_33, output_4_2, output_3_33;
mixer gate_output_3_33(.a(output_4_33), .b(output_4_2), .y(output_3_33));
wire output_1_34, output_1_3, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_3), .y(output_0_34));
wire output_2_34, output_2_3, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_3), .y(output_1_34));
wire output_3_34, output_3_3, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_3), .y(output_2_34));
wire output_4_34, output_4_3, output_3_34;
mixer gate_output_3_34(.a(output_4_34), .b(output_4_3), .y(output_3_34));
wire output_1_35, output_1_0, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_0), .y(output_0_35));
wire output_2_35, output_2_0, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_0), .y(output_1_35));
wire output_3_35, output_3_0, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_0), .y(output_2_35));
wire output_4_35, output_4_0, output_3_35;
mixer gate_output_3_35(.a(output_4_35), .b(output_4_0), .y(output_3_35));
wire output_1_36, output_1_1, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_1), .y(output_0_36));
wire output_2_36, output_2_1, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_1), .y(output_1_36));
wire output_3_36, output_3_1, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_1), .y(output_2_36));
wire output_4_36, output_4_1, output_3_36;
mixer gate_output_3_36(.a(output_4_36), .b(output_4_1), .y(output_3_36));
wire output_1_37, output_1_2, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_2), .y(output_0_37));
wire output_2_37, output_2_2, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_2), .y(output_1_37));
wire output_3_37, output_3_2, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_2), .y(output_2_37));
wire output_4_37, output_4_2, output_3_37;
mixer gate_output_3_37(.a(output_4_37), .b(output_4_2), .y(output_3_37));
wire output_1_38, output_1_3, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_3), .y(output_0_38));
wire output_2_38, output_2_3, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_3), .y(output_1_38));
wire output_3_38, output_3_3, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_3), .y(output_2_38));
wire output_4_38, output_4_3, output_3_38;
mixer gate_output_3_38(.a(output_4_38), .b(output_4_3), .y(output_3_38));
wire output_1_39, output_1_0, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_0), .y(output_0_39));
wire output_2_39, output_2_0, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_0), .y(output_1_39));
wire output_3_39, output_3_0, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_0), .y(output_2_39));
wire output_4_39, output_4_0, output_3_39;
mixer gate_output_3_39(.a(output_4_39), .b(output_4_0), .y(output_3_39));
wire output_1_40, output_1_1, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_1), .y(output_0_40));
wire output_2_40, output_2_1, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_1), .y(output_1_40));
wire output_3_40, output_3_1, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_1), .y(output_2_40));
wire output_4_40, output_4_1, output_3_40;
mixer gate_output_3_40(.a(output_4_40), .b(output_4_1), .y(output_3_40));
wire output_1_41, output_1_2, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_2), .y(output_0_41));
wire output_2_41, output_2_2, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_2), .y(output_1_41));
wire output_3_41, output_3_2, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_2), .y(output_2_41));
wire output_4_41, output_4_2, output_3_41;
mixer gate_output_3_41(.a(output_4_41), .b(output_4_2), .y(output_3_41));
wire output_1_42, output_1_3, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_3), .y(output_0_42));
wire output_2_42, output_2_3, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_3), .y(output_1_42));
wire output_3_42, output_3_3, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_3), .y(output_2_42));
wire output_4_42, output_4_3, output_3_42;
mixer gate_output_3_42(.a(output_4_42), .b(output_4_3), .y(output_3_42));
wire output_1_43, output_1_0, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_0), .y(output_0_43));
wire output_2_43, output_2_0, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_0), .y(output_1_43));
wire output_3_43, output_3_0, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_0), .y(output_2_43));
wire output_4_43, output_4_0, output_3_43;
mixer gate_output_3_43(.a(output_4_43), .b(output_4_0), .y(output_3_43));
wire output_1_44, output_1_1, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_1), .y(output_0_44));
wire output_2_44, output_2_1, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_1), .y(output_1_44));
wire output_3_44, output_3_1, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_1), .y(output_2_44));
wire output_4_44, output_4_1, output_3_44;
mixer gate_output_3_44(.a(output_4_44), .b(output_4_1), .y(output_3_44));
wire output_1_45, output_1_2, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_2), .y(output_0_45));
wire output_2_45, output_2_2, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_2), .y(output_1_45));
wire output_3_45, output_3_2, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_2), .y(output_2_45));
wire output_4_45, output_4_2, output_3_45;
mixer gate_output_3_45(.a(output_4_45), .b(output_4_2), .y(output_3_45));
wire output_1_46, output_1_3, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_3), .y(output_0_46));
wire output_2_46, output_2_3, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_3), .y(output_1_46));
wire output_3_46, output_3_3, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_3), .y(output_2_46));
wire output_4_46, output_4_3, output_3_46;
mixer gate_output_3_46(.a(output_4_46), .b(output_4_3), .y(output_3_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_4_47, output_4_0, output_3_47;
mixer gate_output_3_47(.a(output_4_47), .b(output_4_0), .y(output_3_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_4_48, output_4_1, output_3_48;
mixer gate_output_3_48(.a(output_4_48), .b(output_4_1), .y(output_3_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_4_49, output_4_2, output_3_49;
mixer gate_output_3_49(.a(output_4_49), .b(output_4_2), .y(output_3_49));
wire output_1_50, output_1_3, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_3), .y(output_0_50));
wire output_2_50, output_2_3, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_3), .y(output_1_50));
wire output_3_50, output_3_3, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_3), .y(output_2_50));
wire output_4_50, output_4_3, output_3_50;
mixer gate_output_3_50(.a(output_4_50), .b(output_4_3), .y(output_3_50));
wire output_1_51, output_1_0, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_0), .y(output_0_51));
wire output_2_51, output_2_0, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_0), .y(output_1_51));
wire output_3_51, output_3_0, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_0), .y(output_2_51));
wire output_4_51, output_4_0, output_3_51;
mixer gate_output_3_51(.a(output_4_51), .b(output_4_0), .y(output_3_51));
wire output_1_52, output_1_1, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_1), .y(output_0_52));
wire output_2_52, output_2_1, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_1), .y(output_1_52));
wire output_3_52, output_3_1, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_1), .y(output_2_52));
wire output_4_52, output_4_1, output_3_52;
mixer gate_output_3_52(.a(output_4_52), .b(output_4_1), .y(output_3_52));
wire output_1_53, output_1_2, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_2), .y(output_0_53));
wire output_2_53, output_2_2, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_2), .y(output_1_53));
wire output_3_53, output_3_2, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_2), .y(output_2_53));
wire output_4_53, output_4_2, output_3_53;
mixer gate_output_3_53(.a(output_4_53), .b(output_4_2), .y(output_3_53));
wire output_1_54, output_1_3, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_3), .y(output_0_54));
wire output_2_54, output_2_3, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_3), .y(output_1_54));
wire output_3_54, output_3_3, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_3), .y(output_2_54));
wire output_4_54, output_4_3, output_3_54;
mixer gate_output_3_54(.a(output_4_54), .b(output_4_3), .y(output_3_54));
wire output_1_55, output_1_0, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_0), .y(output_0_55));
wire output_2_55, output_2_0, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_0), .y(output_1_55));
wire output_3_55, output_3_0, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_0), .y(output_2_55));
wire output_4_55, output_4_0, output_3_55;
mixer gate_output_3_55(.a(output_4_55), .b(output_4_0), .y(output_3_55));
wire output_1_56, output_1_1, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_1), .y(output_0_56));
wire output_2_56, output_2_1, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_1), .y(output_1_56));
wire output_3_56, output_3_1, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_1), .y(output_2_56));
wire output_4_56, output_4_1, output_3_56;
mixer gate_output_3_56(.a(output_4_56), .b(output_4_1), .y(output_3_56));
wire output_1_57, output_1_2, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_2), .y(output_0_57));
wire output_2_57, output_2_2, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_2), .y(output_1_57));
wire output_3_57, output_3_2, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_2), .y(output_2_57));
wire output_4_57, output_4_2, output_3_57;
mixer gate_output_3_57(.a(output_4_57), .b(output_4_2), .y(output_3_57));
wire output_1_58, output_1_3, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_3), .y(output_0_58));
wire output_2_58, output_2_3, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_3), .y(output_1_58));
wire output_3_58, output_3_3, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_3), .y(output_2_58));
wire output_4_58, output_4_3, output_3_58;
mixer gate_output_3_58(.a(output_4_58), .b(output_4_3), .y(output_3_58));
wire output_1_59, output_1_0, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_0), .y(output_0_59));
wire output_2_59, output_2_0, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_0), .y(output_1_59));
wire output_3_59, output_3_0, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_0), .y(output_2_59));
wire output_4_59, output_4_0, output_3_59;
mixer gate_output_3_59(.a(output_4_59), .b(output_4_0), .y(output_3_59));
wire output_1_60, output_1_1, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_1), .y(output_0_60));
wire output_2_60, output_2_1, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_1), .y(output_1_60));
wire output_3_60, output_3_1, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_1), .y(output_2_60));
wire output_4_60, output_4_1, output_3_60;
mixer gate_output_3_60(.a(output_4_60), .b(output_4_1), .y(output_3_60));
wire output_1_61, output_1_2, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_2), .y(output_0_61));
wire output_2_61, output_2_2, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_2), .y(output_1_61));
wire output_3_61, output_3_2, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_2), .y(output_2_61));
wire output_4_61, output_4_2, output_3_61;
mixer gate_output_3_61(.a(output_4_61), .b(output_4_2), .y(output_3_61));
wire output_1_62, output_1_3, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_3), .y(output_0_62));
wire output_2_62, output_2_3, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_3), .y(output_1_62));
wire output_3_62, output_3_3, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_3), .y(output_2_62));
wire output_4_62, output_4_3, output_3_62;
mixer gate_output_3_62(.a(output_4_62), .b(output_4_3), .y(output_3_62));
wire output_1_63, output_1_0, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_0), .y(output_0_63));
wire output_2_63, output_2_0, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_0), .y(output_1_63));
wire output_3_63, output_3_0, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_0), .y(output_2_63));
wire output_4_63, output_4_0, output_3_63;
mixer gate_output_3_63(.a(output_4_63), .b(output_4_0), .y(output_3_63));
wire output_1_64, output_1_1, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_1), .y(output_0_64));
wire output_2_64, output_2_1, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_1), .y(output_1_64));
wire output_3_64, output_3_1, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_1), .y(output_2_64));
wire output_4_64, output_4_1, output_3_64;
mixer gate_output_3_64(.a(output_4_64), .b(output_4_1), .y(output_3_64));
wire output_1_65, output_1_2, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_2), .y(output_0_65));
wire output_2_65, output_2_2, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_2), .y(output_1_65));
wire output_3_65, output_3_2, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_2), .y(output_2_65));
wire output_4_65, output_4_2, output_3_65;
mixer gate_output_3_65(.a(output_4_65), .b(output_4_2), .y(output_3_65));
wire output_1_66, output_1_3, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_3), .y(output_0_66));
wire output_2_66, output_2_3, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_3), .y(output_1_66));
wire output_3_66, output_3_3, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_3), .y(output_2_66));
wire output_4_66, output_4_3, output_3_66;
mixer gate_output_3_66(.a(output_4_66), .b(output_4_3), .y(output_3_66));
wire output_1_67, output_1_0, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_0), .y(output_0_67));
wire output_2_67, output_2_0, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_0), .y(output_1_67));
wire output_3_67, output_3_0, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_0), .y(output_2_67));
wire output_4_67, output_4_0, output_3_67;
mixer gate_output_3_67(.a(output_4_67), .b(output_4_0), .y(output_3_67));
wire output_1_68, output_1_1, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_1), .y(output_0_68));
wire output_2_68, output_2_1, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_1), .y(output_1_68));
wire output_3_68, output_3_1, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_1), .y(output_2_68));
wire output_4_68, output_4_1, output_3_68;
mixer gate_output_3_68(.a(output_4_68), .b(output_4_1), .y(output_3_68));
wire output_1_69, output_1_2, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_2), .y(output_0_69));
wire output_2_69, output_2_2, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_2), .y(output_1_69));
wire output_3_69, output_3_2, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_2), .y(output_2_69));
wire output_4_69, output_4_2, output_3_69;
mixer gate_output_3_69(.a(output_4_69), .b(output_4_2), .y(output_3_69));
wire output_1_70, output_1_3, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_3), .y(output_0_70));
wire output_2_70, output_2_3, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_3), .y(output_1_70));
wire output_3_70, output_3_3, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_3), .y(output_2_70));
wire output_4_70, output_4_3, output_3_70;
mixer gate_output_3_70(.a(output_4_70), .b(output_4_3), .y(output_3_70));
wire output_1_71, output_1_0, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_0), .y(output_0_71));
wire output_2_71, output_2_0, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_0), .y(output_1_71));
wire output_3_71, output_3_0, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_0), .y(output_2_71));
wire output_4_71, output_4_0, output_3_71;
mixer gate_output_3_71(.a(output_4_71), .b(output_4_0), .y(output_3_71));
wire output_1_72, output_1_1, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_1), .y(output_0_72));
wire output_2_72, output_2_1, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_1), .y(output_1_72));
wire output_3_72, output_3_1, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_1), .y(output_2_72));
wire output_4_72, output_4_1, output_3_72;
mixer gate_output_3_72(.a(output_4_72), .b(output_4_1), .y(output_3_72));
wire output_1_73, output_1_2, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_2), .y(output_0_73));
wire output_2_73, output_2_2, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_2), .y(output_1_73));
wire output_3_73, output_3_2, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_2), .y(output_2_73));
wire output_4_73, output_4_2, output_3_73;
mixer gate_output_3_73(.a(output_4_73), .b(output_4_2), .y(output_3_73));
wire output_1_74, output_1_3, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_3), .y(output_0_74));
wire output_2_74, output_2_3, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_3), .y(output_1_74));
wire output_3_74, output_3_3, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_3), .y(output_2_74));
wire output_4_74, output_4_3, output_3_74;
mixer gate_output_3_74(.a(output_4_74), .b(output_4_3), .y(output_3_74));
wire output_1_75, output_1_0, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_0), .y(output_0_75));
wire output_2_75, output_2_0, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_0), .y(output_1_75));
wire output_3_75, output_3_0, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_0), .y(output_2_75));
wire output_4_75, output_4_0, output_3_75;
mixer gate_output_3_75(.a(output_4_75), .b(output_4_0), .y(output_3_75));
wire output_1_76, output_1_1, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_1), .y(output_0_76));
wire output_2_76, output_2_1, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_1), .y(output_1_76));
wire output_3_76, output_3_1, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_1), .y(output_2_76));
wire output_4_76, output_4_1, output_3_76;
mixer gate_output_3_76(.a(output_4_76), .b(output_4_1), .y(output_3_76));
wire output_1_77, output_1_2, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_2), .y(output_0_77));
wire output_2_77, output_2_2, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_2), .y(output_1_77));
wire output_3_77, output_3_2, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_2), .y(output_2_77));
wire output_4_77, output_4_2, output_3_77;
mixer gate_output_3_77(.a(output_4_77), .b(output_4_2), .y(output_3_77));
wire output_1_78, output_1_3, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_3), .y(output_0_78));
wire output_2_78, output_2_3, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_3), .y(output_1_78));
wire output_3_78, output_3_3, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_3), .y(output_2_78));
wire output_4_78, output_4_3, output_3_78;
mixer gate_output_3_78(.a(output_4_78), .b(output_4_3), .y(output_3_78));
wire output_1_79, output_1_0, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_0), .y(output_0_79));
wire output_2_79, output_2_0, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_0), .y(output_1_79));
wire output_3_79, output_3_0, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_0), .y(output_2_79));
wire output_4_79, output_4_0, output_3_79;
mixer gate_output_3_79(.a(output_4_79), .b(output_4_0), .y(output_3_79));
wire output_1_80, output_1_1, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_1), .y(output_0_80));
wire output_2_80, output_2_1, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_1), .y(output_1_80));
wire output_3_80, output_3_1, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_1), .y(output_2_80));
wire output_4_80, output_4_1, output_3_80;
mixer gate_output_3_80(.a(output_4_80), .b(output_4_1), .y(output_3_80));
wire output_1_81, output_1_2, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_2), .y(output_0_81));
wire output_2_81, output_2_2, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_2), .y(output_1_81));
wire output_3_81, output_3_2, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_2), .y(output_2_81));
wire output_4_81, output_4_2, output_3_81;
mixer gate_output_3_81(.a(output_4_81), .b(output_4_2), .y(output_3_81));
wire output_1_82, output_1_3, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_3), .y(output_0_82));
wire output_2_82, output_2_3, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_3), .y(output_1_82));
wire output_3_82, output_3_3, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_3), .y(output_2_82));
wire output_4_82, output_4_3, output_3_82;
mixer gate_output_3_82(.a(output_4_82), .b(output_4_3), .y(output_3_82));
wire output_1_83, output_1_0, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_0), .y(output_0_83));
wire output_2_83, output_2_0, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_0), .y(output_1_83));
wire output_3_83, output_3_0, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_0), .y(output_2_83));
wire output_4_83, output_4_0, output_3_83;
mixer gate_output_3_83(.a(output_4_83), .b(output_4_0), .y(output_3_83));
wire output_1_84, output_1_1, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_1), .y(output_0_84));
wire output_2_84, output_2_1, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_1), .y(output_1_84));
wire output_3_84, output_3_1, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_1), .y(output_2_84));
wire output_4_84, output_4_1, output_3_84;
mixer gate_output_3_84(.a(output_4_84), .b(output_4_1), .y(output_3_84));
wire output_1_85, output_1_2, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_2), .y(output_0_85));
wire output_2_85, output_2_2, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_2), .y(output_1_85));
wire output_3_85, output_3_2, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_2), .y(output_2_85));
wire output_4_85, output_4_2, output_3_85;
mixer gate_output_3_85(.a(output_4_85), .b(output_4_2), .y(output_3_85));
wire output_1_86, output_1_3, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_3), .y(output_0_86));
wire output_2_86, output_2_3, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_3), .y(output_1_86));
wire output_3_86, output_3_3, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_3), .y(output_2_86));
wire output_4_86, output_4_3, output_3_86;
mixer gate_output_3_86(.a(output_4_86), .b(output_4_3), .y(output_3_86));
wire output_1_87, output_1_0, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_0), .y(output_0_87));
wire output_2_87, output_2_0, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_0), .y(output_1_87));
wire output_3_87, output_3_0, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_0), .y(output_2_87));
wire output_4_87, output_4_0, output_3_87;
mixer gate_output_3_87(.a(output_4_87), .b(output_4_0), .y(output_3_87));
wire output_1_88, output_1_1, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_1), .y(output_0_88));
wire output_2_88, output_2_1, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_1), .y(output_1_88));
wire output_3_88, output_3_1, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_1), .y(output_2_88));
wire output_4_88, output_4_1, output_3_88;
mixer gate_output_3_88(.a(output_4_88), .b(output_4_1), .y(output_3_88));
wire output_1_89, output_1_2, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_2), .y(output_0_89));
wire output_2_89, output_2_2, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_2), .y(output_1_89));
wire output_3_89, output_3_2, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_2), .y(output_2_89));
wire output_4_89, output_4_2, output_3_89;
mixer gate_output_3_89(.a(output_4_89), .b(output_4_2), .y(output_3_89));
wire output_1_90, output_1_3, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_3), .y(output_0_90));
wire output_2_90, output_2_3, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_3), .y(output_1_90));
wire output_3_90, output_3_3, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_3), .y(output_2_90));
wire output_4_90, output_4_3, output_3_90;
mixer gate_output_3_90(.a(output_4_90), .b(output_4_3), .y(output_3_90));
wire output_1_91, output_1_0, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_0), .y(output_0_91));
wire output_2_91, output_2_0, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_0), .y(output_1_91));
wire output_3_91, output_3_0, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_0), .y(output_2_91));
wire output_4_91, output_4_0, output_3_91;
mixer gate_output_3_91(.a(output_4_91), .b(output_4_0), .y(output_3_91));
wire output_1_92, output_1_1, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_1), .y(output_0_92));
wire output_2_92, output_2_1, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_1), .y(output_1_92));
wire output_3_92, output_3_1, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_1), .y(output_2_92));
wire output_4_92, output_4_1, output_3_92;
mixer gate_output_3_92(.a(output_4_92), .b(output_4_1), .y(output_3_92));
wire output_1_93, output_1_2, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_2), .y(output_0_93));
wire output_2_93, output_2_2, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_2), .y(output_1_93));
wire output_3_93, output_3_2, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_2), .y(output_2_93));
wire output_4_93, output_4_2, output_3_93;
mixer gate_output_3_93(.a(output_4_93), .b(output_4_2), .y(output_3_93));
wire output_1_94, output_1_3, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_3), .y(output_0_94));
wire output_2_94, output_2_3, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_3), .y(output_1_94));
wire output_3_94, output_3_3, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_3), .y(output_2_94));
wire output_4_94, output_4_3, output_3_94;
mixer gate_output_3_94(.a(output_4_94), .b(output_4_3), .y(output_3_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_4_95, output_4_0, output_3_95;
mixer gate_output_3_95(.a(output_4_95), .b(output_4_0), .y(output_3_95));
wire output_1_96, output_1_1, output_0_96;
mixer gate_output_0_96(.a(output_1_96), .b(output_1_1), .y(output_0_96));
wire output_2_96, output_2_1, output_1_96;
mixer gate_output_1_96(.a(output_2_96), .b(output_2_1), .y(output_1_96));
wire output_3_96, output_3_1, output_2_96;
mixer gate_output_2_96(.a(output_3_96), .b(output_3_1), .y(output_2_96));
wire output_4_96, output_4_1, output_3_96;
mixer gate_output_3_96(.a(output_4_96), .b(output_4_1), .y(output_3_96));
wire output_1_97, output_1_2, output_0_97;
mixer gate_output_0_97(.a(output_1_97), .b(output_1_2), .y(output_0_97));
wire output_2_97, output_2_2, output_1_97;
mixer gate_output_1_97(.a(output_2_97), .b(output_2_2), .y(output_1_97));
wire output_3_97, output_3_2, output_2_97;
mixer gate_output_2_97(.a(output_3_97), .b(output_3_2), .y(output_2_97));
wire output_4_97, output_4_2, output_3_97;
mixer gate_output_3_97(.a(output_4_97), .b(output_4_2), .y(output_3_97));
wire output_1_98, output_1_3, output_0_98;
mixer gate_output_0_98(.a(output_1_98), .b(output_1_3), .y(output_0_98));
wire output_2_98, output_2_3, output_1_98;
mixer gate_output_1_98(.a(output_2_98), .b(output_2_3), .y(output_1_98));
wire output_3_98, output_3_3, output_2_98;
mixer gate_output_2_98(.a(output_3_98), .b(output_3_3), .y(output_2_98));
wire output_4_98, output_4_3, output_3_98;
mixer gate_output_3_98(.a(output_4_98), .b(output_4_3), .y(output_3_98));
wire output_1_99, output_1_0, output_0_99;
mixer gate_output_0_99(.a(output_1_99), .b(output_1_0), .y(output_0_99));
wire output_2_99, output_2_0, output_1_99;
mixer gate_output_1_99(.a(output_2_99), .b(output_2_0), .y(output_1_99));
wire output_3_99, output_3_0, output_2_99;
mixer gate_output_2_99(.a(output_3_99), .b(output_3_0), .y(output_2_99));
wire output_4_99, output_4_0, output_3_99;
mixer gate_output_3_99(.a(output_4_99), .b(output_4_0), .y(output_3_99));
wire output_1_100, output_1_1, output_0_100;
mixer gate_output_0_100(.a(output_1_100), .b(output_1_1), .y(output_0_100));
wire output_2_100, output_2_1, output_1_100;
mixer gate_output_1_100(.a(output_2_100), .b(output_2_1), .y(output_1_100));
wire output_3_100, output_3_1, output_2_100;
mixer gate_output_2_100(.a(output_3_100), .b(output_3_1), .y(output_2_100));
wire output_4_100, output_4_1, output_3_100;
mixer gate_output_3_100(.a(output_4_100), .b(output_4_1), .y(output_3_100));
wire output_1_101, output_1_2, output_0_101;
mixer gate_output_0_101(.a(output_1_101), .b(output_1_2), .y(output_0_101));
wire output_2_101, output_2_2, output_1_101;
mixer gate_output_1_101(.a(output_2_101), .b(output_2_2), .y(output_1_101));
wire output_3_101, output_3_2, output_2_101;
mixer gate_output_2_101(.a(output_3_101), .b(output_3_2), .y(output_2_101));
wire output_4_101, output_4_2, output_3_101;
mixer gate_output_3_101(.a(output_4_101), .b(output_4_2), .y(output_3_101));
wire output_1_102, output_1_3, output_0_102;
mixer gate_output_0_102(.a(output_1_102), .b(output_1_3), .y(output_0_102));
wire output_2_102, output_2_3, output_1_102;
mixer gate_output_1_102(.a(output_2_102), .b(output_2_3), .y(output_1_102));
wire output_3_102, output_3_3, output_2_102;
mixer gate_output_2_102(.a(output_3_102), .b(output_3_3), .y(output_2_102));
wire output_4_102, output_4_3, output_3_102;
mixer gate_output_3_102(.a(output_4_102), .b(output_4_3), .y(output_3_102));
wire output_1_103, output_1_0, output_0_103;
mixer gate_output_0_103(.a(output_1_103), .b(output_1_0), .y(output_0_103));
wire output_2_103, output_2_0, output_1_103;
mixer gate_output_1_103(.a(output_2_103), .b(output_2_0), .y(output_1_103));
wire output_3_103, output_3_0, output_2_103;
mixer gate_output_2_103(.a(output_3_103), .b(output_3_0), .y(output_2_103));
wire output_4_103, output_4_0, output_3_103;
mixer gate_output_3_103(.a(output_4_103), .b(output_4_0), .y(output_3_103));
wire output_1_104, output_1_1, output_0_104;
mixer gate_output_0_104(.a(output_1_104), .b(output_1_1), .y(output_0_104));
wire output_2_104, output_2_1, output_1_104;
mixer gate_output_1_104(.a(output_2_104), .b(output_2_1), .y(output_1_104));
wire output_3_104, output_3_1, output_2_104;
mixer gate_output_2_104(.a(output_3_104), .b(output_3_1), .y(output_2_104));
wire output_4_104, output_4_1, output_3_104;
mixer gate_output_3_104(.a(output_4_104), .b(output_4_1), .y(output_3_104));
wire output_1_105, output_1_2, output_0_105;
mixer gate_output_0_105(.a(output_1_105), .b(output_1_2), .y(output_0_105));
wire output_2_105, output_2_2, output_1_105;
mixer gate_output_1_105(.a(output_2_105), .b(output_2_2), .y(output_1_105));
wire output_3_105, output_3_2, output_2_105;
mixer gate_output_2_105(.a(output_3_105), .b(output_3_2), .y(output_2_105));
wire output_4_105, output_4_2, output_3_105;
mixer gate_output_3_105(.a(output_4_105), .b(output_4_2), .y(output_3_105));
wire output_1_106, output_1_3, output_0_106;
mixer gate_output_0_106(.a(output_1_106), .b(output_1_3), .y(output_0_106));
wire output_2_106, output_2_3, output_1_106;
mixer gate_output_1_106(.a(output_2_106), .b(output_2_3), .y(output_1_106));
wire output_3_106, output_3_3, output_2_106;
mixer gate_output_2_106(.a(output_3_106), .b(output_3_3), .y(output_2_106));
wire output_4_106, output_4_3, output_3_106;
mixer gate_output_3_106(.a(output_4_106), .b(output_4_3), .y(output_3_106));
wire output_1_107, output_1_0, output_0_107;
mixer gate_output_0_107(.a(output_1_107), .b(output_1_0), .y(output_0_107));
wire output_2_107, output_2_0, output_1_107;
mixer gate_output_1_107(.a(output_2_107), .b(output_2_0), .y(output_1_107));
wire output_3_107, output_3_0, output_2_107;
mixer gate_output_2_107(.a(output_3_107), .b(output_3_0), .y(output_2_107));
wire output_4_107, output_4_0, output_3_107;
mixer gate_output_3_107(.a(output_4_107), .b(output_4_0), .y(output_3_107));
wire output_1_108, output_1_1, output_0_108;
mixer gate_output_0_108(.a(output_1_108), .b(output_1_1), .y(output_0_108));
wire output_2_108, output_2_1, output_1_108;
mixer gate_output_1_108(.a(output_2_108), .b(output_2_1), .y(output_1_108));
wire output_3_108, output_3_1, output_2_108;
mixer gate_output_2_108(.a(output_3_108), .b(output_3_1), .y(output_2_108));
wire output_4_108, output_4_1, output_3_108;
mixer gate_output_3_108(.a(output_4_108), .b(output_4_1), .y(output_3_108));
wire output_1_109, output_1_2, output_0_109;
mixer gate_output_0_109(.a(output_1_109), .b(output_1_2), .y(output_0_109));
wire output_2_109, output_2_2, output_1_109;
mixer gate_output_1_109(.a(output_2_109), .b(output_2_2), .y(output_1_109));
wire output_3_109, output_3_2, output_2_109;
mixer gate_output_2_109(.a(output_3_109), .b(output_3_2), .y(output_2_109));
wire output_4_109, output_4_2, output_3_109;
mixer gate_output_3_109(.a(output_4_109), .b(output_4_2), .y(output_3_109));
wire output_1_110, output_1_3, output_0_110;
mixer gate_output_0_110(.a(output_1_110), .b(output_1_3), .y(output_0_110));
wire output_2_110, output_2_3, output_1_110;
mixer gate_output_1_110(.a(output_2_110), .b(output_2_3), .y(output_1_110));
wire output_3_110, output_3_3, output_2_110;
mixer gate_output_2_110(.a(output_3_110), .b(output_3_3), .y(output_2_110));
wire output_4_110, output_4_3, output_3_110;
mixer gate_output_3_110(.a(output_4_110), .b(output_4_3), .y(output_3_110));
wire output_1_111, output_1_0, output_0_111;
mixer gate_output_0_111(.a(output_1_111), .b(output_1_0), .y(output_0_111));
wire output_2_111, output_2_0, output_1_111;
mixer gate_output_1_111(.a(output_2_111), .b(output_2_0), .y(output_1_111));
wire output_3_111, output_3_0, output_2_111;
mixer gate_output_2_111(.a(output_3_111), .b(output_3_0), .y(output_2_111));
wire output_4_111, output_4_0, output_3_111;
mixer gate_output_3_111(.a(output_4_111), .b(output_4_0), .y(output_3_111));
wire output_1_112, output_1_1, output_0_112;
mixer gate_output_0_112(.a(output_1_112), .b(output_1_1), .y(output_0_112));
wire output_2_112, output_2_1, output_1_112;
mixer gate_output_1_112(.a(output_2_112), .b(output_2_1), .y(output_1_112));
wire output_3_112, output_3_1, output_2_112;
mixer gate_output_2_112(.a(output_3_112), .b(output_3_1), .y(output_2_112));
wire output_4_112, output_4_1, output_3_112;
mixer gate_output_3_112(.a(output_4_112), .b(output_4_1), .y(output_3_112));
wire output_1_113, output_1_2, output_0_113;
mixer gate_output_0_113(.a(output_1_113), .b(output_1_2), .y(output_0_113));
wire output_2_113, output_2_2, output_1_113;
mixer gate_output_1_113(.a(output_2_113), .b(output_2_2), .y(output_1_113));
wire output_3_113, output_3_2, output_2_113;
mixer gate_output_2_113(.a(output_3_113), .b(output_3_2), .y(output_2_113));
wire output_4_113, output_4_2, output_3_113;
mixer gate_output_3_113(.a(output_4_113), .b(output_4_2), .y(output_3_113));
wire output_1_114, output_1_3, output_0_114;
mixer gate_output_0_114(.a(output_1_114), .b(output_1_3), .y(output_0_114));
wire output_2_114, output_2_3, output_1_114;
mixer gate_output_1_114(.a(output_2_114), .b(output_2_3), .y(output_1_114));
wire output_3_114, output_3_3, output_2_114;
mixer gate_output_2_114(.a(output_3_114), .b(output_3_3), .y(output_2_114));
wire output_4_114, output_4_3, output_3_114;
mixer gate_output_3_114(.a(output_4_114), .b(output_4_3), .y(output_3_114));
wire output_1_115, output_1_0, output_0_115;
mixer gate_output_0_115(.a(output_1_115), .b(output_1_0), .y(output_0_115));
wire output_2_115, output_2_0, output_1_115;
mixer gate_output_1_115(.a(output_2_115), .b(output_2_0), .y(output_1_115));
wire output_3_115, output_3_0, output_2_115;
mixer gate_output_2_115(.a(output_3_115), .b(output_3_0), .y(output_2_115));
wire output_4_115, output_4_0, output_3_115;
mixer gate_output_3_115(.a(output_4_115), .b(output_4_0), .y(output_3_115));
wire output_1_116, output_1_1, output_0_116;
mixer gate_output_0_116(.a(output_1_116), .b(output_1_1), .y(output_0_116));
wire output_2_116, output_2_1, output_1_116;
mixer gate_output_1_116(.a(output_2_116), .b(output_2_1), .y(output_1_116));
wire output_3_116, output_3_1, output_2_116;
mixer gate_output_2_116(.a(output_3_116), .b(output_3_1), .y(output_2_116));
wire output_4_116, output_4_1, output_3_116;
mixer gate_output_3_116(.a(output_4_116), .b(output_4_1), .y(output_3_116));
wire output_1_117, output_1_2, output_0_117;
mixer gate_output_0_117(.a(output_1_117), .b(output_1_2), .y(output_0_117));
wire output_2_117, output_2_2, output_1_117;
mixer gate_output_1_117(.a(output_2_117), .b(output_2_2), .y(output_1_117));
wire output_3_117, output_3_2, output_2_117;
mixer gate_output_2_117(.a(output_3_117), .b(output_3_2), .y(output_2_117));
wire output_4_117, output_4_2, output_3_117;
mixer gate_output_3_117(.a(output_4_117), .b(output_4_2), .y(output_3_117));
wire output_1_118, output_1_3, output_0_118;
mixer gate_output_0_118(.a(output_1_118), .b(output_1_3), .y(output_0_118));
wire output_2_118, output_2_3, output_1_118;
mixer gate_output_1_118(.a(output_2_118), .b(output_2_3), .y(output_1_118));
wire output_3_118, output_3_3, output_2_118;
mixer gate_output_2_118(.a(output_3_118), .b(output_3_3), .y(output_2_118));
wire output_4_118, output_4_3, output_3_118;
mixer gate_output_3_118(.a(output_4_118), .b(output_4_3), .y(output_3_118));
wire output_1_119, output_1_0, output_0_119;
mixer gate_output_0_119(.a(output_1_119), .b(output_1_0), .y(output_0_119));
wire output_2_119, output_2_0, output_1_119;
mixer gate_output_1_119(.a(output_2_119), .b(output_2_0), .y(output_1_119));
wire output_3_119, output_3_0, output_2_119;
mixer gate_output_2_119(.a(output_3_119), .b(output_3_0), .y(output_2_119));
wire output_4_119, output_4_0, output_3_119;
mixer gate_output_3_119(.a(output_4_119), .b(output_4_0), .y(output_3_119));
wire output_1_120, output_1_1, output_0_120;
mixer gate_output_0_120(.a(output_1_120), .b(output_1_1), .y(output_0_120));
wire output_2_120, output_2_1, output_1_120;
mixer gate_output_1_120(.a(output_2_120), .b(output_2_1), .y(output_1_120));
wire output_3_120, output_3_1, output_2_120;
mixer gate_output_2_120(.a(output_3_120), .b(output_3_1), .y(output_2_120));
wire output_4_120, output_4_1, output_3_120;
mixer gate_output_3_120(.a(output_4_120), .b(output_4_1), .y(output_3_120));
wire output_1_121, output_1_2, output_0_121;
mixer gate_output_0_121(.a(output_1_121), .b(output_1_2), .y(output_0_121));
wire output_2_121, output_2_2, output_1_121;
mixer gate_output_1_121(.a(output_2_121), .b(output_2_2), .y(output_1_121));
wire output_3_121, output_3_2, output_2_121;
mixer gate_output_2_121(.a(output_3_121), .b(output_3_2), .y(output_2_121));
wire output_4_121, output_4_2, output_3_121;
mixer gate_output_3_121(.a(output_4_121), .b(output_4_2), .y(output_3_121));
wire output_1_122, output_1_3, output_0_122;
mixer gate_output_0_122(.a(output_1_122), .b(output_1_3), .y(output_0_122));
wire output_2_122, output_2_3, output_1_122;
mixer gate_output_1_122(.a(output_2_122), .b(output_2_3), .y(output_1_122));
wire output_3_122, output_3_3, output_2_122;
mixer gate_output_2_122(.a(output_3_122), .b(output_3_3), .y(output_2_122));
wire output_4_122, output_4_3, output_3_122;
mixer gate_output_3_122(.a(output_4_122), .b(output_4_3), .y(output_3_122));
wire output_1_123, output_1_0, output_0_123;
mixer gate_output_0_123(.a(output_1_123), .b(output_1_0), .y(output_0_123));
wire output_2_123, output_2_0, output_1_123;
mixer gate_output_1_123(.a(output_2_123), .b(output_2_0), .y(output_1_123));
wire output_3_123, output_3_0, output_2_123;
mixer gate_output_2_123(.a(output_3_123), .b(output_3_0), .y(output_2_123));
wire output_4_123, output_4_0, output_3_123;
mixer gate_output_3_123(.a(output_4_123), .b(output_4_0), .y(output_3_123));
wire output_1_124, output_1_1, output_0_124;
mixer gate_output_0_124(.a(output_1_124), .b(output_1_1), .y(output_0_124));
wire output_2_124, output_2_1, output_1_124;
mixer gate_output_1_124(.a(output_2_124), .b(output_2_1), .y(output_1_124));
wire output_3_124, output_3_1, output_2_124;
mixer gate_output_2_124(.a(output_3_124), .b(output_3_1), .y(output_2_124));
wire output_4_124, output_4_1, output_3_124;
mixer gate_output_3_124(.a(output_4_124), .b(output_4_1), .y(output_3_124));
wire output_1_125, output_1_2, output_0_125;
mixer gate_output_0_125(.a(output_1_125), .b(output_1_2), .y(output_0_125));
wire output_2_125, output_2_2, output_1_125;
mixer gate_output_1_125(.a(output_2_125), .b(output_2_2), .y(output_1_125));
wire output_3_125, output_3_2, output_2_125;
mixer gate_output_2_125(.a(output_3_125), .b(output_3_2), .y(output_2_125));
wire output_4_125, output_4_2, output_3_125;
mixer gate_output_3_125(.a(output_4_125), .b(output_4_2), .y(output_3_125));
wire output_1_126, output_1_3, output_0_126;
mixer gate_output_0_126(.a(output_1_126), .b(output_1_3), .y(output_0_126));
wire output_2_126, output_2_3, output_1_126;
mixer gate_output_1_126(.a(output_2_126), .b(output_2_3), .y(output_1_126));
wire output_3_126, output_3_3, output_2_126;
mixer gate_output_2_126(.a(output_3_126), .b(output_3_3), .y(output_2_126));
wire output_4_126, output_4_3, output_3_126;
mixer gate_output_3_126(.a(output_4_126), .b(output_4_3), .y(output_3_126));
wire output_1_127, output_1_0, output_0_127;
mixer gate_output_0_127(.a(output_1_127), .b(output_1_0), .y(output_0_127));
wire output_2_127, output_2_0, output_1_127;
mixer gate_output_1_127(.a(output_2_127), .b(output_2_0), .y(output_1_127));
wire output_3_127, output_3_0, output_2_127;
mixer gate_output_2_127(.a(output_3_127), .b(output_3_0), .y(output_2_127));
wire output_4_127, output_4_0, output_3_127;
mixer gate_output_3_127(.a(output_4_127), .b(output_4_0), .y(output_3_127));
wire output_1_128, output_1_1, output_0_128;
mixer gate_output_0_128(.a(output_1_128), .b(output_1_1), .y(output_0_128));
wire output_2_128, output_2_1, output_1_128;
mixer gate_output_1_128(.a(output_2_128), .b(output_2_1), .y(output_1_128));
wire output_3_128, output_3_1, output_2_128;
mixer gate_output_2_128(.a(output_3_128), .b(output_3_1), .y(output_2_128));
wire output_4_128, output_4_1, output_3_128;
mixer gate_output_3_128(.a(output_4_128), .b(output_4_1), .y(output_3_128));
wire output_1_129, output_1_2, output_0_129;
mixer gate_output_0_129(.a(output_1_129), .b(output_1_2), .y(output_0_129));
wire output_2_129, output_2_2, output_1_129;
mixer gate_output_1_129(.a(output_2_129), .b(output_2_2), .y(output_1_129));
wire output_3_129, output_3_2, output_2_129;
mixer gate_output_2_129(.a(output_3_129), .b(output_3_2), .y(output_2_129));
wire output_4_129, output_4_2, output_3_129;
mixer gate_output_3_129(.a(output_4_129), .b(output_4_2), .y(output_3_129));
wire output_1_130, output_1_3, output_0_130;
mixer gate_output_0_130(.a(output_1_130), .b(output_1_3), .y(output_0_130));
wire output_2_130, output_2_3, output_1_130;
mixer gate_output_1_130(.a(output_2_130), .b(output_2_3), .y(output_1_130));
wire output_3_130, output_3_3, output_2_130;
mixer gate_output_2_130(.a(output_3_130), .b(output_3_3), .y(output_2_130));
wire output_4_130, output_4_3, output_3_130;
mixer gate_output_3_130(.a(output_4_130), .b(output_4_3), .y(output_3_130));
wire output_1_131, output_1_0, output_0_131;
mixer gate_output_0_131(.a(output_1_131), .b(output_1_0), .y(output_0_131));
wire output_2_131, output_2_0, output_1_131;
mixer gate_output_1_131(.a(output_2_131), .b(output_2_0), .y(output_1_131));
wire output_3_131, output_3_0, output_2_131;
mixer gate_output_2_131(.a(output_3_131), .b(output_3_0), .y(output_2_131));
wire output_4_131, output_4_0, output_3_131;
mixer gate_output_3_131(.a(output_4_131), .b(output_4_0), .y(output_3_131));
wire output_1_132, output_1_1, output_0_132;
mixer gate_output_0_132(.a(output_1_132), .b(output_1_1), .y(output_0_132));
wire output_2_132, output_2_1, output_1_132;
mixer gate_output_1_132(.a(output_2_132), .b(output_2_1), .y(output_1_132));
wire output_3_132, output_3_1, output_2_132;
mixer gate_output_2_132(.a(output_3_132), .b(output_3_1), .y(output_2_132));
wire output_4_132, output_4_1, output_3_132;
mixer gate_output_3_132(.a(output_4_132), .b(output_4_1), .y(output_3_132));
wire output_1_133, output_1_2, output_0_133;
mixer gate_output_0_133(.a(output_1_133), .b(output_1_2), .y(output_0_133));
wire output_2_133, output_2_2, output_1_133;
mixer gate_output_1_133(.a(output_2_133), .b(output_2_2), .y(output_1_133));
wire output_3_133, output_3_2, output_2_133;
mixer gate_output_2_133(.a(output_3_133), .b(output_3_2), .y(output_2_133));
wire output_4_133, output_4_2, output_3_133;
mixer gate_output_3_133(.a(output_4_133), .b(output_4_2), .y(output_3_133));
wire output_1_134, output_1_3, output_0_134;
mixer gate_output_0_134(.a(output_1_134), .b(output_1_3), .y(output_0_134));
wire output_2_134, output_2_3, output_1_134;
mixer gate_output_1_134(.a(output_2_134), .b(output_2_3), .y(output_1_134));
wire output_3_134, output_3_3, output_2_134;
mixer gate_output_2_134(.a(output_3_134), .b(output_3_3), .y(output_2_134));
wire output_4_134, output_4_3, output_3_134;
mixer gate_output_3_134(.a(output_4_134), .b(output_4_3), .y(output_3_134));
wire output_1_135, output_1_0, output_0_135;
mixer gate_output_0_135(.a(output_1_135), .b(output_1_0), .y(output_0_135));
wire output_2_135, output_2_0, output_1_135;
mixer gate_output_1_135(.a(output_2_135), .b(output_2_0), .y(output_1_135));
wire output_3_135, output_3_0, output_2_135;
mixer gate_output_2_135(.a(output_3_135), .b(output_3_0), .y(output_2_135));
wire output_4_135, output_4_0, output_3_135;
mixer gate_output_3_135(.a(output_4_135), .b(output_4_0), .y(output_3_135));
wire output_1_136, output_1_1, output_0_136;
mixer gate_output_0_136(.a(output_1_136), .b(output_1_1), .y(output_0_136));
wire output_2_136, output_2_1, output_1_136;
mixer gate_output_1_136(.a(output_2_136), .b(output_2_1), .y(output_1_136));
wire output_3_136, output_3_1, output_2_136;
mixer gate_output_2_136(.a(output_3_136), .b(output_3_1), .y(output_2_136));
wire output_4_136, output_4_1, output_3_136;
mixer gate_output_3_136(.a(output_4_136), .b(output_4_1), .y(output_3_136));
wire output_1_137, output_1_2, output_0_137;
mixer gate_output_0_137(.a(output_1_137), .b(output_1_2), .y(output_0_137));
wire output_2_137, output_2_2, output_1_137;
mixer gate_output_1_137(.a(output_2_137), .b(output_2_2), .y(output_1_137));
wire output_3_137, output_3_2, output_2_137;
mixer gate_output_2_137(.a(output_3_137), .b(output_3_2), .y(output_2_137));
wire output_4_137, output_4_2, output_3_137;
mixer gate_output_3_137(.a(output_4_137), .b(output_4_2), .y(output_3_137));
wire output_1_138, output_1_3, output_0_138;
mixer gate_output_0_138(.a(output_1_138), .b(output_1_3), .y(output_0_138));
wire output_2_138, output_2_3, output_1_138;
mixer gate_output_1_138(.a(output_2_138), .b(output_2_3), .y(output_1_138));
wire output_3_138, output_3_3, output_2_138;
mixer gate_output_2_138(.a(output_3_138), .b(output_3_3), .y(output_2_138));
wire output_4_138, output_4_3, output_3_138;
mixer gate_output_3_138(.a(output_4_138), .b(output_4_3), .y(output_3_138));
wire output_1_139, output_1_0, output_0_139;
mixer gate_output_0_139(.a(output_1_139), .b(output_1_0), .y(output_0_139));
wire output_2_139, output_2_0, output_1_139;
mixer gate_output_1_139(.a(output_2_139), .b(output_2_0), .y(output_1_139));
wire output_3_139, output_3_0, output_2_139;
mixer gate_output_2_139(.a(output_3_139), .b(output_3_0), .y(output_2_139));
wire output_4_139, output_4_0, output_3_139;
mixer gate_output_3_139(.a(output_4_139), .b(output_4_0), .y(output_3_139));
wire output_1_140, output_1_1, output_0_140;
mixer gate_output_0_140(.a(output_1_140), .b(output_1_1), .y(output_0_140));
wire output_2_140, output_2_1, output_1_140;
mixer gate_output_1_140(.a(output_2_140), .b(output_2_1), .y(output_1_140));
wire output_3_140, output_3_1, output_2_140;
mixer gate_output_2_140(.a(output_3_140), .b(output_3_1), .y(output_2_140));
wire output_4_140, output_4_1, output_3_140;
mixer gate_output_3_140(.a(output_4_140), .b(output_4_1), .y(output_3_140));
wire output_1_141, output_1_2, output_0_141;
mixer gate_output_0_141(.a(output_1_141), .b(output_1_2), .y(output_0_141));
wire output_2_141, output_2_2, output_1_141;
mixer gate_output_1_141(.a(output_2_141), .b(output_2_2), .y(output_1_141));
wire output_3_141, output_3_2, output_2_141;
mixer gate_output_2_141(.a(output_3_141), .b(output_3_2), .y(output_2_141));
wire output_4_141, output_4_2, output_3_141;
mixer gate_output_3_141(.a(output_4_141), .b(output_4_2), .y(output_3_141));
wire output_1_142, output_1_3, output_0_142;
mixer gate_output_0_142(.a(output_1_142), .b(output_1_3), .y(output_0_142));
wire output_2_142, output_2_3, output_1_142;
mixer gate_output_1_142(.a(output_2_142), .b(output_2_3), .y(output_1_142));
wire output_3_142, output_3_3, output_2_142;
mixer gate_output_2_142(.a(output_3_142), .b(output_3_3), .y(output_2_142));
wire output_4_142, output_4_3, output_3_142;
mixer gate_output_3_142(.a(output_4_142), .b(output_4_3), .y(output_3_142));
wire output_1_143, output_1_0, output_0_143;
mixer gate_output_0_143(.a(output_1_143), .b(output_1_0), .y(output_0_143));
wire output_2_143, output_2_0, output_1_143;
mixer gate_output_1_143(.a(output_2_143), .b(output_2_0), .y(output_1_143));
wire output_3_143, output_3_0, output_2_143;
mixer gate_output_2_143(.a(output_3_143), .b(output_3_0), .y(output_2_143));
wire output_4_143, output_4_0, output_3_143;
mixer gate_output_3_143(.a(output_4_143), .b(output_4_0), .y(output_3_143));
wire output_1_144, output_1_1, output_0_144;
mixer gate_output_0_144(.a(output_1_144), .b(output_1_1), .y(output_0_144));
wire output_2_144, output_2_1, output_1_144;
mixer gate_output_1_144(.a(output_2_144), .b(output_2_1), .y(output_1_144));
wire output_3_144, output_3_1, output_2_144;
mixer gate_output_2_144(.a(output_3_144), .b(output_3_1), .y(output_2_144));
wire output_4_144, output_4_1, output_3_144;
mixer gate_output_3_144(.a(output_4_144), .b(output_4_1), .y(output_3_144));
wire output_1_145, output_1_2, output_0_145;
mixer gate_output_0_145(.a(output_1_145), .b(output_1_2), .y(output_0_145));
wire output_2_145, output_2_2, output_1_145;
mixer gate_output_1_145(.a(output_2_145), .b(output_2_2), .y(output_1_145));
wire output_3_145, output_3_2, output_2_145;
mixer gate_output_2_145(.a(output_3_145), .b(output_3_2), .y(output_2_145));
wire output_4_145, output_4_2, output_3_145;
mixer gate_output_3_145(.a(output_4_145), .b(output_4_2), .y(output_3_145));
wire output_1_146, output_1_3, output_0_146;
mixer gate_output_0_146(.a(output_1_146), .b(output_1_3), .y(output_0_146));
wire output_2_146, output_2_3, output_1_146;
mixer gate_output_1_146(.a(output_2_146), .b(output_2_3), .y(output_1_146));
wire output_3_146, output_3_3, output_2_146;
mixer gate_output_2_146(.a(output_3_146), .b(output_3_3), .y(output_2_146));
wire output_4_146, output_4_3, output_3_146;
mixer gate_output_3_146(.a(output_4_146), .b(output_4_3), .y(output_3_146));
wire output_1_147, output_1_0, output_0_147;
mixer gate_output_0_147(.a(output_1_147), .b(output_1_0), .y(output_0_147));
wire output_2_147, output_2_0, output_1_147;
mixer gate_output_1_147(.a(output_2_147), .b(output_2_0), .y(output_1_147));
wire output_3_147, output_3_0, output_2_147;
mixer gate_output_2_147(.a(output_3_147), .b(output_3_0), .y(output_2_147));
wire output_4_147, output_4_0, output_3_147;
mixer gate_output_3_147(.a(output_4_147), .b(output_4_0), .y(output_3_147));
wire output_1_148, output_1_1, output_0_148;
mixer gate_output_0_148(.a(output_1_148), .b(output_1_1), .y(output_0_148));
wire output_2_148, output_2_1, output_1_148;
mixer gate_output_1_148(.a(output_2_148), .b(output_2_1), .y(output_1_148));
wire output_3_148, output_3_1, output_2_148;
mixer gate_output_2_148(.a(output_3_148), .b(output_3_1), .y(output_2_148));
wire output_4_148, output_4_1, output_3_148;
mixer gate_output_3_148(.a(output_4_148), .b(output_4_1), .y(output_3_148));
wire output_1_149, output_1_2, output_0_149;
mixer gate_output_0_149(.a(output_1_149), .b(output_1_2), .y(output_0_149));
wire output_2_149, output_2_2, output_1_149;
mixer gate_output_1_149(.a(output_2_149), .b(output_2_2), .y(output_1_149));
wire output_3_149, output_3_2, output_2_149;
mixer gate_output_2_149(.a(output_3_149), .b(output_3_2), .y(output_2_149));
wire output_4_149, output_4_2, output_3_149;
mixer gate_output_3_149(.a(output_4_149), .b(output_4_2), .y(output_3_149));
wire output_1_150, output_1_3, output_0_150;
mixer gate_output_0_150(.a(output_1_150), .b(output_1_3), .y(output_0_150));
wire output_2_150, output_2_3, output_1_150;
mixer gate_output_1_150(.a(output_2_150), .b(output_2_3), .y(output_1_150));
wire output_3_150, output_3_3, output_2_150;
mixer gate_output_2_150(.a(output_3_150), .b(output_3_3), .y(output_2_150));
wire output_4_150, output_4_3, output_3_150;
mixer gate_output_3_150(.a(output_4_150), .b(output_4_3), .y(output_3_150));
wire output_1_151, output_1_0, output_0_151;
mixer gate_output_0_151(.a(output_1_151), .b(output_1_0), .y(output_0_151));
wire output_2_151, output_2_0, output_1_151;
mixer gate_output_1_151(.a(output_2_151), .b(output_2_0), .y(output_1_151));
wire output_3_151, output_3_0, output_2_151;
mixer gate_output_2_151(.a(output_3_151), .b(output_3_0), .y(output_2_151));
wire output_4_151, output_4_0, output_3_151;
mixer gate_output_3_151(.a(output_4_151), .b(output_4_0), .y(output_3_151));
wire output_1_152, output_1_1, output_0_152;
mixer gate_output_0_152(.a(output_1_152), .b(output_1_1), .y(output_0_152));
wire output_2_152, output_2_1, output_1_152;
mixer gate_output_1_152(.a(output_2_152), .b(output_2_1), .y(output_1_152));
wire output_3_152, output_3_1, output_2_152;
mixer gate_output_2_152(.a(output_3_152), .b(output_3_1), .y(output_2_152));
wire output_4_152, output_4_1, output_3_152;
mixer gate_output_3_152(.a(output_4_152), .b(output_4_1), .y(output_3_152));
wire output_1_153, output_1_2, output_0_153;
mixer gate_output_0_153(.a(output_1_153), .b(output_1_2), .y(output_0_153));
wire output_2_153, output_2_2, output_1_153;
mixer gate_output_1_153(.a(output_2_153), .b(output_2_2), .y(output_1_153));
wire output_3_153, output_3_2, output_2_153;
mixer gate_output_2_153(.a(output_3_153), .b(output_3_2), .y(output_2_153));
wire output_4_153, output_4_2, output_3_153;
mixer gate_output_3_153(.a(output_4_153), .b(output_4_2), .y(output_3_153));
wire output_1_154, output_1_3, output_0_154;
mixer gate_output_0_154(.a(output_1_154), .b(output_1_3), .y(output_0_154));
wire output_2_154, output_2_3, output_1_154;
mixer gate_output_1_154(.a(output_2_154), .b(output_2_3), .y(output_1_154));
wire output_3_154, output_3_3, output_2_154;
mixer gate_output_2_154(.a(output_3_154), .b(output_3_3), .y(output_2_154));
wire output_4_154, output_4_3, output_3_154;
mixer gate_output_3_154(.a(output_4_154), .b(output_4_3), .y(output_3_154));
wire output_1_155, output_1_0, output_0_155;
mixer gate_output_0_155(.a(output_1_155), .b(output_1_0), .y(output_0_155));
wire output_2_155, output_2_0, output_1_155;
mixer gate_output_1_155(.a(output_2_155), .b(output_2_0), .y(output_1_155));
wire output_3_155, output_3_0, output_2_155;
mixer gate_output_2_155(.a(output_3_155), .b(output_3_0), .y(output_2_155));
wire output_4_155, output_4_0, output_3_155;
mixer gate_output_3_155(.a(output_4_155), .b(output_4_0), .y(output_3_155));
wire output_1_156, output_1_1, output_0_156;
mixer gate_output_0_156(.a(output_1_156), .b(output_1_1), .y(output_0_156));
wire output_2_156, output_2_1, output_1_156;
mixer gate_output_1_156(.a(output_2_156), .b(output_2_1), .y(output_1_156));
wire output_3_156, output_3_1, output_2_156;
mixer gate_output_2_156(.a(output_3_156), .b(output_3_1), .y(output_2_156));
wire output_4_156, output_4_1, output_3_156;
mixer gate_output_3_156(.a(output_4_156), .b(output_4_1), .y(output_3_156));
wire output_1_157, output_1_2, output_0_157;
mixer gate_output_0_157(.a(output_1_157), .b(output_1_2), .y(output_0_157));
wire output_2_157, output_2_2, output_1_157;
mixer gate_output_1_157(.a(output_2_157), .b(output_2_2), .y(output_1_157));
wire output_3_157, output_3_2, output_2_157;
mixer gate_output_2_157(.a(output_3_157), .b(output_3_2), .y(output_2_157));
wire output_4_157, output_4_2, output_3_157;
mixer gate_output_3_157(.a(output_4_157), .b(output_4_2), .y(output_3_157));
wire output_1_158, output_1_3, output_0_158;
mixer gate_output_0_158(.a(output_1_158), .b(output_1_3), .y(output_0_158));
wire output_2_158, output_2_3, output_1_158;
mixer gate_output_1_158(.a(output_2_158), .b(output_2_3), .y(output_1_158));
wire output_3_158, output_3_3, output_2_158;
mixer gate_output_2_158(.a(output_3_158), .b(output_3_3), .y(output_2_158));
wire output_4_158, output_4_3, output_3_158;
mixer gate_output_3_158(.a(output_4_158), .b(output_4_3), .y(output_3_158));
wire output_1_159, output_1_0, output_0_159;
mixer gate_output_0_159(.a(output_1_159), .b(output_1_0), .y(output_0_159));
wire output_2_159, output_2_0, output_1_159;
mixer gate_output_1_159(.a(output_2_159), .b(output_2_0), .y(output_1_159));
wire output_3_159, output_3_0, output_2_159;
mixer gate_output_2_159(.a(output_3_159), .b(output_3_0), .y(output_2_159));
wire output_4_159, output_4_0, output_3_159;
mixer gate_output_3_159(.a(output_4_159), .b(output_4_0), .y(output_3_159));
wire output_1_160, output_1_1, output_0_160;
mixer gate_output_0_160(.a(output_1_160), .b(output_1_1), .y(output_0_160));
wire output_2_160, output_2_1, output_1_160;
mixer gate_output_1_160(.a(output_2_160), .b(output_2_1), .y(output_1_160));
wire output_3_160, output_3_1, output_2_160;
mixer gate_output_2_160(.a(output_3_160), .b(output_3_1), .y(output_2_160));
wire output_4_160, output_4_1, output_3_160;
mixer gate_output_3_160(.a(output_4_160), .b(output_4_1), .y(output_3_160));
wire output_1_161, output_1_2, output_0_161;
mixer gate_output_0_161(.a(output_1_161), .b(output_1_2), .y(output_0_161));
wire output_2_161, output_2_2, output_1_161;
mixer gate_output_1_161(.a(output_2_161), .b(output_2_2), .y(output_1_161));
wire output_3_161, output_3_2, output_2_161;
mixer gate_output_2_161(.a(output_3_161), .b(output_3_2), .y(output_2_161));
wire output_4_161, output_4_2, output_3_161;
mixer gate_output_3_161(.a(output_4_161), .b(output_4_2), .y(output_3_161));
wire output_1_162, output_1_3, output_0_162;
mixer gate_output_0_162(.a(output_1_162), .b(output_1_3), .y(output_0_162));
wire output_2_162, output_2_3, output_1_162;
mixer gate_output_1_162(.a(output_2_162), .b(output_2_3), .y(output_1_162));
wire output_3_162, output_3_3, output_2_162;
mixer gate_output_2_162(.a(output_3_162), .b(output_3_3), .y(output_2_162));
wire output_4_162, output_4_3, output_3_162;
mixer gate_output_3_162(.a(output_4_162), .b(output_4_3), .y(output_3_162));
wire output_1_163, output_1_0, output_0_163;
mixer gate_output_0_163(.a(output_1_163), .b(output_1_0), .y(output_0_163));
wire output_2_163, output_2_0, output_1_163;
mixer gate_output_1_163(.a(output_2_163), .b(output_2_0), .y(output_1_163));
wire output_3_163, output_3_0, output_2_163;
mixer gate_output_2_163(.a(output_3_163), .b(output_3_0), .y(output_2_163));
wire output_4_163, output_4_0, output_3_163;
mixer gate_output_3_163(.a(output_4_163), .b(output_4_0), .y(output_3_163));
wire output_1_164, output_1_1, output_0_164;
mixer gate_output_0_164(.a(output_1_164), .b(output_1_1), .y(output_0_164));
wire output_2_164, output_2_1, output_1_164;
mixer gate_output_1_164(.a(output_2_164), .b(output_2_1), .y(output_1_164));
wire output_3_164, output_3_1, output_2_164;
mixer gate_output_2_164(.a(output_3_164), .b(output_3_1), .y(output_2_164));
wire output_4_164, output_4_1, output_3_164;
mixer gate_output_3_164(.a(output_4_164), .b(output_4_1), .y(output_3_164));
wire output_1_165, output_1_2, output_0_165;
mixer gate_output_0_165(.a(output_1_165), .b(output_1_2), .y(output_0_165));
wire output_2_165, output_2_2, output_1_165;
mixer gate_output_1_165(.a(output_2_165), .b(output_2_2), .y(output_1_165));
wire output_3_165, output_3_2, output_2_165;
mixer gate_output_2_165(.a(output_3_165), .b(output_3_2), .y(output_2_165));
wire output_4_165, output_4_2, output_3_165;
mixer gate_output_3_165(.a(output_4_165), .b(output_4_2), .y(output_3_165));
wire output_1_166, output_1_3, output_0_166;
mixer gate_output_0_166(.a(output_1_166), .b(output_1_3), .y(output_0_166));
wire output_2_166, output_2_3, output_1_166;
mixer gate_output_1_166(.a(output_2_166), .b(output_2_3), .y(output_1_166));
wire output_3_166, output_3_3, output_2_166;
mixer gate_output_2_166(.a(output_3_166), .b(output_3_3), .y(output_2_166));
wire output_4_166, output_4_3, output_3_166;
mixer gate_output_3_166(.a(output_4_166), .b(output_4_3), .y(output_3_166));
wire output_1_167, output_1_0, output_0_167;
mixer gate_output_0_167(.a(output_1_167), .b(output_1_0), .y(output_0_167));
wire output_2_167, output_2_0, output_1_167;
mixer gate_output_1_167(.a(output_2_167), .b(output_2_0), .y(output_1_167));
wire output_3_167, output_3_0, output_2_167;
mixer gate_output_2_167(.a(output_3_167), .b(output_3_0), .y(output_2_167));
wire output_4_167, output_4_0, output_3_167;
mixer gate_output_3_167(.a(output_4_167), .b(output_4_0), .y(output_3_167));
wire output_1_168, output_1_1, output_0_168;
mixer gate_output_0_168(.a(output_1_168), .b(output_1_1), .y(output_0_168));
wire output_2_168, output_2_1, output_1_168;
mixer gate_output_1_168(.a(output_2_168), .b(output_2_1), .y(output_1_168));
wire output_3_168, output_3_1, output_2_168;
mixer gate_output_2_168(.a(output_3_168), .b(output_3_1), .y(output_2_168));
wire output_4_168, output_4_1, output_3_168;
mixer gate_output_3_168(.a(output_4_168), .b(output_4_1), .y(output_3_168));
wire output_1_169, output_1_2, output_0_169;
mixer gate_output_0_169(.a(output_1_169), .b(output_1_2), .y(output_0_169));
wire output_2_169, output_2_2, output_1_169;
mixer gate_output_1_169(.a(output_2_169), .b(output_2_2), .y(output_1_169));
wire output_3_169, output_3_2, output_2_169;
mixer gate_output_2_169(.a(output_3_169), .b(output_3_2), .y(output_2_169));
wire output_4_169, output_4_2, output_3_169;
mixer gate_output_3_169(.a(output_4_169), .b(output_4_2), .y(output_3_169));
wire output_1_170, output_1_3, output_0_170;
mixer gate_output_0_170(.a(output_1_170), .b(output_1_3), .y(output_0_170));
wire output_2_170, output_2_3, output_1_170;
mixer gate_output_1_170(.a(output_2_170), .b(output_2_3), .y(output_1_170));
wire output_3_170, output_3_3, output_2_170;
mixer gate_output_2_170(.a(output_3_170), .b(output_3_3), .y(output_2_170));
wire output_4_170, output_4_3, output_3_170;
mixer gate_output_3_170(.a(output_4_170), .b(output_4_3), .y(output_3_170));
wire output_1_171, output_1_0, output_0_171;
mixer gate_output_0_171(.a(output_1_171), .b(output_1_0), .y(output_0_171));
wire output_2_171, output_2_0, output_1_171;
mixer gate_output_1_171(.a(output_2_171), .b(output_2_0), .y(output_1_171));
wire output_3_171, output_3_0, output_2_171;
mixer gate_output_2_171(.a(output_3_171), .b(output_3_0), .y(output_2_171));
wire output_4_171, output_4_0, output_3_171;
mixer gate_output_3_171(.a(output_4_171), .b(output_4_0), .y(output_3_171));
wire output_1_172, output_1_1, output_0_172;
mixer gate_output_0_172(.a(output_1_172), .b(output_1_1), .y(output_0_172));
wire output_2_172, output_2_1, output_1_172;
mixer gate_output_1_172(.a(output_2_172), .b(output_2_1), .y(output_1_172));
wire output_3_172, output_3_1, output_2_172;
mixer gate_output_2_172(.a(output_3_172), .b(output_3_1), .y(output_2_172));
wire output_4_172, output_4_1, output_3_172;
mixer gate_output_3_172(.a(output_4_172), .b(output_4_1), .y(output_3_172));
wire output_1_173, output_1_2, output_0_173;
mixer gate_output_0_173(.a(output_1_173), .b(output_1_2), .y(output_0_173));
wire output_2_173, output_2_2, output_1_173;
mixer gate_output_1_173(.a(output_2_173), .b(output_2_2), .y(output_1_173));
wire output_3_173, output_3_2, output_2_173;
mixer gate_output_2_173(.a(output_3_173), .b(output_3_2), .y(output_2_173));
wire output_4_173, output_4_2, output_3_173;
mixer gate_output_3_173(.a(output_4_173), .b(output_4_2), .y(output_3_173));
wire output_1_174, output_1_3, output_0_174;
mixer gate_output_0_174(.a(output_1_174), .b(output_1_3), .y(output_0_174));
wire output_2_174, output_2_3, output_1_174;
mixer gate_output_1_174(.a(output_2_174), .b(output_2_3), .y(output_1_174));
wire output_3_174, output_3_3, output_2_174;
mixer gate_output_2_174(.a(output_3_174), .b(output_3_3), .y(output_2_174));
wire output_4_174, output_4_3, output_3_174;
mixer gate_output_3_174(.a(output_4_174), .b(output_4_3), .y(output_3_174));
wire output_1_175, output_1_0, output_0_175;
mixer gate_output_0_175(.a(output_1_175), .b(output_1_0), .y(output_0_175));
wire output_2_175, output_2_0, output_1_175;
mixer gate_output_1_175(.a(output_2_175), .b(output_2_0), .y(output_1_175));
wire output_3_175, output_3_0, output_2_175;
mixer gate_output_2_175(.a(output_3_175), .b(output_3_0), .y(output_2_175));
wire output_4_175, output_4_0, output_3_175;
mixer gate_output_3_175(.a(output_4_175), .b(output_4_0), .y(output_3_175));
wire output_1_176, output_1_1, output_0_176;
mixer gate_output_0_176(.a(output_1_176), .b(output_1_1), .y(output_0_176));
wire output_2_176, output_2_1, output_1_176;
mixer gate_output_1_176(.a(output_2_176), .b(output_2_1), .y(output_1_176));
wire output_3_176, output_3_1, output_2_176;
mixer gate_output_2_176(.a(output_3_176), .b(output_3_1), .y(output_2_176));
wire output_4_176, output_4_1, output_3_176;
mixer gate_output_3_176(.a(output_4_176), .b(output_4_1), .y(output_3_176));
wire output_1_177, output_1_2, output_0_177;
mixer gate_output_0_177(.a(output_1_177), .b(output_1_2), .y(output_0_177));
wire output_2_177, output_2_2, output_1_177;
mixer gate_output_1_177(.a(output_2_177), .b(output_2_2), .y(output_1_177));
wire output_3_177, output_3_2, output_2_177;
mixer gate_output_2_177(.a(output_3_177), .b(output_3_2), .y(output_2_177));
wire output_4_177, output_4_2, output_3_177;
mixer gate_output_3_177(.a(output_4_177), .b(output_4_2), .y(output_3_177));
wire output_1_178, output_1_3, output_0_178;
mixer gate_output_0_178(.a(output_1_178), .b(output_1_3), .y(output_0_178));
wire output_2_178, output_2_3, output_1_178;
mixer gate_output_1_178(.a(output_2_178), .b(output_2_3), .y(output_1_178));
wire output_3_178, output_3_3, output_2_178;
mixer gate_output_2_178(.a(output_3_178), .b(output_3_3), .y(output_2_178));
wire output_4_178, output_4_3, output_3_178;
mixer gate_output_3_178(.a(output_4_178), .b(output_4_3), .y(output_3_178));
wire output_1_179, output_1_0, output_0_179;
mixer gate_output_0_179(.a(output_1_179), .b(output_1_0), .y(output_0_179));
wire output_2_179, output_2_0, output_1_179;
mixer gate_output_1_179(.a(output_2_179), .b(output_2_0), .y(output_1_179));
wire output_3_179, output_3_0, output_2_179;
mixer gate_output_2_179(.a(output_3_179), .b(output_3_0), .y(output_2_179));
wire output_4_179, output_4_0, output_3_179;
mixer gate_output_3_179(.a(output_4_179), .b(output_4_0), .y(output_3_179));
wire output_1_180, output_1_1, output_0_180;
mixer gate_output_0_180(.a(output_1_180), .b(output_1_1), .y(output_0_180));
wire output_2_180, output_2_1, output_1_180;
mixer gate_output_1_180(.a(output_2_180), .b(output_2_1), .y(output_1_180));
wire output_3_180, output_3_1, output_2_180;
mixer gate_output_2_180(.a(output_3_180), .b(output_3_1), .y(output_2_180));
wire output_4_180, output_4_1, output_3_180;
mixer gate_output_3_180(.a(output_4_180), .b(output_4_1), .y(output_3_180));
wire output_1_181, output_1_2, output_0_181;
mixer gate_output_0_181(.a(output_1_181), .b(output_1_2), .y(output_0_181));
wire output_2_181, output_2_2, output_1_181;
mixer gate_output_1_181(.a(output_2_181), .b(output_2_2), .y(output_1_181));
wire output_3_181, output_3_2, output_2_181;
mixer gate_output_2_181(.a(output_3_181), .b(output_3_2), .y(output_2_181));
wire output_4_181, output_4_2, output_3_181;
mixer gate_output_3_181(.a(output_4_181), .b(output_4_2), .y(output_3_181));
wire output_1_182, output_1_3, output_0_182;
mixer gate_output_0_182(.a(output_1_182), .b(output_1_3), .y(output_0_182));
wire output_2_182, output_2_3, output_1_182;
mixer gate_output_1_182(.a(output_2_182), .b(output_2_3), .y(output_1_182));
wire output_3_182, output_3_3, output_2_182;
mixer gate_output_2_182(.a(output_3_182), .b(output_3_3), .y(output_2_182));
wire output_4_182, output_4_3, output_3_182;
mixer gate_output_3_182(.a(output_4_182), .b(output_4_3), .y(output_3_182));
wire output_1_183, output_1_0, output_0_183;
mixer gate_output_0_183(.a(output_1_183), .b(output_1_0), .y(output_0_183));
wire output_2_183, output_2_0, output_1_183;
mixer gate_output_1_183(.a(output_2_183), .b(output_2_0), .y(output_1_183));
wire output_3_183, output_3_0, output_2_183;
mixer gate_output_2_183(.a(output_3_183), .b(output_3_0), .y(output_2_183));
wire output_4_183, output_4_0, output_3_183;
mixer gate_output_3_183(.a(output_4_183), .b(output_4_0), .y(output_3_183));
wire output_1_184, output_1_1, output_0_184;
mixer gate_output_0_184(.a(output_1_184), .b(output_1_1), .y(output_0_184));
wire output_2_184, output_2_1, output_1_184;
mixer gate_output_1_184(.a(output_2_184), .b(output_2_1), .y(output_1_184));
wire output_3_184, output_3_1, output_2_184;
mixer gate_output_2_184(.a(output_3_184), .b(output_3_1), .y(output_2_184));
wire output_4_184, output_4_1, output_3_184;
mixer gate_output_3_184(.a(output_4_184), .b(output_4_1), .y(output_3_184));
wire output_1_185, output_1_2, output_0_185;
mixer gate_output_0_185(.a(output_1_185), .b(output_1_2), .y(output_0_185));
wire output_2_185, output_2_2, output_1_185;
mixer gate_output_1_185(.a(output_2_185), .b(output_2_2), .y(output_1_185));
wire output_3_185, output_3_2, output_2_185;
mixer gate_output_2_185(.a(output_3_185), .b(output_3_2), .y(output_2_185));
wire output_4_185, output_4_2, output_3_185;
mixer gate_output_3_185(.a(output_4_185), .b(output_4_2), .y(output_3_185));
wire output_1_186, output_1_3, output_0_186;
mixer gate_output_0_186(.a(output_1_186), .b(output_1_3), .y(output_0_186));
wire output_2_186, output_2_3, output_1_186;
mixer gate_output_1_186(.a(output_2_186), .b(output_2_3), .y(output_1_186));
wire output_3_186, output_3_3, output_2_186;
mixer gate_output_2_186(.a(output_3_186), .b(output_3_3), .y(output_2_186));
wire output_4_186, output_4_3, output_3_186;
mixer gate_output_3_186(.a(output_4_186), .b(output_4_3), .y(output_3_186));
wire output_1_187, output_1_0, output_0_187;
mixer gate_output_0_187(.a(output_1_187), .b(output_1_0), .y(output_0_187));
wire output_2_187, output_2_0, output_1_187;
mixer gate_output_1_187(.a(output_2_187), .b(output_2_0), .y(output_1_187));
wire output_3_187, output_3_0, output_2_187;
mixer gate_output_2_187(.a(output_3_187), .b(output_3_0), .y(output_2_187));
wire output_4_187, output_4_0, output_3_187;
mixer gate_output_3_187(.a(output_4_187), .b(output_4_0), .y(output_3_187));
wire output_1_188, output_1_1, output_0_188;
mixer gate_output_0_188(.a(output_1_188), .b(output_1_1), .y(output_0_188));
wire output_2_188, output_2_1, output_1_188;
mixer gate_output_1_188(.a(output_2_188), .b(output_2_1), .y(output_1_188));
wire output_3_188, output_3_1, output_2_188;
mixer gate_output_2_188(.a(output_3_188), .b(output_3_1), .y(output_2_188));
wire output_4_188, output_4_1, output_3_188;
mixer gate_output_3_188(.a(output_4_188), .b(output_4_1), .y(output_3_188));
wire output_1_189, output_1_2, output_0_189;
mixer gate_output_0_189(.a(output_1_189), .b(output_1_2), .y(output_0_189));
wire output_2_189, output_2_2, output_1_189;
mixer gate_output_1_189(.a(output_2_189), .b(output_2_2), .y(output_1_189));
wire output_3_189, output_3_2, output_2_189;
mixer gate_output_2_189(.a(output_3_189), .b(output_3_2), .y(output_2_189));
wire output_4_189, output_4_2, output_3_189;
mixer gate_output_3_189(.a(output_4_189), .b(output_4_2), .y(output_3_189));
wire output_1_190, output_1_3, output_0_190;
mixer gate_output_0_190(.a(output_1_190), .b(output_1_3), .y(output_0_190));
wire output_2_190, output_2_3, output_1_190;
mixer gate_output_1_190(.a(output_2_190), .b(output_2_3), .y(output_1_190));
wire output_3_190, output_3_3, output_2_190;
mixer gate_output_2_190(.a(output_3_190), .b(output_3_3), .y(output_2_190));
wire output_4_190, output_4_3, output_3_190;
mixer gate_output_3_190(.a(output_4_190), .b(output_4_3), .y(output_3_190));
wire output_1_191, output_1_0, output_0_191;
mixer gate_output_0_191(.a(output_1_191), .b(output_1_0), .y(output_0_191));
wire output_2_191, output_2_0, output_1_191;
mixer gate_output_1_191(.a(output_2_191), .b(output_2_0), .y(output_1_191));
wire output_3_191, output_3_0, output_2_191;
mixer gate_output_2_191(.a(output_3_191), .b(output_3_0), .y(output_2_191));
wire output_4_191, output_4_0, output_3_191;
mixer gate_output_3_191(.a(output_4_191), .b(output_4_0), .y(output_3_191));
wire output_1_192, output_1_1, output_0_192;
mixer gate_output_0_192(.a(output_1_192), .b(output_1_1), .y(output_0_192));
wire output_2_192, output_2_1, output_1_192;
mixer gate_output_1_192(.a(output_2_192), .b(output_2_1), .y(output_1_192));
wire output_3_192, output_3_1, output_2_192;
mixer gate_output_2_192(.a(output_3_192), .b(output_3_1), .y(output_2_192));
wire output_4_192, output_4_1, output_3_192;
mixer gate_output_3_192(.a(output_4_192), .b(output_4_1), .y(output_3_192));
wire output_1_193, output_1_2, output_0_193;
mixer gate_output_0_193(.a(output_1_193), .b(output_1_2), .y(output_0_193));
wire output_2_193, output_2_2, output_1_193;
mixer gate_output_1_193(.a(output_2_193), .b(output_2_2), .y(output_1_193));
wire output_3_193, output_3_2, output_2_193;
mixer gate_output_2_193(.a(output_3_193), .b(output_3_2), .y(output_2_193));
wire output_4_193, output_4_2, output_3_193;
mixer gate_output_3_193(.a(output_4_193), .b(output_4_2), .y(output_3_193));
wire output_1_194, output_1_3, output_0_194;
mixer gate_output_0_194(.a(output_1_194), .b(output_1_3), .y(output_0_194));
wire output_2_194, output_2_3, output_1_194;
mixer gate_output_1_194(.a(output_2_194), .b(output_2_3), .y(output_1_194));
wire output_3_194, output_3_3, output_2_194;
mixer gate_output_2_194(.a(output_3_194), .b(output_3_3), .y(output_2_194));
wire output_4_194, output_4_3, output_3_194;
mixer gate_output_3_194(.a(output_4_194), .b(output_4_3), .y(output_3_194));
wire output_1_195, output_1_0, output_0_195;
mixer gate_output_0_195(.a(output_1_195), .b(output_1_0), .y(output_0_195));
wire output_2_195, output_2_0, output_1_195;
mixer gate_output_1_195(.a(output_2_195), .b(output_2_0), .y(output_1_195));
wire output_3_195, output_3_0, output_2_195;
mixer gate_output_2_195(.a(output_3_195), .b(output_3_0), .y(output_2_195));
wire output_4_195, output_4_0, output_3_195;
mixer gate_output_3_195(.a(output_4_195), .b(output_4_0), .y(output_3_195));
wire output_1_196, output_1_1, output_0_196;
mixer gate_output_0_196(.a(output_1_196), .b(output_1_1), .y(output_0_196));
wire output_2_196, output_2_1, output_1_196;
mixer gate_output_1_196(.a(output_2_196), .b(output_2_1), .y(output_1_196));
wire output_3_196, output_3_1, output_2_196;
mixer gate_output_2_196(.a(output_3_196), .b(output_3_1), .y(output_2_196));
wire output_4_196, output_4_1, output_3_196;
mixer gate_output_3_196(.a(output_4_196), .b(output_4_1), .y(output_3_196));
wire output_1_197, output_1_2, output_0_197;
mixer gate_output_0_197(.a(output_1_197), .b(output_1_2), .y(output_0_197));
wire output_2_197, output_2_2, output_1_197;
mixer gate_output_1_197(.a(output_2_197), .b(output_2_2), .y(output_1_197));
wire output_3_197, output_3_2, output_2_197;
mixer gate_output_2_197(.a(output_3_197), .b(output_3_2), .y(output_2_197));
wire output_4_197, output_4_2, output_3_197;
mixer gate_output_3_197(.a(output_4_197), .b(output_4_2), .y(output_3_197));
wire output_1_198, output_1_3, output_0_198;
mixer gate_output_0_198(.a(output_1_198), .b(output_1_3), .y(output_0_198));
wire output_2_198, output_2_3, output_1_198;
mixer gate_output_1_198(.a(output_2_198), .b(output_2_3), .y(output_1_198));
wire output_3_198, output_3_3, output_2_198;
mixer gate_output_2_198(.a(output_3_198), .b(output_3_3), .y(output_2_198));
wire output_4_198, output_4_3, output_3_198;
mixer gate_output_3_198(.a(output_4_198), .b(output_4_3), .y(output_3_198));
wire output_1_199, output_1_0, output_0_199;
mixer gate_output_0_199(.a(output_1_199), .b(output_1_0), .y(output_0_199));
wire output_2_199, output_2_0, output_1_199;
mixer gate_output_1_199(.a(output_2_199), .b(output_2_0), .y(output_1_199));
wire output_3_199, output_3_0, output_2_199;
mixer gate_output_2_199(.a(output_3_199), .b(output_3_0), .y(output_2_199));
wire output_4_199, output_4_0, output_3_199;
mixer gate_output_3_199(.a(output_4_199), .b(output_4_0), .y(output_3_199));
wire output_1_200, output_1_1, output_0_200;
mixer gate_output_0_200(.a(output_1_200), .b(output_1_1), .y(output_0_200));
wire output_2_200, output_2_1, output_1_200;
mixer gate_output_1_200(.a(output_2_200), .b(output_2_1), .y(output_1_200));
wire output_3_200, output_3_1, output_2_200;
mixer gate_output_2_200(.a(output_3_200), .b(output_3_1), .y(output_2_200));
wire output_4_200, output_4_1, output_3_200;
mixer gate_output_3_200(.a(output_4_200), .b(output_4_1), .y(output_3_200));
wire output_1_201, output_1_2, output_0_201;
mixer gate_output_0_201(.a(output_1_201), .b(output_1_2), .y(output_0_201));
wire output_2_201, output_2_2, output_1_201;
mixer gate_output_1_201(.a(output_2_201), .b(output_2_2), .y(output_1_201));
wire output_3_201, output_3_2, output_2_201;
mixer gate_output_2_201(.a(output_3_201), .b(output_3_2), .y(output_2_201));
wire output_4_201, output_4_2, output_3_201;
mixer gate_output_3_201(.a(output_4_201), .b(output_4_2), .y(output_3_201));
wire output_1_202, output_1_3, output_0_202;
mixer gate_output_0_202(.a(output_1_202), .b(output_1_3), .y(output_0_202));
wire output_2_202, output_2_3, output_1_202;
mixer gate_output_1_202(.a(output_2_202), .b(output_2_3), .y(output_1_202));
wire output_3_202, output_3_3, output_2_202;
mixer gate_output_2_202(.a(output_3_202), .b(output_3_3), .y(output_2_202));
wire output_4_202, output_4_3, output_3_202;
mixer gate_output_3_202(.a(output_4_202), .b(output_4_3), .y(output_3_202));
wire output_1_203, output_1_0, output_0_203;
mixer gate_output_0_203(.a(output_1_203), .b(output_1_0), .y(output_0_203));
wire output_2_203, output_2_0, output_1_203;
mixer gate_output_1_203(.a(output_2_203), .b(output_2_0), .y(output_1_203));
wire output_3_203, output_3_0, output_2_203;
mixer gate_output_2_203(.a(output_3_203), .b(output_3_0), .y(output_2_203));
wire output_4_203, output_4_0, output_3_203;
mixer gate_output_3_203(.a(output_4_203), .b(output_4_0), .y(output_3_203));
wire output_1_204, output_1_1, output_0_204;
mixer gate_output_0_204(.a(output_1_204), .b(output_1_1), .y(output_0_204));
wire output_2_204, output_2_1, output_1_204;
mixer gate_output_1_204(.a(output_2_204), .b(output_2_1), .y(output_1_204));
wire output_3_204, output_3_1, output_2_204;
mixer gate_output_2_204(.a(output_3_204), .b(output_3_1), .y(output_2_204));
wire output_4_204, output_4_1, output_3_204;
mixer gate_output_3_204(.a(output_4_204), .b(output_4_1), .y(output_3_204));
wire output_1_205, output_1_2, output_0_205;
mixer gate_output_0_205(.a(output_1_205), .b(output_1_2), .y(output_0_205));
wire output_2_205, output_2_2, output_1_205;
mixer gate_output_1_205(.a(output_2_205), .b(output_2_2), .y(output_1_205));
wire output_3_205, output_3_2, output_2_205;
mixer gate_output_2_205(.a(output_3_205), .b(output_3_2), .y(output_2_205));
wire output_4_205, output_4_2, output_3_205;
mixer gate_output_3_205(.a(output_4_205), .b(output_4_2), .y(output_3_205));
wire output_1_206, output_1_3, output_0_206;
mixer gate_output_0_206(.a(output_1_206), .b(output_1_3), .y(output_0_206));
wire output_2_206, output_2_3, output_1_206;
mixer gate_output_1_206(.a(output_2_206), .b(output_2_3), .y(output_1_206));
wire output_3_206, output_3_3, output_2_206;
mixer gate_output_2_206(.a(output_3_206), .b(output_3_3), .y(output_2_206));
wire output_4_206, output_4_3, output_3_206;
mixer gate_output_3_206(.a(output_4_206), .b(output_4_3), .y(output_3_206));
wire output_1_207, output_1_0, output_0_207;
mixer gate_output_0_207(.a(output_1_207), .b(output_1_0), .y(output_0_207));
wire output_2_207, output_2_0, output_1_207;
mixer gate_output_1_207(.a(output_2_207), .b(output_2_0), .y(output_1_207));
wire output_3_207, output_3_0, output_2_207;
mixer gate_output_2_207(.a(output_3_207), .b(output_3_0), .y(output_2_207));
wire output_4_207, output_4_0, output_3_207;
mixer gate_output_3_207(.a(output_4_207), .b(output_4_0), .y(output_3_207));
wire output_1_208, output_1_1, output_0_208;
mixer gate_output_0_208(.a(output_1_208), .b(output_1_1), .y(output_0_208));
wire output_2_208, output_2_1, output_1_208;
mixer gate_output_1_208(.a(output_2_208), .b(output_2_1), .y(output_1_208));
wire output_3_208, output_3_1, output_2_208;
mixer gate_output_2_208(.a(output_3_208), .b(output_3_1), .y(output_2_208));
wire output_4_208, output_4_1, output_3_208;
mixer gate_output_3_208(.a(output_4_208), .b(output_4_1), .y(output_3_208));
wire output_1_209, output_1_2, output_0_209;
mixer gate_output_0_209(.a(output_1_209), .b(output_1_2), .y(output_0_209));
wire output_2_209, output_2_2, output_1_209;
mixer gate_output_1_209(.a(output_2_209), .b(output_2_2), .y(output_1_209));
wire output_3_209, output_3_2, output_2_209;
mixer gate_output_2_209(.a(output_3_209), .b(output_3_2), .y(output_2_209));
wire output_4_209, output_4_2, output_3_209;
mixer gate_output_3_209(.a(output_4_209), .b(output_4_2), .y(output_3_209));
wire output_1_210, output_1_3, output_0_210;
mixer gate_output_0_210(.a(output_1_210), .b(output_1_3), .y(output_0_210));
wire output_2_210, output_2_3, output_1_210;
mixer gate_output_1_210(.a(output_2_210), .b(output_2_3), .y(output_1_210));
wire output_3_210, output_3_3, output_2_210;
mixer gate_output_2_210(.a(output_3_210), .b(output_3_3), .y(output_2_210));
wire output_4_210, output_4_3, output_3_210;
mixer gate_output_3_210(.a(output_4_210), .b(output_4_3), .y(output_3_210));
wire output_1_211, output_1_0, output_0_211;
mixer gate_output_0_211(.a(output_1_211), .b(output_1_0), .y(output_0_211));
wire output_2_211, output_2_0, output_1_211;
mixer gate_output_1_211(.a(output_2_211), .b(output_2_0), .y(output_1_211));
wire output_3_211, output_3_0, output_2_211;
mixer gate_output_2_211(.a(output_3_211), .b(output_3_0), .y(output_2_211));
wire output_4_211, output_4_0, output_3_211;
mixer gate_output_3_211(.a(output_4_211), .b(output_4_0), .y(output_3_211));
wire output_1_212, output_1_1, output_0_212;
mixer gate_output_0_212(.a(output_1_212), .b(output_1_1), .y(output_0_212));
wire output_2_212, output_2_1, output_1_212;
mixer gate_output_1_212(.a(output_2_212), .b(output_2_1), .y(output_1_212));
wire output_3_212, output_3_1, output_2_212;
mixer gate_output_2_212(.a(output_3_212), .b(output_3_1), .y(output_2_212));
wire output_4_212, output_4_1, output_3_212;
mixer gate_output_3_212(.a(output_4_212), .b(output_4_1), .y(output_3_212));
wire output_1_213, output_1_2, output_0_213;
mixer gate_output_0_213(.a(output_1_213), .b(output_1_2), .y(output_0_213));
wire output_2_213, output_2_2, output_1_213;
mixer gate_output_1_213(.a(output_2_213), .b(output_2_2), .y(output_1_213));
wire output_3_213, output_3_2, output_2_213;
mixer gate_output_2_213(.a(output_3_213), .b(output_3_2), .y(output_2_213));
wire output_4_213, output_4_2, output_3_213;
mixer gate_output_3_213(.a(output_4_213), .b(output_4_2), .y(output_3_213));
wire output_1_214, output_1_3, output_0_214;
mixer gate_output_0_214(.a(output_1_214), .b(output_1_3), .y(output_0_214));
wire output_2_214, output_2_3, output_1_214;
mixer gate_output_1_214(.a(output_2_214), .b(output_2_3), .y(output_1_214));
wire output_3_214, output_3_3, output_2_214;
mixer gate_output_2_214(.a(output_3_214), .b(output_3_3), .y(output_2_214));
wire output_4_214, output_4_3, output_3_214;
mixer gate_output_3_214(.a(output_4_214), .b(output_4_3), .y(output_3_214));
wire output_1_215, output_1_0, output_0_215;
mixer gate_output_0_215(.a(output_1_215), .b(output_1_0), .y(output_0_215));
wire output_2_215, output_2_0, output_1_215;
mixer gate_output_1_215(.a(output_2_215), .b(output_2_0), .y(output_1_215));
wire output_3_215, output_3_0, output_2_215;
mixer gate_output_2_215(.a(output_3_215), .b(output_3_0), .y(output_2_215));
wire output_4_215, output_4_0, output_3_215;
mixer gate_output_3_215(.a(output_4_215), .b(output_4_0), .y(output_3_215));
wire output_1_216, output_1_1, output_0_216;
mixer gate_output_0_216(.a(output_1_216), .b(output_1_1), .y(output_0_216));
wire output_2_216, output_2_1, output_1_216;
mixer gate_output_1_216(.a(output_2_216), .b(output_2_1), .y(output_1_216));
wire output_3_216, output_3_1, output_2_216;
mixer gate_output_2_216(.a(output_3_216), .b(output_3_1), .y(output_2_216));
wire output_4_216, output_4_1, output_3_216;
mixer gate_output_3_216(.a(output_4_216), .b(output_4_1), .y(output_3_216));
wire output_1_217, output_1_2, output_0_217;
mixer gate_output_0_217(.a(output_1_217), .b(output_1_2), .y(output_0_217));
wire output_2_217, output_2_2, output_1_217;
mixer gate_output_1_217(.a(output_2_217), .b(output_2_2), .y(output_1_217));
wire output_3_217, output_3_2, output_2_217;
mixer gate_output_2_217(.a(output_3_217), .b(output_3_2), .y(output_2_217));
wire output_4_217, output_4_2, output_3_217;
mixer gate_output_3_217(.a(output_4_217), .b(output_4_2), .y(output_3_217));
wire output_1_218, output_1_3, output_0_218;
mixer gate_output_0_218(.a(output_1_218), .b(output_1_3), .y(output_0_218));
wire output_2_218, output_2_3, output_1_218;
mixer gate_output_1_218(.a(output_2_218), .b(output_2_3), .y(output_1_218));
wire output_3_218, output_3_3, output_2_218;
mixer gate_output_2_218(.a(output_3_218), .b(output_3_3), .y(output_2_218));
wire output_4_218, output_4_3, output_3_218;
mixer gate_output_3_218(.a(output_4_218), .b(output_4_3), .y(output_3_218));
wire output_1_219, output_1_0, output_0_219;
mixer gate_output_0_219(.a(output_1_219), .b(output_1_0), .y(output_0_219));
wire output_2_219, output_2_0, output_1_219;
mixer gate_output_1_219(.a(output_2_219), .b(output_2_0), .y(output_1_219));
wire output_3_219, output_3_0, output_2_219;
mixer gate_output_2_219(.a(output_3_219), .b(output_3_0), .y(output_2_219));
wire output_4_219, output_4_0, output_3_219;
mixer gate_output_3_219(.a(output_4_219), .b(output_4_0), .y(output_3_219));
wire output_1_220, output_1_1, output_0_220;
mixer gate_output_0_220(.a(output_1_220), .b(output_1_1), .y(output_0_220));
wire output_2_220, output_2_1, output_1_220;
mixer gate_output_1_220(.a(output_2_220), .b(output_2_1), .y(output_1_220));
wire output_3_220, output_3_1, output_2_220;
mixer gate_output_2_220(.a(output_3_220), .b(output_3_1), .y(output_2_220));
wire output_4_220, output_4_1, output_3_220;
mixer gate_output_3_220(.a(output_4_220), .b(output_4_1), .y(output_3_220));
wire output_1_221, output_1_2, output_0_221;
mixer gate_output_0_221(.a(output_1_221), .b(output_1_2), .y(output_0_221));
wire output_2_221, output_2_2, output_1_221;
mixer gate_output_1_221(.a(output_2_221), .b(output_2_2), .y(output_1_221));
wire output_3_221, output_3_2, output_2_221;
mixer gate_output_2_221(.a(output_3_221), .b(output_3_2), .y(output_2_221));
wire output_4_221, output_4_2, output_3_221;
mixer gate_output_3_221(.a(output_4_221), .b(output_4_2), .y(output_3_221));
wire output_1_222, output_1_3, output_0_222;
mixer gate_output_0_222(.a(output_1_222), .b(output_1_3), .y(output_0_222));
wire output_2_222, output_2_3, output_1_222;
mixer gate_output_1_222(.a(output_2_222), .b(output_2_3), .y(output_1_222));
wire output_3_222, output_3_3, output_2_222;
mixer gate_output_2_222(.a(output_3_222), .b(output_3_3), .y(output_2_222));
wire output_4_222, output_4_3, output_3_222;
mixer gate_output_3_222(.a(output_4_222), .b(output_4_3), .y(output_3_222));
wire output_1_223, output_1_0, output_0_223;
mixer gate_output_0_223(.a(output_1_223), .b(output_1_0), .y(output_0_223));
wire output_2_223, output_2_0, output_1_223;
mixer gate_output_1_223(.a(output_2_223), .b(output_2_0), .y(output_1_223));
wire output_3_223, output_3_0, output_2_223;
mixer gate_output_2_223(.a(output_3_223), .b(output_3_0), .y(output_2_223));
wire output_4_223, output_4_0, output_3_223;
mixer gate_output_3_223(.a(output_4_223), .b(output_4_0), .y(output_3_223));
wire output_1_224, output_1_1, output_0_224;
mixer gate_output_0_224(.a(output_1_224), .b(output_1_1), .y(output_0_224));
wire output_2_224, output_2_1, output_1_224;
mixer gate_output_1_224(.a(output_2_224), .b(output_2_1), .y(output_1_224));
wire output_3_224, output_3_1, output_2_224;
mixer gate_output_2_224(.a(output_3_224), .b(output_3_1), .y(output_2_224));
wire output_4_224, output_4_1, output_3_224;
mixer gate_output_3_224(.a(output_4_224), .b(output_4_1), .y(output_3_224));
wire output_1_225, output_1_2, output_0_225;
mixer gate_output_0_225(.a(output_1_225), .b(output_1_2), .y(output_0_225));
wire output_2_225, output_2_2, output_1_225;
mixer gate_output_1_225(.a(output_2_225), .b(output_2_2), .y(output_1_225));
wire output_3_225, output_3_2, output_2_225;
mixer gate_output_2_225(.a(output_3_225), .b(output_3_2), .y(output_2_225));
wire output_4_225, output_4_2, output_3_225;
mixer gate_output_3_225(.a(output_4_225), .b(output_4_2), .y(output_3_225));
wire output_1_226, output_1_3, output_0_226;
mixer gate_output_0_226(.a(output_1_226), .b(output_1_3), .y(output_0_226));
wire output_2_226, output_2_3, output_1_226;
mixer gate_output_1_226(.a(output_2_226), .b(output_2_3), .y(output_1_226));
wire output_3_226, output_3_3, output_2_226;
mixer gate_output_2_226(.a(output_3_226), .b(output_3_3), .y(output_2_226));
wire output_4_226, output_4_3, output_3_226;
mixer gate_output_3_226(.a(output_4_226), .b(output_4_3), .y(output_3_226));
wire output_1_227, output_1_0, output_0_227;
mixer gate_output_0_227(.a(output_1_227), .b(output_1_0), .y(output_0_227));
wire output_2_227, output_2_0, output_1_227;
mixer gate_output_1_227(.a(output_2_227), .b(output_2_0), .y(output_1_227));
wire output_3_227, output_3_0, output_2_227;
mixer gate_output_2_227(.a(output_3_227), .b(output_3_0), .y(output_2_227));
wire output_4_227, output_4_0, output_3_227;
mixer gate_output_3_227(.a(output_4_227), .b(output_4_0), .y(output_3_227));
wire output_1_228, output_1_1, output_0_228;
mixer gate_output_0_228(.a(output_1_228), .b(output_1_1), .y(output_0_228));
wire output_2_228, output_2_1, output_1_228;
mixer gate_output_1_228(.a(output_2_228), .b(output_2_1), .y(output_1_228));
wire output_3_228, output_3_1, output_2_228;
mixer gate_output_2_228(.a(output_3_228), .b(output_3_1), .y(output_2_228));
wire output_4_228, output_4_1, output_3_228;
mixer gate_output_3_228(.a(output_4_228), .b(output_4_1), .y(output_3_228));
wire output_1_229, output_1_2, output_0_229;
mixer gate_output_0_229(.a(output_1_229), .b(output_1_2), .y(output_0_229));
wire output_2_229, output_2_2, output_1_229;
mixer gate_output_1_229(.a(output_2_229), .b(output_2_2), .y(output_1_229));
wire output_3_229, output_3_2, output_2_229;
mixer gate_output_2_229(.a(output_3_229), .b(output_3_2), .y(output_2_229));
wire output_4_229, output_4_2, output_3_229;
mixer gate_output_3_229(.a(output_4_229), .b(output_4_2), .y(output_3_229));
wire output_1_230, output_1_3, output_0_230;
mixer gate_output_0_230(.a(output_1_230), .b(output_1_3), .y(output_0_230));
wire output_2_230, output_2_3, output_1_230;
mixer gate_output_1_230(.a(output_2_230), .b(output_2_3), .y(output_1_230));
wire output_3_230, output_3_3, output_2_230;
mixer gate_output_2_230(.a(output_3_230), .b(output_3_3), .y(output_2_230));
wire output_4_230, output_4_3, output_3_230;
mixer gate_output_3_230(.a(output_4_230), .b(output_4_3), .y(output_3_230));
wire output_1_231, output_1_0, output_0_231;
mixer gate_output_0_231(.a(output_1_231), .b(output_1_0), .y(output_0_231));
wire output_2_231, output_2_0, output_1_231;
mixer gate_output_1_231(.a(output_2_231), .b(output_2_0), .y(output_1_231));
wire output_3_231, output_3_0, output_2_231;
mixer gate_output_2_231(.a(output_3_231), .b(output_3_0), .y(output_2_231));
wire output_4_231, output_4_0, output_3_231;
mixer gate_output_3_231(.a(output_4_231), .b(output_4_0), .y(output_3_231));
wire output_1_232, output_1_1, output_0_232;
mixer gate_output_0_232(.a(output_1_232), .b(output_1_1), .y(output_0_232));
wire output_2_232, output_2_1, output_1_232;
mixer gate_output_1_232(.a(output_2_232), .b(output_2_1), .y(output_1_232));
wire output_3_232, output_3_1, output_2_232;
mixer gate_output_2_232(.a(output_3_232), .b(output_3_1), .y(output_2_232));
wire output_4_232, output_4_1, output_3_232;
mixer gate_output_3_232(.a(output_4_232), .b(output_4_1), .y(output_3_232));
wire output_1_233, output_1_2, output_0_233;
mixer gate_output_0_233(.a(output_1_233), .b(output_1_2), .y(output_0_233));
wire output_2_233, output_2_2, output_1_233;
mixer gate_output_1_233(.a(output_2_233), .b(output_2_2), .y(output_1_233));
wire output_3_233, output_3_2, output_2_233;
mixer gate_output_2_233(.a(output_3_233), .b(output_3_2), .y(output_2_233));
wire output_4_233, output_4_2, output_3_233;
mixer gate_output_3_233(.a(output_4_233), .b(output_4_2), .y(output_3_233));
wire output_1_234, output_1_3, output_0_234;
mixer gate_output_0_234(.a(output_1_234), .b(output_1_3), .y(output_0_234));
wire output_2_234, output_2_3, output_1_234;
mixer gate_output_1_234(.a(output_2_234), .b(output_2_3), .y(output_1_234));
wire output_3_234, output_3_3, output_2_234;
mixer gate_output_2_234(.a(output_3_234), .b(output_3_3), .y(output_2_234));
wire output_4_234, output_4_3, output_3_234;
mixer gate_output_3_234(.a(output_4_234), .b(output_4_3), .y(output_3_234));
wire output_1_235, output_1_0, output_0_235;
mixer gate_output_0_235(.a(output_1_235), .b(output_1_0), .y(output_0_235));
wire output_2_235, output_2_0, output_1_235;
mixer gate_output_1_235(.a(output_2_235), .b(output_2_0), .y(output_1_235));
wire output_3_235, output_3_0, output_2_235;
mixer gate_output_2_235(.a(output_3_235), .b(output_3_0), .y(output_2_235));
wire output_4_235, output_4_0, output_3_235;
mixer gate_output_3_235(.a(output_4_235), .b(output_4_0), .y(output_3_235));
wire output_1_236, output_1_1, output_0_236;
mixer gate_output_0_236(.a(output_1_236), .b(output_1_1), .y(output_0_236));
wire output_2_236, output_2_1, output_1_236;
mixer gate_output_1_236(.a(output_2_236), .b(output_2_1), .y(output_1_236));
wire output_3_236, output_3_1, output_2_236;
mixer gate_output_2_236(.a(output_3_236), .b(output_3_1), .y(output_2_236));
wire output_4_236, output_4_1, output_3_236;
mixer gate_output_3_236(.a(output_4_236), .b(output_4_1), .y(output_3_236));
wire output_1_237, output_1_2, output_0_237;
mixer gate_output_0_237(.a(output_1_237), .b(output_1_2), .y(output_0_237));
wire output_2_237, output_2_2, output_1_237;
mixer gate_output_1_237(.a(output_2_237), .b(output_2_2), .y(output_1_237));
wire output_3_237, output_3_2, output_2_237;
mixer gate_output_2_237(.a(output_3_237), .b(output_3_2), .y(output_2_237));
wire output_4_237, output_4_2, output_3_237;
mixer gate_output_3_237(.a(output_4_237), .b(output_4_2), .y(output_3_237));
wire output_1_238, output_1_3, output_0_238;
mixer gate_output_0_238(.a(output_1_238), .b(output_1_3), .y(output_0_238));
wire output_2_238, output_2_3, output_1_238;
mixer gate_output_1_238(.a(output_2_238), .b(output_2_3), .y(output_1_238));
wire output_3_238, output_3_3, output_2_238;
mixer gate_output_2_238(.a(output_3_238), .b(output_3_3), .y(output_2_238));
wire output_4_238, output_4_3, output_3_238;
mixer gate_output_3_238(.a(output_4_238), .b(output_4_3), .y(output_3_238));
wire output_1_239, output_1_0, output_0_239;
mixer gate_output_0_239(.a(output_1_239), .b(output_1_0), .y(output_0_239));
wire output_2_239, output_2_0, output_1_239;
mixer gate_output_1_239(.a(output_2_239), .b(output_2_0), .y(output_1_239));
wire output_3_239, output_3_0, output_2_239;
mixer gate_output_2_239(.a(output_3_239), .b(output_3_0), .y(output_2_239));
wire output_4_239, output_4_0, output_3_239;
mixer gate_output_3_239(.a(output_4_239), .b(output_4_0), .y(output_3_239));
wire output_1_240, output_1_1, output_0_240;
mixer gate_output_0_240(.a(output_1_240), .b(output_1_1), .y(output_0_240));
wire output_2_240, output_2_1, output_1_240;
mixer gate_output_1_240(.a(output_2_240), .b(output_2_1), .y(output_1_240));
wire output_3_240, output_3_1, output_2_240;
mixer gate_output_2_240(.a(output_3_240), .b(output_3_1), .y(output_2_240));
wire output_4_240, output_4_1, output_3_240;
mixer gate_output_3_240(.a(output_4_240), .b(output_4_1), .y(output_3_240));
wire output_1_241, output_1_2, output_0_241;
mixer gate_output_0_241(.a(output_1_241), .b(output_1_2), .y(output_0_241));
wire output_2_241, output_2_2, output_1_241;
mixer gate_output_1_241(.a(output_2_241), .b(output_2_2), .y(output_1_241));
wire output_3_241, output_3_2, output_2_241;
mixer gate_output_2_241(.a(output_3_241), .b(output_3_2), .y(output_2_241));
wire output_4_241, output_4_2, output_3_241;
mixer gate_output_3_241(.a(output_4_241), .b(output_4_2), .y(output_3_241));
wire output_1_242, output_1_3, output_0_242;
mixer gate_output_0_242(.a(output_1_242), .b(output_1_3), .y(output_0_242));
wire output_2_242, output_2_3, output_1_242;
mixer gate_output_1_242(.a(output_2_242), .b(output_2_3), .y(output_1_242));
wire output_3_242, output_3_3, output_2_242;
mixer gate_output_2_242(.a(output_3_242), .b(output_3_3), .y(output_2_242));
wire output_4_242, output_4_3, output_3_242;
mixer gate_output_3_242(.a(output_4_242), .b(output_4_3), .y(output_3_242));
wire output_1_243, output_1_0, output_0_243;
mixer gate_output_0_243(.a(output_1_243), .b(output_1_0), .y(output_0_243));
wire output_2_243, output_2_0, output_1_243;
mixer gate_output_1_243(.a(output_2_243), .b(output_2_0), .y(output_1_243));
wire output_3_243, output_3_0, output_2_243;
mixer gate_output_2_243(.a(output_3_243), .b(output_3_0), .y(output_2_243));
wire output_4_243, output_4_0, output_3_243;
mixer gate_output_3_243(.a(output_4_243), .b(output_4_0), .y(output_3_243));
wire output_1_244, output_1_1, output_0_244;
mixer gate_output_0_244(.a(output_1_244), .b(output_1_1), .y(output_0_244));
wire output_2_244, output_2_1, output_1_244;
mixer gate_output_1_244(.a(output_2_244), .b(output_2_1), .y(output_1_244));
wire output_3_244, output_3_1, output_2_244;
mixer gate_output_2_244(.a(output_3_244), .b(output_3_1), .y(output_2_244));
wire output_4_244, output_4_1, output_3_244;
mixer gate_output_3_244(.a(output_4_244), .b(output_4_1), .y(output_3_244));
wire output_1_245, output_1_2, output_0_245;
mixer gate_output_0_245(.a(output_1_245), .b(output_1_2), .y(output_0_245));
wire output_2_245, output_2_2, output_1_245;
mixer gate_output_1_245(.a(output_2_245), .b(output_2_2), .y(output_1_245));
wire output_3_245, output_3_2, output_2_245;
mixer gate_output_2_245(.a(output_3_245), .b(output_3_2), .y(output_2_245));
wire output_4_245, output_4_2, output_3_245;
mixer gate_output_3_245(.a(output_4_245), .b(output_4_2), .y(output_3_245));
wire output_1_246, output_1_3, output_0_246;
mixer gate_output_0_246(.a(output_1_246), .b(output_1_3), .y(output_0_246));
wire output_2_246, output_2_3, output_1_246;
mixer gate_output_1_246(.a(output_2_246), .b(output_2_3), .y(output_1_246));
wire output_3_246, output_3_3, output_2_246;
mixer gate_output_2_246(.a(output_3_246), .b(output_3_3), .y(output_2_246));
wire output_4_246, output_4_3, output_3_246;
mixer gate_output_3_246(.a(output_4_246), .b(output_4_3), .y(output_3_246));
wire output_1_247, output_1_0, output_0_247;
mixer gate_output_0_247(.a(output_1_247), .b(output_1_0), .y(output_0_247));
wire output_2_247, output_2_0, output_1_247;
mixer gate_output_1_247(.a(output_2_247), .b(output_2_0), .y(output_1_247));
wire output_3_247, output_3_0, output_2_247;
mixer gate_output_2_247(.a(output_3_247), .b(output_3_0), .y(output_2_247));
wire output_4_247, output_4_0, output_3_247;
mixer gate_output_3_247(.a(output_4_247), .b(output_4_0), .y(output_3_247));
wire output_1_248, output_1_1, output_0_248;
mixer gate_output_0_248(.a(output_1_248), .b(output_1_1), .y(output_0_248));
wire output_2_248, output_2_1, output_1_248;
mixer gate_output_1_248(.a(output_2_248), .b(output_2_1), .y(output_1_248));
wire output_3_248, output_3_1, output_2_248;
mixer gate_output_2_248(.a(output_3_248), .b(output_3_1), .y(output_2_248));
wire output_4_248, output_4_1, output_3_248;
mixer gate_output_3_248(.a(output_4_248), .b(output_4_1), .y(output_3_248));
wire output_1_249, output_1_2, output_0_249;
mixer gate_output_0_249(.a(output_1_249), .b(output_1_2), .y(output_0_249));
wire output_2_249, output_2_2, output_1_249;
mixer gate_output_1_249(.a(output_2_249), .b(output_2_2), .y(output_1_249));
wire output_3_249, output_3_2, output_2_249;
mixer gate_output_2_249(.a(output_3_249), .b(output_3_2), .y(output_2_249));
wire output_4_249, output_4_2, output_3_249;
mixer gate_output_3_249(.a(output_4_249), .b(output_4_2), .y(output_3_249));
wire output_1_250, output_1_3, output_0_250;
mixer gate_output_0_250(.a(output_1_250), .b(output_1_3), .y(output_0_250));
wire output_2_250, output_2_3, output_1_250;
mixer gate_output_1_250(.a(output_2_250), .b(output_2_3), .y(output_1_250));
wire output_3_250, output_3_3, output_2_250;
mixer gate_output_2_250(.a(output_3_250), .b(output_3_3), .y(output_2_250));
wire output_4_250, output_4_3, output_3_250;
mixer gate_output_3_250(.a(output_4_250), .b(output_4_3), .y(output_3_250));
wire output_1_251, output_1_0, output_0_251;
mixer gate_output_0_251(.a(output_1_251), .b(output_1_0), .y(output_0_251));
wire output_2_251, output_2_0, output_1_251;
mixer gate_output_1_251(.a(output_2_251), .b(output_2_0), .y(output_1_251));
wire output_3_251, output_3_0, output_2_251;
mixer gate_output_2_251(.a(output_3_251), .b(output_3_0), .y(output_2_251));
wire output_4_251, output_4_0, output_3_251;
mixer gate_output_3_251(.a(output_4_251), .b(output_4_0), .y(output_3_251));
wire output_1_252, output_1_1, output_0_252;
mixer gate_output_0_252(.a(output_1_252), .b(output_1_1), .y(output_0_252));
wire output_2_252, output_2_1, output_1_252;
mixer gate_output_1_252(.a(output_2_252), .b(output_2_1), .y(output_1_252));
wire output_3_252, output_3_1, output_2_252;
mixer gate_output_2_252(.a(output_3_252), .b(output_3_1), .y(output_2_252));
wire output_4_252, output_4_1, output_3_252;
mixer gate_output_3_252(.a(output_4_252), .b(output_4_1), .y(output_3_252));
wire output_1_253, output_1_2, output_0_253;
mixer gate_output_0_253(.a(output_1_253), .b(output_1_2), .y(output_0_253));
wire output_2_253, output_2_2, output_1_253;
mixer gate_output_1_253(.a(output_2_253), .b(output_2_2), .y(output_1_253));
wire output_3_253, output_3_2, output_2_253;
mixer gate_output_2_253(.a(output_3_253), .b(output_3_2), .y(output_2_253));
wire output_4_253, output_4_2, output_3_253;
mixer gate_output_3_253(.a(output_4_253), .b(output_4_2), .y(output_3_253));
wire output_1_254, output_1_3, output_0_254;
mixer gate_output_0_254(.a(output_1_254), .b(output_1_3), .y(output_0_254));
wire output_2_254, output_2_3, output_1_254;
mixer gate_output_1_254(.a(output_2_254), .b(output_2_3), .y(output_1_254));
wire output_3_254, output_3_3, output_2_254;
mixer gate_output_2_254(.a(output_3_254), .b(output_3_3), .y(output_2_254));
wire output_4_254, output_4_3, output_3_254;
mixer gate_output_3_254(.a(output_4_254), .b(output_4_3), .y(output_3_254));
wire output_1_255, output_1_0, output_0_255;
mixer gate_output_0_255(.a(output_1_255), .b(output_1_0), .y(output_0_255));
wire output_2_255, output_2_0, output_1_255;
mixer gate_output_1_255(.a(output_2_255), .b(output_2_0), .y(output_1_255));
wire output_3_255, output_3_0, output_2_255;
mixer gate_output_2_255(.a(output_3_255), .b(output_3_0), .y(output_2_255));
wire output_4_255, output_4_0, output_3_255;
mixer gate_output_3_255(.a(output_4_255), .b(output_4_0), .y(output_3_255));
assign output_0 = output_0_0;
wire output_0_256;
assign output_0_256 = input_0;
assign output_1 = output_1_0;
wire output_1_256;
assign output_1_256 = input_1;
assign output_2 = output_2_0;
wire output_2_256;
assign output_2_256 = input_2;
assign output_3 = output_3_0;
wire output_3_256;
assign output_3_256 = input_3;
endmodule
