module fanout2_braid_3_1024 (
output output_0,output output_1,output output_2,input input_0,input input_1,input input_2
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_1_2, output_1_0, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_0), .y(output_0_2));
wire output_2_2, output_2_0, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_0), .y(output_1_2));
wire output_3_2, output_3_0, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_0), .y(output_2_2));
wire output_1_3, output_1_1, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_1), .y(output_0_3));
wire output_2_3, output_2_1, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_1), .y(output_1_3));
wire output_3_3, output_3_1, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_1), .y(output_2_3));
wire output_1_4, output_1_2, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_2), .y(output_0_4));
wire output_2_4, output_2_2, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_2), .y(output_1_4));
wire output_3_4, output_3_2, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_2), .y(output_2_4));
wire output_1_5, output_1_0, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_0), .y(output_0_5));
wire output_2_5, output_2_0, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_0), .y(output_1_5));
wire output_3_5, output_3_0, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_0), .y(output_2_5));
wire output_1_6, output_1_1, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_1), .y(output_0_6));
wire output_2_6, output_2_1, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_1), .y(output_1_6));
wire output_3_6, output_3_1, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_1), .y(output_2_6));
wire output_1_7, output_1_2, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_2), .y(output_0_7));
wire output_2_7, output_2_2, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_2), .y(output_1_7));
wire output_3_7, output_3_2, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_2), .y(output_2_7));
wire output_1_8, output_1_0, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_0), .y(output_0_8));
wire output_2_8, output_2_0, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_0), .y(output_1_8));
wire output_3_8, output_3_0, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_0), .y(output_2_8));
wire output_1_9, output_1_1, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_1), .y(output_0_9));
wire output_2_9, output_2_1, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_1), .y(output_1_9));
wire output_3_9, output_3_1, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_1), .y(output_2_9));
wire output_1_10, output_1_2, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_2), .y(output_0_10));
wire output_2_10, output_2_2, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_2), .y(output_1_10));
wire output_3_10, output_3_2, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_2), .y(output_2_10));
wire output_1_11, output_1_0, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_0), .y(output_0_11));
wire output_2_11, output_2_0, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_0), .y(output_1_11));
wire output_3_11, output_3_0, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_0), .y(output_2_11));
wire output_1_12, output_1_1, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_1), .y(output_0_12));
wire output_2_12, output_2_1, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_1), .y(output_1_12));
wire output_3_12, output_3_1, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_1), .y(output_2_12));
wire output_1_13, output_1_2, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_2), .y(output_0_13));
wire output_2_13, output_2_2, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_2), .y(output_1_13));
wire output_3_13, output_3_2, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_2), .y(output_2_13));
wire output_1_14, output_1_0, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_0), .y(output_0_14));
wire output_2_14, output_2_0, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_0), .y(output_1_14));
wire output_3_14, output_3_0, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_0), .y(output_2_14));
wire output_1_15, output_1_1, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_1), .y(output_0_15));
wire output_2_15, output_2_1, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_1), .y(output_1_15));
wire output_3_15, output_3_1, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_1), .y(output_2_15));
wire output_1_16, output_1_2, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_2), .y(output_0_16));
wire output_2_16, output_2_2, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_2), .y(output_1_16));
wire output_3_16, output_3_2, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_2), .y(output_2_16));
wire output_1_17, output_1_0, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_0), .y(output_0_17));
wire output_2_17, output_2_0, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_0), .y(output_1_17));
wire output_3_17, output_3_0, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_0), .y(output_2_17));
wire output_1_18, output_1_1, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_1), .y(output_0_18));
wire output_2_18, output_2_1, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_1), .y(output_1_18));
wire output_3_18, output_3_1, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_1), .y(output_2_18));
wire output_1_19, output_1_2, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_2), .y(output_0_19));
wire output_2_19, output_2_2, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_2), .y(output_1_19));
wire output_3_19, output_3_2, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_2), .y(output_2_19));
wire output_1_20, output_1_0, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_0), .y(output_0_20));
wire output_2_20, output_2_0, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_0), .y(output_1_20));
wire output_3_20, output_3_0, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_0), .y(output_2_20));
wire output_1_21, output_1_1, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_1), .y(output_0_21));
wire output_2_21, output_2_1, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_1), .y(output_1_21));
wire output_3_21, output_3_1, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_1), .y(output_2_21));
wire output_1_22, output_1_2, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_2), .y(output_0_22));
wire output_2_22, output_2_2, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_2), .y(output_1_22));
wire output_3_22, output_3_2, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_2), .y(output_2_22));
wire output_1_23, output_1_0, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_0), .y(output_0_23));
wire output_2_23, output_2_0, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_0), .y(output_1_23));
wire output_3_23, output_3_0, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_0), .y(output_2_23));
wire output_1_24, output_1_1, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_1), .y(output_0_24));
wire output_2_24, output_2_1, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_1), .y(output_1_24));
wire output_3_24, output_3_1, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_1), .y(output_2_24));
wire output_1_25, output_1_2, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_2), .y(output_0_25));
wire output_2_25, output_2_2, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_2), .y(output_1_25));
wire output_3_25, output_3_2, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_2), .y(output_2_25));
wire output_1_26, output_1_0, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_0), .y(output_0_26));
wire output_2_26, output_2_0, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_0), .y(output_1_26));
wire output_3_26, output_3_0, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_0), .y(output_2_26));
wire output_1_27, output_1_1, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_1), .y(output_0_27));
wire output_2_27, output_2_1, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_1), .y(output_1_27));
wire output_3_27, output_3_1, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_1), .y(output_2_27));
wire output_1_28, output_1_2, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_2), .y(output_0_28));
wire output_2_28, output_2_2, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_2), .y(output_1_28));
wire output_3_28, output_3_2, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_2), .y(output_2_28));
wire output_1_29, output_1_0, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_0), .y(output_0_29));
wire output_2_29, output_2_0, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_0), .y(output_1_29));
wire output_3_29, output_3_0, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_0), .y(output_2_29));
wire output_1_30, output_1_1, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_1), .y(output_0_30));
wire output_2_30, output_2_1, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_1), .y(output_1_30));
wire output_3_30, output_3_1, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_1), .y(output_2_30));
wire output_1_31, output_1_2, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_2), .y(output_0_31));
wire output_2_31, output_2_2, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_2), .y(output_1_31));
wire output_3_31, output_3_2, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_2), .y(output_2_31));
wire output_1_32, output_1_0, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_0), .y(output_0_32));
wire output_2_32, output_2_0, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_0), .y(output_1_32));
wire output_3_32, output_3_0, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_0), .y(output_2_32));
wire output_1_33, output_1_1, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_1), .y(output_0_33));
wire output_2_33, output_2_1, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_1), .y(output_1_33));
wire output_3_33, output_3_1, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_1), .y(output_2_33));
wire output_1_34, output_1_2, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_2), .y(output_0_34));
wire output_2_34, output_2_2, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_2), .y(output_1_34));
wire output_3_34, output_3_2, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_2), .y(output_2_34));
wire output_1_35, output_1_0, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_0), .y(output_0_35));
wire output_2_35, output_2_0, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_0), .y(output_1_35));
wire output_3_35, output_3_0, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_0), .y(output_2_35));
wire output_1_36, output_1_1, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_1), .y(output_0_36));
wire output_2_36, output_2_1, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_1), .y(output_1_36));
wire output_3_36, output_3_1, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_1), .y(output_2_36));
wire output_1_37, output_1_2, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_2), .y(output_0_37));
wire output_2_37, output_2_2, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_2), .y(output_1_37));
wire output_3_37, output_3_2, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_2), .y(output_2_37));
wire output_1_38, output_1_0, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_0), .y(output_0_38));
wire output_2_38, output_2_0, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_0), .y(output_1_38));
wire output_3_38, output_3_0, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_0), .y(output_2_38));
wire output_1_39, output_1_1, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_1), .y(output_0_39));
wire output_2_39, output_2_1, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_1), .y(output_1_39));
wire output_3_39, output_3_1, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_1), .y(output_2_39));
wire output_1_40, output_1_2, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_2), .y(output_0_40));
wire output_2_40, output_2_2, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_2), .y(output_1_40));
wire output_3_40, output_3_2, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_2), .y(output_2_40));
wire output_1_41, output_1_0, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_0), .y(output_0_41));
wire output_2_41, output_2_0, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_0), .y(output_1_41));
wire output_3_41, output_3_0, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_0), .y(output_2_41));
wire output_1_42, output_1_1, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_1), .y(output_0_42));
wire output_2_42, output_2_1, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_1), .y(output_1_42));
wire output_3_42, output_3_1, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_1), .y(output_2_42));
wire output_1_43, output_1_2, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_2), .y(output_0_43));
wire output_2_43, output_2_2, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_2), .y(output_1_43));
wire output_3_43, output_3_2, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_2), .y(output_2_43));
wire output_1_44, output_1_0, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_0), .y(output_0_44));
wire output_2_44, output_2_0, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_0), .y(output_1_44));
wire output_3_44, output_3_0, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_0), .y(output_2_44));
wire output_1_45, output_1_1, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_1), .y(output_0_45));
wire output_2_45, output_2_1, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_1), .y(output_1_45));
wire output_3_45, output_3_1, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_1), .y(output_2_45));
wire output_1_46, output_1_2, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_2), .y(output_0_46));
wire output_2_46, output_2_2, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_2), .y(output_1_46));
wire output_3_46, output_3_2, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_2), .y(output_2_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_1_50, output_1_0, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_0), .y(output_0_50));
wire output_2_50, output_2_0, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_0), .y(output_1_50));
wire output_3_50, output_3_0, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_0), .y(output_2_50));
wire output_1_51, output_1_1, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_1), .y(output_0_51));
wire output_2_51, output_2_1, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_1), .y(output_1_51));
wire output_3_51, output_3_1, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_1), .y(output_2_51));
wire output_1_52, output_1_2, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_2), .y(output_0_52));
wire output_2_52, output_2_2, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_2), .y(output_1_52));
wire output_3_52, output_3_2, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_2), .y(output_2_52));
wire output_1_53, output_1_0, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_0), .y(output_0_53));
wire output_2_53, output_2_0, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_0), .y(output_1_53));
wire output_3_53, output_3_0, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_0), .y(output_2_53));
wire output_1_54, output_1_1, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_1), .y(output_0_54));
wire output_2_54, output_2_1, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_1), .y(output_1_54));
wire output_3_54, output_3_1, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_1), .y(output_2_54));
wire output_1_55, output_1_2, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_2), .y(output_0_55));
wire output_2_55, output_2_2, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_2), .y(output_1_55));
wire output_3_55, output_3_2, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_2), .y(output_2_55));
wire output_1_56, output_1_0, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_0), .y(output_0_56));
wire output_2_56, output_2_0, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_0), .y(output_1_56));
wire output_3_56, output_3_0, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_0), .y(output_2_56));
wire output_1_57, output_1_1, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_1), .y(output_0_57));
wire output_2_57, output_2_1, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_1), .y(output_1_57));
wire output_3_57, output_3_1, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_1), .y(output_2_57));
wire output_1_58, output_1_2, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_2), .y(output_0_58));
wire output_2_58, output_2_2, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_2), .y(output_1_58));
wire output_3_58, output_3_2, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_2), .y(output_2_58));
wire output_1_59, output_1_0, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_0), .y(output_0_59));
wire output_2_59, output_2_0, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_0), .y(output_1_59));
wire output_3_59, output_3_0, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_0), .y(output_2_59));
wire output_1_60, output_1_1, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_1), .y(output_0_60));
wire output_2_60, output_2_1, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_1), .y(output_1_60));
wire output_3_60, output_3_1, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_1), .y(output_2_60));
wire output_1_61, output_1_2, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_2), .y(output_0_61));
wire output_2_61, output_2_2, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_2), .y(output_1_61));
wire output_3_61, output_3_2, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_2), .y(output_2_61));
wire output_1_62, output_1_0, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_0), .y(output_0_62));
wire output_2_62, output_2_0, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_0), .y(output_1_62));
wire output_3_62, output_3_0, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_0), .y(output_2_62));
wire output_1_63, output_1_1, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_1), .y(output_0_63));
wire output_2_63, output_2_1, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_1), .y(output_1_63));
wire output_3_63, output_3_1, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_1), .y(output_2_63));
wire output_1_64, output_1_2, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_2), .y(output_0_64));
wire output_2_64, output_2_2, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_2), .y(output_1_64));
wire output_3_64, output_3_2, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_2), .y(output_2_64));
wire output_1_65, output_1_0, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_0), .y(output_0_65));
wire output_2_65, output_2_0, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_0), .y(output_1_65));
wire output_3_65, output_3_0, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_0), .y(output_2_65));
wire output_1_66, output_1_1, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_1), .y(output_0_66));
wire output_2_66, output_2_1, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_1), .y(output_1_66));
wire output_3_66, output_3_1, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_1), .y(output_2_66));
wire output_1_67, output_1_2, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_2), .y(output_0_67));
wire output_2_67, output_2_2, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_2), .y(output_1_67));
wire output_3_67, output_3_2, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_2), .y(output_2_67));
wire output_1_68, output_1_0, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_0), .y(output_0_68));
wire output_2_68, output_2_0, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_0), .y(output_1_68));
wire output_3_68, output_3_0, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_0), .y(output_2_68));
wire output_1_69, output_1_1, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_1), .y(output_0_69));
wire output_2_69, output_2_1, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_1), .y(output_1_69));
wire output_3_69, output_3_1, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_1), .y(output_2_69));
wire output_1_70, output_1_2, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_2), .y(output_0_70));
wire output_2_70, output_2_2, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_2), .y(output_1_70));
wire output_3_70, output_3_2, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_2), .y(output_2_70));
wire output_1_71, output_1_0, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_0), .y(output_0_71));
wire output_2_71, output_2_0, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_0), .y(output_1_71));
wire output_3_71, output_3_0, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_0), .y(output_2_71));
wire output_1_72, output_1_1, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_1), .y(output_0_72));
wire output_2_72, output_2_1, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_1), .y(output_1_72));
wire output_3_72, output_3_1, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_1), .y(output_2_72));
wire output_1_73, output_1_2, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_2), .y(output_0_73));
wire output_2_73, output_2_2, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_2), .y(output_1_73));
wire output_3_73, output_3_2, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_2), .y(output_2_73));
wire output_1_74, output_1_0, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_0), .y(output_0_74));
wire output_2_74, output_2_0, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_0), .y(output_1_74));
wire output_3_74, output_3_0, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_0), .y(output_2_74));
wire output_1_75, output_1_1, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_1), .y(output_0_75));
wire output_2_75, output_2_1, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_1), .y(output_1_75));
wire output_3_75, output_3_1, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_1), .y(output_2_75));
wire output_1_76, output_1_2, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_2), .y(output_0_76));
wire output_2_76, output_2_2, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_2), .y(output_1_76));
wire output_3_76, output_3_2, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_2), .y(output_2_76));
wire output_1_77, output_1_0, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_0), .y(output_0_77));
wire output_2_77, output_2_0, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_0), .y(output_1_77));
wire output_3_77, output_3_0, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_0), .y(output_2_77));
wire output_1_78, output_1_1, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_1), .y(output_0_78));
wire output_2_78, output_2_1, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_1), .y(output_1_78));
wire output_3_78, output_3_1, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_1), .y(output_2_78));
wire output_1_79, output_1_2, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_2), .y(output_0_79));
wire output_2_79, output_2_2, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_2), .y(output_1_79));
wire output_3_79, output_3_2, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_2), .y(output_2_79));
wire output_1_80, output_1_0, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_0), .y(output_0_80));
wire output_2_80, output_2_0, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_0), .y(output_1_80));
wire output_3_80, output_3_0, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_0), .y(output_2_80));
wire output_1_81, output_1_1, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_1), .y(output_0_81));
wire output_2_81, output_2_1, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_1), .y(output_1_81));
wire output_3_81, output_3_1, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_1), .y(output_2_81));
wire output_1_82, output_1_2, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_2), .y(output_0_82));
wire output_2_82, output_2_2, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_2), .y(output_1_82));
wire output_3_82, output_3_2, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_2), .y(output_2_82));
wire output_1_83, output_1_0, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_0), .y(output_0_83));
wire output_2_83, output_2_0, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_0), .y(output_1_83));
wire output_3_83, output_3_0, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_0), .y(output_2_83));
wire output_1_84, output_1_1, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_1), .y(output_0_84));
wire output_2_84, output_2_1, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_1), .y(output_1_84));
wire output_3_84, output_3_1, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_1), .y(output_2_84));
wire output_1_85, output_1_2, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_2), .y(output_0_85));
wire output_2_85, output_2_2, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_2), .y(output_1_85));
wire output_3_85, output_3_2, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_2), .y(output_2_85));
wire output_1_86, output_1_0, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_0), .y(output_0_86));
wire output_2_86, output_2_0, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_0), .y(output_1_86));
wire output_3_86, output_3_0, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_0), .y(output_2_86));
wire output_1_87, output_1_1, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_1), .y(output_0_87));
wire output_2_87, output_2_1, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_1), .y(output_1_87));
wire output_3_87, output_3_1, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_1), .y(output_2_87));
wire output_1_88, output_1_2, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_2), .y(output_0_88));
wire output_2_88, output_2_2, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_2), .y(output_1_88));
wire output_3_88, output_3_2, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_2), .y(output_2_88));
wire output_1_89, output_1_0, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_0), .y(output_0_89));
wire output_2_89, output_2_0, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_0), .y(output_1_89));
wire output_3_89, output_3_0, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_0), .y(output_2_89));
wire output_1_90, output_1_1, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_1), .y(output_0_90));
wire output_2_90, output_2_1, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_1), .y(output_1_90));
wire output_3_90, output_3_1, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_1), .y(output_2_90));
wire output_1_91, output_1_2, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_2), .y(output_0_91));
wire output_2_91, output_2_2, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_2), .y(output_1_91));
wire output_3_91, output_3_2, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_2), .y(output_2_91));
wire output_1_92, output_1_0, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_0), .y(output_0_92));
wire output_2_92, output_2_0, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_0), .y(output_1_92));
wire output_3_92, output_3_0, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_0), .y(output_2_92));
wire output_1_93, output_1_1, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_1), .y(output_0_93));
wire output_2_93, output_2_1, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_1), .y(output_1_93));
wire output_3_93, output_3_1, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_1), .y(output_2_93));
wire output_1_94, output_1_2, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_2), .y(output_0_94));
wire output_2_94, output_2_2, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_2), .y(output_1_94));
wire output_3_94, output_3_2, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_2), .y(output_2_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_1_96, output_1_1, output_0_96;
mixer gate_output_0_96(.a(output_1_96), .b(output_1_1), .y(output_0_96));
wire output_2_96, output_2_1, output_1_96;
mixer gate_output_1_96(.a(output_2_96), .b(output_2_1), .y(output_1_96));
wire output_3_96, output_3_1, output_2_96;
mixer gate_output_2_96(.a(output_3_96), .b(output_3_1), .y(output_2_96));
wire output_1_97, output_1_2, output_0_97;
mixer gate_output_0_97(.a(output_1_97), .b(output_1_2), .y(output_0_97));
wire output_2_97, output_2_2, output_1_97;
mixer gate_output_1_97(.a(output_2_97), .b(output_2_2), .y(output_1_97));
wire output_3_97, output_3_2, output_2_97;
mixer gate_output_2_97(.a(output_3_97), .b(output_3_2), .y(output_2_97));
wire output_1_98, output_1_0, output_0_98;
mixer gate_output_0_98(.a(output_1_98), .b(output_1_0), .y(output_0_98));
wire output_2_98, output_2_0, output_1_98;
mixer gate_output_1_98(.a(output_2_98), .b(output_2_0), .y(output_1_98));
wire output_3_98, output_3_0, output_2_98;
mixer gate_output_2_98(.a(output_3_98), .b(output_3_0), .y(output_2_98));
wire output_1_99, output_1_1, output_0_99;
mixer gate_output_0_99(.a(output_1_99), .b(output_1_1), .y(output_0_99));
wire output_2_99, output_2_1, output_1_99;
mixer gate_output_1_99(.a(output_2_99), .b(output_2_1), .y(output_1_99));
wire output_3_99, output_3_1, output_2_99;
mixer gate_output_2_99(.a(output_3_99), .b(output_3_1), .y(output_2_99));
wire output_1_100, output_1_2, output_0_100;
mixer gate_output_0_100(.a(output_1_100), .b(output_1_2), .y(output_0_100));
wire output_2_100, output_2_2, output_1_100;
mixer gate_output_1_100(.a(output_2_100), .b(output_2_2), .y(output_1_100));
wire output_3_100, output_3_2, output_2_100;
mixer gate_output_2_100(.a(output_3_100), .b(output_3_2), .y(output_2_100));
wire output_1_101, output_1_0, output_0_101;
mixer gate_output_0_101(.a(output_1_101), .b(output_1_0), .y(output_0_101));
wire output_2_101, output_2_0, output_1_101;
mixer gate_output_1_101(.a(output_2_101), .b(output_2_0), .y(output_1_101));
wire output_3_101, output_3_0, output_2_101;
mixer gate_output_2_101(.a(output_3_101), .b(output_3_0), .y(output_2_101));
wire output_1_102, output_1_1, output_0_102;
mixer gate_output_0_102(.a(output_1_102), .b(output_1_1), .y(output_0_102));
wire output_2_102, output_2_1, output_1_102;
mixer gate_output_1_102(.a(output_2_102), .b(output_2_1), .y(output_1_102));
wire output_3_102, output_3_1, output_2_102;
mixer gate_output_2_102(.a(output_3_102), .b(output_3_1), .y(output_2_102));
wire output_1_103, output_1_2, output_0_103;
mixer gate_output_0_103(.a(output_1_103), .b(output_1_2), .y(output_0_103));
wire output_2_103, output_2_2, output_1_103;
mixer gate_output_1_103(.a(output_2_103), .b(output_2_2), .y(output_1_103));
wire output_3_103, output_3_2, output_2_103;
mixer gate_output_2_103(.a(output_3_103), .b(output_3_2), .y(output_2_103));
wire output_1_104, output_1_0, output_0_104;
mixer gate_output_0_104(.a(output_1_104), .b(output_1_0), .y(output_0_104));
wire output_2_104, output_2_0, output_1_104;
mixer gate_output_1_104(.a(output_2_104), .b(output_2_0), .y(output_1_104));
wire output_3_104, output_3_0, output_2_104;
mixer gate_output_2_104(.a(output_3_104), .b(output_3_0), .y(output_2_104));
wire output_1_105, output_1_1, output_0_105;
mixer gate_output_0_105(.a(output_1_105), .b(output_1_1), .y(output_0_105));
wire output_2_105, output_2_1, output_1_105;
mixer gate_output_1_105(.a(output_2_105), .b(output_2_1), .y(output_1_105));
wire output_3_105, output_3_1, output_2_105;
mixer gate_output_2_105(.a(output_3_105), .b(output_3_1), .y(output_2_105));
wire output_1_106, output_1_2, output_0_106;
mixer gate_output_0_106(.a(output_1_106), .b(output_1_2), .y(output_0_106));
wire output_2_106, output_2_2, output_1_106;
mixer gate_output_1_106(.a(output_2_106), .b(output_2_2), .y(output_1_106));
wire output_3_106, output_3_2, output_2_106;
mixer gate_output_2_106(.a(output_3_106), .b(output_3_2), .y(output_2_106));
wire output_1_107, output_1_0, output_0_107;
mixer gate_output_0_107(.a(output_1_107), .b(output_1_0), .y(output_0_107));
wire output_2_107, output_2_0, output_1_107;
mixer gate_output_1_107(.a(output_2_107), .b(output_2_0), .y(output_1_107));
wire output_3_107, output_3_0, output_2_107;
mixer gate_output_2_107(.a(output_3_107), .b(output_3_0), .y(output_2_107));
wire output_1_108, output_1_1, output_0_108;
mixer gate_output_0_108(.a(output_1_108), .b(output_1_1), .y(output_0_108));
wire output_2_108, output_2_1, output_1_108;
mixer gate_output_1_108(.a(output_2_108), .b(output_2_1), .y(output_1_108));
wire output_3_108, output_3_1, output_2_108;
mixer gate_output_2_108(.a(output_3_108), .b(output_3_1), .y(output_2_108));
wire output_1_109, output_1_2, output_0_109;
mixer gate_output_0_109(.a(output_1_109), .b(output_1_2), .y(output_0_109));
wire output_2_109, output_2_2, output_1_109;
mixer gate_output_1_109(.a(output_2_109), .b(output_2_2), .y(output_1_109));
wire output_3_109, output_3_2, output_2_109;
mixer gate_output_2_109(.a(output_3_109), .b(output_3_2), .y(output_2_109));
wire output_1_110, output_1_0, output_0_110;
mixer gate_output_0_110(.a(output_1_110), .b(output_1_0), .y(output_0_110));
wire output_2_110, output_2_0, output_1_110;
mixer gate_output_1_110(.a(output_2_110), .b(output_2_0), .y(output_1_110));
wire output_3_110, output_3_0, output_2_110;
mixer gate_output_2_110(.a(output_3_110), .b(output_3_0), .y(output_2_110));
wire output_1_111, output_1_1, output_0_111;
mixer gate_output_0_111(.a(output_1_111), .b(output_1_1), .y(output_0_111));
wire output_2_111, output_2_1, output_1_111;
mixer gate_output_1_111(.a(output_2_111), .b(output_2_1), .y(output_1_111));
wire output_3_111, output_3_1, output_2_111;
mixer gate_output_2_111(.a(output_3_111), .b(output_3_1), .y(output_2_111));
wire output_1_112, output_1_2, output_0_112;
mixer gate_output_0_112(.a(output_1_112), .b(output_1_2), .y(output_0_112));
wire output_2_112, output_2_2, output_1_112;
mixer gate_output_1_112(.a(output_2_112), .b(output_2_2), .y(output_1_112));
wire output_3_112, output_3_2, output_2_112;
mixer gate_output_2_112(.a(output_3_112), .b(output_3_2), .y(output_2_112));
wire output_1_113, output_1_0, output_0_113;
mixer gate_output_0_113(.a(output_1_113), .b(output_1_0), .y(output_0_113));
wire output_2_113, output_2_0, output_1_113;
mixer gate_output_1_113(.a(output_2_113), .b(output_2_0), .y(output_1_113));
wire output_3_113, output_3_0, output_2_113;
mixer gate_output_2_113(.a(output_3_113), .b(output_3_0), .y(output_2_113));
wire output_1_114, output_1_1, output_0_114;
mixer gate_output_0_114(.a(output_1_114), .b(output_1_1), .y(output_0_114));
wire output_2_114, output_2_1, output_1_114;
mixer gate_output_1_114(.a(output_2_114), .b(output_2_1), .y(output_1_114));
wire output_3_114, output_3_1, output_2_114;
mixer gate_output_2_114(.a(output_3_114), .b(output_3_1), .y(output_2_114));
wire output_1_115, output_1_2, output_0_115;
mixer gate_output_0_115(.a(output_1_115), .b(output_1_2), .y(output_0_115));
wire output_2_115, output_2_2, output_1_115;
mixer gate_output_1_115(.a(output_2_115), .b(output_2_2), .y(output_1_115));
wire output_3_115, output_3_2, output_2_115;
mixer gate_output_2_115(.a(output_3_115), .b(output_3_2), .y(output_2_115));
wire output_1_116, output_1_0, output_0_116;
mixer gate_output_0_116(.a(output_1_116), .b(output_1_0), .y(output_0_116));
wire output_2_116, output_2_0, output_1_116;
mixer gate_output_1_116(.a(output_2_116), .b(output_2_0), .y(output_1_116));
wire output_3_116, output_3_0, output_2_116;
mixer gate_output_2_116(.a(output_3_116), .b(output_3_0), .y(output_2_116));
wire output_1_117, output_1_1, output_0_117;
mixer gate_output_0_117(.a(output_1_117), .b(output_1_1), .y(output_0_117));
wire output_2_117, output_2_1, output_1_117;
mixer gate_output_1_117(.a(output_2_117), .b(output_2_1), .y(output_1_117));
wire output_3_117, output_3_1, output_2_117;
mixer gate_output_2_117(.a(output_3_117), .b(output_3_1), .y(output_2_117));
wire output_1_118, output_1_2, output_0_118;
mixer gate_output_0_118(.a(output_1_118), .b(output_1_2), .y(output_0_118));
wire output_2_118, output_2_2, output_1_118;
mixer gate_output_1_118(.a(output_2_118), .b(output_2_2), .y(output_1_118));
wire output_3_118, output_3_2, output_2_118;
mixer gate_output_2_118(.a(output_3_118), .b(output_3_2), .y(output_2_118));
wire output_1_119, output_1_0, output_0_119;
mixer gate_output_0_119(.a(output_1_119), .b(output_1_0), .y(output_0_119));
wire output_2_119, output_2_0, output_1_119;
mixer gate_output_1_119(.a(output_2_119), .b(output_2_0), .y(output_1_119));
wire output_3_119, output_3_0, output_2_119;
mixer gate_output_2_119(.a(output_3_119), .b(output_3_0), .y(output_2_119));
wire output_1_120, output_1_1, output_0_120;
mixer gate_output_0_120(.a(output_1_120), .b(output_1_1), .y(output_0_120));
wire output_2_120, output_2_1, output_1_120;
mixer gate_output_1_120(.a(output_2_120), .b(output_2_1), .y(output_1_120));
wire output_3_120, output_3_1, output_2_120;
mixer gate_output_2_120(.a(output_3_120), .b(output_3_1), .y(output_2_120));
wire output_1_121, output_1_2, output_0_121;
mixer gate_output_0_121(.a(output_1_121), .b(output_1_2), .y(output_0_121));
wire output_2_121, output_2_2, output_1_121;
mixer gate_output_1_121(.a(output_2_121), .b(output_2_2), .y(output_1_121));
wire output_3_121, output_3_2, output_2_121;
mixer gate_output_2_121(.a(output_3_121), .b(output_3_2), .y(output_2_121));
wire output_1_122, output_1_0, output_0_122;
mixer gate_output_0_122(.a(output_1_122), .b(output_1_0), .y(output_0_122));
wire output_2_122, output_2_0, output_1_122;
mixer gate_output_1_122(.a(output_2_122), .b(output_2_0), .y(output_1_122));
wire output_3_122, output_3_0, output_2_122;
mixer gate_output_2_122(.a(output_3_122), .b(output_3_0), .y(output_2_122));
wire output_1_123, output_1_1, output_0_123;
mixer gate_output_0_123(.a(output_1_123), .b(output_1_1), .y(output_0_123));
wire output_2_123, output_2_1, output_1_123;
mixer gate_output_1_123(.a(output_2_123), .b(output_2_1), .y(output_1_123));
wire output_3_123, output_3_1, output_2_123;
mixer gate_output_2_123(.a(output_3_123), .b(output_3_1), .y(output_2_123));
wire output_1_124, output_1_2, output_0_124;
mixer gate_output_0_124(.a(output_1_124), .b(output_1_2), .y(output_0_124));
wire output_2_124, output_2_2, output_1_124;
mixer gate_output_1_124(.a(output_2_124), .b(output_2_2), .y(output_1_124));
wire output_3_124, output_3_2, output_2_124;
mixer gate_output_2_124(.a(output_3_124), .b(output_3_2), .y(output_2_124));
wire output_1_125, output_1_0, output_0_125;
mixer gate_output_0_125(.a(output_1_125), .b(output_1_0), .y(output_0_125));
wire output_2_125, output_2_0, output_1_125;
mixer gate_output_1_125(.a(output_2_125), .b(output_2_0), .y(output_1_125));
wire output_3_125, output_3_0, output_2_125;
mixer gate_output_2_125(.a(output_3_125), .b(output_3_0), .y(output_2_125));
wire output_1_126, output_1_1, output_0_126;
mixer gate_output_0_126(.a(output_1_126), .b(output_1_1), .y(output_0_126));
wire output_2_126, output_2_1, output_1_126;
mixer gate_output_1_126(.a(output_2_126), .b(output_2_1), .y(output_1_126));
wire output_3_126, output_3_1, output_2_126;
mixer gate_output_2_126(.a(output_3_126), .b(output_3_1), .y(output_2_126));
wire output_1_127, output_1_2, output_0_127;
mixer gate_output_0_127(.a(output_1_127), .b(output_1_2), .y(output_0_127));
wire output_2_127, output_2_2, output_1_127;
mixer gate_output_1_127(.a(output_2_127), .b(output_2_2), .y(output_1_127));
wire output_3_127, output_3_2, output_2_127;
mixer gate_output_2_127(.a(output_3_127), .b(output_3_2), .y(output_2_127));
wire output_1_128, output_1_0, output_0_128;
mixer gate_output_0_128(.a(output_1_128), .b(output_1_0), .y(output_0_128));
wire output_2_128, output_2_0, output_1_128;
mixer gate_output_1_128(.a(output_2_128), .b(output_2_0), .y(output_1_128));
wire output_3_128, output_3_0, output_2_128;
mixer gate_output_2_128(.a(output_3_128), .b(output_3_0), .y(output_2_128));
wire output_1_129, output_1_1, output_0_129;
mixer gate_output_0_129(.a(output_1_129), .b(output_1_1), .y(output_0_129));
wire output_2_129, output_2_1, output_1_129;
mixer gate_output_1_129(.a(output_2_129), .b(output_2_1), .y(output_1_129));
wire output_3_129, output_3_1, output_2_129;
mixer gate_output_2_129(.a(output_3_129), .b(output_3_1), .y(output_2_129));
wire output_1_130, output_1_2, output_0_130;
mixer gate_output_0_130(.a(output_1_130), .b(output_1_2), .y(output_0_130));
wire output_2_130, output_2_2, output_1_130;
mixer gate_output_1_130(.a(output_2_130), .b(output_2_2), .y(output_1_130));
wire output_3_130, output_3_2, output_2_130;
mixer gate_output_2_130(.a(output_3_130), .b(output_3_2), .y(output_2_130));
wire output_1_131, output_1_0, output_0_131;
mixer gate_output_0_131(.a(output_1_131), .b(output_1_0), .y(output_0_131));
wire output_2_131, output_2_0, output_1_131;
mixer gate_output_1_131(.a(output_2_131), .b(output_2_0), .y(output_1_131));
wire output_3_131, output_3_0, output_2_131;
mixer gate_output_2_131(.a(output_3_131), .b(output_3_0), .y(output_2_131));
wire output_1_132, output_1_1, output_0_132;
mixer gate_output_0_132(.a(output_1_132), .b(output_1_1), .y(output_0_132));
wire output_2_132, output_2_1, output_1_132;
mixer gate_output_1_132(.a(output_2_132), .b(output_2_1), .y(output_1_132));
wire output_3_132, output_3_1, output_2_132;
mixer gate_output_2_132(.a(output_3_132), .b(output_3_1), .y(output_2_132));
wire output_1_133, output_1_2, output_0_133;
mixer gate_output_0_133(.a(output_1_133), .b(output_1_2), .y(output_0_133));
wire output_2_133, output_2_2, output_1_133;
mixer gate_output_1_133(.a(output_2_133), .b(output_2_2), .y(output_1_133));
wire output_3_133, output_3_2, output_2_133;
mixer gate_output_2_133(.a(output_3_133), .b(output_3_2), .y(output_2_133));
wire output_1_134, output_1_0, output_0_134;
mixer gate_output_0_134(.a(output_1_134), .b(output_1_0), .y(output_0_134));
wire output_2_134, output_2_0, output_1_134;
mixer gate_output_1_134(.a(output_2_134), .b(output_2_0), .y(output_1_134));
wire output_3_134, output_3_0, output_2_134;
mixer gate_output_2_134(.a(output_3_134), .b(output_3_0), .y(output_2_134));
wire output_1_135, output_1_1, output_0_135;
mixer gate_output_0_135(.a(output_1_135), .b(output_1_1), .y(output_0_135));
wire output_2_135, output_2_1, output_1_135;
mixer gate_output_1_135(.a(output_2_135), .b(output_2_1), .y(output_1_135));
wire output_3_135, output_3_1, output_2_135;
mixer gate_output_2_135(.a(output_3_135), .b(output_3_1), .y(output_2_135));
wire output_1_136, output_1_2, output_0_136;
mixer gate_output_0_136(.a(output_1_136), .b(output_1_2), .y(output_0_136));
wire output_2_136, output_2_2, output_1_136;
mixer gate_output_1_136(.a(output_2_136), .b(output_2_2), .y(output_1_136));
wire output_3_136, output_3_2, output_2_136;
mixer gate_output_2_136(.a(output_3_136), .b(output_3_2), .y(output_2_136));
wire output_1_137, output_1_0, output_0_137;
mixer gate_output_0_137(.a(output_1_137), .b(output_1_0), .y(output_0_137));
wire output_2_137, output_2_0, output_1_137;
mixer gate_output_1_137(.a(output_2_137), .b(output_2_0), .y(output_1_137));
wire output_3_137, output_3_0, output_2_137;
mixer gate_output_2_137(.a(output_3_137), .b(output_3_0), .y(output_2_137));
wire output_1_138, output_1_1, output_0_138;
mixer gate_output_0_138(.a(output_1_138), .b(output_1_1), .y(output_0_138));
wire output_2_138, output_2_1, output_1_138;
mixer gate_output_1_138(.a(output_2_138), .b(output_2_1), .y(output_1_138));
wire output_3_138, output_3_1, output_2_138;
mixer gate_output_2_138(.a(output_3_138), .b(output_3_1), .y(output_2_138));
wire output_1_139, output_1_2, output_0_139;
mixer gate_output_0_139(.a(output_1_139), .b(output_1_2), .y(output_0_139));
wire output_2_139, output_2_2, output_1_139;
mixer gate_output_1_139(.a(output_2_139), .b(output_2_2), .y(output_1_139));
wire output_3_139, output_3_2, output_2_139;
mixer gate_output_2_139(.a(output_3_139), .b(output_3_2), .y(output_2_139));
wire output_1_140, output_1_0, output_0_140;
mixer gate_output_0_140(.a(output_1_140), .b(output_1_0), .y(output_0_140));
wire output_2_140, output_2_0, output_1_140;
mixer gate_output_1_140(.a(output_2_140), .b(output_2_0), .y(output_1_140));
wire output_3_140, output_3_0, output_2_140;
mixer gate_output_2_140(.a(output_3_140), .b(output_3_0), .y(output_2_140));
wire output_1_141, output_1_1, output_0_141;
mixer gate_output_0_141(.a(output_1_141), .b(output_1_1), .y(output_0_141));
wire output_2_141, output_2_1, output_1_141;
mixer gate_output_1_141(.a(output_2_141), .b(output_2_1), .y(output_1_141));
wire output_3_141, output_3_1, output_2_141;
mixer gate_output_2_141(.a(output_3_141), .b(output_3_1), .y(output_2_141));
wire output_1_142, output_1_2, output_0_142;
mixer gate_output_0_142(.a(output_1_142), .b(output_1_2), .y(output_0_142));
wire output_2_142, output_2_2, output_1_142;
mixer gate_output_1_142(.a(output_2_142), .b(output_2_2), .y(output_1_142));
wire output_3_142, output_3_2, output_2_142;
mixer gate_output_2_142(.a(output_3_142), .b(output_3_2), .y(output_2_142));
wire output_1_143, output_1_0, output_0_143;
mixer gate_output_0_143(.a(output_1_143), .b(output_1_0), .y(output_0_143));
wire output_2_143, output_2_0, output_1_143;
mixer gate_output_1_143(.a(output_2_143), .b(output_2_0), .y(output_1_143));
wire output_3_143, output_3_0, output_2_143;
mixer gate_output_2_143(.a(output_3_143), .b(output_3_0), .y(output_2_143));
wire output_1_144, output_1_1, output_0_144;
mixer gate_output_0_144(.a(output_1_144), .b(output_1_1), .y(output_0_144));
wire output_2_144, output_2_1, output_1_144;
mixer gate_output_1_144(.a(output_2_144), .b(output_2_1), .y(output_1_144));
wire output_3_144, output_3_1, output_2_144;
mixer gate_output_2_144(.a(output_3_144), .b(output_3_1), .y(output_2_144));
wire output_1_145, output_1_2, output_0_145;
mixer gate_output_0_145(.a(output_1_145), .b(output_1_2), .y(output_0_145));
wire output_2_145, output_2_2, output_1_145;
mixer gate_output_1_145(.a(output_2_145), .b(output_2_2), .y(output_1_145));
wire output_3_145, output_3_2, output_2_145;
mixer gate_output_2_145(.a(output_3_145), .b(output_3_2), .y(output_2_145));
wire output_1_146, output_1_0, output_0_146;
mixer gate_output_0_146(.a(output_1_146), .b(output_1_0), .y(output_0_146));
wire output_2_146, output_2_0, output_1_146;
mixer gate_output_1_146(.a(output_2_146), .b(output_2_0), .y(output_1_146));
wire output_3_146, output_3_0, output_2_146;
mixer gate_output_2_146(.a(output_3_146), .b(output_3_0), .y(output_2_146));
wire output_1_147, output_1_1, output_0_147;
mixer gate_output_0_147(.a(output_1_147), .b(output_1_1), .y(output_0_147));
wire output_2_147, output_2_1, output_1_147;
mixer gate_output_1_147(.a(output_2_147), .b(output_2_1), .y(output_1_147));
wire output_3_147, output_3_1, output_2_147;
mixer gate_output_2_147(.a(output_3_147), .b(output_3_1), .y(output_2_147));
wire output_1_148, output_1_2, output_0_148;
mixer gate_output_0_148(.a(output_1_148), .b(output_1_2), .y(output_0_148));
wire output_2_148, output_2_2, output_1_148;
mixer gate_output_1_148(.a(output_2_148), .b(output_2_2), .y(output_1_148));
wire output_3_148, output_3_2, output_2_148;
mixer gate_output_2_148(.a(output_3_148), .b(output_3_2), .y(output_2_148));
wire output_1_149, output_1_0, output_0_149;
mixer gate_output_0_149(.a(output_1_149), .b(output_1_0), .y(output_0_149));
wire output_2_149, output_2_0, output_1_149;
mixer gate_output_1_149(.a(output_2_149), .b(output_2_0), .y(output_1_149));
wire output_3_149, output_3_0, output_2_149;
mixer gate_output_2_149(.a(output_3_149), .b(output_3_0), .y(output_2_149));
wire output_1_150, output_1_1, output_0_150;
mixer gate_output_0_150(.a(output_1_150), .b(output_1_1), .y(output_0_150));
wire output_2_150, output_2_1, output_1_150;
mixer gate_output_1_150(.a(output_2_150), .b(output_2_1), .y(output_1_150));
wire output_3_150, output_3_1, output_2_150;
mixer gate_output_2_150(.a(output_3_150), .b(output_3_1), .y(output_2_150));
wire output_1_151, output_1_2, output_0_151;
mixer gate_output_0_151(.a(output_1_151), .b(output_1_2), .y(output_0_151));
wire output_2_151, output_2_2, output_1_151;
mixer gate_output_1_151(.a(output_2_151), .b(output_2_2), .y(output_1_151));
wire output_3_151, output_3_2, output_2_151;
mixer gate_output_2_151(.a(output_3_151), .b(output_3_2), .y(output_2_151));
wire output_1_152, output_1_0, output_0_152;
mixer gate_output_0_152(.a(output_1_152), .b(output_1_0), .y(output_0_152));
wire output_2_152, output_2_0, output_1_152;
mixer gate_output_1_152(.a(output_2_152), .b(output_2_0), .y(output_1_152));
wire output_3_152, output_3_0, output_2_152;
mixer gate_output_2_152(.a(output_3_152), .b(output_3_0), .y(output_2_152));
wire output_1_153, output_1_1, output_0_153;
mixer gate_output_0_153(.a(output_1_153), .b(output_1_1), .y(output_0_153));
wire output_2_153, output_2_1, output_1_153;
mixer gate_output_1_153(.a(output_2_153), .b(output_2_1), .y(output_1_153));
wire output_3_153, output_3_1, output_2_153;
mixer gate_output_2_153(.a(output_3_153), .b(output_3_1), .y(output_2_153));
wire output_1_154, output_1_2, output_0_154;
mixer gate_output_0_154(.a(output_1_154), .b(output_1_2), .y(output_0_154));
wire output_2_154, output_2_2, output_1_154;
mixer gate_output_1_154(.a(output_2_154), .b(output_2_2), .y(output_1_154));
wire output_3_154, output_3_2, output_2_154;
mixer gate_output_2_154(.a(output_3_154), .b(output_3_2), .y(output_2_154));
wire output_1_155, output_1_0, output_0_155;
mixer gate_output_0_155(.a(output_1_155), .b(output_1_0), .y(output_0_155));
wire output_2_155, output_2_0, output_1_155;
mixer gate_output_1_155(.a(output_2_155), .b(output_2_0), .y(output_1_155));
wire output_3_155, output_3_0, output_2_155;
mixer gate_output_2_155(.a(output_3_155), .b(output_3_0), .y(output_2_155));
wire output_1_156, output_1_1, output_0_156;
mixer gate_output_0_156(.a(output_1_156), .b(output_1_1), .y(output_0_156));
wire output_2_156, output_2_1, output_1_156;
mixer gate_output_1_156(.a(output_2_156), .b(output_2_1), .y(output_1_156));
wire output_3_156, output_3_1, output_2_156;
mixer gate_output_2_156(.a(output_3_156), .b(output_3_1), .y(output_2_156));
wire output_1_157, output_1_2, output_0_157;
mixer gate_output_0_157(.a(output_1_157), .b(output_1_2), .y(output_0_157));
wire output_2_157, output_2_2, output_1_157;
mixer gate_output_1_157(.a(output_2_157), .b(output_2_2), .y(output_1_157));
wire output_3_157, output_3_2, output_2_157;
mixer gate_output_2_157(.a(output_3_157), .b(output_3_2), .y(output_2_157));
wire output_1_158, output_1_0, output_0_158;
mixer gate_output_0_158(.a(output_1_158), .b(output_1_0), .y(output_0_158));
wire output_2_158, output_2_0, output_1_158;
mixer gate_output_1_158(.a(output_2_158), .b(output_2_0), .y(output_1_158));
wire output_3_158, output_3_0, output_2_158;
mixer gate_output_2_158(.a(output_3_158), .b(output_3_0), .y(output_2_158));
wire output_1_159, output_1_1, output_0_159;
mixer gate_output_0_159(.a(output_1_159), .b(output_1_1), .y(output_0_159));
wire output_2_159, output_2_1, output_1_159;
mixer gate_output_1_159(.a(output_2_159), .b(output_2_1), .y(output_1_159));
wire output_3_159, output_3_1, output_2_159;
mixer gate_output_2_159(.a(output_3_159), .b(output_3_1), .y(output_2_159));
wire output_1_160, output_1_2, output_0_160;
mixer gate_output_0_160(.a(output_1_160), .b(output_1_2), .y(output_0_160));
wire output_2_160, output_2_2, output_1_160;
mixer gate_output_1_160(.a(output_2_160), .b(output_2_2), .y(output_1_160));
wire output_3_160, output_3_2, output_2_160;
mixer gate_output_2_160(.a(output_3_160), .b(output_3_2), .y(output_2_160));
wire output_1_161, output_1_0, output_0_161;
mixer gate_output_0_161(.a(output_1_161), .b(output_1_0), .y(output_0_161));
wire output_2_161, output_2_0, output_1_161;
mixer gate_output_1_161(.a(output_2_161), .b(output_2_0), .y(output_1_161));
wire output_3_161, output_3_0, output_2_161;
mixer gate_output_2_161(.a(output_3_161), .b(output_3_0), .y(output_2_161));
wire output_1_162, output_1_1, output_0_162;
mixer gate_output_0_162(.a(output_1_162), .b(output_1_1), .y(output_0_162));
wire output_2_162, output_2_1, output_1_162;
mixer gate_output_1_162(.a(output_2_162), .b(output_2_1), .y(output_1_162));
wire output_3_162, output_3_1, output_2_162;
mixer gate_output_2_162(.a(output_3_162), .b(output_3_1), .y(output_2_162));
wire output_1_163, output_1_2, output_0_163;
mixer gate_output_0_163(.a(output_1_163), .b(output_1_2), .y(output_0_163));
wire output_2_163, output_2_2, output_1_163;
mixer gate_output_1_163(.a(output_2_163), .b(output_2_2), .y(output_1_163));
wire output_3_163, output_3_2, output_2_163;
mixer gate_output_2_163(.a(output_3_163), .b(output_3_2), .y(output_2_163));
wire output_1_164, output_1_0, output_0_164;
mixer gate_output_0_164(.a(output_1_164), .b(output_1_0), .y(output_0_164));
wire output_2_164, output_2_0, output_1_164;
mixer gate_output_1_164(.a(output_2_164), .b(output_2_0), .y(output_1_164));
wire output_3_164, output_3_0, output_2_164;
mixer gate_output_2_164(.a(output_3_164), .b(output_3_0), .y(output_2_164));
wire output_1_165, output_1_1, output_0_165;
mixer gate_output_0_165(.a(output_1_165), .b(output_1_1), .y(output_0_165));
wire output_2_165, output_2_1, output_1_165;
mixer gate_output_1_165(.a(output_2_165), .b(output_2_1), .y(output_1_165));
wire output_3_165, output_3_1, output_2_165;
mixer gate_output_2_165(.a(output_3_165), .b(output_3_1), .y(output_2_165));
wire output_1_166, output_1_2, output_0_166;
mixer gate_output_0_166(.a(output_1_166), .b(output_1_2), .y(output_0_166));
wire output_2_166, output_2_2, output_1_166;
mixer gate_output_1_166(.a(output_2_166), .b(output_2_2), .y(output_1_166));
wire output_3_166, output_3_2, output_2_166;
mixer gate_output_2_166(.a(output_3_166), .b(output_3_2), .y(output_2_166));
wire output_1_167, output_1_0, output_0_167;
mixer gate_output_0_167(.a(output_1_167), .b(output_1_0), .y(output_0_167));
wire output_2_167, output_2_0, output_1_167;
mixer gate_output_1_167(.a(output_2_167), .b(output_2_0), .y(output_1_167));
wire output_3_167, output_3_0, output_2_167;
mixer gate_output_2_167(.a(output_3_167), .b(output_3_0), .y(output_2_167));
wire output_1_168, output_1_1, output_0_168;
mixer gate_output_0_168(.a(output_1_168), .b(output_1_1), .y(output_0_168));
wire output_2_168, output_2_1, output_1_168;
mixer gate_output_1_168(.a(output_2_168), .b(output_2_1), .y(output_1_168));
wire output_3_168, output_3_1, output_2_168;
mixer gate_output_2_168(.a(output_3_168), .b(output_3_1), .y(output_2_168));
wire output_1_169, output_1_2, output_0_169;
mixer gate_output_0_169(.a(output_1_169), .b(output_1_2), .y(output_0_169));
wire output_2_169, output_2_2, output_1_169;
mixer gate_output_1_169(.a(output_2_169), .b(output_2_2), .y(output_1_169));
wire output_3_169, output_3_2, output_2_169;
mixer gate_output_2_169(.a(output_3_169), .b(output_3_2), .y(output_2_169));
wire output_1_170, output_1_0, output_0_170;
mixer gate_output_0_170(.a(output_1_170), .b(output_1_0), .y(output_0_170));
wire output_2_170, output_2_0, output_1_170;
mixer gate_output_1_170(.a(output_2_170), .b(output_2_0), .y(output_1_170));
wire output_3_170, output_3_0, output_2_170;
mixer gate_output_2_170(.a(output_3_170), .b(output_3_0), .y(output_2_170));
wire output_1_171, output_1_1, output_0_171;
mixer gate_output_0_171(.a(output_1_171), .b(output_1_1), .y(output_0_171));
wire output_2_171, output_2_1, output_1_171;
mixer gate_output_1_171(.a(output_2_171), .b(output_2_1), .y(output_1_171));
wire output_3_171, output_3_1, output_2_171;
mixer gate_output_2_171(.a(output_3_171), .b(output_3_1), .y(output_2_171));
wire output_1_172, output_1_2, output_0_172;
mixer gate_output_0_172(.a(output_1_172), .b(output_1_2), .y(output_0_172));
wire output_2_172, output_2_2, output_1_172;
mixer gate_output_1_172(.a(output_2_172), .b(output_2_2), .y(output_1_172));
wire output_3_172, output_3_2, output_2_172;
mixer gate_output_2_172(.a(output_3_172), .b(output_3_2), .y(output_2_172));
wire output_1_173, output_1_0, output_0_173;
mixer gate_output_0_173(.a(output_1_173), .b(output_1_0), .y(output_0_173));
wire output_2_173, output_2_0, output_1_173;
mixer gate_output_1_173(.a(output_2_173), .b(output_2_0), .y(output_1_173));
wire output_3_173, output_3_0, output_2_173;
mixer gate_output_2_173(.a(output_3_173), .b(output_3_0), .y(output_2_173));
wire output_1_174, output_1_1, output_0_174;
mixer gate_output_0_174(.a(output_1_174), .b(output_1_1), .y(output_0_174));
wire output_2_174, output_2_1, output_1_174;
mixer gate_output_1_174(.a(output_2_174), .b(output_2_1), .y(output_1_174));
wire output_3_174, output_3_1, output_2_174;
mixer gate_output_2_174(.a(output_3_174), .b(output_3_1), .y(output_2_174));
wire output_1_175, output_1_2, output_0_175;
mixer gate_output_0_175(.a(output_1_175), .b(output_1_2), .y(output_0_175));
wire output_2_175, output_2_2, output_1_175;
mixer gate_output_1_175(.a(output_2_175), .b(output_2_2), .y(output_1_175));
wire output_3_175, output_3_2, output_2_175;
mixer gate_output_2_175(.a(output_3_175), .b(output_3_2), .y(output_2_175));
wire output_1_176, output_1_0, output_0_176;
mixer gate_output_0_176(.a(output_1_176), .b(output_1_0), .y(output_0_176));
wire output_2_176, output_2_0, output_1_176;
mixer gate_output_1_176(.a(output_2_176), .b(output_2_0), .y(output_1_176));
wire output_3_176, output_3_0, output_2_176;
mixer gate_output_2_176(.a(output_3_176), .b(output_3_0), .y(output_2_176));
wire output_1_177, output_1_1, output_0_177;
mixer gate_output_0_177(.a(output_1_177), .b(output_1_1), .y(output_0_177));
wire output_2_177, output_2_1, output_1_177;
mixer gate_output_1_177(.a(output_2_177), .b(output_2_1), .y(output_1_177));
wire output_3_177, output_3_1, output_2_177;
mixer gate_output_2_177(.a(output_3_177), .b(output_3_1), .y(output_2_177));
wire output_1_178, output_1_2, output_0_178;
mixer gate_output_0_178(.a(output_1_178), .b(output_1_2), .y(output_0_178));
wire output_2_178, output_2_2, output_1_178;
mixer gate_output_1_178(.a(output_2_178), .b(output_2_2), .y(output_1_178));
wire output_3_178, output_3_2, output_2_178;
mixer gate_output_2_178(.a(output_3_178), .b(output_3_2), .y(output_2_178));
wire output_1_179, output_1_0, output_0_179;
mixer gate_output_0_179(.a(output_1_179), .b(output_1_0), .y(output_0_179));
wire output_2_179, output_2_0, output_1_179;
mixer gate_output_1_179(.a(output_2_179), .b(output_2_0), .y(output_1_179));
wire output_3_179, output_3_0, output_2_179;
mixer gate_output_2_179(.a(output_3_179), .b(output_3_0), .y(output_2_179));
wire output_1_180, output_1_1, output_0_180;
mixer gate_output_0_180(.a(output_1_180), .b(output_1_1), .y(output_0_180));
wire output_2_180, output_2_1, output_1_180;
mixer gate_output_1_180(.a(output_2_180), .b(output_2_1), .y(output_1_180));
wire output_3_180, output_3_1, output_2_180;
mixer gate_output_2_180(.a(output_3_180), .b(output_3_1), .y(output_2_180));
wire output_1_181, output_1_2, output_0_181;
mixer gate_output_0_181(.a(output_1_181), .b(output_1_2), .y(output_0_181));
wire output_2_181, output_2_2, output_1_181;
mixer gate_output_1_181(.a(output_2_181), .b(output_2_2), .y(output_1_181));
wire output_3_181, output_3_2, output_2_181;
mixer gate_output_2_181(.a(output_3_181), .b(output_3_2), .y(output_2_181));
wire output_1_182, output_1_0, output_0_182;
mixer gate_output_0_182(.a(output_1_182), .b(output_1_0), .y(output_0_182));
wire output_2_182, output_2_0, output_1_182;
mixer gate_output_1_182(.a(output_2_182), .b(output_2_0), .y(output_1_182));
wire output_3_182, output_3_0, output_2_182;
mixer gate_output_2_182(.a(output_3_182), .b(output_3_0), .y(output_2_182));
wire output_1_183, output_1_1, output_0_183;
mixer gate_output_0_183(.a(output_1_183), .b(output_1_1), .y(output_0_183));
wire output_2_183, output_2_1, output_1_183;
mixer gate_output_1_183(.a(output_2_183), .b(output_2_1), .y(output_1_183));
wire output_3_183, output_3_1, output_2_183;
mixer gate_output_2_183(.a(output_3_183), .b(output_3_1), .y(output_2_183));
wire output_1_184, output_1_2, output_0_184;
mixer gate_output_0_184(.a(output_1_184), .b(output_1_2), .y(output_0_184));
wire output_2_184, output_2_2, output_1_184;
mixer gate_output_1_184(.a(output_2_184), .b(output_2_2), .y(output_1_184));
wire output_3_184, output_3_2, output_2_184;
mixer gate_output_2_184(.a(output_3_184), .b(output_3_2), .y(output_2_184));
wire output_1_185, output_1_0, output_0_185;
mixer gate_output_0_185(.a(output_1_185), .b(output_1_0), .y(output_0_185));
wire output_2_185, output_2_0, output_1_185;
mixer gate_output_1_185(.a(output_2_185), .b(output_2_0), .y(output_1_185));
wire output_3_185, output_3_0, output_2_185;
mixer gate_output_2_185(.a(output_3_185), .b(output_3_0), .y(output_2_185));
wire output_1_186, output_1_1, output_0_186;
mixer gate_output_0_186(.a(output_1_186), .b(output_1_1), .y(output_0_186));
wire output_2_186, output_2_1, output_1_186;
mixer gate_output_1_186(.a(output_2_186), .b(output_2_1), .y(output_1_186));
wire output_3_186, output_3_1, output_2_186;
mixer gate_output_2_186(.a(output_3_186), .b(output_3_1), .y(output_2_186));
wire output_1_187, output_1_2, output_0_187;
mixer gate_output_0_187(.a(output_1_187), .b(output_1_2), .y(output_0_187));
wire output_2_187, output_2_2, output_1_187;
mixer gate_output_1_187(.a(output_2_187), .b(output_2_2), .y(output_1_187));
wire output_3_187, output_3_2, output_2_187;
mixer gate_output_2_187(.a(output_3_187), .b(output_3_2), .y(output_2_187));
wire output_1_188, output_1_0, output_0_188;
mixer gate_output_0_188(.a(output_1_188), .b(output_1_0), .y(output_0_188));
wire output_2_188, output_2_0, output_1_188;
mixer gate_output_1_188(.a(output_2_188), .b(output_2_0), .y(output_1_188));
wire output_3_188, output_3_0, output_2_188;
mixer gate_output_2_188(.a(output_3_188), .b(output_3_0), .y(output_2_188));
wire output_1_189, output_1_1, output_0_189;
mixer gate_output_0_189(.a(output_1_189), .b(output_1_1), .y(output_0_189));
wire output_2_189, output_2_1, output_1_189;
mixer gate_output_1_189(.a(output_2_189), .b(output_2_1), .y(output_1_189));
wire output_3_189, output_3_1, output_2_189;
mixer gate_output_2_189(.a(output_3_189), .b(output_3_1), .y(output_2_189));
wire output_1_190, output_1_2, output_0_190;
mixer gate_output_0_190(.a(output_1_190), .b(output_1_2), .y(output_0_190));
wire output_2_190, output_2_2, output_1_190;
mixer gate_output_1_190(.a(output_2_190), .b(output_2_2), .y(output_1_190));
wire output_3_190, output_3_2, output_2_190;
mixer gate_output_2_190(.a(output_3_190), .b(output_3_2), .y(output_2_190));
wire output_1_191, output_1_0, output_0_191;
mixer gate_output_0_191(.a(output_1_191), .b(output_1_0), .y(output_0_191));
wire output_2_191, output_2_0, output_1_191;
mixer gate_output_1_191(.a(output_2_191), .b(output_2_0), .y(output_1_191));
wire output_3_191, output_3_0, output_2_191;
mixer gate_output_2_191(.a(output_3_191), .b(output_3_0), .y(output_2_191));
wire output_1_192, output_1_1, output_0_192;
mixer gate_output_0_192(.a(output_1_192), .b(output_1_1), .y(output_0_192));
wire output_2_192, output_2_1, output_1_192;
mixer gate_output_1_192(.a(output_2_192), .b(output_2_1), .y(output_1_192));
wire output_3_192, output_3_1, output_2_192;
mixer gate_output_2_192(.a(output_3_192), .b(output_3_1), .y(output_2_192));
wire output_1_193, output_1_2, output_0_193;
mixer gate_output_0_193(.a(output_1_193), .b(output_1_2), .y(output_0_193));
wire output_2_193, output_2_2, output_1_193;
mixer gate_output_1_193(.a(output_2_193), .b(output_2_2), .y(output_1_193));
wire output_3_193, output_3_2, output_2_193;
mixer gate_output_2_193(.a(output_3_193), .b(output_3_2), .y(output_2_193));
wire output_1_194, output_1_0, output_0_194;
mixer gate_output_0_194(.a(output_1_194), .b(output_1_0), .y(output_0_194));
wire output_2_194, output_2_0, output_1_194;
mixer gate_output_1_194(.a(output_2_194), .b(output_2_0), .y(output_1_194));
wire output_3_194, output_3_0, output_2_194;
mixer gate_output_2_194(.a(output_3_194), .b(output_3_0), .y(output_2_194));
wire output_1_195, output_1_1, output_0_195;
mixer gate_output_0_195(.a(output_1_195), .b(output_1_1), .y(output_0_195));
wire output_2_195, output_2_1, output_1_195;
mixer gate_output_1_195(.a(output_2_195), .b(output_2_1), .y(output_1_195));
wire output_3_195, output_3_1, output_2_195;
mixer gate_output_2_195(.a(output_3_195), .b(output_3_1), .y(output_2_195));
wire output_1_196, output_1_2, output_0_196;
mixer gate_output_0_196(.a(output_1_196), .b(output_1_2), .y(output_0_196));
wire output_2_196, output_2_2, output_1_196;
mixer gate_output_1_196(.a(output_2_196), .b(output_2_2), .y(output_1_196));
wire output_3_196, output_3_2, output_2_196;
mixer gate_output_2_196(.a(output_3_196), .b(output_3_2), .y(output_2_196));
wire output_1_197, output_1_0, output_0_197;
mixer gate_output_0_197(.a(output_1_197), .b(output_1_0), .y(output_0_197));
wire output_2_197, output_2_0, output_1_197;
mixer gate_output_1_197(.a(output_2_197), .b(output_2_0), .y(output_1_197));
wire output_3_197, output_3_0, output_2_197;
mixer gate_output_2_197(.a(output_3_197), .b(output_3_0), .y(output_2_197));
wire output_1_198, output_1_1, output_0_198;
mixer gate_output_0_198(.a(output_1_198), .b(output_1_1), .y(output_0_198));
wire output_2_198, output_2_1, output_1_198;
mixer gate_output_1_198(.a(output_2_198), .b(output_2_1), .y(output_1_198));
wire output_3_198, output_3_1, output_2_198;
mixer gate_output_2_198(.a(output_3_198), .b(output_3_1), .y(output_2_198));
wire output_1_199, output_1_2, output_0_199;
mixer gate_output_0_199(.a(output_1_199), .b(output_1_2), .y(output_0_199));
wire output_2_199, output_2_2, output_1_199;
mixer gate_output_1_199(.a(output_2_199), .b(output_2_2), .y(output_1_199));
wire output_3_199, output_3_2, output_2_199;
mixer gate_output_2_199(.a(output_3_199), .b(output_3_2), .y(output_2_199));
wire output_1_200, output_1_0, output_0_200;
mixer gate_output_0_200(.a(output_1_200), .b(output_1_0), .y(output_0_200));
wire output_2_200, output_2_0, output_1_200;
mixer gate_output_1_200(.a(output_2_200), .b(output_2_0), .y(output_1_200));
wire output_3_200, output_3_0, output_2_200;
mixer gate_output_2_200(.a(output_3_200), .b(output_3_0), .y(output_2_200));
wire output_1_201, output_1_1, output_0_201;
mixer gate_output_0_201(.a(output_1_201), .b(output_1_1), .y(output_0_201));
wire output_2_201, output_2_1, output_1_201;
mixer gate_output_1_201(.a(output_2_201), .b(output_2_1), .y(output_1_201));
wire output_3_201, output_3_1, output_2_201;
mixer gate_output_2_201(.a(output_3_201), .b(output_3_1), .y(output_2_201));
wire output_1_202, output_1_2, output_0_202;
mixer gate_output_0_202(.a(output_1_202), .b(output_1_2), .y(output_0_202));
wire output_2_202, output_2_2, output_1_202;
mixer gate_output_1_202(.a(output_2_202), .b(output_2_2), .y(output_1_202));
wire output_3_202, output_3_2, output_2_202;
mixer gate_output_2_202(.a(output_3_202), .b(output_3_2), .y(output_2_202));
wire output_1_203, output_1_0, output_0_203;
mixer gate_output_0_203(.a(output_1_203), .b(output_1_0), .y(output_0_203));
wire output_2_203, output_2_0, output_1_203;
mixer gate_output_1_203(.a(output_2_203), .b(output_2_0), .y(output_1_203));
wire output_3_203, output_3_0, output_2_203;
mixer gate_output_2_203(.a(output_3_203), .b(output_3_0), .y(output_2_203));
wire output_1_204, output_1_1, output_0_204;
mixer gate_output_0_204(.a(output_1_204), .b(output_1_1), .y(output_0_204));
wire output_2_204, output_2_1, output_1_204;
mixer gate_output_1_204(.a(output_2_204), .b(output_2_1), .y(output_1_204));
wire output_3_204, output_3_1, output_2_204;
mixer gate_output_2_204(.a(output_3_204), .b(output_3_1), .y(output_2_204));
wire output_1_205, output_1_2, output_0_205;
mixer gate_output_0_205(.a(output_1_205), .b(output_1_2), .y(output_0_205));
wire output_2_205, output_2_2, output_1_205;
mixer gate_output_1_205(.a(output_2_205), .b(output_2_2), .y(output_1_205));
wire output_3_205, output_3_2, output_2_205;
mixer gate_output_2_205(.a(output_3_205), .b(output_3_2), .y(output_2_205));
wire output_1_206, output_1_0, output_0_206;
mixer gate_output_0_206(.a(output_1_206), .b(output_1_0), .y(output_0_206));
wire output_2_206, output_2_0, output_1_206;
mixer gate_output_1_206(.a(output_2_206), .b(output_2_0), .y(output_1_206));
wire output_3_206, output_3_0, output_2_206;
mixer gate_output_2_206(.a(output_3_206), .b(output_3_0), .y(output_2_206));
wire output_1_207, output_1_1, output_0_207;
mixer gate_output_0_207(.a(output_1_207), .b(output_1_1), .y(output_0_207));
wire output_2_207, output_2_1, output_1_207;
mixer gate_output_1_207(.a(output_2_207), .b(output_2_1), .y(output_1_207));
wire output_3_207, output_3_1, output_2_207;
mixer gate_output_2_207(.a(output_3_207), .b(output_3_1), .y(output_2_207));
wire output_1_208, output_1_2, output_0_208;
mixer gate_output_0_208(.a(output_1_208), .b(output_1_2), .y(output_0_208));
wire output_2_208, output_2_2, output_1_208;
mixer gate_output_1_208(.a(output_2_208), .b(output_2_2), .y(output_1_208));
wire output_3_208, output_3_2, output_2_208;
mixer gate_output_2_208(.a(output_3_208), .b(output_3_2), .y(output_2_208));
wire output_1_209, output_1_0, output_0_209;
mixer gate_output_0_209(.a(output_1_209), .b(output_1_0), .y(output_0_209));
wire output_2_209, output_2_0, output_1_209;
mixer gate_output_1_209(.a(output_2_209), .b(output_2_0), .y(output_1_209));
wire output_3_209, output_3_0, output_2_209;
mixer gate_output_2_209(.a(output_3_209), .b(output_3_0), .y(output_2_209));
wire output_1_210, output_1_1, output_0_210;
mixer gate_output_0_210(.a(output_1_210), .b(output_1_1), .y(output_0_210));
wire output_2_210, output_2_1, output_1_210;
mixer gate_output_1_210(.a(output_2_210), .b(output_2_1), .y(output_1_210));
wire output_3_210, output_3_1, output_2_210;
mixer gate_output_2_210(.a(output_3_210), .b(output_3_1), .y(output_2_210));
wire output_1_211, output_1_2, output_0_211;
mixer gate_output_0_211(.a(output_1_211), .b(output_1_2), .y(output_0_211));
wire output_2_211, output_2_2, output_1_211;
mixer gate_output_1_211(.a(output_2_211), .b(output_2_2), .y(output_1_211));
wire output_3_211, output_3_2, output_2_211;
mixer gate_output_2_211(.a(output_3_211), .b(output_3_2), .y(output_2_211));
wire output_1_212, output_1_0, output_0_212;
mixer gate_output_0_212(.a(output_1_212), .b(output_1_0), .y(output_0_212));
wire output_2_212, output_2_0, output_1_212;
mixer gate_output_1_212(.a(output_2_212), .b(output_2_0), .y(output_1_212));
wire output_3_212, output_3_0, output_2_212;
mixer gate_output_2_212(.a(output_3_212), .b(output_3_0), .y(output_2_212));
wire output_1_213, output_1_1, output_0_213;
mixer gate_output_0_213(.a(output_1_213), .b(output_1_1), .y(output_0_213));
wire output_2_213, output_2_1, output_1_213;
mixer gate_output_1_213(.a(output_2_213), .b(output_2_1), .y(output_1_213));
wire output_3_213, output_3_1, output_2_213;
mixer gate_output_2_213(.a(output_3_213), .b(output_3_1), .y(output_2_213));
wire output_1_214, output_1_2, output_0_214;
mixer gate_output_0_214(.a(output_1_214), .b(output_1_2), .y(output_0_214));
wire output_2_214, output_2_2, output_1_214;
mixer gate_output_1_214(.a(output_2_214), .b(output_2_2), .y(output_1_214));
wire output_3_214, output_3_2, output_2_214;
mixer gate_output_2_214(.a(output_3_214), .b(output_3_2), .y(output_2_214));
wire output_1_215, output_1_0, output_0_215;
mixer gate_output_0_215(.a(output_1_215), .b(output_1_0), .y(output_0_215));
wire output_2_215, output_2_0, output_1_215;
mixer gate_output_1_215(.a(output_2_215), .b(output_2_0), .y(output_1_215));
wire output_3_215, output_3_0, output_2_215;
mixer gate_output_2_215(.a(output_3_215), .b(output_3_0), .y(output_2_215));
wire output_1_216, output_1_1, output_0_216;
mixer gate_output_0_216(.a(output_1_216), .b(output_1_1), .y(output_0_216));
wire output_2_216, output_2_1, output_1_216;
mixer gate_output_1_216(.a(output_2_216), .b(output_2_1), .y(output_1_216));
wire output_3_216, output_3_1, output_2_216;
mixer gate_output_2_216(.a(output_3_216), .b(output_3_1), .y(output_2_216));
wire output_1_217, output_1_2, output_0_217;
mixer gate_output_0_217(.a(output_1_217), .b(output_1_2), .y(output_0_217));
wire output_2_217, output_2_2, output_1_217;
mixer gate_output_1_217(.a(output_2_217), .b(output_2_2), .y(output_1_217));
wire output_3_217, output_3_2, output_2_217;
mixer gate_output_2_217(.a(output_3_217), .b(output_3_2), .y(output_2_217));
wire output_1_218, output_1_0, output_0_218;
mixer gate_output_0_218(.a(output_1_218), .b(output_1_0), .y(output_0_218));
wire output_2_218, output_2_0, output_1_218;
mixer gate_output_1_218(.a(output_2_218), .b(output_2_0), .y(output_1_218));
wire output_3_218, output_3_0, output_2_218;
mixer gate_output_2_218(.a(output_3_218), .b(output_3_0), .y(output_2_218));
wire output_1_219, output_1_1, output_0_219;
mixer gate_output_0_219(.a(output_1_219), .b(output_1_1), .y(output_0_219));
wire output_2_219, output_2_1, output_1_219;
mixer gate_output_1_219(.a(output_2_219), .b(output_2_1), .y(output_1_219));
wire output_3_219, output_3_1, output_2_219;
mixer gate_output_2_219(.a(output_3_219), .b(output_3_1), .y(output_2_219));
wire output_1_220, output_1_2, output_0_220;
mixer gate_output_0_220(.a(output_1_220), .b(output_1_2), .y(output_0_220));
wire output_2_220, output_2_2, output_1_220;
mixer gate_output_1_220(.a(output_2_220), .b(output_2_2), .y(output_1_220));
wire output_3_220, output_3_2, output_2_220;
mixer gate_output_2_220(.a(output_3_220), .b(output_3_2), .y(output_2_220));
wire output_1_221, output_1_0, output_0_221;
mixer gate_output_0_221(.a(output_1_221), .b(output_1_0), .y(output_0_221));
wire output_2_221, output_2_0, output_1_221;
mixer gate_output_1_221(.a(output_2_221), .b(output_2_0), .y(output_1_221));
wire output_3_221, output_3_0, output_2_221;
mixer gate_output_2_221(.a(output_3_221), .b(output_3_0), .y(output_2_221));
wire output_1_222, output_1_1, output_0_222;
mixer gate_output_0_222(.a(output_1_222), .b(output_1_1), .y(output_0_222));
wire output_2_222, output_2_1, output_1_222;
mixer gate_output_1_222(.a(output_2_222), .b(output_2_1), .y(output_1_222));
wire output_3_222, output_3_1, output_2_222;
mixer gate_output_2_222(.a(output_3_222), .b(output_3_1), .y(output_2_222));
wire output_1_223, output_1_2, output_0_223;
mixer gate_output_0_223(.a(output_1_223), .b(output_1_2), .y(output_0_223));
wire output_2_223, output_2_2, output_1_223;
mixer gate_output_1_223(.a(output_2_223), .b(output_2_2), .y(output_1_223));
wire output_3_223, output_3_2, output_2_223;
mixer gate_output_2_223(.a(output_3_223), .b(output_3_2), .y(output_2_223));
wire output_1_224, output_1_0, output_0_224;
mixer gate_output_0_224(.a(output_1_224), .b(output_1_0), .y(output_0_224));
wire output_2_224, output_2_0, output_1_224;
mixer gate_output_1_224(.a(output_2_224), .b(output_2_0), .y(output_1_224));
wire output_3_224, output_3_0, output_2_224;
mixer gate_output_2_224(.a(output_3_224), .b(output_3_0), .y(output_2_224));
wire output_1_225, output_1_1, output_0_225;
mixer gate_output_0_225(.a(output_1_225), .b(output_1_1), .y(output_0_225));
wire output_2_225, output_2_1, output_1_225;
mixer gate_output_1_225(.a(output_2_225), .b(output_2_1), .y(output_1_225));
wire output_3_225, output_3_1, output_2_225;
mixer gate_output_2_225(.a(output_3_225), .b(output_3_1), .y(output_2_225));
wire output_1_226, output_1_2, output_0_226;
mixer gate_output_0_226(.a(output_1_226), .b(output_1_2), .y(output_0_226));
wire output_2_226, output_2_2, output_1_226;
mixer gate_output_1_226(.a(output_2_226), .b(output_2_2), .y(output_1_226));
wire output_3_226, output_3_2, output_2_226;
mixer gate_output_2_226(.a(output_3_226), .b(output_3_2), .y(output_2_226));
wire output_1_227, output_1_0, output_0_227;
mixer gate_output_0_227(.a(output_1_227), .b(output_1_0), .y(output_0_227));
wire output_2_227, output_2_0, output_1_227;
mixer gate_output_1_227(.a(output_2_227), .b(output_2_0), .y(output_1_227));
wire output_3_227, output_3_0, output_2_227;
mixer gate_output_2_227(.a(output_3_227), .b(output_3_0), .y(output_2_227));
wire output_1_228, output_1_1, output_0_228;
mixer gate_output_0_228(.a(output_1_228), .b(output_1_1), .y(output_0_228));
wire output_2_228, output_2_1, output_1_228;
mixer gate_output_1_228(.a(output_2_228), .b(output_2_1), .y(output_1_228));
wire output_3_228, output_3_1, output_2_228;
mixer gate_output_2_228(.a(output_3_228), .b(output_3_1), .y(output_2_228));
wire output_1_229, output_1_2, output_0_229;
mixer gate_output_0_229(.a(output_1_229), .b(output_1_2), .y(output_0_229));
wire output_2_229, output_2_2, output_1_229;
mixer gate_output_1_229(.a(output_2_229), .b(output_2_2), .y(output_1_229));
wire output_3_229, output_3_2, output_2_229;
mixer gate_output_2_229(.a(output_3_229), .b(output_3_2), .y(output_2_229));
wire output_1_230, output_1_0, output_0_230;
mixer gate_output_0_230(.a(output_1_230), .b(output_1_0), .y(output_0_230));
wire output_2_230, output_2_0, output_1_230;
mixer gate_output_1_230(.a(output_2_230), .b(output_2_0), .y(output_1_230));
wire output_3_230, output_3_0, output_2_230;
mixer gate_output_2_230(.a(output_3_230), .b(output_3_0), .y(output_2_230));
wire output_1_231, output_1_1, output_0_231;
mixer gate_output_0_231(.a(output_1_231), .b(output_1_1), .y(output_0_231));
wire output_2_231, output_2_1, output_1_231;
mixer gate_output_1_231(.a(output_2_231), .b(output_2_1), .y(output_1_231));
wire output_3_231, output_3_1, output_2_231;
mixer gate_output_2_231(.a(output_3_231), .b(output_3_1), .y(output_2_231));
wire output_1_232, output_1_2, output_0_232;
mixer gate_output_0_232(.a(output_1_232), .b(output_1_2), .y(output_0_232));
wire output_2_232, output_2_2, output_1_232;
mixer gate_output_1_232(.a(output_2_232), .b(output_2_2), .y(output_1_232));
wire output_3_232, output_3_2, output_2_232;
mixer gate_output_2_232(.a(output_3_232), .b(output_3_2), .y(output_2_232));
wire output_1_233, output_1_0, output_0_233;
mixer gate_output_0_233(.a(output_1_233), .b(output_1_0), .y(output_0_233));
wire output_2_233, output_2_0, output_1_233;
mixer gate_output_1_233(.a(output_2_233), .b(output_2_0), .y(output_1_233));
wire output_3_233, output_3_0, output_2_233;
mixer gate_output_2_233(.a(output_3_233), .b(output_3_0), .y(output_2_233));
wire output_1_234, output_1_1, output_0_234;
mixer gate_output_0_234(.a(output_1_234), .b(output_1_1), .y(output_0_234));
wire output_2_234, output_2_1, output_1_234;
mixer gate_output_1_234(.a(output_2_234), .b(output_2_1), .y(output_1_234));
wire output_3_234, output_3_1, output_2_234;
mixer gate_output_2_234(.a(output_3_234), .b(output_3_1), .y(output_2_234));
wire output_1_235, output_1_2, output_0_235;
mixer gate_output_0_235(.a(output_1_235), .b(output_1_2), .y(output_0_235));
wire output_2_235, output_2_2, output_1_235;
mixer gate_output_1_235(.a(output_2_235), .b(output_2_2), .y(output_1_235));
wire output_3_235, output_3_2, output_2_235;
mixer gate_output_2_235(.a(output_3_235), .b(output_3_2), .y(output_2_235));
wire output_1_236, output_1_0, output_0_236;
mixer gate_output_0_236(.a(output_1_236), .b(output_1_0), .y(output_0_236));
wire output_2_236, output_2_0, output_1_236;
mixer gate_output_1_236(.a(output_2_236), .b(output_2_0), .y(output_1_236));
wire output_3_236, output_3_0, output_2_236;
mixer gate_output_2_236(.a(output_3_236), .b(output_3_0), .y(output_2_236));
wire output_1_237, output_1_1, output_0_237;
mixer gate_output_0_237(.a(output_1_237), .b(output_1_1), .y(output_0_237));
wire output_2_237, output_2_1, output_1_237;
mixer gate_output_1_237(.a(output_2_237), .b(output_2_1), .y(output_1_237));
wire output_3_237, output_3_1, output_2_237;
mixer gate_output_2_237(.a(output_3_237), .b(output_3_1), .y(output_2_237));
wire output_1_238, output_1_2, output_0_238;
mixer gate_output_0_238(.a(output_1_238), .b(output_1_2), .y(output_0_238));
wire output_2_238, output_2_2, output_1_238;
mixer gate_output_1_238(.a(output_2_238), .b(output_2_2), .y(output_1_238));
wire output_3_238, output_3_2, output_2_238;
mixer gate_output_2_238(.a(output_3_238), .b(output_3_2), .y(output_2_238));
wire output_1_239, output_1_0, output_0_239;
mixer gate_output_0_239(.a(output_1_239), .b(output_1_0), .y(output_0_239));
wire output_2_239, output_2_0, output_1_239;
mixer gate_output_1_239(.a(output_2_239), .b(output_2_0), .y(output_1_239));
wire output_3_239, output_3_0, output_2_239;
mixer gate_output_2_239(.a(output_3_239), .b(output_3_0), .y(output_2_239));
wire output_1_240, output_1_1, output_0_240;
mixer gate_output_0_240(.a(output_1_240), .b(output_1_1), .y(output_0_240));
wire output_2_240, output_2_1, output_1_240;
mixer gate_output_1_240(.a(output_2_240), .b(output_2_1), .y(output_1_240));
wire output_3_240, output_3_1, output_2_240;
mixer gate_output_2_240(.a(output_3_240), .b(output_3_1), .y(output_2_240));
wire output_1_241, output_1_2, output_0_241;
mixer gate_output_0_241(.a(output_1_241), .b(output_1_2), .y(output_0_241));
wire output_2_241, output_2_2, output_1_241;
mixer gate_output_1_241(.a(output_2_241), .b(output_2_2), .y(output_1_241));
wire output_3_241, output_3_2, output_2_241;
mixer gate_output_2_241(.a(output_3_241), .b(output_3_2), .y(output_2_241));
wire output_1_242, output_1_0, output_0_242;
mixer gate_output_0_242(.a(output_1_242), .b(output_1_0), .y(output_0_242));
wire output_2_242, output_2_0, output_1_242;
mixer gate_output_1_242(.a(output_2_242), .b(output_2_0), .y(output_1_242));
wire output_3_242, output_3_0, output_2_242;
mixer gate_output_2_242(.a(output_3_242), .b(output_3_0), .y(output_2_242));
wire output_1_243, output_1_1, output_0_243;
mixer gate_output_0_243(.a(output_1_243), .b(output_1_1), .y(output_0_243));
wire output_2_243, output_2_1, output_1_243;
mixer gate_output_1_243(.a(output_2_243), .b(output_2_1), .y(output_1_243));
wire output_3_243, output_3_1, output_2_243;
mixer gate_output_2_243(.a(output_3_243), .b(output_3_1), .y(output_2_243));
wire output_1_244, output_1_2, output_0_244;
mixer gate_output_0_244(.a(output_1_244), .b(output_1_2), .y(output_0_244));
wire output_2_244, output_2_2, output_1_244;
mixer gate_output_1_244(.a(output_2_244), .b(output_2_2), .y(output_1_244));
wire output_3_244, output_3_2, output_2_244;
mixer gate_output_2_244(.a(output_3_244), .b(output_3_2), .y(output_2_244));
wire output_1_245, output_1_0, output_0_245;
mixer gate_output_0_245(.a(output_1_245), .b(output_1_0), .y(output_0_245));
wire output_2_245, output_2_0, output_1_245;
mixer gate_output_1_245(.a(output_2_245), .b(output_2_0), .y(output_1_245));
wire output_3_245, output_3_0, output_2_245;
mixer gate_output_2_245(.a(output_3_245), .b(output_3_0), .y(output_2_245));
wire output_1_246, output_1_1, output_0_246;
mixer gate_output_0_246(.a(output_1_246), .b(output_1_1), .y(output_0_246));
wire output_2_246, output_2_1, output_1_246;
mixer gate_output_1_246(.a(output_2_246), .b(output_2_1), .y(output_1_246));
wire output_3_246, output_3_1, output_2_246;
mixer gate_output_2_246(.a(output_3_246), .b(output_3_1), .y(output_2_246));
wire output_1_247, output_1_2, output_0_247;
mixer gate_output_0_247(.a(output_1_247), .b(output_1_2), .y(output_0_247));
wire output_2_247, output_2_2, output_1_247;
mixer gate_output_1_247(.a(output_2_247), .b(output_2_2), .y(output_1_247));
wire output_3_247, output_3_2, output_2_247;
mixer gate_output_2_247(.a(output_3_247), .b(output_3_2), .y(output_2_247));
wire output_1_248, output_1_0, output_0_248;
mixer gate_output_0_248(.a(output_1_248), .b(output_1_0), .y(output_0_248));
wire output_2_248, output_2_0, output_1_248;
mixer gate_output_1_248(.a(output_2_248), .b(output_2_0), .y(output_1_248));
wire output_3_248, output_3_0, output_2_248;
mixer gate_output_2_248(.a(output_3_248), .b(output_3_0), .y(output_2_248));
wire output_1_249, output_1_1, output_0_249;
mixer gate_output_0_249(.a(output_1_249), .b(output_1_1), .y(output_0_249));
wire output_2_249, output_2_1, output_1_249;
mixer gate_output_1_249(.a(output_2_249), .b(output_2_1), .y(output_1_249));
wire output_3_249, output_3_1, output_2_249;
mixer gate_output_2_249(.a(output_3_249), .b(output_3_1), .y(output_2_249));
wire output_1_250, output_1_2, output_0_250;
mixer gate_output_0_250(.a(output_1_250), .b(output_1_2), .y(output_0_250));
wire output_2_250, output_2_2, output_1_250;
mixer gate_output_1_250(.a(output_2_250), .b(output_2_2), .y(output_1_250));
wire output_3_250, output_3_2, output_2_250;
mixer gate_output_2_250(.a(output_3_250), .b(output_3_2), .y(output_2_250));
wire output_1_251, output_1_0, output_0_251;
mixer gate_output_0_251(.a(output_1_251), .b(output_1_0), .y(output_0_251));
wire output_2_251, output_2_0, output_1_251;
mixer gate_output_1_251(.a(output_2_251), .b(output_2_0), .y(output_1_251));
wire output_3_251, output_3_0, output_2_251;
mixer gate_output_2_251(.a(output_3_251), .b(output_3_0), .y(output_2_251));
wire output_1_252, output_1_1, output_0_252;
mixer gate_output_0_252(.a(output_1_252), .b(output_1_1), .y(output_0_252));
wire output_2_252, output_2_1, output_1_252;
mixer gate_output_1_252(.a(output_2_252), .b(output_2_1), .y(output_1_252));
wire output_3_252, output_3_1, output_2_252;
mixer gate_output_2_252(.a(output_3_252), .b(output_3_1), .y(output_2_252));
wire output_1_253, output_1_2, output_0_253;
mixer gate_output_0_253(.a(output_1_253), .b(output_1_2), .y(output_0_253));
wire output_2_253, output_2_2, output_1_253;
mixer gate_output_1_253(.a(output_2_253), .b(output_2_2), .y(output_1_253));
wire output_3_253, output_3_2, output_2_253;
mixer gate_output_2_253(.a(output_3_253), .b(output_3_2), .y(output_2_253));
wire output_1_254, output_1_0, output_0_254;
mixer gate_output_0_254(.a(output_1_254), .b(output_1_0), .y(output_0_254));
wire output_2_254, output_2_0, output_1_254;
mixer gate_output_1_254(.a(output_2_254), .b(output_2_0), .y(output_1_254));
wire output_3_254, output_3_0, output_2_254;
mixer gate_output_2_254(.a(output_3_254), .b(output_3_0), .y(output_2_254));
wire output_1_255, output_1_1, output_0_255;
mixer gate_output_0_255(.a(output_1_255), .b(output_1_1), .y(output_0_255));
wire output_2_255, output_2_1, output_1_255;
mixer gate_output_1_255(.a(output_2_255), .b(output_2_1), .y(output_1_255));
wire output_3_255, output_3_1, output_2_255;
mixer gate_output_2_255(.a(output_3_255), .b(output_3_1), .y(output_2_255));
wire output_1_256, output_1_2, output_0_256;
mixer gate_output_0_256(.a(output_1_256), .b(output_1_2), .y(output_0_256));
wire output_2_256, output_2_2, output_1_256;
mixer gate_output_1_256(.a(output_2_256), .b(output_2_2), .y(output_1_256));
wire output_3_256, output_3_2, output_2_256;
mixer gate_output_2_256(.a(output_3_256), .b(output_3_2), .y(output_2_256));
wire output_1_257, output_1_0, output_0_257;
mixer gate_output_0_257(.a(output_1_257), .b(output_1_0), .y(output_0_257));
wire output_2_257, output_2_0, output_1_257;
mixer gate_output_1_257(.a(output_2_257), .b(output_2_0), .y(output_1_257));
wire output_3_257, output_3_0, output_2_257;
mixer gate_output_2_257(.a(output_3_257), .b(output_3_0), .y(output_2_257));
wire output_1_258, output_1_1, output_0_258;
mixer gate_output_0_258(.a(output_1_258), .b(output_1_1), .y(output_0_258));
wire output_2_258, output_2_1, output_1_258;
mixer gate_output_1_258(.a(output_2_258), .b(output_2_1), .y(output_1_258));
wire output_3_258, output_3_1, output_2_258;
mixer gate_output_2_258(.a(output_3_258), .b(output_3_1), .y(output_2_258));
wire output_1_259, output_1_2, output_0_259;
mixer gate_output_0_259(.a(output_1_259), .b(output_1_2), .y(output_0_259));
wire output_2_259, output_2_2, output_1_259;
mixer gate_output_1_259(.a(output_2_259), .b(output_2_2), .y(output_1_259));
wire output_3_259, output_3_2, output_2_259;
mixer gate_output_2_259(.a(output_3_259), .b(output_3_2), .y(output_2_259));
wire output_1_260, output_1_0, output_0_260;
mixer gate_output_0_260(.a(output_1_260), .b(output_1_0), .y(output_0_260));
wire output_2_260, output_2_0, output_1_260;
mixer gate_output_1_260(.a(output_2_260), .b(output_2_0), .y(output_1_260));
wire output_3_260, output_3_0, output_2_260;
mixer gate_output_2_260(.a(output_3_260), .b(output_3_0), .y(output_2_260));
wire output_1_261, output_1_1, output_0_261;
mixer gate_output_0_261(.a(output_1_261), .b(output_1_1), .y(output_0_261));
wire output_2_261, output_2_1, output_1_261;
mixer gate_output_1_261(.a(output_2_261), .b(output_2_1), .y(output_1_261));
wire output_3_261, output_3_1, output_2_261;
mixer gate_output_2_261(.a(output_3_261), .b(output_3_1), .y(output_2_261));
wire output_1_262, output_1_2, output_0_262;
mixer gate_output_0_262(.a(output_1_262), .b(output_1_2), .y(output_0_262));
wire output_2_262, output_2_2, output_1_262;
mixer gate_output_1_262(.a(output_2_262), .b(output_2_2), .y(output_1_262));
wire output_3_262, output_3_2, output_2_262;
mixer gate_output_2_262(.a(output_3_262), .b(output_3_2), .y(output_2_262));
wire output_1_263, output_1_0, output_0_263;
mixer gate_output_0_263(.a(output_1_263), .b(output_1_0), .y(output_0_263));
wire output_2_263, output_2_0, output_1_263;
mixer gate_output_1_263(.a(output_2_263), .b(output_2_0), .y(output_1_263));
wire output_3_263, output_3_0, output_2_263;
mixer gate_output_2_263(.a(output_3_263), .b(output_3_0), .y(output_2_263));
wire output_1_264, output_1_1, output_0_264;
mixer gate_output_0_264(.a(output_1_264), .b(output_1_1), .y(output_0_264));
wire output_2_264, output_2_1, output_1_264;
mixer gate_output_1_264(.a(output_2_264), .b(output_2_1), .y(output_1_264));
wire output_3_264, output_3_1, output_2_264;
mixer gate_output_2_264(.a(output_3_264), .b(output_3_1), .y(output_2_264));
wire output_1_265, output_1_2, output_0_265;
mixer gate_output_0_265(.a(output_1_265), .b(output_1_2), .y(output_0_265));
wire output_2_265, output_2_2, output_1_265;
mixer gate_output_1_265(.a(output_2_265), .b(output_2_2), .y(output_1_265));
wire output_3_265, output_3_2, output_2_265;
mixer gate_output_2_265(.a(output_3_265), .b(output_3_2), .y(output_2_265));
wire output_1_266, output_1_0, output_0_266;
mixer gate_output_0_266(.a(output_1_266), .b(output_1_0), .y(output_0_266));
wire output_2_266, output_2_0, output_1_266;
mixer gate_output_1_266(.a(output_2_266), .b(output_2_0), .y(output_1_266));
wire output_3_266, output_3_0, output_2_266;
mixer gate_output_2_266(.a(output_3_266), .b(output_3_0), .y(output_2_266));
wire output_1_267, output_1_1, output_0_267;
mixer gate_output_0_267(.a(output_1_267), .b(output_1_1), .y(output_0_267));
wire output_2_267, output_2_1, output_1_267;
mixer gate_output_1_267(.a(output_2_267), .b(output_2_1), .y(output_1_267));
wire output_3_267, output_3_1, output_2_267;
mixer gate_output_2_267(.a(output_3_267), .b(output_3_1), .y(output_2_267));
wire output_1_268, output_1_2, output_0_268;
mixer gate_output_0_268(.a(output_1_268), .b(output_1_2), .y(output_0_268));
wire output_2_268, output_2_2, output_1_268;
mixer gate_output_1_268(.a(output_2_268), .b(output_2_2), .y(output_1_268));
wire output_3_268, output_3_2, output_2_268;
mixer gate_output_2_268(.a(output_3_268), .b(output_3_2), .y(output_2_268));
wire output_1_269, output_1_0, output_0_269;
mixer gate_output_0_269(.a(output_1_269), .b(output_1_0), .y(output_0_269));
wire output_2_269, output_2_0, output_1_269;
mixer gate_output_1_269(.a(output_2_269), .b(output_2_0), .y(output_1_269));
wire output_3_269, output_3_0, output_2_269;
mixer gate_output_2_269(.a(output_3_269), .b(output_3_0), .y(output_2_269));
wire output_1_270, output_1_1, output_0_270;
mixer gate_output_0_270(.a(output_1_270), .b(output_1_1), .y(output_0_270));
wire output_2_270, output_2_1, output_1_270;
mixer gate_output_1_270(.a(output_2_270), .b(output_2_1), .y(output_1_270));
wire output_3_270, output_3_1, output_2_270;
mixer gate_output_2_270(.a(output_3_270), .b(output_3_1), .y(output_2_270));
wire output_1_271, output_1_2, output_0_271;
mixer gate_output_0_271(.a(output_1_271), .b(output_1_2), .y(output_0_271));
wire output_2_271, output_2_2, output_1_271;
mixer gate_output_1_271(.a(output_2_271), .b(output_2_2), .y(output_1_271));
wire output_3_271, output_3_2, output_2_271;
mixer gate_output_2_271(.a(output_3_271), .b(output_3_2), .y(output_2_271));
wire output_1_272, output_1_0, output_0_272;
mixer gate_output_0_272(.a(output_1_272), .b(output_1_0), .y(output_0_272));
wire output_2_272, output_2_0, output_1_272;
mixer gate_output_1_272(.a(output_2_272), .b(output_2_0), .y(output_1_272));
wire output_3_272, output_3_0, output_2_272;
mixer gate_output_2_272(.a(output_3_272), .b(output_3_0), .y(output_2_272));
wire output_1_273, output_1_1, output_0_273;
mixer gate_output_0_273(.a(output_1_273), .b(output_1_1), .y(output_0_273));
wire output_2_273, output_2_1, output_1_273;
mixer gate_output_1_273(.a(output_2_273), .b(output_2_1), .y(output_1_273));
wire output_3_273, output_3_1, output_2_273;
mixer gate_output_2_273(.a(output_3_273), .b(output_3_1), .y(output_2_273));
wire output_1_274, output_1_2, output_0_274;
mixer gate_output_0_274(.a(output_1_274), .b(output_1_2), .y(output_0_274));
wire output_2_274, output_2_2, output_1_274;
mixer gate_output_1_274(.a(output_2_274), .b(output_2_2), .y(output_1_274));
wire output_3_274, output_3_2, output_2_274;
mixer gate_output_2_274(.a(output_3_274), .b(output_3_2), .y(output_2_274));
wire output_1_275, output_1_0, output_0_275;
mixer gate_output_0_275(.a(output_1_275), .b(output_1_0), .y(output_0_275));
wire output_2_275, output_2_0, output_1_275;
mixer gate_output_1_275(.a(output_2_275), .b(output_2_0), .y(output_1_275));
wire output_3_275, output_3_0, output_2_275;
mixer gate_output_2_275(.a(output_3_275), .b(output_3_0), .y(output_2_275));
wire output_1_276, output_1_1, output_0_276;
mixer gate_output_0_276(.a(output_1_276), .b(output_1_1), .y(output_0_276));
wire output_2_276, output_2_1, output_1_276;
mixer gate_output_1_276(.a(output_2_276), .b(output_2_1), .y(output_1_276));
wire output_3_276, output_3_1, output_2_276;
mixer gate_output_2_276(.a(output_3_276), .b(output_3_1), .y(output_2_276));
wire output_1_277, output_1_2, output_0_277;
mixer gate_output_0_277(.a(output_1_277), .b(output_1_2), .y(output_0_277));
wire output_2_277, output_2_2, output_1_277;
mixer gate_output_1_277(.a(output_2_277), .b(output_2_2), .y(output_1_277));
wire output_3_277, output_3_2, output_2_277;
mixer gate_output_2_277(.a(output_3_277), .b(output_3_2), .y(output_2_277));
wire output_1_278, output_1_0, output_0_278;
mixer gate_output_0_278(.a(output_1_278), .b(output_1_0), .y(output_0_278));
wire output_2_278, output_2_0, output_1_278;
mixer gate_output_1_278(.a(output_2_278), .b(output_2_0), .y(output_1_278));
wire output_3_278, output_3_0, output_2_278;
mixer gate_output_2_278(.a(output_3_278), .b(output_3_0), .y(output_2_278));
wire output_1_279, output_1_1, output_0_279;
mixer gate_output_0_279(.a(output_1_279), .b(output_1_1), .y(output_0_279));
wire output_2_279, output_2_1, output_1_279;
mixer gate_output_1_279(.a(output_2_279), .b(output_2_1), .y(output_1_279));
wire output_3_279, output_3_1, output_2_279;
mixer gate_output_2_279(.a(output_3_279), .b(output_3_1), .y(output_2_279));
wire output_1_280, output_1_2, output_0_280;
mixer gate_output_0_280(.a(output_1_280), .b(output_1_2), .y(output_0_280));
wire output_2_280, output_2_2, output_1_280;
mixer gate_output_1_280(.a(output_2_280), .b(output_2_2), .y(output_1_280));
wire output_3_280, output_3_2, output_2_280;
mixer gate_output_2_280(.a(output_3_280), .b(output_3_2), .y(output_2_280));
wire output_1_281, output_1_0, output_0_281;
mixer gate_output_0_281(.a(output_1_281), .b(output_1_0), .y(output_0_281));
wire output_2_281, output_2_0, output_1_281;
mixer gate_output_1_281(.a(output_2_281), .b(output_2_0), .y(output_1_281));
wire output_3_281, output_3_0, output_2_281;
mixer gate_output_2_281(.a(output_3_281), .b(output_3_0), .y(output_2_281));
wire output_1_282, output_1_1, output_0_282;
mixer gate_output_0_282(.a(output_1_282), .b(output_1_1), .y(output_0_282));
wire output_2_282, output_2_1, output_1_282;
mixer gate_output_1_282(.a(output_2_282), .b(output_2_1), .y(output_1_282));
wire output_3_282, output_3_1, output_2_282;
mixer gate_output_2_282(.a(output_3_282), .b(output_3_1), .y(output_2_282));
wire output_1_283, output_1_2, output_0_283;
mixer gate_output_0_283(.a(output_1_283), .b(output_1_2), .y(output_0_283));
wire output_2_283, output_2_2, output_1_283;
mixer gate_output_1_283(.a(output_2_283), .b(output_2_2), .y(output_1_283));
wire output_3_283, output_3_2, output_2_283;
mixer gate_output_2_283(.a(output_3_283), .b(output_3_2), .y(output_2_283));
wire output_1_284, output_1_0, output_0_284;
mixer gate_output_0_284(.a(output_1_284), .b(output_1_0), .y(output_0_284));
wire output_2_284, output_2_0, output_1_284;
mixer gate_output_1_284(.a(output_2_284), .b(output_2_0), .y(output_1_284));
wire output_3_284, output_3_0, output_2_284;
mixer gate_output_2_284(.a(output_3_284), .b(output_3_0), .y(output_2_284));
wire output_1_285, output_1_1, output_0_285;
mixer gate_output_0_285(.a(output_1_285), .b(output_1_1), .y(output_0_285));
wire output_2_285, output_2_1, output_1_285;
mixer gate_output_1_285(.a(output_2_285), .b(output_2_1), .y(output_1_285));
wire output_3_285, output_3_1, output_2_285;
mixer gate_output_2_285(.a(output_3_285), .b(output_3_1), .y(output_2_285));
wire output_1_286, output_1_2, output_0_286;
mixer gate_output_0_286(.a(output_1_286), .b(output_1_2), .y(output_0_286));
wire output_2_286, output_2_2, output_1_286;
mixer gate_output_1_286(.a(output_2_286), .b(output_2_2), .y(output_1_286));
wire output_3_286, output_3_2, output_2_286;
mixer gate_output_2_286(.a(output_3_286), .b(output_3_2), .y(output_2_286));
wire output_1_287, output_1_0, output_0_287;
mixer gate_output_0_287(.a(output_1_287), .b(output_1_0), .y(output_0_287));
wire output_2_287, output_2_0, output_1_287;
mixer gate_output_1_287(.a(output_2_287), .b(output_2_0), .y(output_1_287));
wire output_3_287, output_3_0, output_2_287;
mixer gate_output_2_287(.a(output_3_287), .b(output_3_0), .y(output_2_287));
wire output_1_288, output_1_1, output_0_288;
mixer gate_output_0_288(.a(output_1_288), .b(output_1_1), .y(output_0_288));
wire output_2_288, output_2_1, output_1_288;
mixer gate_output_1_288(.a(output_2_288), .b(output_2_1), .y(output_1_288));
wire output_3_288, output_3_1, output_2_288;
mixer gate_output_2_288(.a(output_3_288), .b(output_3_1), .y(output_2_288));
wire output_1_289, output_1_2, output_0_289;
mixer gate_output_0_289(.a(output_1_289), .b(output_1_2), .y(output_0_289));
wire output_2_289, output_2_2, output_1_289;
mixer gate_output_1_289(.a(output_2_289), .b(output_2_2), .y(output_1_289));
wire output_3_289, output_3_2, output_2_289;
mixer gate_output_2_289(.a(output_3_289), .b(output_3_2), .y(output_2_289));
wire output_1_290, output_1_0, output_0_290;
mixer gate_output_0_290(.a(output_1_290), .b(output_1_0), .y(output_0_290));
wire output_2_290, output_2_0, output_1_290;
mixer gate_output_1_290(.a(output_2_290), .b(output_2_0), .y(output_1_290));
wire output_3_290, output_3_0, output_2_290;
mixer gate_output_2_290(.a(output_3_290), .b(output_3_0), .y(output_2_290));
wire output_1_291, output_1_1, output_0_291;
mixer gate_output_0_291(.a(output_1_291), .b(output_1_1), .y(output_0_291));
wire output_2_291, output_2_1, output_1_291;
mixer gate_output_1_291(.a(output_2_291), .b(output_2_1), .y(output_1_291));
wire output_3_291, output_3_1, output_2_291;
mixer gate_output_2_291(.a(output_3_291), .b(output_3_1), .y(output_2_291));
wire output_1_292, output_1_2, output_0_292;
mixer gate_output_0_292(.a(output_1_292), .b(output_1_2), .y(output_0_292));
wire output_2_292, output_2_2, output_1_292;
mixer gate_output_1_292(.a(output_2_292), .b(output_2_2), .y(output_1_292));
wire output_3_292, output_3_2, output_2_292;
mixer gate_output_2_292(.a(output_3_292), .b(output_3_2), .y(output_2_292));
wire output_1_293, output_1_0, output_0_293;
mixer gate_output_0_293(.a(output_1_293), .b(output_1_0), .y(output_0_293));
wire output_2_293, output_2_0, output_1_293;
mixer gate_output_1_293(.a(output_2_293), .b(output_2_0), .y(output_1_293));
wire output_3_293, output_3_0, output_2_293;
mixer gate_output_2_293(.a(output_3_293), .b(output_3_0), .y(output_2_293));
wire output_1_294, output_1_1, output_0_294;
mixer gate_output_0_294(.a(output_1_294), .b(output_1_1), .y(output_0_294));
wire output_2_294, output_2_1, output_1_294;
mixer gate_output_1_294(.a(output_2_294), .b(output_2_1), .y(output_1_294));
wire output_3_294, output_3_1, output_2_294;
mixer gate_output_2_294(.a(output_3_294), .b(output_3_1), .y(output_2_294));
wire output_1_295, output_1_2, output_0_295;
mixer gate_output_0_295(.a(output_1_295), .b(output_1_2), .y(output_0_295));
wire output_2_295, output_2_2, output_1_295;
mixer gate_output_1_295(.a(output_2_295), .b(output_2_2), .y(output_1_295));
wire output_3_295, output_3_2, output_2_295;
mixer gate_output_2_295(.a(output_3_295), .b(output_3_2), .y(output_2_295));
wire output_1_296, output_1_0, output_0_296;
mixer gate_output_0_296(.a(output_1_296), .b(output_1_0), .y(output_0_296));
wire output_2_296, output_2_0, output_1_296;
mixer gate_output_1_296(.a(output_2_296), .b(output_2_0), .y(output_1_296));
wire output_3_296, output_3_0, output_2_296;
mixer gate_output_2_296(.a(output_3_296), .b(output_3_0), .y(output_2_296));
wire output_1_297, output_1_1, output_0_297;
mixer gate_output_0_297(.a(output_1_297), .b(output_1_1), .y(output_0_297));
wire output_2_297, output_2_1, output_1_297;
mixer gate_output_1_297(.a(output_2_297), .b(output_2_1), .y(output_1_297));
wire output_3_297, output_3_1, output_2_297;
mixer gate_output_2_297(.a(output_3_297), .b(output_3_1), .y(output_2_297));
wire output_1_298, output_1_2, output_0_298;
mixer gate_output_0_298(.a(output_1_298), .b(output_1_2), .y(output_0_298));
wire output_2_298, output_2_2, output_1_298;
mixer gate_output_1_298(.a(output_2_298), .b(output_2_2), .y(output_1_298));
wire output_3_298, output_3_2, output_2_298;
mixer gate_output_2_298(.a(output_3_298), .b(output_3_2), .y(output_2_298));
wire output_1_299, output_1_0, output_0_299;
mixer gate_output_0_299(.a(output_1_299), .b(output_1_0), .y(output_0_299));
wire output_2_299, output_2_0, output_1_299;
mixer gate_output_1_299(.a(output_2_299), .b(output_2_0), .y(output_1_299));
wire output_3_299, output_3_0, output_2_299;
mixer gate_output_2_299(.a(output_3_299), .b(output_3_0), .y(output_2_299));
wire output_1_300, output_1_1, output_0_300;
mixer gate_output_0_300(.a(output_1_300), .b(output_1_1), .y(output_0_300));
wire output_2_300, output_2_1, output_1_300;
mixer gate_output_1_300(.a(output_2_300), .b(output_2_1), .y(output_1_300));
wire output_3_300, output_3_1, output_2_300;
mixer gate_output_2_300(.a(output_3_300), .b(output_3_1), .y(output_2_300));
wire output_1_301, output_1_2, output_0_301;
mixer gate_output_0_301(.a(output_1_301), .b(output_1_2), .y(output_0_301));
wire output_2_301, output_2_2, output_1_301;
mixer gate_output_1_301(.a(output_2_301), .b(output_2_2), .y(output_1_301));
wire output_3_301, output_3_2, output_2_301;
mixer gate_output_2_301(.a(output_3_301), .b(output_3_2), .y(output_2_301));
wire output_1_302, output_1_0, output_0_302;
mixer gate_output_0_302(.a(output_1_302), .b(output_1_0), .y(output_0_302));
wire output_2_302, output_2_0, output_1_302;
mixer gate_output_1_302(.a(output_2_302), .b(output_2_0), .y(output_1_302));
wire output_3_302, output_3_0, output_2_302;
mixer gate_output_2_302(.a(output_3_302), .b(output_3_0), .y(output_2_302));
wire output_1_303, output_1_1, output_0_303;
mixer gate_output_0_303(.a(output_1_303), .b(output_1_1), .y(output_0_303));
wire output_2_303, output_2_1, output_1_303;
mixer gate_output_1_303(.a(output_2_303), .b(output_2_1), .y(output_1_303));
wire output_3_303, output_3_1, output_2_303;
mixer gate_output_2_303(.a(output_3_303), .b(output_3_1), .y(output_2_303));
wire output_1_304, output_1_2, output_0_304;
mixer gate_output_0_304(.a(output_1_304), .b(output_1_2), .y(output_0_304));
wire output_2_304, output_2_2, output_1_304;
mixer gate_output_1_304(.a(output_2_304), .b(output_2_2), .y(output_1_304));
wire output_3_304, output_3_2, output_2_304;
mixer gate_output_2_304(.a(output_3_304), .b(output_3_2), .y(output_2_304));
wire output_1_305, output_1_0, output_0_305;
mixer gate_output_0_305(.a(output_1_305), .b(output_1_0), .y(output_0_305));
wire output_2_305, output_2_0, output_1_305;
mixer gate_output_1_305(.a(output_2_305), .b(output_2_0), .y(output_1_305));
wire output_3_305, output_3_0, output_2_305;
mixer gate_output_2_305(.a(output_3_305), .b(output_3_0), .y(output_2_305));
wire output_1_306, output_1_1, output_0_306;
mixer gate_output_0_306(.a(output_1_306), .b(output_1_1), .y(output_0_306));
wire output_2_306, output_2_1, output_1_306;
mixer gate_output_1_306(.a(output_2_306), .b(output_2_1), .y(output_1_306));
wire output_3_306, output_3_1, output_2_306;
mixer gate_output_2_306(.a(output_3_306), .b(output_3_1), .y(output_2_306));
wire output_1_307, output_1_2, output_0_307;
mixer gate_output_0_307(.a(output_1_307), .b(output_1_2), .y(output_0_307));
wire output_2_307, output_2_2, output_1_307;
mixer gate_output_1_307(.a(output_2_307), .b(output_2_2), .y(output_1_307));
wire output_3_307, output_3_2, output_2_307;
mixer gate_output_2_307(.a(output_3_307), .b(output_3_2), .y(output_2_307));
wire output_1_308, output_1_0, output_0_308;
mixer gate_output_0_308(.a(output_1_308), .b(output_1_0), .y(output_0_308));
wire output_2_308, output_2_0, output_1_308;
mixer gate_output_1_308(.a(output_2_308), .b(output_2_0), .y(output_1_308));
wire output_3_308, output_3_0, output_2_308;
mixer gate_output_2_308(.a(output_3_308), .b(output_3_0), .y(output_2_308));
wire output_1_309, output_1_1, output_0_309;
mixer gate_output_0_309(.a(output_1_309), .b(output_1_1), .y(output_0_309));
wire output_2_309, output_2_1, output_1_309;
mixer gate_output_1_309(.a(output_2_309), .b(output_2_1), .y(output_1_309));
wire output_3_309, output_3_1, output_2_309;
mixer gate_output_2_309(.a(output_3_309), .b(output_3_1), .y(output_2_309));
wire output_1_310, output_1_2, output_0_310;
mixer gate_output_0_310(.a(output_1_310), .b(output_1_2), .y(output_0_310));
wire output_2_310, output_2_2, output_1_310;
mixer gate_output_1_310(.a(output_2_310), .b(output_2_2), .y(output_1_310));
wire output_3_310, output_3_2, output_2_310;
mixer gate_output_2_310(.a(output_3_310), .b(output_3_2), .y(output_2_310));
wire output_1_311, output_1_0, output_0_311;
mixer gate_output_0_311(.a(output_1_311), .b(output_1_0), .y(output_0_311));
wire output_2_311, output_2_0, output_1_311;
mixer gate_output_1_311(.a(output_2_311), .b(output_2_0), .y(output_1_311));
wire output_3_311, output_3_0, output_2_311;
mixer gate_output_2_311(.a(output_3_311), .b(output_3_0), .y(output_2_311));
wire output_1_312, output_1_1, output_0_312;
mixer gate_output_0_312(.a(output_1_312), .b(output_1_1), .y(output_0_312));
wire output_2_312, output_2_1, output_1_312;
mixer gate_output_1_312(.a(output_2_312), .b(output_2_1), .y(output_1_312));
wire output_3_312, output_3_1, output_2_312;
mixer gate_output_2_312(.a(output_3_312), .b(output_3_1), .y(output_2_312));
wire output_1_313, output_1_2, output_0_313;
mixer gate_output_0_313(.a(output_1_313), .b(output_1_2), .y(output_0_313));
wire output_2_313, output_2_2, output_1_313;
mixer gate_output_1_313(.a(output_2_313), .b(output_2_2), .y(output_1_313));
wire output_3_313, output_3_2, output_2_313;
mixer gate_output_2_313(.a(output_3_313), .b(output_3_2), .y(output_2_313));
wire output_1_314, output_1_0, output_0_314;
mixer gate_output_0_314(.a(output_1_314), .b(output_1_0), .y(output_0_314));
wire output_2_314, output_2_0, output_1_314;
mixer gate_output_1_314(.a(output_2_314), .b(output_2_0), .y(output_1_314));
wire output_3_314, output_3_0, output_2_314;
mixer gate_output_2_314(.a(output_3_314), .b(output_3_0), .y(output_2_314));
wire output_1_315, output_1_1, output_0_315;
mixer gate_output_0_315(.a(output_1_315), .b(output_1_1), .y(output_0_315));
wire output_2_315, output_2_1, output_1_315;
mixer gate_output_1_315(.a(output_2_315), .b(output_2_1), .y(output_1_315));
wire output_3_315, output_3_1, output_2_315;
mixer gate_output_2_315(.a(output_3_315), .b(output_3_1), .y(output_2_315));
wire output_1_316, output_1_2, output_0_316;
mixer gate_output_0_316(.a(output_1_316), .b(output_1_2), .y(output_0_316));
wire output_2_316, output_2_2, output_1_316;
mixer gate_output_1_316(.a(output_2_316), .b(output_2_2), .y(output_1_316));
wire output_3_316, output_3_2, output_2_316;
mixer gate_output_2_316(.a(output_3_316), .b(output_3_2), .y(output_2_316));
wire output_1_317, output_1_0, output_0_317;
mixer gate_output_0_317(.a(output_1_317), .b(output_1_0), .y(output_0_317));
wire output_2_317, output_2_0, output_1_317;
mixer gate_output_1_317(.a(output_2_317), .b(output_2_0), .y(output_1_317));
wire output_3_317, output_3_0, output_2_317;
mixer gate_output_2_317(.a(output_3_317), .b(output_3_0), .y(output_2_317));
wire output_1_318, output_1_1, output_0_318;
mixer gate_output_0_318(.a(output_1_318), .b(output_1_1), .y(output_0_318));
wire output_2_318, output_2_1, output_1_318;
mixer gate_output_1_318(.a(output_2_318), .b(output_2_1), .y(output_1_318));
wire output_3_318, output_3_1, output_2_318;
mixer gate_output_2_318(.a(output_3_318), .b(output_3_1), .y(output_2_318));
wire output_1_319, output_1_2, output_0_319;
mixer gate_output_0_319(.a(output_1_319), .b(output_1_2), .y(output_0_319));
wire output_2_319, output_2_2, output_1_319;
mixer gate_output_1_319(.a(output_2_319), .b(output_2_2), .y(output_1_319));
wire output_3_319, output_3_2, output_2_319;
mixer gate_output_2_319(.a(output_3_319), .b(output_3_2), .y(output_2_319));
wire output_1_320, output_1_0, output_0_320;
mixer gate_output_0_320(.a(output_1_320), .b(output_1_0), .y(output_0_320));
wire output_2_320, output_2_0, output_1_320;
mixer gate_output_1_320(.a(output_2_320), .b(output_2_0), .y(output_1_320));
wire output_3_320, output_3_0, output_2_320;
mixer gate_output_2_320(.a(output_3_320), .b(output_3_0), .y(output_2_320));
wire output_1_321, output_1_1, output_0_321;
mixer gate_output_0_321(.a(output_1_321), .b(output_1_1), .y(output_0_321));
wire output_2_321, output_2_1, output_1_321;
mixer gate_output_1_321(.a(output_2_321), .b(output_2_1), .y(output_1_321));
wire output_3_321, output_3_1, output_2_321;
mixer gate_output_2_321(.a(output_3_321), .b(output_3_1), .y(output_2_321));
wire output_1_322, output_1_2, output_0_322;
mixer gate_output_0_322(.a(output_1_322), .b(output_1_2), .y(output_0_322));
wire output_2_322, output_2_2, output_1_322;
mixer gate_output_1_322(.a(output_2_322), .b(output_2_2), .y(output_1_322));
wire output_3_322, output_3_2, output_2_322;
mixer gate_output_2_322(.a(output_3_322), .b(output_3_2), .y(output_2_322));
wire output_1_323, output_1_0, output_0_323;
mixer gate_output_0_323(.a(output_1_323), .b(output_1_0), .y(output_0_323));
wire output_2_323, output_2_0, output_1_323;
mixer gate_output_1_323(.a(output_2_323), .b(output_2_0), .y(output_1_323));
wire output_3_323, output_3_0, output_2_323;
mixer gate_output_2_323(.a(output_3_323), .b(output_3_0), .y(output_2_323));
wire output_1_324, output_1_1, output_0_324;
mixer gate_output_0_324(.a(output_1_324), .b(output_1_1), .y(output_0_324));
wire output_2_324, output_2_1, output_1_324;
mixer gate_output_1_324(.a(output_2_324), .b(output_2_1), .y(output_1_324));
wire output_3_324, output_3_1, output_2_324;
mixer gate_output_2_324(.a(output_3_324), .b(output_3_1), .y(output_2_324));
wire output_1_325, output_1_2, output_0_325;
mixer gate_output_0_325(.a(output_1_325), .b(output_1_2), .y(output_0_325));
wire output_2_325, output_2_2, output_1_325;
mixer gate_output_1_325(.a(output_2_325), .b(output_2_2), .y(output_1_325));
wire output_3_325, output_3_2, output_2_325;
mixer gate_output_2_325(.a(output_3_325), .b(output_3_2), .y(output_2_325));
wire output_1_326, output_1_0, output_0_326;
mixer gate_output_0_326(.a(output_1_326), .b(output_1_0), .y(output_0_326));
wire output_2_326, output_2_0, output_1_326;
mixer gate_output_1_326(.a(output_2_326), .b(output_2_0), .y(output_1_326));
wire output_3_326, output_3_0, output_2_326;
mixer gate_output_2_326(.a(output_3_326), .b(output_3_0), .y(output_2_326));
wire output_1_327, output_1_1, output_0_327;
mixer gate_output_0_327(.a(output_1_327), .b(output_1_1), .y(output_0_327));
wire output_2_327, output_2_1, output_1_327;
mixer gate_output_1_327(.a(output_2_327), .b(output_2_1), .y(output_1_327));
wire output_3_327, output_3_1, output_2_327;
mixer gate_output_2_327(.a(output_3_327), .b(output_3_1), .y(output_2_327));
wire output_1_328, output_1_2, output_0_328;
mixer gate_output_0_328(.a(output_1_328), .b(output_1_2), .y(output_0_328));
wire output_2_328, output_2_2, output_1_328;
mixer gate_output_1_328(.a(output_2_328), .b(output_2_2), .y(output_1_328));
wire output_3_328, output_3_2, output_2_328;
mixer gate_output_2_328(.a(output_3_328), .b(output_3_2), .y(output_2_328));
wire output_1_329, output_1_0, output_0_329;
mixer gate_output_0_329(.a(output_1_329), .b(output_1_0), .y(output_0_329));
wire output_2_329, output_2_0, output_1_329;
mixer gate_output_1_329(.a(output_2_329), .b(output_2_0), .y(output_1_329));
wire output_3_329, output_3_0, output_2_329;
mixer gate_output_2_329(.a(output_3_329), .b(output_3_0), .y(output_2_329));
wire output_1_330, output_1_1, output_0_330;
mixer gate_output_0_330(.a(output_1_330), .b(output_1_1), .y(output_0_330));
wire output_2_330, output_2_1, output_1_330;
mixer gate_output_1_330(.a(output_2_330), .b(output_2_1), .y(output_1_330));
wire output_3_330, output_3_1, output_2_330;
mixer gate_output_2_330(.a(output_3_330), .b(output_3_1), .y(output_2_330));
wire output_1_331, output_1_2, output_0_331;
mixer gate_output_0_331(.a(output_1_331), .b(output_1_2), .y(output_0_331));
wire output_2_331, output_2_2, output_1_331;
mixer gate_output_1_331(.a(output_2_331), .b(output_2_2), .y(output_1_331));
wire output_3_331, output_3_2, output_2_331;
mixer gate_output_2_331(.a(output_3_331), .b(output_3_2), .y(output_2_331));
wire output_1_332, output_1_0, output_0_332;
mixer gate_output_0_332(.a(output_1_332), .b(output_1_0), .y(output_0_332));
wire output_2_332, output_2_0, output_1_332;
mixer gate_output_1_332(.a(output_2_332), .b(output_2_0), .y(output_1_332));
wire output_3_332, output_3_0, output_2_332;
mixer gate_output_2_332(.a(output_3_332), .b(output_3_0), .y(output_2_332));
wire output_1_333, output_1_1, output_0_333;
mixer gate_output_0_333(.a(output_1_333), .b(output_1_1), .y(output_0_333));
wire output_2_333, output_2_1, output_1_333;
mixer gate_output_1_333(.a(output_2_333), .b(output_2_1), .y(output_1_333));
wire output_3_333, output_3_1, output_2_333;
mixer gate_output_2_333(.a(output_3_333), .b(output_3_1), .y(output_2_333));
wire output_1_334, output_1_2, output_0_334;
mixer gate_output_0_334(.a(output_1_334), .b(output_1_2), .y(output_0_334));
wire output_2_334, output_2_2, output_1_334;
mixer gate_output_1_334(.a(output_2_334), .b(output_2_2), .y(output_1_334));
wire output_3_334, output_3_2, output_2_334;
mixer gate_output_2_334(.a(output_3_334), .b(output_3_2), .y(output_2_334));
wire output_1_335, output_1_0, output_0_335;
mixer gate_output_0_335(.a(output_1_335), .b(output_1_0), .y(output_0_335));
wire output_2_335, output_2_0, output_1_335;
mixer gate_output_1_335(.a(output_2_335), .b(output_2_0), .y(output_1_335));
wire output_3_335, output_3_0, output_2_335;
mixer gate_output_2_335(.a(output_3_335), .b(output_3_0), .y(output_2_335));
wire output_1_336, output_1_1, output_0_336;
mixer gate_output_0_336(.a(output_1_336), .b(output_1_1), .y(output_0_336));
wire output_2_336, output_2_1, output_1_336;
mixer gate_output_1_336(.a(output_2_336), .b(output_2_1), .y(output_1_336));
wire output_3_336, output_3_1, output_2_336;
mixer gate_output_2_336(.a(output_3_336), .b(output_3_1), .y(output_2_336));
wire output_1_337, output_1_2, output_0_337;
mixer gate_output_0_337(.a(output_1_337), .b(output_1_2), .y(output_0_337));
wire output_2_337, output_2_2, output_1_337;
mixer gate_output_1_337(.a(output_2_337), .b(output_2_2), .y(output_1_337));
wire output_3_337, output_3_2, output_2_337;
mixer gate_output_2_337(.a(output_3_337), .b(output_3_2), .y(output_2_337));
wire output_1_338, output_1_0, output_0_338;
mixer gate_output_0_338(.a(output_1_338), .b(output_1_0), .y(output_0_338));
wire output_2_338, output_2_0, output_1_338;
mixer gate_output_1_338(.a(output_2_338), .b(output_2_0), .y(output_1_338));
wire output_3_338, output_3_0, output_2_338;
mixer gate_output_2_338(.a(output_3_338), .b(output_3_0), .y(output_2_338));
wire output_1_339, output_1_1, output_0_339;
mixer gate_output_0_339(.a(output_1_339), .b(output_1_1), .y(output_0_339));
wire output_2_339, output_2_1, output_1_339;
mixer gate_output_1_339(.a(output_2_339), .b(output_2_1), .y(output_1_339));
wire output_3_339, output_3_1, output_2_339;
mixer gate_output_2_339(.a(output_3_339), .b(output_3_1), .y(output_2_339));
wire output_1_340, output_1_2, output_0_340;
mixer gate_output_0_340(.a(output_1_340), .b(output_1_2), .y(output_0_340));
wire output_2_340, output_2_2, output_1_340;
mixer gate_output_1_340(.a(output_2_340), .b(output_2_2), .y(output_1_340));
wire output_3_340, output_3_2, output_2_340;
mixer gate_output_2_340(.a(output_3_340), .b(output_3_2), .y(output_2_340));
wire output_1_341, output_1_0, output_0_341;
mixer gate_output_0_341(.a(output_1_341), .b(output_1_0), .y(output_0_341));
wire output_2_341, output_2_0, output_1_341;
mixer gate_output_1_341(.a(output_2_341), .b(output_2_0), .y(output_1_341));
wire output_3_341, output_3_0, output_2_341;
mixer gate_output_2_341(.a(output_3_341), .b(output_3_0), .y(output_2_341));
wire output_1_342, output_1_1, output_0_342;
mixer gate_output_0_342(.a(output_1_342), .b(output_1_1), .y(output_0_342));
wire output_2_342, output_2_1, output_1_342;
mixer gate_output_1_342(.a(output_2_342), .b(output_2_1), .y(output_1_342));
wire output_3_342, output_3_1, output_2_342;
mixer gate_output_2_342(.a(output_3_342), .b(output_3_1), .y(output_2_342));
wire output_1_343, output_1_2, output_0_343;
mixer gate_output_0_343(.a(output_1_343), .b(output_1_2), .y(output_0_343));
wire output_2_343, output_2_2, output_1_343;
mixer gate_output_1_343(.a(output_2_343), .b(output_2_2), .y(output_1_343));
wire output_3_343, output_3_2, output_2_343;
mixer gate_output_2_343(.a(output_3_343), .b(output_3_2), .y(output_2_343));
wire output_1_344, output_1_0, output_0_344;
mixer gate_output_0_344(.a(output_1_344), .b(output_1_0), .y(output_0_344));
wire output_2_344, output_2_0, output_1_344;
mixer gate_output_1_344(.a(output_2_344), .b(output_2_0), .y(output_1_344));
wire output_3_344, output_3_0, output_2_344;
mixer gate_output_2_344(.a(output_3_344), .b(output_3_0), .y(output_2_344));
wire output_1_345, output_1_1, output_0_345;
mixer gate_output_0_345(.a(output_1_345), .b(output_1_1), .y(output_0_345));
wire output_2_345, output_2_1, output_1_345;
mixer gate_output_1_345(.a(output_2_345), .b(output_2_1), .y(output_1_345));
wire output_3_345, output_3_1, output_2_345;
mixer gate_output_2_345(.a(output_3_345), .b(output_3_1), .y(output_2_345));
wire output_1_346, output_1_2, output_0_346;
mixer gate_output_0_346(.a(output_1_346), .b(output_1_2), .y(output_0_346));
wire output_2_346, output_2_2, output_1_346;
mixer gate_output_1_346(.a(output_2_346), .b(output_2_2), .y(output_1_346));
wire output_3_346, output_3_2, output_2_346;
mixer gate_output_2_346(.a(output_3_346), .b(output_3_2), .y(output_2_346));
wire output_1_347, output_1_0, output_0_347;
mixer gate_output_0_347(.a(output_1_347), .b(output_1_0), .y(output_0_347));
wire output_2_347, output_2_0, output_1_347;
mixer gate_output_1_347(.a(output_2_347), .b(output_2_0), .y(output_1_347));
wire output_3_347, output_3_0, output_2_347;
mixer gate_output_2_347(.a(output_3_347), .b(output_3_0), .y(output_2_347));
wire output_1_348, output_1_1, output_0_348;
mixer gate_output_0_348(.a(output_1_348), .b(output_1_1), .y(output_0_348));
wire output_2_348, output_2_1, output_1_348;
mixer gate_output_1_348(.a(output_2_348), .b(output_2_1), .y(output_1_348));
wire output_3_348, output_3_1, output_2_348;
mixer gate_output_2_348(.a(output_3_348), .b(output_3_1), .y(output_2_348));
wire output_1_349, output_1_2, output_0_349;
mixer gate_output_0_349(.a(output_1_349), .b(output_1_2), .y(output_0_349));
wire output_2_349, output_2_2, output_1_349;
mixer gate_output_1_349(.a(output_2_349), .b(output_2_2), .y(output_1_349));
wire output_3_349, output_3_2, output_2_349;
mixer gate_output_2_349(.a(output_3_349), .b(output_3_2), .y(output_2_349));
wire output_1_350, output_1_0, output_0_350;
mixer gate_output_0_350(.a(output_1_350), .b(output_1_0), .y(output_0_350));
wire output_2_350, output_2_0, output_1_350;
mixer gate_output_1_350(.a(output_2_350), .b(output_2_0), .y(output_1_350));
wire output_3_350, output_3_0, output_2_350;
mixer gate_output_2_350(.a(output_3_350), .b(output_3_0), .y(output_2_350));
wire output_1_351, output_1_1, output_0_351;
mixer gate_output_0_351(.a(output_1_351), .b(output_1_1), .y(output_0_351));
wire output_2_351, output_2_1, output_1_351;
mixer gate_output_1_351(.a(output_2_351), .b(output_2_1), .y(output_1_351));
wire output_3_351, output_3_1, output_2_351;
mixer gate_output_2_351(.a(output_3_351), .b(output_3_1), .y(output_2_351));
wire output_1_352, output_1_2, output_0_352;
mixer gate_output_0_352(.a(output_1_352), .b(output_1_2), .y(output_0_352));
wire output_2_352, output_2_2, output_1_352;
mixer gate_output_1_352(.a(output_2_352), .b(output_2_2), .y(output_1_352));
wire output_3_352, output_3_2, output_2_352;
mixer gate_output_2_352(.a(output_3_352), .b(output_3_2), .y(output_2_352));
wire output_1_353, output_1_0, output_0_353;
mixer gate_output_0_353(.a(output_1_353), .b(output_1_0), .y(output_0_353));
wire output_2_353, output_2_0, output_1_353;
mixer gate_output_1_353(.a(output_2_353), .b(output_2_0), .y(output_1_353));
wire output_3_353, output_3_0, output_2_353;
mixer gate_output_2_353(.a(output_3_353), .b(output_3_0), .y(output_2_353));
wire output_1_354, output_1_1, output_0_354;
mixer gate_output_0_354(.a(output_1_354), .b(output_1_1), .y(output_0_354));
wire output_2_354, output_2_1, output_1_354;
mixer gate_output_1_354(.a(output_2_354), .b(output_2_1), .y(output_1_354));
wire output_3_354, output_3_1, output_2_354;
mixer gate_output_2_354(.a(output_3_354), .b(output_3_1), .y(output_2_354));
wire output_1_355, output_1_2, output_0_355;
mixer gate_output_0_355(.a(output_1_355), .b(output_1_2), .y(output_0_355));
wire output_2_355, output_2_2, output_1_355;
mixer gate_output_1_355(.a(output_2_355), .b(output_2_2), .y(output_1_355));
wire output_3_355, output_3_2, output_2_355;
mixer gate_output_2_355(.a(output_3_355), .b(output_3_2), .y(output_2_355));
wire output_1_356, output_1_0, output_0_356;
mixer gate_output_0_356(.a(output_1_356), .b(output_1_0), .y(output_0_356));
wire output_2_356, output_2_0, output_1_356;
mixer gate_output_1_356(.a(output_2_356), .b(output_2_0), .y(output_1_356));
wire output_3_356, output_3_0, output_2_356;
mixer gate_output_2_356(.a(output_3_356), .b(output_3_0), .y(output_2_356));
wire output_1_357, output_1_1, output_0_357;
mixer gate_output_0_357(.a(output_1_357), .b(output_1_1), .y(output_0_357));
wire output_2_357, output_2_1, output_1_357;
mixer gate_output_1_357(.a(output_2_357), .b(output_2_1), .y(output_1_357));
wire output_3_357, output_3_1, output_2_357;
mixer gate_output_2_357(.a(output_3_357), .b(output_3_1), .y(output_2_357));
wire output_1_358, output_1_2, output_0_358;
mixer gate_output_0_358(.a(output_1_358), .b(output_1_2), .y(output_0_358));
wire output_2_358, output_2_2, output_1_358;
mixer gate_output_1_358(.a(output_2_358), .b(output_2_2), .y(output_1_358));
wire output_3_358, output_3_2, output_2_358;
mixer gate_output_2_358(.a(output_3_358), .b(output_3_2), .y(output_2_358));
wire output_1_359, output_1_0, output_0_359;
mixer gate_output_0_359(.a(output_1_359), .b(output_1_0), .y(output_0_359));
wire output_2_359, output_2_0, output_1_359;
mixer gate_output_1_359(.a(output_2_359), .b(output_2_0), .y(output_1_359));
wire output_3_359, output_3_0, output_2_359;
mixer gate_output_2_359(.a(output_3_359), .b(output_3_0), .y(output_2_359));
wire output_1_360, output_1_1, output_0_360;
mixer gate_output_0_360(.a(output_1_360), .b(output_1_1), .y(output_0_360));
wire output_2_360, output_2_1, output_1_360;
mixer gate_output_1_360(.a(output_2_360), .b(output_2_1), .y(output_1_360));
wire output_3_360, output_3_1, output_2_360;
mixer gate_output_2_360(.a(output_3_360), .b(output_3_1), .y(output_2_360));
wire output_1_361, output_1_2, output_0_361;
mixer gate_output_0_361(.a(output_1_361), .b(output_1_2), .y(output_0_361));
wire output_2_361, output_2_2, output_1_361;
mixer gate_output_1_361(.a(output_2_361), .b(output_2_2), .y(output_1_361));
wire output_3_361, output_3_2, output_2_361;
mixer gate_output_2_361(.a(output_3_361), .b(output_3_2), .y(output_2_361));
wire output_1_362, output_1_0, output_0_362;
mixer gate_output_0_362(.a(output_1_362), .b(output_1_0), .y(output_0_362));
wire output_2_362, output_2_0, output_1_362;
mixer gate_output_1_362(.a(output_2_362), .b(output_2_0), .y(output_1_362));
wire output_3_362, output_3_0, output_2_362;
mixer gate_output_2_362(.a(output_3_362), .b(output_3_0), .y(output_2_362));
wire output_1_363, output_1_1, output_0_363;
mixer gate_output_0_363(.a(output_1_363), .b(output_1_1), .y(output_0_363));
wire output_2_363, output_2_1, output_1_363;
mixer gate_output_1_363(.a(output_2_363), .b(output_2_1), .y(output_1_363));
wire output_3_363, output_3_1, output_2_363;
mixer gate_output_2_363(.a(output_3_363), .b(output_3_1), .y(output_2_363));
wire output_1_364, output_1_2, output_0_364;
mixer gate_output_0_364(.a(output_1_364), .b(output_1_2), .y(output_0_364));
wire output_2_364, output_2_2, output_1_364;
mixer gate_output_1_364(.a(output_2_364), .b(output_2_2), .y(output_1_364));
wire output_3_364, output_3_2, output_2_364;
mixer gate_output_2_364(.a(output_3_364), .b(output_3_2), .y(output_2_364));
wire output_1_365, output_1_0, output_0_365;
mixer gate_output_0_365(.a(output_1_365), .b(output_1_0), .y(output_0_365));
wire output_2_365, output_2_0, output_1_365;
mixer gate_output_1_365(.a(output_2_365), .b(output_2_0), .y(output_1_365));
wire output_3_365, output_3_0, output_2_365;
mixer gate_output_2_365(.a(output_3_365), .b(output_3_0), .y(output_2_365));
wire output_1_366, output_1_1, output_0_366;
mixer gate_output_0_366(.a(output_1_366), .b(output_1_1), .y(output_0_366));
wire output_2_366, output_2_1, output_1_366;
mixer gate_output_1_366(.a(output_2_366), .b(output_2_1), .y(output_1_366));
wire output_3_366, output_3_1, output_2_366;
mixer gate_output_2_366(.a(output_3_366), .b(output_3_1), .y(output_2_366));
wire output_1_367, output_1_2, output_0_367;
mixer gate_output_0_367(.a(output_1_367), .b(output_1_2), .y(output_0_367));
wire output_2_367, output_2_2, output_1_367;
mixer gate_output_1_367(.a(output_2_367), .b(output_2_2), .y(output_1_367));
wire output_3_367, output_3_2, output_2_367;
mixer gate_output_2_367(.a(output_3_367), .b(output_3_2), .y(output_2_367));
wire output_1_368, output_1_0, output_0_368;
mixer gate_output_0_368(.a(output_1_368), .b(output_1_0), .y(output_0_368));
wire output_2_368, output_2_0, output_1_368;
mixer gate_output_1_368(.a(output_2_368), .b(output_2_0), .y(output_1_368));
wire output_3_368, output_3_0, output_2_368;
mixer gate_output_2_368(.a(output_3_368), .b(output_3_0), .y(output_2_368));
wire output_1_369, output_1_1, output_0_369;
mixer gate_output_0_369(.a(output_1_369), .b(output_1_1), .y(output_0_369));
wire output_2_369, output_2_1, output_1_369;
mixer gate_output_1_369(.a(output_2_369), .b(output_2_1), .y(output_1_369));
wire output_3_369, output_3_1, output_2_369;
mixer gate_output_2_369(.a(output_3_369), .b(output_3_1), .y(output_2_369));
wire output_1_370, output_1_2, output_0_370;
mixer gate_output_0_370(.a(output_1_370), .b(output_1_2), .y(output_0_370));
wire output_2_370, output_2_2, output_1_370;
mixer gate_output_1_370(.a(output_2_370), .b(output_2_2), .y(output_1_370));
wire output_3_370, output_3_2, output_2_370;
mixer gate_output_2_370(.a(output_3_370), .b(output_3_2), .y(output_2_370));
wire output_1_371, output_1_0, output_0_371;
mixer gate_output_0_371(.a(output_1_371), .b(output_1_0), .y(output_0_371));
wire output_2_371, output_2_0, output_1_371;
mixer gate_output_1_371(.a(output_2_371), .b(output_2_0), .y(output_1_371));
wire output_3_371, output_3_0, output_2_371;
mixer gate_output_2_371(.a(output_3_371), .b(output_3_0), .y(output_2_371));
wire output_1_372, output_1_1, output_0_372;
mixer gate_output_0_372(.a(output_1_372), .b(output_1_1), .y(output_0_372));
wire output_2_372, output_2_1, output_1_372;
mixer gate_output_1_372(.a(output_2_372), .b(output_2_1), .y(output_1_372));
wire output_3_372, output_3_1, output_2_372;
mixer gate_output_2_372(.a(output_3_372), .b(output_3_1), .y(output_2_372));
wire output_1_373, output_1_2, output_0_373;
mixer gate_output_0_373(.a(output_1_373), .b(output_1_2), .y(output_0_373));
wire output_2_373, output_2_2, output_1_373;
mixer gate_output_1_373(.a(output_2_373), .b(output_2_2), .y(output_1_373));
wire output_3_373, output_3_2, output_2_373;
mixer gate_output_2_373(.a(output_3_373), .b(output_3_2), .y(output_2_373));
wire output_1_374, output_1_0, output_0_374;
mixer gate_output_0_374(.a(output_1_374), .b(output_1_0), .y(output_0_374));
wire output_2_374, output_2_0, output_1_374;
mixer gate_output_1_374(.a(output_2_374), .b(output_2_0), .y(output_1_374));
wire output_3_374, output_3_0, output_2_374;
mixer gate_output_2_374(.a(output_3_374), .b(output_3_0), .y(output_2_374));
wire output_1_375, output_1_1, output_0_375;
mixer gate_output_0_375(.a(output_1_375), .b(output_1_1), .y(output_0_375));
wire output_2_375, output_2_1, output_1_375;
mixer gate_output_1_375(.a(output_2_375), .b(output_2_1), .y(output_1_375));
wire output_3_375, output_3_1, output_2_375;
mixer gate_output_2_375(.a(output_3_375), .b(output_3_1), .y(output_2_375));
wire output_1_376, output_1_2, output_0_376;
mixer gate_output_0_376(.a(output_1_376), .b(output_1_2), .y(output_0_376));
wire output_2_376, output_2_2, output_1_376;
mixer gate_output_1_376(.a(output_2_376), .b(output_2_2), .y(output_1_376));
wire output_3_376, output_3_2, output_2_376;
mixer gate_output_2_376(.a(output_3_376), .b(output_3_2), .y(output_2_376));
wire output_1_377, output_1_0, output_0_377;
mixer gate_output_0_377(.a(output_1_377), .b(output_1_0), .y(output_0_377));
wire output_2_377, output_2_0, output_1_377;
mixer gate_output_1_377(.a(output_2_377), .b(output_2_0), .y(output_1_377));
wire output_3_377, output_3_0, output_2_377;
mixer gate_output_2_377(.a(output_3_377), .b(output_3_0), .y(output_2_377));
wire output_1_378, output_1_1, output_0_378;
mixer gate_output_0_378(.a(output_1_378), .b(output_1_1), .y(output_0_378));
wire output_2_378, output_2_1, output_1_378;
mixer gate_output_1_378(.a(output_2_378), .b(output_2_1), .y(output_1_378));
wire output_3_378, output_3_1, output_2_378;
mixer gate_output_2_378(.a(output_3_378), .b(output_3_1), .y(output_2_378));
wire output_1_379, output_1_2, output_0_379;
mixer gate_output_0_379(.a(output_1_379), .b(output_1_2), .y(output_0_379));
wire output_2_379, output_2_2, output_1_379;
mixer gate_output_1_379(.a(output_2_379), .b(output_2_2), .y(output_1_379));
wire output_3_379, output_3_2, output_2_379;
mixer gate_output_2_379(.a(output_3_379), .b(output_3_2), .y(output_2_379));
wire output_1_380, output_1_0, output_0_380;
mixer gate_output_0_380(.a(output_1_380), .b(output_1_0), .y(output_0_380));
wire output_2_380, output_2_0, output_1_380;
mixer gate_output_1_380(.a(output_2_380), .b(output_2_0), .y(output_1_380));
wire output_3_380, output_3_0, output_2_380;
mixer gate_output_2_380(.a(output_3_380), .b(output_3_0), .y(output_2_380));
wire output_1_381, output_1_1, output_0_381;
mixer gate_output_0_381(.a(output_1_381), .b(output_1_1), .y(output_0_381));
wire output_2_381, output_2_1, output_1_381;
mixer gate_output_1_381(.a(output_2_381), .b(output_2_1), .y(output_1_381));
wire output_3_381, output_3_1, output_2_381;
mixer gate_output_2_381(.a(output_3_381), .b(output_3_1), .y(output_2_381));
wire output_1_382, output_1_2, output_0_382;
mixer gate_output_0_382(.a(output_1_382), .b(output_1_2), .y(output_0_382));
wire output_2_382, output_2_2, output_1_382;
mixer gate_output_1_382(.a(output_2_382), .b(output_2_2), .y(output_1_382));
wire output_3_382, output_3_2, output_2_382;
mixer gate_output_2_382(.a(output_3_382), .b(output_3_2), .y(output_2_382));
wire output_1_383, output_1_0, output_0_383;
mixer gate_output_0_383(.a(output_1_383), .b(output_1_0), .y(output_0_383));
wire output_2_383, output_2_0, output_1_383;
mixer gate_output_1_383(.a(output_2_383), .b(output_2_0), .y(output_1_383));
wire output_3_383, output_3_0, output_2_383;
mixer gate_output_2_383(.a(output_3_383), .b(output_3_0), .y(output_2_383));
wire output_1_384, output_1_1, output_0_384;
mixer gate_output_0_384(.a(output_1_384), .b(output_1_1), .y(output_0_384));
wire output_2_384, output_2_1, output_1_384;
mixer gate_output_1_384(.a(output_2_384), .b(output_2_1), .y(output_1_384));
wire output_3_384, output_3_1, output_2_384;
mixer gate_output_2_384(.a(output_3_384), .b(output_3_1), .y(output_2_384));
wire output_1_385, output_1_2, output_0_385;
mixer gate_output_0_385(.a(output_1_385), .b(output_1_2), .y(output_0_385));
wire output_2_385, output_2_2, output_1_385;
mixer gate_output_1_385(.a(output_2_385), .b(output_2_2), .y(output_1_385));
wire output_3_385, output_3_2, output_2_385;
mixer gate_output_2_385(.a(output_3_385), .b(output_3_2), .y(output_2_385));
wire output_1_386, output_1_0, output_0_386;
mixer gate_output_0_386(.a(output_1_386), .b(output_1_0), .y(output_0_386));
wire output_2_386, output_2_0, output_1_386;
mixer gate_output_1_386(.a(output_2_386), .b(output_2_0), .y(output_1_386));
wire output_3_386, output_3_0, output_2_386;
mixer gate_output_2_386(.a(output_3_386), .b(output_3_0), .y(output_2_386));
wire output_1_387, output_1_1, output_0_387;
mixer gate_output_0_387(.a(output_1_387), .b(output_1_1), .y(output_0_387));
wire output_2_387, output_2_1, output_1_387;
mixer gate_output_1_387(.a(output_2_387), .b(output_2_1), .y(output_1_387));
wire output_3_387, output_3_1, output_2_387;
mixer gate_output_2_387(.a(output_3_387), .b(output_3_1), .y(output_2_387));
wire output_1_388, output_1_2, output_0_388;
mixer gate_output_0_388(.a(output_1_388), .b(output_1_2), .y(output_0_388));
wire output_2_388, output_2_2, output_1_388;
mixer gate_output_1_388(.a(output_2_388), .b(output_2_2), .y(output_1_388));
wire output_3_388, output_3_2, output_2_388;
mixer gate_output_2_388(.a(output_3_388), .b(output_3_2), .y(output_2_388));
wire output_1_389, output_1_0, output_0_389;
mixer gate_output_0_389(.a(output_1_389), .b(output_1_0), .y(output_0_389));
wire output_2_389, output_2_0, output_1_389;
mixer gate_output_1_389(.a(output_2_389), .b(output_2_0), .y(output_1_389));
wire output_3_389, output_3_0, output_2_389;
mixer gate_output_2_389(.a(output_3_389), .b(output_3_0), .y(output_2_389));
wire output_1_390, output_1_1, output_0_390;
mixer gate_output_0_390(.a(output_1_390), .b(output_1_1), .y(output_0_390));
wire output_2_390, output_2_1, output_1_390;
mixer gate_output_1_390(.a(output_2_390), .b(output_2_1), .y(output_1_390));
wire output_3_390, output_3_1, output_2_390;
mixer gate_output_2_390(.a(output_3_390), .b(output_3_1), .y(output_2_390));
wire output_1_391, output_1_2, output_0_391;
mixer gate_output_0_391(.a(output_1_391), .b(output_1_2), .y(output_0_391));
wire output_2_391, output_2_2, output_1_391;
mixer gate_output_1_391(.a(output_2_391), .b(output_2_2), .y(output_1_391));
wire output_3_391, output_3_2, output_2_391;
mixer gate_output_2_391(.a(output_3_391), .b(output_3_2), .y(output_2_391));
wire output_1_392, output_1_0, output_0_392;
mixer gate_output_0_392(.a(output_1_392), .b(output_1_0), .y(output_0_392));
wire output_2_392, output_2_0, output_1_392;
mixer gate_output_1_392(.a(output_2_392), .b(output_2_0), .y(output_1_392));
wire output_3_392, output_3_0, output_2_392;
mixer gate_output_2_392(.a(output_3_392), .b(output_3_0), .y(output_2_392));
wire output_1_393, output_1_1, output_0_393;
mixer gate_output_0_393(.a(output_1_393), .b(output_1_1), .y(output_0_393));
wire output_2_393, output_2_1, output_1_393;
mixer gate_output_1_393(.a(output_2_393), .b(output_2_1), .y(output_1_393));
wire output_3_393, output_3_1, output_2_393;
mixer gate_output_2_393(.a(output_3_393), .b(output_3_1), .y(output_2_393));
wire output_1_394, output_1_2, output_0_394;
mixer gate_output_0_394(.a(output_1_394), .b(output_1_2), .y(output_0_394));
wire output_2_394, output_2_2, output_1_394;
mixer gate_output_1_394(.a(output_2_394), .b(output_2_2), .y(output_1_394));
wire output_3_394, output_3_2, output_2_394;
mixer gate_output_2_394(.a(output_3_394), .b(output_3_2), .y(output_2_394));
wire output_1_395, output_1_0, output_0_395;
mixer gate_output_0_395(.a(output_1_395), .b(output_1_0), .y(output_0_395));
wire output_2_395, output_2_0, output_1_395;
mixer gate_output_1_395(.a(output_2_395), .b(output_2_0), .y(output_1_395));
wire output_3_395, output_3_0, output_2_395;
mixer gate_output_2_395(.a(output_3_395), .b(output_3_0), .y(output_2_395));
wire output_1_396, output_1_1, output_0_396;
mixer gate_output_0_396(.a(output_1_396), .b(output_1_1), .y(output_0_396));
wire output_2_396, output_2_1, output_1_396;
mixer gate_output_1_396(.a(output_2_396), .b(output_2_1), .y(output_1_396));
wire output_3_396, output_3_1, output_2_396;
mixer gate_output_2_396(.a(output_3_396), .b(output_3_1), .y(output_2_396));
wire output_1_397, output_1_2, output_0_397;
mixer gate_output_0_397(.a(output_1_397), .b(output_1_2), .y(output_0_397));
wire output_2_397, output_2_2, output_1_397;
mixer gate_output_1_397(.a(output_2_397), .b(output_2_2), .y(output_1_397));
wire output_3_397, output_3_2, output_2_397;
mixer gate_output_2_397(.a(output_3_397), .b(output_3_2), .y(output_2_397));
wire output_1_398, output_1_0, output_0_398;
mixer gate_output_0_398(.a(output_1_398), .b(output_1_0), .y(output_0_398));
wire output_2_398, output_2_0, output_1_398;
mixer gate_output_1_398(.a(output_2_398), .b(output_2_0), .y(output_1_398));
wire output_3_398, output_3_0, output_2_398;
mixer gate_output_2_398(.a(output_3_398), .b(output_3_0), .y(output_2_398));
wire output_1_399, output_1_1, output_0_399;
mixer gate_output_0_399(.a(output_1_399), .b(output_1_1), .y(output_0_399));
wire output_2_399, output_2_1, output_1_399;
mixer gate_output_1_399(.a(output_2_399), .b(output_2_1), .y(output_1_399));
wire output_3_399, output_3_1, output_2_399;
mixer gate_output_2_399(.a(output_3_399), .b(output_3_1), .y(output_2_399));
wire output_1_400, output_1_2, output_0_400;
mixer gate_output_0_400(.a(output_1_400), .b(output_1_2), .y(output_0_400));
wire output_2_400, output_2_2, output_1_400;
mixer gate_output_1_400(.a(output_2_400), .b(output_2_2), .y(output_1_400));
wire output_3_400, output_3_2, output_2_400;
mixer gate_output_2_400(.a(output_3_400), .b(output_3_2), .y(output_2_400));
wire output_1_401, output_1_0, output_0_401;
mixer gate_output_0_401(.a(output_1_401), .b(output_1_0), .y(output_0_401));
wire output_2_401, output_2_0, output_1_401;
mixer gate_output_1_401(.a(output_2_401), .b(output_2_0), .y(output_1_401));
wire output_3_401, output_3_0, output_2_401;
mixer gate_output_2_401(.a(output_3_401), .b(output_3_0), .y(output_2_401));
wire output_1_402, output_1_1, output_0_402;
mixer gate_output_0_402(.a(output_1_402), .b(output_1_1), .y(output_0_402));
wire output_2_402, output_2_1, output_1_402;
mixer gate_output_1_402(.a(output_2_402), .b(output_2_1), .y(output_1_402));
wire output_3_402, output_3_1, output_2_402;
mixer gate_output_2_402(.a(output_3_402), .b(output_3_1), .y(output_2_402));
wire output_1_403, output_1_2, output_0_403;
mixer gate_output_0_403(.a(output_1_403), .b(output_1_2), .y(output_0_403));
wire output_2_403, output_2_2, output_1_403;
mixer gate_output_1_403(.a(output_2_403), .b(output_2_2), .y(output_1_403));
wire output_3_403, output_3_2, output_2_403;
mixer gate_output_2_403(.a(output_3_403), .b(output_3_2), .y(output_2_403));
wire output_1_404, output_1_0, output_0_404;
mixer gate_output_0_404(.a(output_1_404), .b(output_1_0), .y(output_0_404));
wire output_2_404, output_2_0, output_1_404;
mixer gate_output_1_404(.a(output_2_404), .b(output_2_0), .y(output_1_404));
wire output_3_404, output_3_0, output_2_404;
mixer gate_output_2_404(.a(output_3_404), .b(output_3_0), .y(output_2_404));
wire output_1_405, output_1_1, output_0_405;
mixer gate_output_0_405(.a(output_1_405), .b(output_1_1), .y(output_0_405));
wire output_2_405, output_2_1, output_1_405;
mixer gate_output_1_405(.a(output_2_405), .b(output_2_1), .y(output_1_405));
wire output_3_405, output_3_1, output_2_405;
mixer gate_output_2_405(.a(output_3_405), .b(output_3_1), .y(output_2_405));
wire output_1_406, output_1_2, output_0_406;
mixer gate_output_0_406(.a(output_1_406), .b(output_1_2), .y(output_0_406));
wire output_2_406, output_2_2, output_1_406;
mixer gate_output_1_406(.a(output_2_406), .b(output_2_2), .y(output_1_406));
wire output_3_406, output_3_2, output_2_406;
mixer gate_output_2_406(.a(output_3_406), .b(output_3_2), .y(output_2_406));
wire output_1_407, output_1_0, output_0_407;
mixer gate_output_0_407(.a(output_1_407), .b(output_1_0), .y(output_0_407));
wire output_2_407, output_2_0, output_1_407;
mixer gate_output_1_407(.a(output_2_407), .b(output_2_0), .y(output_1_407));
wire output_3_407, output_3_0, output_2_407;
mixer gate_output_2_407(.a(output_3_407), .b(output_3_0), .y(output_2_407));
wire output_1_408, output_1_1, output_0_408;
mixer gate_output_0_408(.a(output_1_408), .b(output_1_1), .y(output_0_408));
wire output_2_408, output_2_1, output_1_408;
mixer gate_output_1_408(.a(output_2_408), .b(output_2_1), .y(output_1_408));
wire output_3_408, output_3_1, output_2_408;
mixer gate_output_2_408(.a(output_3_408), .b(output_3_1), .y(output_2_408));
wire output_1_409, output_1_2, output_0_409;
mixer gate_output_0_409(.a(output_1_409), .b(output_1_2), .y(output_0_409));
wire output_2_409, output_2_2, output_1_409;
mixer gate_output_1_409(.a(output_2_409), .b(output_2_2), .y(output_1_409));
wire output_3_409, output_3_2, output_2_409;
mixer gate_output_2_409(.a(output_3_409), .b(output_3_2), .y(output_2_409));
wire output_1_410, output_1_0, output_0_410;
mixer gate_output_0_410(.a(output_1_410), .b(output_1_0), .y(output_0_410));
wire output_2_410, output_2_0, output_1_410;
mixer gate_output_1_410(.a(output_2_410), .b(output_2_0), .y(output_1_410));
wire output_3_410, output_3_0, output_2_410;
mixer gate_output_2_410(.a(output_3_410), .b(output_3_0), .y(output_2_410));
wire output_1_411, output_1_1, output_0_411;
mixer gate_output_0_411(.a(output_1_411), .b(output_1_1), .y(output_0_411));
wire output_2_411, output_2_1, output_1_411;
mixer gate_output_1_411(.a(output_2_411), .b(output_2_1), .y(output_1_411));
wire output_3_411, output_3_1, output_2_411;
mixer gate_output_2_411(.a(output_3_411), .b(output_3_1), .y(output_2_411));
wire output_1_412, output_1_2, output_0_412;
mixer gate_output_0_412(.a(output_1_412), .b(output_1_2), .y(output_0_412));
wire output_2_412, output_2_2, output_1_412;
mixer gate_output_1_412(.a(output_2_412), .b(output_2_2), .y(output_1_412));
wire output_3_412, output_3_2, output_2_412;
mixer gate_output_2_412(.a(output_3_412), .b(output_3_2), .y(output_2_412));
wire output_1_413, output_1_0, output_0_413;
mixer gate_output_0_413(.a(output_1_413), .b(output_1_0), .y(output_0_413));
wire output_2_413, output_2_0, output_1_413;
mixer gate_output_1_413(.a(output_2_413), .b(output_2_0), .y(output_1_413));
wire output_3_413, output_3_0, output_2_413;
mixer gate_output_2_413(.a(output_3_413), .b(output_3_0), .y(output_2_413));
wire output_1_414, output_1_1, output_0_414;
mixer gate_output_0_414(.a(output_1_414), .b(output_1_1), .y(output_0_414));
wire output_2_414, output_2_1, output_1_414;
mixer gate_output_1_414(.a(output_2_414), .b(output_2_1), .y(output_1_414));
wire output_3_414, output_3_1, output_2_414;
mixer gate_output_2_414(.a(output_3_414), .b(output_3_1), .y(output_2_414));
wire output_1_415, output_1_2, output_0_415;
mixer gate_output_0_415(.a(output_1_415), .b(output_1_2), .y(output_0_415));
wire output_2_415, output_2_2, output_1_415;
mixer gate_output_1_415(.a(output_2_415), .b(output_2_2), .y(output_1_415));
wire output_3_415, output_3_2, output_2_415;
mixer gate_output_2_415(.a(output_3_415), .b(output_3_2), .y(output_2_415));
wire output_1_416, output_1_0, output_0_416;
mixer gate_output_0_416(.a(output_1_416), .b(output_1_0), .y(output_0_416));
wire output_2_416, output_2_0, output_1_416;
mixer gate_output_1_416(.a(output_2_416), .b(output_2_0), .y(output_1_416));
wire output_3_416, output_3_0, output_2_416;
mixer gate_output_2_416(.a(output_3_416), .b(output_3_0), .y(output_2_416));
wire output_1_417, output_1_1, output_0_417;
mixer gate_output_0_417(.a(output_1_417), .b(output_1_1), .y(output_0_417));
wire output_2_417, output_2_1, output_1_417;
mixer gate_output_1_417(.a(output_2_417), .b(output_2_1), .y(output_1_417));
wire output_3_417, output_3_1, output_2_417;
mixer gate_output_2_417(.a(output_3_417), .b(output_3_1), .y(output_2_417));
wire output_1_418, output_1_2, output_0_418;
mixer gate_output_0_418(.a(output_1_418), .b(output_1_2), .y(output_0_418));
wire output_2_418, output_2_2, output_1_418;
mixer gate_output_1_418(.a(output_2_418), .b(output_2_2), .y(output_1_418));
wire output_3_418, output_3_2, output_2_418;
mixer gate_output_2_418(.a(output_3_418), .b(output_3_2), .y(output_2_418));
wire output_1_419, output_1_0, output_0_419;
mixer gate_output_0_419(.a(output_1_419), .b(output_1_0), .y(output_0_419));
wire output_2_419, output_2_0, output_1_419;
mixer gate_output_1_419(.a(output_2_419), .b(output_2_0), .y(output_1_419));
wire output_3_419, output_3_0, output_2_419;
mixer gate_output_2_419(.a(output_3_419), .b(output_3_0), .y(output_2_419));
wire output_1_420, output_1_1, output_0_420;
mixer gate_output_0_420(.a(output_1_420), .b(output_1_1), .y(output_0_420));
wire output_2_420, output_2_1, output_1_420;
mixer gate_output_1_420(.a(output_2_420), .b(output_2_1), .y(output_1_420));
wire output_3_420, output_3_1, output_2_420;
mixer gate_output_2_420(.a(output_3_420), .b(output_3_1), .y(output_2_420));
wire output_1_421, output_1_2, output_0_421;
mixer gate_output_0_421(.a(output_1_421), .b(output_1_2), .y(output_0_421));
wire output_2_421, output_2_2, output_1_421;
mixer gate_output_1_421(.a(output_2_421), .b(output_2_2), .y(output_1_421));
wire output_3_421, output_3_2, output_2_421;
mixer gate_output_2_421(.a(output_3_421), .b(output_3_2), .y(output_2_421));
wire output_1_422, output_1_0, output_0_422;
mixer gate_output_0_422(.a(output_1_422), .b(output_1_0), .y(output_0_422));
wire output_2_422, output_2_0, output_1_422;
mixer gate_output_1_422(.a(output_2_422), .b(output_2_0), .y(output_1_422));
wire output_3_422, output_3_0, output_2_422;
mixer gate_output_2_422(.a(output_3_422), .b(output_3_0), .y(output_2_422));
wire output_1_423, output_1_1, output_0_423;
mixer gate_output_0_423(.a(output_1_423), .b(output_1_1), .y(output_0_423));
wire output_2_423, output_2_1, output_1_423;
mixer gate_output_1_423(.a(output_2_423), .b(output_2_1), .y(output_1_423));
wire output_3_423, output_3_1, output_2_423;
mixer gate_output_2_423(.a(output_3_423), .b(output_3_1), .y(output_2_423));
wire output_1_424, output_1_2, output_0_424;
mixer gate_output_0_424(.a(output_1_424), .b(output_1_2), .y(output_0_424));
wire output_2_424, output_2_2, output_1_424;
mixer gate_output_1_424(.a(output_2_424), .b(output_2_2), .y(output_1_424));
wire output_3_424, output_3_2, output_2_424;
mixer gate_output_2_424(.a(output_3_424), .b(output_3_2), .y(output_2_424));
wire output_1_425, output_1_0, output_0_425;
mixer gate_output_0_425(.a(output_1_425), .b(output_1_0), .y(output_0_425));
wire output_2_425, output_2_0, output_1_425;
mixer gate_output_1_425(.a(output_2_425), .b(output_2_0), .y(output_1_425));
wire output_3_425, output_3_0, output_2_425;
mixer gate_output_2_425(.a(output_3_425), .b(output_3_0), .y(output_2_425));
wire output_1_426, output_1_1, output_0_426;
mixer gate_output_0_426(.a(output_1_426), .b(output_1_1), .y(output_0_426));
wire output_2_426, output_2_1, output_1_426;
mixer gate_output_1_426(.a(output_2_426), .b(output_2_1), .y(output_1_426));
wire output_3_426, output_3_1, output_2_426;
mixer gate_output_2_426(.a(output_3_426), .b(output_3_1), .y(output_2_426));
wire output_1_427, output_1_2, output_0_427;
mixer gate_output_0_427(.a(output_1_427), .b(output_1_2), .y(output_0_427));
wire output_2_427, output_2_2, output_1_427;
mixer gate_output_1_427(.a(output_2_427), .b(output_2_2), .y(output_1_427));
wire output_3_427, output_3_2, output_2_427;
mixer gate_output_2_427(.a(output_3_427), .b(output_3_2), .y(output_2_427));
wire output_1_428, output_1_0, output_0_428;
mixer gate_output_0_428(.a(output_1_428), .b(output_1_0), .y(output_0_428));
wire output_2_428, output_2_0, output_1_428;
mixer gate_output_1_428(.a(output_2_428), .b(output_2_0), .y(output_1_428));
wire output_3_428, output_3_0, output_2_428;
mixer gate_output_2_428(.a(output_3_428), .b(output_3_0), .y(output_2_428));
wire output_1_429, output_1_1, output_0_429;
mixer gate_output_0_429(.a(output_1_429), .b(output_1_1), .y(output_0_429));
wire output_2_429, output_2_1, output_1_429;
mixer gate_output_1_429(.a(output_2_429), .b(output_2_1), .y(output_1_429));
wire output_3_429, output_3_1, output_2_429;
mixer gate_output_2_429(.a(output_3_429), .b(output_3_1), .y(output_2_429));
wire output_1_430, output_1_2, output_0_430;
mixer gate_output_0_430(.a(output_1_430), .b(output_1_2), .y(output_0_430));
wire output_2_430, output_2_2, output_1_430;
mixer gate_output_1_430(.a(output_2_430), .b(output_2_2), .y(output_1_430));
wire output_3_430, output_3_2, output_2_430;
mixer gate_output_2_430(.a(output_3_430), .b(output_3_2), .y(output_2_430));
wire output_1_431, output_1_0, output_0_431;
mixer gate_output_0_431(.a(output_1_431), .b(output_1_0), .y(output_0_431));
wire output_2_431, output_2_0, output_1_431;
mixer gate_output_1_431(.a(output_2_431), .b(output_2_0), .y(output_1_431));
wire output_3_431, output_3_0, output_2_431;
mixer gate_output_2_431(.a(output_3_431), .b(output_3_0), .y(output_2_431));
wire output_1_432, output_1_1, output_0_432;
mixer gate_output_0_432(.a(output_1_432), .b(output_1_1), .y(output_0_432));
wire output_2_432, output_2_1, output_1_432;
mixer gate_output_1_432(.a(output_2_432), .b(output_2_1), .y(output_1_432));
wire output_3_432, output_3_1, output_2_432;
mixer gate_output_2_432(.a(output_3_432), .b(output_3_1), .y(output_2_432));
wire output_1_433, output_1_2, output_0_433;
mixer gate_output_0_433(.a(output_1_433), .b(output_1_2), .y(output_0_433));
wire output_2_433, output_2_2, output_1_433;
mixer gate_output_1_433(.a(output_2_433), .b(output_2_2), .y(output_1_433));
wire output_3_433, output_3_2, output_2_433;
mixer gate_output_2_433(.a(output_3_433), .b(output_3_2), .y(output_2_433));
wire output_1_434, output_1_0, output_0_434;
mixer gate_output_0_434(.a(output_1_434), .b(output_1_0), .y(output_0_434));
wire output_2_434, output_2_0, output_1_434;
mixer gate_output_1_434(.a(output_2_434), .b(output_2_0), .y(output_1_434));
wire output_3_434, output_3_0, output_2_434;
mixer gate_output_2_434(.a(output_3_434), .b(output_3_0), .y(output_2_434));
wire output_1_435, output_1_1, output_0_435;
mixer gate_output_0_435(.a(output_1_435), .b(output_1_1), .y(output_0_435));
wire output_2_435, output_2_1, output_1_435;
mixer gate_output_1_435(.a(output_2_435), .b(output_2_1), .y(output_1_435));
wire output_3_435, output_3_1, output_2_435;
mixer gate_output_2_435(.a(output_3_435), .b(output_3_1), .y(output_2_435));
wire output_1_436, output_1_2, output_0_436;
mixer gate_output_0_436(.a(output_1_436), .b(output_1_2), .y(output_0_436));
wire output_2_436, output_2_2, output_1_436;
mixer gate_output_1_436(.a(output_2_436), .b(output_2_2), .y(output_1_436));
wire output_3_436, output_3_2, output_2_436;
mixer gate_output_2_436(.a(output_3_436), .b(output_3_2), .y(output_2_436));
wire output_1_437, output_1_0, output_0_437;
mixer gate_output_0_437(.a(output_1_437), .b(output_1_0), .y(output_0_437));
wire output_2_437, output_2_0, output_1_437;
mixer gate_output_1_437(.a(output_2_437), .b(output_2_0), .y(output_1_437));
wire output_3_437, output_3_0, output_2_437;
mixer gate_output_2_437(.a(output_3_437), .b(output_3_0), .y(output_2_437));
wire output_1_438, output_1_1, output_0_438;
mixer gate_output_0_438(.a(output_1_438), .b(output_1_1), .y(output_0_438));
wire output_2_438, output_2_1, output_1_438;
mixer gate_output_1_438(.a(output_2_438), .b(output_2_1), .y(output_1_438));
wire output_3_438, output_3_1, output_2_438;
mixer gate_output_2_438(.a(output_3_438), .b(output_3_1), .y(output_2_438));
wire output_1_439, output_1_2, output_0_439;
mixer gate_output_0_439(.a(output_1_439), .b(output_1_2), .y(output_0_439));
wire output_2_439, output_2_2, output_1_439;
mixer gate_output_1_439(.a(output_2_439), .b(output_2_2), .y(output_1_439));
wire output_3_439, output_3_2, output_2_439;
mixer gate_output_2_439(.a(output_3_439), .b(output_3_2), .y(output_2_439));
wire output_1_440, output_1_0, output_0_440;
mixer gate_output_0_440(.a(output_1_440), .b(output_1_0), .y(output_0_440));
wire output_2_440, output_2_0, output_1_440;
mixer gate_output_1_440(.a(output_2_440), .b(output_2_0), .y(output_1_440));
wire output_3_440, output_3_0, output_2_440;
mixer gate_output_2_440(.a(output_3_440), .b(output_3_0), .y(output_2_440));
wire output_1_441, output_1_1, output_0_441;
mixer gate_output_0_441(.a(output_1_441), .b(output_1_1), .y(output_0_441));
wire output_2_441, output_2_1, output_1_441;
mixer gate_output_1_441(.a(output_2_441), .b(output_2_1), .y(output_1_441));
wire output_3_441, output_3_1, output_2_441;
mixer gate_output_2_441(.a(output_3_441), .b(output_3_1), .y(output_2_441));
wire output_1_442, output_1_2, output_0_442;
mixer gate_output_0_442(.a(output_1_442), .b(output_1_2), .y(output_0_442));
wire output_2_442, output_2_2, output_1_442;
mixer gate_output_1_442(.a(output_2_442), .b(output_2_2), .y(output_1_442));
wire output_3_442, output_3_2, output_2_442;
mixer gate_output_2_442(.a(output_3_442), .b(output_3_2), .y(output_2_442));
wire output_1_443, output_1_0, output_0_443;
mixer gate_output_0_443(.a(output_1_443), .b(output_1_0), .y(output_0_443));
wire output_2_443, output_2_0, output_1_443;
mixer gate_output_1_443(.a(output_2_443), .b(output_2_0), .y(output_1_443));
wire output_3_443, output_3_0, output_2_443;
mixer gate_output_2_443(.a(output_3_443), .b(output_3_0), .y(output_2_443));
wire output_1_444, output_1_1, output_0_444;
mixer gate_output_0_444(.a(output_1_444), .b(output_1_1), .y(output_0_444));
wire output_2_444, output_2_1, output_1_444;
mixer gate_output_1_444(.a(output_2_444), .b(output_2_1), .y(output_1_444));
wire output_3_444, output_3_1, output_2_444;
mixer gate_output_2_444(.a(output_3_444), .b(output_3_1), .y(output_2_444));
wire output_1_445, output_1_2, output_0_445;
mixer gate_output_0_445(.a(output_1_445), .b(output_1_2), .y(output_0_445));
wire output_2_445, output_2_2, output_1_445;
mixer gate_output_1_445(.a(output_2_445), .b(output_2_2), .y(output_1_445));
wire output_3_445, output_3_2, output_2_445;
mixer gate_output_2_445(.a(output_3_445), .b(output_3_2), .y(output_2_445));
wire output_1_446, output_1_0, output_0_446;
mixer gate_output_0_446(.a(output_1_446), .b(output_1_0), .y(output_0_446));
wire output_2_446, output_2_0, output_1_446;
mixer gate_output_1_446(.a(output_2_446), .b(output_2_0), .y(output_1_446));
wire output_3_446, output_3_0, output_2_446;
mixer gate_output_2_446(.a(output_3_446), .b(output_3_0), .y(output_2_446));
wire output_1_447, output_1_1, output_0_447;
mixer gate_output_0_447(.a(output_1_447), .b(output_1_1), .y(output_0_447));
wire output_2_447, output_2_1, output_1_447;
mixer gate_output_1_447(.a(output_2_447), .b(output_2_1), .y(output_1_447));
wire output_3_447, output_3_1, output_2_447;
mixer gate_output_2_447(.a(output_3_447), .b(output_3_1), .y(output_2_447));
wire output_1_448, output_1_2, output_0_448;
mixer gate_output_0_448(.a(output_1_448), .b(output_1_2), .y(output_0_448));
wire output_2_448, output_2_2, output_1_448;
mixer gate_output_1_448(.a(output_2_448), .b(output_2_2), .y(output_1_448));
wire output_3_448, output_3_2, output_2_448;
mixer gate_output_2_448(.a(output_3_448), .b(output_3_2), .y(output_2_448));
wire output_1_449, output_1_0, output_0_449;
mixer gate_output_0_449(.a(output_1_449), .b(output_1_0), .y(output_0_449));
wire output_2_449, output_2_0, output_1_449;
mixer gate_output_1_449(.a(output_2_449), .b(output_2_0), .y(output_1_449));
wire output_3_449, output_3_0, output_2_449;
mixer gate_output_2_449(.a(output_3_449), .b(output_3_0), .y(output_2_449));
wire output_1_450, output_1_1, output_0_450;
mixer gate_output_0_450(.a(output_1_450), .b(output_1_1), .y(output_0_450));
wire output_2_450, output_2_1, output_1_450;
mixer gate_output_1_450(.a(output_2_450), .b(output_2_1), .y(output_1_450));
wire output_3_450, output_3_1, output_2_450;
mixer gate_output_2_450(.a(output_3_450), .b(output_3_1), .y(output_2_450));
wire output_1_451, output_1_2, output_0_451;
mixer gate_output_0_451(.a(output_1_451), .b(output_1_2), .y(output_0_451));
wire output_2_451, output_2_2, output_1_451;
mixer gate_output_1_451(.a(output_2_451), .b(output_2_2), .y(output_1_451));
wire output_3_451, output_3_2, output_2_451;
mixer gate_output_2_451(.a(output_3_451), .b(output_3_2), .y(output_2_451));
wire output_1_452, output_1_0, output_0_452;
mixer gate_output_0_452(.a(output_1_452), .b(output_1_0), .y(output_0_452));
wire output_2_452, output_2_0, output_1_452;
mixer gate_output_1_452(.a(output_2_452), .b(output_2_0), .y(output_1_452));
wire output_3_452, output_3_0, output_2_452;
mixer gate_output_2_452(.a(output_3_452), .b(output_3_0), .y(output_2_452));
wire output_1_453, output_1_1, output_0_453;
mixer gate_output_0_453(.a(output_1_453), .b(output_1_1), .y(output_0_453));
wire output_2_453, output_2_1, output_1_453;
mixer gate_output_1_453(.a(output_2_453), .b(output_2_1), .y(output_1_453));
wire output_3_453, output_3_1, output_2_453;
mixer gate_output_2_453(.a(output_3_453), .b(output_3_1), .y(output_2_453));
wire output_1_454, output_1_2, output_0_454;
mixer gate_output_0_454(.a(output_1_454), .b(output_1_2), .y(output_0_454));
wire output_2_454, output_2_2, output_1_454;
mixer gate_output_1_454(.a(output_2_454), .b(output_2_2), .y(output_1_454));
wire output_3_454, output_3_2, output_2_454;
mixer gate_output_2_454(.a(output_3_454), .b(output_3_2), .y(output_2_454));
wire output_1_455, output_1_0, output_0_455;
mixer gate_output_0_455(.a(output_1_455), .b(output_1_0), .y(output_0_455));
wire output_2_455, output_2_0, output_1_455;
mixer gate_output_1_455(.a(output_2_455), .b(output_2_0), .y(output_1_455));
wire output_3_455, output_3_0, output_2_455;
mixer gate_output_2_455(.a(output_3_455), .b(output_3_0), .y(output_2_455));
wire output_1_456, output_1_1, output_0_456;
mixer gate_output_0_456(.a(output_1_456), .b(output_1_1), .y(output_0_456));
wire output_2_456, output_2_1, output_1_456;
mixer gate_output_1_456(.a(output_2_456), .b(output_2_1), .y(output_1_456));
wire output_3_456, output_3_1, output_2_456;
mixer gate_output_2_456(.a(output_3_456), .b(output_3_1), .y(output_2_456));
wire output_1_457, output_1_2, output_0_457;
mixer gate_output_0_457(.a(output_1_457), .b(output_1_2), .y(output_0_457));
wire output_2_457, output_2_2, output_1_457;
mixer gate_output_1_457(.a(output_2_457), .b(output_2_2), .y(output_1_457));
wire output_3_457, output_3_2, output_2_457;
mixer gate_output_2_457(.a(output_3_457), .b(output_3_2), .y(output_2_457));
wire output_1_458, output_1_0, output_0_458;
mixer gate_output_0_458(.a(output_1_458), .b(output_1_0), .y(output_0_458));
wire output_2_458, output_2_0, output_1_458;
mixer gate_output_1_458(.a(output_2_458), .b(output_2_0), .y(output_1_458));
wire output_3_458, output_3_0, output_2_458;
mixer gate_output_2_458(.a(output_3_458), .b(output_3_0), .y(output_2_458));
wire output_1_459, output_1_1, output_0_459;
mixer gate_output_0_459(.a(output_1_459), .b(output_1_1), .y(output_0_459));
wire output_2_459, output_2_1, output_1_459;
mixer gate_output_1_459(.a(output_2_459), .b(output_2_1), .y(output_1_459));
wire output_3_459, output_3_1, output_2_459;
mixer gate_output_2_459(.a(output_3_459), .b(output_3_1), .y(output_2_459));
wire output_1_460, output_1_2, output_0_460;
mixer gate_output_0_460(.a(output_1_460), .b(output_1_2), .y(output_0_460));
wire output_2_460, output_2_2, output_1_460;
mixer gate_output_1_460(.a(output_2_460), .b(output_2_2), .y(output_1_460));
wire output_3_460, output_3_2, output_2_460;
mixer gate_output_2_460(.a(output_3_460), .b(output_3_2), .y(output_2_460));
wire output_1_461, output_1_0, output_0_461;
mixer gate_output_0_461(.a(output_1_461), .b(output_1_0), .y(output_0_461));
wire output_2_461, output_2_0, output_1_461;
mixer gate_output_1_461(.a(output_2_461), .b(output_2_0), .y(output_1_461));
wire output_3_461, output_3_0, output_2_461;
mixer gate_output_2_461(.a(output_3_461), .b(output_3_0), .y(output_2_461));
wire output_1_462, output_1_1, output_0_462;
mixer gate_output_0_462(.a(output_1_462), .b(output_1_1), .y(output_0_462));
wire output_2_462, output_2_1, output_1_462;
mixer gate_output_1_462(.a(output_2_462), .b(output_2_1), .y(output_1_462));
wire output_3_462, output_3_1, output_2_462;
mixer gate_output_2_462(.a(output_3_462), .b(output_3_1), .y(output_2_462));
wire output_1_463, output_1_2, output_0_463;
mixer gate_output_0_463(.a(output_1_463), .b(output_1_2), .y(output_0_463));
wire output_2_463, output_2_2, output_1_463;
mixer gate_output_1_463(.a(output_2_463), .b(output_2_2), .y(output_1_463));
wire output_3_463, output_3_2, output_2_463;
mixer gate_output_2_463(.a(output_3_463), .b(output_3_2), .y(output_2_463));
wire output_1_464, output_1_0, output_0_464;
mixer gate_output_0_464(.a(output_1_464), .b(output_1_0), .y(output_0_464));
wire output_2_464, output_2_0, output_1_464;
mixer gate_output_1_464(.a(output_2_464), .b(output_2_0), .y(output_1_464));
wire output_3_464, output_3_0, output_2_464;
mixer gate_output_2_464(.a(output_3_464), .b(output_3_0), .y(output_2_464));
wire output_1_465, output_1_1, output_0_465;
mixer gate_output_0_465(.a(output_1_465), .b(output_1_1), .y(output_0_465));
wire output_2_465, output_2_1, output_1_465;
mixer gate_output_1_465(.a(output_2_465), .b(output_2_1), .y(output_1_465));
wire output_3_465, output_3_1, output_2_465;
mixer gate_output_2_465(.a(output_3_465), .b(output_3_1), .y(output_2_465));
wire output_1_466, output_1_2, output_0_466;
mixer gate_output_0_466(.a(output_1_466), .b(output_1_2), .y(output_0_466));
wire output_2_466, output_2_2, output_1_466;
mixer gate_output_1_466(.a(output_2_466), .b(output_2_2), .y(output_1_466));
wire output_3_466, output_3_2, output_2_466;
mixer gate_output_2_466(.a(output_3_466), .b(output_3_2), .y(output_2_466));
wire output_1_467, output_1_0, output_0_467;
mixer gate_output_0_467(.a(output_1_467), .b(output_1_0), .y(output_0_467));
wire output_2_467, output_2_0, output_1_467;
mixer gate_output_1_467(.a(output_2_467), .b(output_2_0), .y(output_1_467));
wire output_3_467, output_3_0, output_2_467;
mixer gate_output_2_467(.a(output_3_467), .b(output_3_0), .y(output_2_467));
wire output_1_468, output_1_1, output_0_468;
mixer gate_output_0_468(.a(output_1_468), .b(output_1_1), .y(output_0_468));
wire output_2_468, output_2_1, output_1_468;
mixer gate_output_1_468(.a(output_2_468), .b(output_2_1), .y(output_1_468));
wire output_3_468, output_3_1, output_2_468;
mixer gate_output_2_468(.a(output_3_468), .b(output_3_1), .y(output_2_468));
wire output_1_469, output_1_2, output_0_469;
mixer gate_output_0_469(.a(output_1_469), .b(output_1_2), .y(output_0_469));
wire output_2_469, output_2_2, output_1_469;
mixer gate_output_1_469(.a(output_2_469), .b(output_2_2), .y(output_1_469));
wire output_3_469, output_3_2, output_2_469;
mixer gate_output_2_469(.a(output_3_469), .b(output_3_2), .y(output_2_469));
wire output_1_470, output_1_0, output_0_470;
mixer gate_output_0_470(.a(output_1_470), .b(output_1_0), .y(output_0_470));
wire output_2_470, output_2_0, output_1_470;
mixer gate_output_1_470(.a(output_2_470), .b(output_2_0), .y(output_1_470));
wire output_3_470, output_3_0, output_2_470;
mixer gate_output_2_470(.a(output_3_470), .b(output_3_0), .y(output_2_470));
wire output_1_471, output_1_1, output_0_471;
mixer gate_output_0_471(.a(output_1_471), .b(output_1_1), .y(output_0_471));
wire output_2_471, output_2_1, output_1_471;
mixer gate_output_1_471(.a(output_2_471), .b(output_2_1), .y(output_1_471));
wire output_3_471, output_3_1, output_2_471;
mixer gate_output_2_471(.a(output_3_471), .b(output_3_1), .y(output_2_471));
wire output_1_472, output_1_2, output_0_472;
mixer gate_output_0_472(.a(output_1_472), .b(output_1_2), .y(output_0_472));
wire output_2_472, output_2_2, output_1_472;
mixer gate_output_1_472(.a(output_2_472), .b(output_2_2), .y(output_1_472));
wire output_3_472, output_3_2, output_2_472;
mixer gate_output_2_472(.a(output_3_472), .b(output_3_2), .y(output_2_472));
wire output_1_473, output_1_0, output_0_473;
mixer gate_output_0_473(.a(output_1_473), .b(output_1_0), .y(output_0_473));
wire output_2_473, output_2_0, output_1_473;
mixer gate_output_1_473(.a(output_2_473), .b(output_2_0), .y(output_1_473));
wire output_3_473, output_3_0, output_2_473;
mixer gate_output_2_473(.a(output_3_473), .b(output_3_0), .y(output_2_473));
wire output_1_474, output_1_1, output_0_474;
mixer gate_output_0_474(.a(output_1_474), .b(output_1_1), .y(output_0_474));
wire output_2_474, output_2_1, output_1_474;
mixer gate_output_1_474(.a(output_2_474), .b(output_2_1), .y(output_1_474));
wire output_3_474, output_3_1, output_2_474;
mixer gate_output_2_474(.a(output_3_474), .b(output_3_1), .y(output_2_474));
wire output_1_475, output_1_2, output_0_475;
mixer gate_output_0_475(.a(output_1_475), .b(output_1_2), .y(output_0_475));
wire output_2_475, output_2_2, output_1_475;
mixer gate_output_1_475(.a(output_2_475), .b(output_2_2), .y(output_1_475));
wire output_3_475, output_3_2, output_2_475;
mixer gate_output_2_475(.a(output_3_475), .b(output_3_2), .y(output_2_475));
wire output_1_476, output_1_0, output_0_476;
mixer gate_output_0_476(.a(output_1_476), .b(output_1_0), .y(output_0_476));
wire output_2_476, output_2_0, output_1_476;
mixer gate_output_1_476(.a(output_2_476), .b(output_2_0), .y(output_1_476));
wire output_3_476, output_3_0, output_2_476;
mixer gate_output_2_476(.a(output_3_476), .b(output_3_0), .y(output_2_476));
wire output_1_477, output_1_1, output_0_477;
mixer gate_output_0_477(.a(output_1_477), .b(output_1_1), .y(output_0_477));
wire output_2_477, output_2_1, output_1_477;
mixer gate_output_1_477(.a(output_2_477), .b(output_2_1), .y(output_1_477));
wire output_3_477, output_3_1, output_2_477;
mixer gate_output_2_477(.a(output_3_477), .b(output_3_1), .y(output_2_477));
wire output_1_478, output_1_2, output_0_478;
mixer gate_output_0_478(.a(output_1_478), .b(output_1_2), .y(output_0_478));
wire output_2_478, output_2_2, output_1_478;
mixer gate_output_1_478(.a(output_2_478), .b(output_2_2), .y(output_1_478));
wire output_3_478, output_3_2, output_2_478;
mixer gate_output_2_478(.a(output_3_478), .b(output_3_2), .y(output_2_478));
wire output_1_479, output_1_0, output_0_479;
mixer gate_output_0_479(.a(output_1_479), .b(output_1_0), .y(output_0_479));
wire output_2_479, output_2_0, output_1_479;
mixer gate_output_1_479(.a(output_2_479), .b(output_2_0), .y(output_1_479));
wire output_3_479, output_3_0, output_2_479;
mixer gate_output_2_479(.a(output_3_479), .b(output_3_0), .y(output_2_479));
wire output_1_480, output_1_1, output_0_480;
mixer gate_output_0_480(.a(output_1_480), .b(output_1_1), .y(output_0_480));
wire output_2_480, output_2_1, output_1_480;
mixer gate_output_1_480(.a(output_2_480), .b(output_2_1), .y(output_1_480));
wire output_3_480, output_3_1, output_2_480;
mixer gate_output_2_480(.a(output_3_480), .b(output_3_1), .y(output_2_480));
wire output_1_481, output_1_2, output_0_481;
mixer gate_output_0_481(.a(output_1_481), .b(output_1_2), .y(output_0_481));
wire output_2_481, output_2_2, output_1_481;
mixer gate_output_1_481(.a(output_2_481), .b(output_2_2), .y(output_1_481));
wire output_3_481, output_3_2, output_2_481;
mixer gate_output_2_481(.a(output_3_481), .b(output_3_2), .y(output_2_481));
wire output_1_482, output_1_0, output_0_482;
mixer gate_output_0_482(.a(output_1_482), .b(output_1_0), .y(output_0_482));
wire output_2_482, output_2_0, output_1_482;
mixer gate_output_1_482(.a(output_2_482), .b(output_2_0), .y(output_1_482));
wire output_3_482, output_3_0, output_2_482;
mixer gate_output_2_482(.a(output_3_482), .b(output_3_0), .y(output_2_482));
wire output_1_483, output_1_1, output_0_483;
mixer gate_output_0_483(.a(output_1_483), .b(output_1_1), .y(output_0_483));
wire output_2_483, output_2_1, output_1_483;
mixer gate_output_1_483(.a(output_2_483), .b(output_2_1), .y(output_1_483));
wire output_3_483, output_3_1, output_2_483;
mixer gate_output_2_483(.a(output_3_483), .b(output_3_1), .y(output_2_483));
wire output_1_484, output_1_2, output_0_484;
mixer gate_output_0_484(.a(output_1_484), .b(output_1_2), .y(output_0_484));
wire output_2_484, output_2_2, output_1_484;
mixer gate_output_1_484(.a(output_2_484), .b(output_2_2), .y(output_1_484));
wire output_3_484, output_3_2, output_2_484;
mixer gate_output_2_484(.a(output_3_484), .b(output_3_2), .y(output_2_484));
wire output_1_485, output_1_0, output_0_485;
mixer gate_output_0_485(.a(output_1_485), .b(output_1_0), .y(output_0_485));
wire output_2_485, output_2_0, output_1_485;
mixer gate_output_1_485(.a(output_2_485), .b(output_2_0), .y(output_1_485));
wire output_3_485, output_3_0, output_2_485;
mixer gate_output_2_485(.a(output_3_485), .b(output_3_0), .y(output_2_485));
wire output_1_486, output_1_1, output_0_486;
mixer gate_output_0_486(.a(output_1_486), .b(output_1_1), .y(output_0_486));
wire output_2_486, output_2_1, output_1_486;
mixer gate_output_1_486(.a(output_2_486), .b(output_2_1), .y(output_1_486));
wire output_3_486, output_3_1, output_2_486;
mixer gate_output_2_486(.a(output_3_486), .b(output_3_1), .y(output_2_486));
wire output_1_487, output_1_2, output_0_487;
mixer gate_output_0_487(.a(output_1_487), .b(output_1_2), .y(output_0_487));
wire output_2_487, output_2_2, output_1_487;
mixer gate_output_1_487(.a(output_2_487), .b(output_2_2), .y(output_1_487));
wire output_3_487, output_3_2, output_2_487;
mixer gate_output_2_487(.a(output_3_487), .b(output_3_2), .y(output_2_487));
wire output_1_488, output_1_0, output_0_488;
mixer gate_output_0_488(.a(output_1_488), .b(output_1_0), .y(output_0_488));
wire output_2_488, output_2_0, output_1_488;
mixer gate_output_1_488(.a(output_2_488), .b(output_2_0), .y(output_1_488));
wire output_3_488, output_3_0, output_2_488;
mixer gate_output_2_488(.a(output_3_488), .b(output_3_0), .y(output_2_488));
wire output_1_489, output_1_1, output_0_489;
mixer gate_output_0_489(.a(output_1_489), .b(output_1_1), .y(output_0_489));
wire output_2_489, output_2_1, output_1_489;
mixer gate_output_1_489(.a(output_2_489), .b(output_2_1), .y(output_1_489));
wire output_3_489, output_3_1, output_2_489;
mixer gate_output_2_489(.a(output_3_489), .b(output_3_1), .y(output_2_489));
wire output_1_490, output_1_2, output_0_490;
mixer gate_output_0_490(.a(output_1_490), .b(output_1_2), .y(output_0_490));
wire output_2_490, output_2_2, output_1_490;
mixer gate_output_1_490(.a(output_2_490), .b(output_2_2), .y(output_1_490));
wire output_3_490, output_3_2, output_2_490;
mixer gate_output_2_490(.a(output_3_490), .b(output_3_2), .y(output_2_490));
wire output_1_491, output_1_0, output_0_491;
mixer gate_output_0_491(.a(output_1_491), .b(output_1_0), .y(output_0_491));
wire output_2_491, output_2_0, output_1_491;
mixer gate_output_1_491(.a(output_2_491), .b(output_2_0), .y(output_1_491));
wire output_3_491, output_3_0, output_2_491;
mixer gate_output_2_491(.a(output_3_491), .b(output_3_0), .y(output_2_491));
wire output_1_492, output_1_1, output_0_492;
mixer gate_output_0_492(.a(output_1_492), .b(output_1_1), .y(output_0_492));
wire output_2_492, output_2_1, output_1_492;
mixer gate_output_1_492(.a(output_2_492), .b(output_2_1), .y(output_1_492));
wire output_3_492, output_3_1, output_2_492;
mixer gate_output_2_492(.a(output_3_492), .b(output_3_1), .y(output_2_492));
wire output_1_493, output_1_2, output_0_493;
mixer gate_output_0_493(.a(output_1_493), .b(output_1_2), .y(output_0_493));
wire output_2_493, output_2_2, output_1_493;
mixer gate_output_1_493(.a(output_2_493), .b(output_2_2), .y(output_1_493));
wire output_3_493, output_3_2, output_2_493;
mixer gate_output_2_493(.a(output_3_493), .b(output_3_2), .y(output_2_493));
wire output_1_494, output_1_0, output_0_494;
mixer gate_output_0_494(.a(output_1_494), .b(output_1_0), .y(output_0_494));
wire output_2_494, output_2_0, output_1_494;
mixer gate_output_1_494(.a(output_2_494), .b(output_2_0), .y(output_1_494));
wire output_3_494, output_3_0, output_2_494;
mixer gate_output_2_494(.a(output_3_494), .b(output_3_0), .y(output_2_494));
wire output_1_495, output_1_1, output_0_495;
mixer gate_output_0_495(.a(output_1_495), .b(output_1_1), .y(output_0_495));
wire output_2_495, output_2_1, output_1_495;
mixer gate_output_1_495(.a(output_2_495), .b(output_2_1), .y(output_1_495));
wire output_3_495, output_3_1, output_2_495;
mixer gate_output_2_495(.a(output_3_495), .b(output_3_1), .y(output_2_495));
wire output_1_496, output_1_2, output_0_496;
mixer gate_output_0_496(.a(output_1_496), .b(output_1_2), .y(output_0_496));
wire output_2_496, output_2_2, output_1_496;
mixer gate_output_1_496(.a(output_2_496), .b(output_2_2), .y(output_1_496));
wire output_3_496, output_3_2, output_2_496;
mixer gate_output_2_496(.a(output_3_496), .b(output_3_2), .y(output_2_496));
wire output_1_497, output_1_0, output_0_497;
mixer gate_output_0_497(.a(output_1_497), .b(output_1_0), .y(output_0_497));
wire output_2_497, output_2_0, output_1_497;
mixer gate_output_1_497(.a(output_2_497), .b(output_2_0), .y(output_1_497));
wire output_3_497, output_3_0, output_2_497;
mixer gate_output_2_497(.a(output_3_497), .b(output_3_0), .y(output_2_497));
wire output_1_498, output_1_1, output_0_498;
mixer gate_output_0_498(.a(output_1_498), .b(output_1_1), .y(output_0_498));
wire output_2_498, output_2_1, output_1_498;
mixer gate_output_1_498(.a(output_2_498), .b(output_2_1), .y(output_1_498));
wire output_3_498, output_3_1, output_2_498;
mixer gate_output_2_498(.a(output_3_498), .b(output_3_1), .y(output_2_498));
wire output_1_499, output_1_2, output_0_499;
mixer gate_output_0_499(.a(output_1_499), .b(output_1_2), .y(output_0_499));
wire output_2_499, output_2_2, output_1_499;
mixer gate_output_1_499(.a(output_2_499), .b(output_2_2), .y(output_1_499));
wire output_3_499, output_3_2, output_2_499;
mixer gate_output_2_499(.a(output_3_499), .b(output_3_2), .y(output_2_499));
wire output_1_500, output_1_0, output_0_500;
mixer gate_output_0_500(.a(output_1_500), .b(output_1_0), .y(output_0_500));
wire output_2_500, output_2_0, output_1_500;
mixer gate_output_1_500(.a(output_2_500), .b(output_2_0), .y(output_1_500));
wire output_3_500, output_3_0, output_2_500;
mixer gate_output_2_500(.a(output_3_500), .b(output_3_0), .y(output_2_500));
wire output_1_501, output_1_1, output_0_501;
mixer gate_output_0_501(.a(output_1_501), .b(output_1_1), .y(output_0_501));
wire output_2_501, output_2_1, output_1_501;
mixer gate_output_1_501(.a(output_2_501), .b(output_2_1), .y(output_1_501));
wire output_3_501, output_3_1, output_2_501;
mixer gate_output_2_501(.a(output_3_501), .b(output_3_1), .y(output_2_501));
wire output_1_502, output_1_2, output_0_502;
mixer gate_output_0_502(.a(output_1_502), .b(output_1_2), .y(output_0_502));
wire output_2_502, output_2_2, output_1_502;
mixer gate_output_1_502(.a(output_2_502), .b(output_2_2), .y(output_1_502));
wire output_3_502, output_3_2, output_2_502;
mixer gate_output_2_502(.a(output_3_502), .b(output_3_2), .y(output_2_502));
wire output_1_503, output_1_0, output_0_503;
mixer gate_output_0_503(.a(output_1_503), .b(output_1_0), .y(output_0_503));
wire output_2_503, output_2_0, output_1_503;
mixer gate_output_1_503(.a(output_2_503), .b(output_2_0), .y(output_1_503));
wire output_3_503, output_3_0, output_2_503;
mixer gate_output_2_503(.a(output_3_503), .b(output_3_0), .y(output_2_503));
wire output_1_504, output_1_1, output_0_504;
mixer gate_output_0_504(.a(output_1_504), .b(output_1_1), .y(output_0_504));
wire output_2_504, output_2_1, output_1_504;
mixer gate_output_1_504(.a(output_2_504), .b(output_2_1), .y(output_1_504));
wire output_3_504, output_3_1, output_2_504;
mixer gate_output_2_504(.a(output_3_504), .b(output_3_1), .y(output_2_504));
wire output_1_505, output_1_2, output_0_505;
mixer gate_output_0_505(.a(output_1_505), .b(output_1_2), .y(output_0_505));
wire output_2_505, output_2_2, output_1_505;
mixer gate_output_1_505(.a(output_2_505), .b(output_2_2), .y(output_1_505));
wire output_3_505, output_3_2, output_2_505;
mixer gate_output_2_505(.a(output_3_505), .b(output_3_2), .y(output_2_505));
wire output_1_506, output_1_0, output_0_506;
mixer gate_output_0_506(.a(output_1_506), .b(output_1_0), .y(output_0_506));
wire output_2_506, output_2_0, output_1_506;
mixer gate_output_1_506(.a(output_2_506), .b(output_2_0), .y(output_1_506));
wire output_3_506, output_3_0, output_2_506;
mixer gate_output_2_506(.a(output_3_506), .b(output_3_0), .y(output_2_506));
wire output_1_507, output_1_1, output_0_507;
mixer gate_output_0_507(.a(output_1_507), .b(output_1_1), .y(output_0_507));
wire output_2_507, output_2_1, output_1_507;
mixer gate_output_1_507(.a(output_2_507), .b(output_2_1), .y(output_1_507));
wire output_3_507, output_3_1, output_2_507;
mixer gate_output_2_507(.a(output_3_507), .b(output_3_1), .y(output_2_507));
wire output_1_508, output_1_2, output_0_508;
mixer gate_output_0_508(.a(output_1_508), .b(output_1_2), .y(output_0_508));
wire output_2_508, output_2_2, output_1_508;
mixer gate_output_1_508(.a(output_2_508), .b(output_2_2), .y(output_1_508));
wire output_3_508, output_3_2, output_2_508;
mixer gate_output_2_508(.a(output_3_508), .b(output_3_2), .y(output_2_508));
wire output_1_509, output_1_0, output_0_509;
mixer gate_output_0_509(.a(output_1_509), .b(output_1_0), .y(output_0_509));
wire output_2_509, output_2_0, output_1_509;
mixer gate_output_1_509(.a(output_2_509), .b(output_2_0), .y(output_1_509));
wire output_3_509, output_3_0, output_2_509;
mixer gate_output_2_509(.a(output_3_509), .b(output_3_0), .y(output_2_509));
wire output_1_510, output_1_1, output_0_510;
mixer gate_output_0_510(.a(output_1_510), .b(output_1_1), .y(output_0_510));
wire output_2_510, output_2_1, output_1_510;
mixer gate_output_1_510(.a(output_2_510), .b(output_2_1), .y(output_1_510));
wire output_3_510, output_3_1, output_2_510;
mixer gate_output_2_510(.a(output_3_510), .b(output_3_1), .y(output_2_510));
wire output_1_511, output_1_2, output_0_511;
mixer gate_output_0_511(.a(output_1_511), .b(output_1_2), .y(output_0_511));
wire output_2_511, output_2_2, output_1_511;
mixer gate_output_1_511(.a(output_2_511), .b(output_2_2), .y(output_1_511));
wire output_3_511, output_3_2, output_2_511;
mixer gate_output_2_511(.a(output_3_511), .b(output_3_2), .y(output_2_511));
wire output_1_512, output_1_0, output_0_512;
mixer gate_output_0_512(.a(output_1_512), .b(output_1_0), .y(output_0_512));
wire output_2_512, output_2_0, output_1_512;
mixer gate_output_1_512(.a(output_2_512), .b(output_2_0), .y(output_1_512));
wire output_3_512, output_3_0, output_2_512;
mixer gate_output_2_512(.a(output_3_512), .b(output_3_0), .y(output_2_512));
wire output_1_513, output_1_1, output_0_513;
mixer gate_output_0_513(.a(output_1_513), .b(output_1_1), .y(output_0_513));
wire output_2_513, output_2_1, output_1_513;
mixer gate_output_1_513(.a(output_2_513), .b(output_2_1), .y(output_1_513));
wire output_3_513, output_3_1, output_2_513;
mixer gate_output_2_513(.a(output_3_513), .b(output_3_1), .y(output_2_513));
wire output_1_514, output_1_2, output_0_514;
mixer gate_output_0_514(.a(output_1_514), .b(output_1_2), .y(output_0_514));
wire output_2_514, output_2_2, output_1_514;
mixer gate_output_1_514(.a(output_2_514), .b(output_2_2), .y(output_1_514));
wire output_3_514, output_3_2, output_2_514;
mixer gate_output_2_514(.a(output_3_514), .b(output_3_2), .y(output_2_514));
wire output_1_515, output_1_0, output_0_515;
mixer gate_output_0_515(.a(output_1_515), .b(output_1_0), .y(output_0_515));
wire output_2_515, output_2_0, output_1_515;
mixer gate_output_1_515(.a(output_2_515), .b(output_2_0), .y(output_1_515));
wire output_3_515, output_3_0, output_2_515;
mixer gate_output_2_515(.a(output_3_515), .b(output_3_0), .y(output_2_515));
wire output_1_516, output_1_1, output_0_516;
mixer gate_output_0_516(.a(output_1_516), .b(output_1_1), .y(output_0_516));
wire output_2_516, output_2_1, output_1_516;
mixer gate_output_1_516(.a(output_2_516), .b(output_2_1), .y(output_1_516));
wire output_3_516, output_3_1, output_2_516;
mixer gate_output_2_516(.a(output_3_516), .b(output_3_1), .y(output_2_516));
wire output_1_517, output_1_2, output_0_517;
mixer gate_output_0_517(.a(output_1_517), .b(output_1_2), .y(output_0_517));
wire output_2_517, output_2_2, output_1_517;
mixer gate_output_1_517(.a(output_2_517), .b(output_2_2), .y(output_1_517));
wire output_3_517, output_3_2, output_2_517;
mixer gate_output_2_517(.a(output_3_517), .b(output_3_2), .y(output_2_517));
wire output_1_518, output_1_0, output_0_518;
mixer gate_output_0_518(.a(output_1_518), .b(output_1_0), .y(output_0_518));
wire output_2_518, output_2_0, output_1_518;
mixer gate_output_1_518(.a(output_2_518), .b(output_2_0), .y(output_1_518));
wire output_3_518, output_3_0, output_2_518;
mixer gate_output_2_518(.a(output_3_518), .b(output_3_0), .y(output_2_518));
wire output_1_519, output_1_1, output_0_519;
mixer gate_output_0_519(.a(output_1_519), .b(output_1_1), .y(output_0_519));
wire output_2_519, output_2_1, output_1_519;
mixer gate_output_1_519(.a(output_2_519), .b(output_2_1), .y(output_1_519));
wire output_3_519, output_3_1, output_2_519;
mixer gate_output_2_519(.a(output_3_519), .b(output_3_1), .y(output_2_519));
wire output_1_520, output_1_2, output_0_520;
mixer gate_output_0_520(.a(output_1_520), .b(output_1_2), .y(output_0_520));
wire output_2_520, output_2_2, output_1_520;
mixer gate_output_1_520(.a(output_2_520), .b(output_2_2), .y(output_1_520));
wire output_3_520, output_3_2, output_2_520;
mixer gate_output_2_520(.a(output_3_520), .b(output_3_2), .y(output_2_520));
wire output_1_521, output_1_0, output_0_521;
mixer gate_output_0_521(.a(output_1_521), .b(output_1_0), .y(output_0_521));
wire output_2_521, output_2_0, output_1_521;
mixer gate_output_1_521(.a(output_2_521), .b(output_2_0), .y(output_1_521));
wire output_3_521, output_3_0, output_2_521;
mixer gate_output_2_521(.a(output_3_521), .b(output_3_0), .y(output_2_521));
wire output_1_522, output_1_1, output_0_522;
mixer gate_output_0_522(.a(output_1_522), .b(output_1_1), .y(output_0_522));
wire output_2_522, output_2_1, output_1_522;
mixer gate_output_1_522(.a(output_2_522), .b(output_2_1), .y(output_1_522));
wire output_3_522, output_3_1, output_2_522;
mixer gate_output_2_522(.a(output_3_522), .b(output_3_1), .y(output_2_522));
wire output_1_523, output_1_2, output_0_523;
mixer gate_output_0_523(.a(output_1_523), .b(output_1_2), .y(output_0_523));
wire output_2_523, output_2_2, output_1_523;
mixer gate_output_1_523(.a(output_2_523), .b(output_2_2), .y(output_1_523));
wire output_3_523, output_3_2, output_2_523;
mixer gate_output_2_523(.a(output_3_523), .b(output_3_2), .y(output_2_523));
wire output_1_524, output_1_0, output_0_524;
mixer gate_output_0_524(.a(output_1_524), .b(output_1_0), .y(output_0_524));
wire output_2_524, output_2_0, output_1_524;
mixer gate_output_1_524(.a(output_2_524), .b(output_2_0), .y(output_1_524));
wire output_3_524, output_3_0, output_2_524;
mixer gate_output_2_524(.a(output_3_524), .b(output_3_0), .y(output_2_524));
wire output_1_525, output_1_1, output_0_525;
mixer gate_output_0_525(.a(output_1_525), .b(output_1_1), .y(output_0_525));
wire output_2_525, output_2_1, output_1_525;
mixer gate_output_1_525(.a(output_2_525), .b(output_2_1), .y(output_1_525));
wire output_3_525, output_3_1, output_2_525;
mixer gate_output_2_525(.a(output_3_525), .b(output_3_1), .y(output_2_525));
wire output_1_526, output_1_2, output_0_526;
mixer gate_output_0_526(.a(output_1_526), .b(output_1_2), .y(output_0_526));
wire output_2_526, output_2_2, output_1_526;
mixer gate_output_1_526(.a(output_2_526), .b(output_2_2), .y(output_1_526));
wire output_3_526, output_3_2, output_2_526;
mixer gate_output_2_526(.a(output_3_526), .b(output_3_2), .y(output_2_526));
wire output_1_527, output_1_0, output_0_527;
mixer gate_output_0_527(.a(output_1_527), .b(output_1_0), .y(output_0_527));
wire output_2_527, output_2_0, output_1_527;
mixer gate_output_1_527(.a(output_2_527), .b(output_2_0), .y(output_1_527));
wire output_3_527, output_3_0, output_2_527;
mixer gate_output_2_527(.a(output_3_527), .b(output_3_0), .y(output_2_527));
wire output_1_528, output_1_1, output_0_528;
mixer gate_output_0_528(.a(output_1_528), .b(output_1_1), .y(output_0_528));
wire output_2_528, output_2_1, output_1_528;
mixer gate_output_1_528(.a(output_2_528), .b(output_2_1), .y(output_1_528));
wire output_3_528, output_3_1, output_2_528;
mixer gate_output_2_528(.a(output_3_528), .b(output_3_1), .y(output_2_528));
wire output_1_529, output_1_2, output_0_529;
mixer gate_output_0_529(.a(output_1_529), .b(output_1_2), .y(output_0_529));
wire output_2_529, output_2_2, output_1_529;
mixer gate_output_1_529(.a(output_2_529), .b(output_2_2), .y(output_1_529));
wire output_3_529, output_3_2, output_2_529;
mixer gate_output_2_529(.a(output_3_529), .b(output_3_2), .y(output_2_529));
wire output_1_530, output_1_0, output_0_530;
mixer gate_output_0_530(.a(output_1_530), .b(output_1_0), .y(output_0_530));
wire output_2_530, output_2_0, output_1_530;
mixer gate_output_1_530(.a(output_2_530), .b(output_2_0), .y(output_1_530));
wire output_3_530, output_3_0, output_2_530;
mixer gate_output_2_530(.a(output_3_530), .b(output_3_0), .y(output_2_530));
wire output_1_531, output_1_1, output_0_531;
mixer gate_output_0_531(.a(output_1_531), .b(output_1_1), .y(output_0_531));
wire output_2_531, output_2_1, output_1_531;
mixer gate_output_1_531(.a(output_2_531), .b(output_2_1), .y(output_1_531));
wire output_3_531, output_3_1, output_2_531;
mixer gate_output_2_531(.a(output_3_531), .b(output_3_1), .y(output_2_531));
wire output_1_532, output_1_2, output_0_532;
mixer gate_output_0_532(.a(output_1_532), .b(output_1_2), .y(output_0_532));
wire output_2_532, output_2_2, output_1_532;
mixer gate_output_1_532(.a(output_2_532), .b(output_2_2), .y(output_1_532));
wire output_3_532, output_3_2, output_2_532;
mixer gate_output_2_532(.a(output_3_532), .b(output_3_2), .y(output_2_532));
wire output_1_533, output_1_0, output_0_533;
mixer gate_output_0_533(.a(output_1_533), .b(output_1_0), .y(output_0_533));
wire output_2_533, output_2_0, output_1_533;
mixer gate_output_1_533(.a(output_2_533), .b(output_2_0), .y(output_1_533));
wire output_3_533, output_3_0, output_2_533;
mixer gate_output_2_533(.a(output_3_533), .b(output_3_0), .y(output_2_533));
wire output_1_534, output_1_1, output_0_534;
mixer gate_output_0_534(.a(output_1_534), .b(output_1_1), .y(output_0_534));
wire output_2_534, output_2_1, output_1_534;
mixer gate_output_1_534(.a(output_2_534), .b(output_2_1), .y(output_1_534));
wire output_3_534, output_3_1, output_2_534;
mixer gate_output_2_534(.a(output_3_534), .b(output_3_1), .y(output_2_534));
wire output_1_535, output_1_2, output_0_535;
mixer gate_output_0_535(.a(output_1_535), .b(output_1_2), .y(output_0_535));
wire output_2_535, output_2_2, output_1_535;
mixer gate_output_1_535(.a(output_2_535), .b(output_2_2), .y(output_1_535));
wire output_3_535, output_3_2, output_2_535;
mixer gate_output_2_535(.a(output_3_535), .b(output_3_2), .y(output_2_535));
wire output_1_536, output_1_0, output_0_536;
mixer gate_output_0_536(.a(output_1_536), .b(output_1_0), .y(output_0_536));
wire output_2_536, output_2_0, output_1_536;
mixer gate_output_1_536(.a(output_2_536), .b(output_2_0), .y(output_1_536));
wire output_3_536, output_3_0, output_2_536;
mixer gate_output_2_536(.a(output_3_536), .b(output_3_0), .y(output_2_536));
wire output_1_537, output_1_1, output_0_537;
mixer gate_output_0_537(.a(output_1_537), .b(output_1_1), .y(output_0_537));
wire output_2_537, output_2_1, output_1_537;
mixer gate_output_1_537(.a(output_2_537), .b(output_2_1), .y(output_1_537));
wire output_3_537, output_3_1, output_2_537;
mixer gate_output_2_537(.a(output_3_537), .b(output_3_1), .y(output_2_537));
wire output_1_538, output_1_2, output_0_538;
mixer gate_output_0_538(.a(output_1_538), .b(output_1_2), .y(output_0_538));
wire output_2_538, output_2_2, output_1_538;
mixer gate_output_1_538(.a(output_2_538), .b(output_2_2), .y(output_1_538));
wire output_3_538, output_3_2, output_2_538;
mixer gate_output_2_538(.a(output_3_538), .b(output_3_2), .y(output_2_538));
wire output_1_539, output_1_0, output_0_539;
mixer gate_output_0_539(.a(output_1_539), .b(output_1_0), .y(output_0_539));
wire output_2_539, output_2_0, output_1_539;
mixer gate_output_1_539(.a(output_2_539), .b(output_2_0), .y(output_1_539));
wire output_3_539, output_3_0, output_2_539;
mixer gate_output_2_539(.a(output_3_539), .b(output_3_0), .y(output_2_539));
wire output_1_540, output_1_1, output_0_540;
mixer gate_output_0_540(.a(output_1_540), .b(output_1_1), .y(output_0_540));
wire output_2_540, output_2_1, output_1_540;
mixer gate_output_1_540(.a(output_2_540), .b(output_2_1), .y(output_1_540));
wire output_3_540, output_3_1, output_2_540;
mixer gate_output_2_540(.a(output_3_540), .b(output_3_1), .y(output_2_540));
wire output_1_541, output_1_2, output_0_541;
mixer gate_output_0_541(.a(output_1_541), .b(output_1_2), .y(output_0_541));
wire output_2_541, output_2_2, output_1_541;
mixer gate_output_1_541(.a(output_2_541), .b(output_2_2), .y(output_1_541));
wire output_3_541, output_3_2, output_2_541;
mixer gate_output_2_541(.a(output_3_541), .b(output_3_2), .y(output_2_541));
wire output_1_542, output_1_0, output_0_542;
mixer gate_output_0_542(.a(output_1_542), .b(output_1_0), .y(output_0_542));
wire output_2_542, output_2_0, output_1_542;
mixer gate_output_1_542(.a(output_2_542), .b(output_2_0), .y(output_1_542));
wire output_3_542, output_3_0, output_2_542;
mixer gate_output_2_542(.a(output_3_542), .b(output_3_0), .y(output_2_542));
wire output_1_543, output_1_1, output_0_543;
mixer gate_output_0_543(.a(output_1_543), .b(output_1_1), .y(output_0_543));
wire output_2_543, output_2_1, output_1_543;
mixer gate_output_1_543(.a(output_2_543), .b(output_2_1), .y(output_1_543));
wire output_3_543, output_3_1, output_2_543;
mixer gate_output_2_543(.a(output_3_543), .b(output_3_1), .y(output_2_543));
wire output_1_544, output_1_2, output_0_544;
mixer gate_output_0_544(.a(output_1_544), .b(output_1_2), .y(output_0_544));
wire output_2_544, output_2_2, output_1_544;
mixer gate_output_1_544(.a(output_2_544), .b(output_2_2), .y(output_1_544));
wire output_3_544, output_3_2, output_2_544;
mixer gate_output_2_544(.a(output_3_544), .b(output_3_2), .y(output_2_544));
wire output_1_545, output_1_0, output_0_545;
mixer gate_output_0_545(.a(output_1_545), .b(output_1_0), .y(output_0_545));
wire output_2_545, output_2_0, output_1_545;
mixer gate_output_1_545(.a(output_2_545), .b(output_2_0), .y(output_1_545));
wire output_3_545, output_3_0, output_2_545;
mixer gate_output_2_545(.a(output_3_545), .b(output_3_0), .y(output_2_545));
wire output_1_546, output_1_1, output_0_546;
mixer gate_output_0_546(.a(output_1_546), .b(output_1_1), .y(output_0_546));
wire output_2_546, output_2_1, output_1_546;
mixer gate_output_1_546(.a(output_2_546), .b(output_2_1), .y(output_1_546));
wire output_3_546, output_3_1, output_2_546;
mixer gate_output_2_546(.a(output_3_546), .b(output_3_1), .y(output_2_546));
wire output_1_547, output_1_2, output_0_547;
mixer gate_output_0_547(.a(output_1_547), .b(output_1_2), .y(output_0_547));
wire output_2_547, output_2_2, output_1_547;
mixer gate_output_1_547(.a(output_2_547), .b(output_2_2), .y(output_1_547));
wire output_3_547, output_3_2, output_2_547;
mixer gate_output_2_547(.a(output_3_547), .b(output_3_2), .y(output_2_547));
wire output_1_548, output_1_0, output_0_548;
mixer gate_output_0_548(.a(output_1_548), .b(output_1_0), .y(output_0_548));
wire output_2_548, output_2_0, output_1_548;
mixer gate_output_1_548(.a(output_2_548), .b(output_2_0), .y(output_1_548));
wire output_3_548, output_3_0, output_2_548;
mixer gate_output_2_548(.a(output_3_548), .b(output_3_0), .y(output_2_548));
wire output_1_549, output_1_1, output_0_549;
mixer gate_output_0_549(.a(output_1_549), .b(output_1_1), .y(output_0_549));
wire output_2_549, output_2_1, output_1_549;
mixer gate_output_1_549(.a(output_2_549), .b(output_2_1), .y(output_1_549));
wire output_3_549, output_3_1, output_2_549;
mixer gate_output_2_549(.a(output_3_549), .b(output_3_1), .y(output_2_549));
wire output_1_550, output_1_2, output_0_550;
mixer gate_output_0_550(.a(output_1_550), .b(output_1_2), .y(output_0_550));
wire output_2_550, output_2_2, output_1_550;
mixer gate_output_1_550(.a(output_2_550), .b(output_2_2), .y(output_1_550));
wire output_3_550, output_3_2, output_2_550;
mixer gate_output_2_550(.a(output_3_550), .b(output_3_2), .y(output_2_550));
wire output_1_551, output_1_0, output_0_551;
mixer gate_output_0_551(.a(output_1_551), .b(output_1_0), .y(output_0_551));
wire output_2_551, output_2_0, output_1_551;
mixer gate_output_1_551(.a(output_2_551), .b(output_2_0), .y(output_1_551));
wire output_3_551, output_3_0, output_2_551;
mixer gate_output_2_551(.a(output_3_551), .b(output_3_0), .y(output_2_551));
wire output_1_552, output_1_1, output_0_552;
mixer gate_output_0_552(.a(output_1_552), .b(output_1_1), .y(output_0_552));
wire output_2_552, output_2_1, output_1_552;
mixer gate_output_1_552(.a(output_2_552), .b(output_2_1), .y(output_1_552));
wire output_3_552, output_3_1, output_2_552;
mixer gate_output_2_552(.a(output_3_552), .b(output_3_1), .y(output_2_552));
wire output_1_553, output_1_2, output_0_553;
mixer gate_output_0_553(.a(output_1_553), .b(output_1_2), .y(output_0_553));
wire output_2_553, output_2_2, output_1_553;
mixer gate_output_1_553(.a(output_2_553), .b(output_2_2), .y(output_1_553));
wire output_3_553, output_3_2, output_2_553;
mixer gate_output_2_553(.a(output_3_553), .b(output_3_2), .y(output_2_553));
wire output_1_554, output_1_0, output_0_554;
mixer gate_output_0_554(.a(output_1_554), .b(output_1_0), .y(output_0_554));
wire output_2_554, output_2_0, output_1_554;
mixer gate_output_1_554(.a(output_2_554), .b(output_2_0), .y(output_1_554));
wire output_3_554, output_3_0, output_2_554;
mixer gate_output_2_554(.a(output_3_554), .b(output_3_0), .y(output_2_554));
wire output_1_555, output_1_1, output_0_555;
mixer gate_output_0_555(.a(output_1_555), .b(output_1_1), .y(output_0_555));
wire output_2_555, output_2_1, output_1_555;
mixer gate_output_1_555(.a(output_2_555), .b(output_2_1), .y(output_1_555));
wire output_3_555, output_3_1, output_2_555;
mixer gate_output_2_555(.a(output_3_555), .b(output_3_1), .y(output_2_555));
wire output_1_556, output_1_2, output_0_556;
mixer gate_output_0_556(.a(output_1_556), .b(output_1_2), .y(output_0_556));
wire output_2_556, output_2_2, output_1_556;
mixer gate_output_1_556(.a(output_2_556), .b(output_2_2), .y(output_1_556));
wire output_3_556, output_3_2, output_2_556;
mixer gate_output_2_556(.a(output_3_556), .b(output_3_2), .y(output_2_556));
wire output_1_557, output_1_0, output_0_557;
mixer gate_output_0_557(.a(output_1_557), .b(output_1_0), .y(output_0_557));
wire output_2_557, output_2_0, output_1_557;
mixer gate_output_1_557(.a(output_2_557), .b(output_2_0), .y(output_1_557));
wire output_3_557, output_3_0, output_2_557;
mixer gate_output_2_557(.a(output_3_557), .b(output_3_0), .y(output_2_557));
wire output_1_558, output_1_1, output_0_558;
mixer gate_output_0_558(.a(output_1_558), .b(output_1_1), .y(output_0_558));
wire output_2_558, output_2_1, output_1_558;
mixer gate_output_1_558(.a(output_2_558), .b(output_2_1), .y(output_1_558));
wire output_3_558, output_3_1, output_2_558;
mixer gate_output_2_558(.a(output_3_558), .b(output_3_1), .y(output_2_558));
wire output_1_559, output_1_2, output_0_559;
mixer gate_output_0_559(.a(output_1_559), .b(output_1_2), .y(output_0_559));
wire output_2_559, output_2_2, output_1_559;
mixer gate_output_1_559(.a(output_2_559), .b(output_2_2), .y(output_1_559));
wire output_3_559, output_3_2, output_2_559;
mixer gate_output_2_559(.a(output_3_559), .b(output_3_2), .y(output_2_559));
wire output_1_560, output_1_0, output_0_560;
mixer gate_output_0_560(.a(output_1_560), .b(output_1_0), .y(output_0_560));
wire output_2_560, output_2_0, output_1_560;
mixer gate_output_1_560(.a(output_2_560), .b(output_2_0), .y(output_1_560));
wire output_3_560, output_3_0, output_2_560;
mixer gate_output_2_560(.a(output_3_560), .b(output_3_0), .y(output_2_560));
wire output_1_561, output_1_1, output_0_561;
mixer gate_output_0_561(.a(output_1_561), .b(output_1_1), .y(output_0_561));
wire output_2_561, output_2_1, output_1_561;
mixer gate_output_1_561(.a(output_2_561), .b(output_2_1), .y(output_1_561));
wire output_3_561, output_3_1, output_2_561;
mixer gate_output_2_561(.a(output_3_561), .b(output_3_1), .y(output_2_561));
wire output_1_562, output_1_2, output_0_562;
mixer gate_output_0_562(.a(output_1_562), .b(output_1_2), .y(output_0_562));
wire output_2_562, output_2_2, output_1_562;
mixer gate_output_1_562(.a(output_2_562), .b(output_2_2), .y(output_1_562));
wire output_3_562, output_3_2, output_2_562;
mixer gate_output_2_562(.a(output_3_562), .b(output_3_2), .y(output_2_562));
wire output_1_563, output_1_0, output_0_563;
mixer gate_output_0_563(.a(output_1_563), .b(output_1_0), .y(output_0_563));
wire output_2_563, output_2_0, output_1_563;
mixer gate_output_1_563(.a(output_2_563), .b(output_2_0), .y(output_1_563));
wire output_3_563, output_3_0, output_2_563;
mixer gate_output_2_563(.a(output_3_563), .b(output_3_0), .y(output_2_563));
wire output_1_564, output_1_1, output_0_564;
mixer gate_output_0_564(.a(output_1_564), .b(output_1_1), .y(output_0_564));
wire output_2_564, output_2_1, output_1_564;
mixer gate_output_1_564(.a(output_2_564), .b(output_2_1), .y(output_1_564));
wire output_3_564, output_3_1, output_2_564;
mixer gate_output_2_564(.a(output_3_564), .b(output_3_1), .y(output_2_564));
wire output_1_565, output_1_2, output_0_565;
mixer gate_output_0_565(.a(output_1_565), .b(output_1_2), .y(output_0_565));
wire output_2_565, output_2_2, output_1_565;
mixer gate_output_1_565(.a(output_2_565), .b(output_2_2), .y(output_1_565));
wire output_3_565, output_3_2, output_2_565;
mixer gate_output_2_565(.a(output_3_565), .b(output_3_2), .y(output_2_565));
wire output_1_566, output_1_0, output_0_566;
mixer gate_output_0_566(.a(output_1_566), .b(output_1_0), .y(output_0_566));
wire output_2_566, output_2_0, output_1_566;
mixer gate_output_1_566(.a(output_2_566), .b(output_2_0), .y(output_1_566));
wire output_3_566, output_3_0, output_2_566;
mixer gate_output_2_566(.a(output_3_566), .b(output_3_0), .y(output_2_566));
wire output_1_567, output_1_1, output_0_567;
mixer gate_output_0_567(.a(output_1_567), .b(output_1_1), .y(output_0_567));
wire output_2_567, output_2_1, output_1_567;
mixer gate_output_1_567(.a(output_2_567), .b(output_2_1), .y(output_1_567));
wire output_3_567, output_3_1, output_2_567;
mixer gate_output_2_567(.a(output_3_567), .b(output_3_1), .y(output_2_567));
wire output_1_568, output_1_2, output_0_568;
mixer gate_output_0_568(.a(output_1_568), .b(output_1_2), .y(output_0_568));
wire output_2_568, output_2_2, output_1_568;
mixer gate_output_1_568(.a(output_2_568), .b(output_2_2), .y(output_1_568));
wire output_3_568, output_3_2, output_2_568;
mixer gate_output_2_568(.a(output_3_568), .b(output_3_2), .y(output_2_568));
wire output_1_569, output_1_0, output_0_569;
mixer gate_output_0_569(.a(output_1_569), .b(output_1_0), .y(output_0_569));
wire output_2_569, output_2_0, output_1_569;
mixer gate_output_1_569(.a(output_2_569), .b(output_2_0), .y(output_1_569));
wire output_3_569, output_3_0, output_2_569;
mixer gate_output_2_569(.a(output_3_569), .b(output_3_0), .y(output_2_569));
wire output_1_570, output_1_1, output_0_570;
mixer gate_output_0_570(.a(output_1_570), .b(output_1_1), .y(output_0_570));
wire output_2_570, output_2_1, output_1_570;
mixer gate_output_1_570(.a(output_2_570), .b(output_2_1), .y(output_1_570));
wire output_3_570, output_3_1, output_2_570;
mixer gate_output_2_570(.a(output_3_570), .b(output_3_1), .y(output_2_570));
wire output_1_571, output_1_2, output_0_571;
mixer gate_output_0_571(.a(output_1_571), .b(output_1_2), .y(output_0_571));
wire output_2_571, output_2_2, output_1_571;
mixer gate_output_1_571(.a(output_2_571), .b(output_2_2), .y(output_1_571));
wire output_3_571, output_3_2, output_2_571;
mixer gate_output_2_571(.a(output_3_571), .b(output_3_2), .y(output_2_571));
wire output_1_572, output_1_0, output_0_572;
mixer gate_output_0_572(.a(output_1_572), .b(output_1_0), .y(output_0_572));
wire output_2_572, output_2_0, output_1_572;
mixer gate_output_1_572(.a(output_2_572), .b(output_2_0), .y(output_1_572));
wire output_3_572, output_3_0, output_2_572;
mixer gate_output_2_572(.a(output_3_572), .b(output_3_0), .y(output_2_572));
wire output_1_573, output_1_1, output_0_573;
mixer gate_output_0_573(.a(output_1_573), .b(output_1_1), .y(output_0_573));
wire output_2_573, output_2_1, output_1_573;
mixer gate_output_1_573(.a(output_2_573), .b(output_2_1), .y(output_1_573));
wire output_3_573, output_3_1, output_2_573;
mixer gate_output_2_573(.a(output_3_573), .b(output_3_1), .y(output_2_573));
wire output_1_574, output_1_2, output_0_574;
mixer gate_output_0_574(.a(output_1_574), .b(output_1_2), .y(output_0_574));
wire output_2_574, output_2_2, output_1_574;
mixer gate_output_1_574(.a(output_2_574), .b(output_2_2), .y(output_1_574));
wire output_3_574, output_3_2, output_2_574;
mixer gate_output_2_574(.a(output_3_574), .b(output_3_2), .y(output_2_574));
wire output_1_575, output_1_0, output_0_575;
mixer gate_output_0_575(.a(output_1_575), .b(output_1_0), .y(output_0_575));
wire output_2_575, output_2_0, output_1_575;
mixer gate_output_1_575(.a(output_2_575), .b(output_2_0), .y(output_1_575));
wire output_3_575, output_3_0, output_2_575;
mixer gate_output_2_575(.a(output_3_575), .b(output_3_0), .y(output_2_575));
wire output_1_576, output_1_1, output_0_576;
mixer gate_output_0_576(.a(output_1_576), .b(output_1_1), .y(output_0_576));
wire output_2_576, output_2_1, output_1_576;
mixer gate_output_1_576(.a(output_2_576), .b(output_2_1), .y(output_1_576));
wire output_3_576, output_3_1, output_2_576;
mixer gate_output_2_576(.a(output_3_576), .b(output_3_1), .y(output_2_576));
wire output_1_577, output_1_2, output_0_577;
mixer gate_output_0_577(.a(output_1_577), .b(output_1_2), .y(output_0_577));
wire output_2_577, output_2_2, output_1_577;
mixer gate_output_1_577(.a(output_2_577), .b(output_2_2), .y(output_1_577));
wire output_3_577, output_3_2, output_2_577;
mixer gate_output_2_577(.a(output_3_577), .b(output_3_2), .y(output_2_577));
wire output_1_578, output_1_0, output_0_578;
mixer gate_output_0_578(.a(output_1_578), .b(output_1_0), .y(output_0_578));
wire output_2_578, output_2_0, output_1_578;
mixer gate_output_1_578(.a(output_2_578), .b(output_2_0), .y(output_1_578));
wire output_3_578, output_3_0, output_2_578;
mixer gate_output_2_578(.a(output_3_578), .b(output_3_0), .y(output_2_578));
wire output_1_579, output_1_1, output_0_579;
mixer gate_output_0_579(.a(output_1_579), .b(output_1_1), .y(output_0_579));
wire output_2_579, output_2_1, output_1_579;
mixer gate_output_1_579(.a(output_2_579), .b(output_2_1), .y(output_1_579));
wire output_3_579, output_3_1, output_2_579;
mixer gate_output_2_579(.a(output_3_579), .b(output_3_1), .y(output_2_579));
wire output_1_580, output_1_2, output_0_580;
mixer gate_output_0_580(.a(output_1_580), .b(output_1_2), .y(output_0_580));
wire output_2_580, output_2_2, output_1_580;
mixer gate_output_1_580(.a(output_2_580), .b(output_2_2), .y(output_1_580));
wire output_3_580, output_3_2, output_2_580;
mixer gate_output_2_580(.a(output_3_580), .b(output_3_2), .y(output_2_580));
wire output_1_581, output_1_0, output_0_581;
mixer gate_output_0_581(.a(output_1_581), .b(output_1_0), .y(output_0_581));
wire output_2_581, output_2_0, output_1_581;
mixer gate_output_1_581(.a(output_2_581), .b(output_2_0), .y(output_1_581));
wire output_3_581, output_3_0, output_2_581;
mixer gate_output_2_581(.a(output_3_581), .b(output_3_0), .y(output_2_581));
wire output_1_582, output_1_1, output_0_582;
mixer gate_output_0_582(.a(output_1_582), .b(output_1_1), .y(output_0_582));
wire output_2_582, output_2_1, output_1_582;
mixer gate_output_1_582(.a(output_2_582), .b(output_2_1), .y(output_1_582));
wire output_3_582, output_3_1, output_2_582;
mixer gate_output_2_582(.a(output_3_582), .b(output_3_1), .y(output_2_582));
wire output_1_583, output_1_2, output_0_583;
mixer gate_output_0_583(.a(output_1_583), .b(output_1_2), .y(output_0_583));
wire output_2_583, output_2_2, output_1_583;
mixer gate_output_1_583(.a(output_2_583), .b(output_2_2), .y(output_1_583));
wire output_3_583, output_3_2, output_2_583;
mixer gate_output_2_583(.a(output_3_583), .b(output_3_2), .y(output_2_583));
wire output_1_584, output_1_0, output_0_584;
mixer gate_output_0_584(.a(output_1_584), .b(output_1_0), .y(output_0_584));
wire output_2_584, output_2_0, output_1_584;
mixer gate_output_1_584(.a(output_2_584), .b(output_2_0), .y(output_1_584));
wire output_3_584, output_3_0, output_2_584;
mixer gate_output_2_584(.a(output_3_584), .b(output_3_0), .y(output_2_584));
wire output_1_585, output_1_1, output_0_585;
mixer gate_output_0_585(.a(output_1_585), .b(output_1_1), .y(output_0_585));
wire output_2_585, output_2_1, output_1_585;
mixer gate_output_1_585(.a(output_2_585), .b(output_2_1), .y(output_1_585));
wire output_3_585, output_3_1, output_2_585;
mixer gate_output_2_585(.a(output_3_585), .b(output_3_1), .y(output_2_585));
wire output_1_586, output_1_2, output_0_586;
mixer gate_output_0_586(.a(output_1_586), .b(output_1_2), .y(output_0_586));
wire output_2_586, output_2_2, output_1_586;
mixer gate_output_1_586(.a(output_2_586), .b(output_2_2), .y(output_1_586));
wire output_3_586, output_3_2, output_2_586;
mixer gate_output_2_586(.a(output_3_586), .b(output_3_2), .y(output_2_586));
wire output_1_587, output_1_0, output_0_587;
mixer gate_output_0_587(.a(output_1_587), .b(output_1_0), .y(output_0_587));
wire output_2_587, output_2_0, output_1_587;
mixer gate_output_1_587(.a(output_2_587), .b(output_2_0), .y(output_1_587));
wire output_3_587, output_3_0, output_2_587;
mixer gate_output_2_587(.a(output_3_587), .b(output_3_0), .y(output_2_587));
wire output_1_588, output_1_1, output_0_588;
mixer gate_output_0_588(.a(output_1_588), .b(output_1_1), .y(output_0_588));
wire output_2_588, output_2_1, output_1_588;
mixer gate_output_1_588(.a(output_2_588), .b(output_2_1), .y(output_1_588));
wire output_3_588, output_3_1, output_2_588;
mixer gate_output_2_588(.a(output_3_588), .b(output_3_1), .y(output_2_588));
wire output_1_589, output_1_2, output_0_589;
mixer gate_output_0_589(.a(output_1_589), .b(output_1_2), .y(output_0_589));
wire output_2_589, output_2_2, output_1_589;
mixer gate_output_1_589(.a(output_2_589), .b(output_2_2), .y(output_1_589));
wire output_3_589, output_3_2, output_2_589;
mixer gate_output_2_589(.a(output_3_589), .b(output_3_2), .y(output_2_589));
wire output_1_590, output_1_0, output_0_590;
mixer gate_output_0_590(.a(output_1_590), .b(output_1_0), .y(output_0_590));
wire output_2_590, output_2_0, output_1_590;
mixer gate_output_1_590(.a(output_2_590), .b(output_2_0), .y(output_1_590));
wire output_3_590, output_3_0, output_2_590;
mixer gate_output_2_590(.a(output_3_590), .b(output_3_0), .y(output_2_590));
wire output_1_591, output_1_1, output_0_591;
mixer gate_output_0_591(.a(output_1_591), .b(output_1_1), .y(output_0_591));
wire output_2_591, output_2_1, output_1_591;
mixer gate_output_1_591(.a(output_2_591), .b(output_2_1), .y(output_1_591));
wire output_3_591, output_3_1, output_2_591;
mixer gate_output_2_591(.a(output_3_591), .b(output_3_1), .y(output_2_591));
wire output_1_592, output_1_2, output_0_592;
mixer gate_output_0_592(.a(output_1_592), .b(output_1_2), .y(output_0_592));
wire output_2_592, output_2_2, output_1_592;
mixer gate_output_1_592(.a(output_2_592), .b(output_2_2), .y(output_1_592));
wire output_3_592, output_3_2, output_2_592;
mixer gate_output_2_592(.a(output_3_592), .b(output_3_2), .y(output_2_592));
wire output_1_593, output_1_0, output_0_593;
mixer gate_output_0_593(.a(output_1_593), .b(output_1_0), .y(output_0_593));
wire output_2_593, output_2_0, output_1_593;
mixer gate_output_1_593(.a(output_2_593), .b(output_2_0), .y(output_1_593));
wire output_3_593, output_3_0, output_2_593;
mixer gate_output_2_593(.a(output_3_593), .b(output_3_0), .y(output_2_593));
wire output_1_594, output_1_1, output_0_594;
mixer gate_output_0_594(.a(output_1_594), .b(output_1_1), .y(output_0_594));
wire output_2_594, output_2_1, output_1_594;
mixer gate_output_1_594(.a(output_2_594), .b(output_2_1), .y(output_1_594));
wire output_3_594, output_3_1, output_2_594;
mixer gate_output_2_594(.a(output_3_594), .b(output_3_1), .y(output_2_594));
wire output_1_595, output_1_2, output_0_595;
mixer gate_output_0_595(.a(output_1_595), .b(output_1_2), .y(output_0_595));
wire output_2_595, output_2_2, output_1_595;
mixer gate_output_1_595(.a(output_2_595), .b(output_2_2), .y(output_1_595));
wire output_3_595, output_3_2, output_2_595;
mixer gate_output_2_595(.a(output_3_595), .b(output_3_2), .y(output_2_595));
wire output_1_596, output_1_0, output_0_596;
mixer gate_output_0_596(.a(output_1_596), .b(output_1_0), .y(output_0_596));
wire output_2_596, output_2_0, output_1_596;
mixer gate_output_1_596(.a(output_2_596), .b(output_2_0), .y(output_1_596));
wire output_3_596, output_3_0, output_2_596;
mixer gate_output_2_596(.a(output_3_596), .b(output_3_0), .y(output_2_596));
wire output_1_597, output_1_1, output_0_597;
mixer gate_output_0_597(.a(output_1_597), .b(output_1_1), .y(output_0_597));
wire output_2_597, output_2_1, output_1_597;
mixer gate_output_1_597(.a(output_2_597), .b(output_2_1), .y(output_1_597));
wire output_3_597, output_3_1, output_2_597;
mixer gate_output_2_597(.a(output_3_597), .b(output_3_1), .y(output_2_597));
wire output_1_598, output_1_2, output_0_598;
mixer gate_output_0_598(.a(output_1_598), .b(output_1_2), .y(output_0_598));
wire output_2_598, output_2_2, output_1_598;
mixer gate_output_1_598(.a(output_2_598), .b(output_2_2), .y(output_1_598));
wire output_3_598, output_3_2, output_2_598;
mixer gate_output_2_598(.a(output_3_598), .b(output_3_2), .y(output_2_598));
wire output_1_599, output_1_0, output_0_599;
mixer gate_output_0_599(.a(output_1_599), .b(output_1_0), .y(output_0_599));
wire output_2_599, output_2_0, output_1_599;
mixer gate_output_1_599(.a(output_2_599), .b(output_2_0), .y(output_1_599));
wire output_3_599, output_3_0, output_2_599;
mixer gate_output_2_599(.a(output_3_599), .b(output_3_0), .y(output_2_599));
wire output_1_600, output_1_1, output_0_600;
mixer gate_output_0_600(.a(output_1_600), .b(output_1_1), .y(output_0_600));
wire output_2_600, output_2_1, output_1_600;
mixer gate_output_1_600(.a(output_2_600), .b(output_2_1), .y(output_1_600));
wire output_3_600, output_3_1, output_2_600;
mixer gate_output_2_600(.a(output_3_600), .b(output_3_1), .y(output_2_600));
wire output_1_601, output_1_2, output_0_601;
mixer gate_output_0_601(.a(output_1_601), .b(output_1_2), .y(output_0_601));
wire output_2_601, output_2_2, output_1_601;
mixer gate_output_1_601(.a(output_2_601), .b(output_2_2), .y(output_1_601));
wire output_3_601, output_3_2, output_2_601;
mixer gate_output_2_601(.a(output_3_601), .b(output_3_2), .y(output_2_601));
wire output_1_602, output_1_0, output_0_602;
mixer gate_output_0_602(.a(output_1_602), .b(output_1_0), .y(output_0_602));
wire output_2_602, output_2_0, output_1_602;
mixer gate_output_1_602(.a(output_2_602), .b(output_2_0), .y(output_1_602));
wire output_3_602, output_3_0, output_2_602;
mixer gate_output_2_602(.a(output_3_602), .b(output_3_0), .y(output_2_602));
wire output_1_603, output_1_1, output_0_603;
mixer gate_output_0_603(.a(output_1_603), .b(output_1_1), .y(output_0_603));
wire output_2_603, output_2_1, output_1_603;
mixer gate_output_1_603(.a(output_2_603), .b(output_2_1), .y(output_1_603));
wire output_3_603, output_3_1, output_2_603;
mixer gate_output_2_603(.a(output_3_603), .b(output_3_1), .y(output_2_603));
wire output_1_604, output_1_2, output_0_604;
mixer gate_output_0_604(.a(output_1_604), .b(output_1_2), .y(output_0_604));
wire output_2_604, output_2_2, output_1_604;
mixer gate_output_1_604(.a(output_2_604), .b(output_2_2), .y(output_1_604));
wire output_3_604, output_3_2, output_2_604;
mixer gate_output_2_604(.a(output_3_604), .b(output_3_2), .y(output_2_604));
wire output_1_605, output_1_0, output_0_605;
mixer gate_output_0_605(.a(output_1_605), .b(output_1_0), .y(output_0_605));
wire output_2_605, output_2_0, output_1_605;
mixer gate_output_1_605(.a(output_2_605), .b(output_2_0), .y(output_1_605));
wire output_3_605, output_3_0, output_2_605;
mixer gate_output_2_605(.a(output_3_605), .b(output_3_0), .y(output_2_605));
wire output_1_606, output_1_1, output_0_606;
mixer gate_output_0_606(.a(output_1_606), .b(output_1_1), .y(output_0_606));
wire output_2_606, output_2_1, output_1_606;
mixer gate_output_1_606(.a(output_2_606), .b(output_2_1), .y(output_1_606));
wire output_3_606, output_3_1, output_2_606;
mixer gate_output_2_606(.a(output_3_606), .b(output_3_1), .y(output_2_606));
wire output_1_607, output_1_2, output_0_607;
mixer gate_output_0_607(.a(output_1_607), .b(output_1_2), .y(output_0_607));
wire output_2_607, output_2_2, output_1_607;
mixer gate_output_1_607(.a(output_2_607), .b(output_2_2), .y(output_1_607));
wire output_3_607, output_3_2, output_2_607;
mixer gate_output_2_607(.a(output_3_607), .b(output_3_2), .y(output_2_607));
wire output_1_608, output_1_0, output_0_608;
mixer gate_output_0_608(.a(output_1_608), .b(output_1_0), .y(output_0_608));
wire output_2_608, output_2_0, output_1_608;
mixer gate_output_1_608(.a(output_2_608), .b(output_2_0), .y(output_1_608));
wire output_3_608, output_3_0, output_2_608;
mixer gate_output_2_608(.a(output_3_608), .b(output_3_0), .y(output_2_608));
wire output_1_609, output_1_1, output_0_609;
mixer gate_output_0_609(.a(output_1_609), .b(output_1_1), .y(output_0_609));
wire output_2_609, output_2_1, output_1_609;
mixer gate_output_1_609(.a(output_2_609), .b(output_2_1), .y(output_1_609));
wire output_3_609, output_3_1, output_2_609;
mixer gate_output_2_609(.a(output_3_609), .b(output_3_1), .y(output_2_609));
wire output_1_610, output_1_2, output_0_610;
mixer gate_output_0_610(.a(output_1_610), .b(output_1_2), .y(output_0_610));
wire output_2_610, output_2_2, output_1_610;
mixer gate_output_1_610(.a(output_2_610), .b(output_2_2), .y(output_1_610));
wire output_3_610, output_3_2, output_2_610;
mixer gate_output_2_610(.a(output_3_610), .b(output_3_2), .y(output_2_610));
wire output_1_611, output_1_0, output_0_611;
mixer gate_output_0_611(.a(output_1_611), .b(output_1_0), .y(output_0_611));
wire output_2_611, output_2_0, output_1_611;
mixer gate_output_1_611(.a(output_2_611), .b(output_2_0), .y(output_1_611));
wire output_3_611, output_3_0, output_2_611;
mixer gate_output_2_611(.a(output_3_611), .b(output_3_0), .y(output_2_611));
wire output_1_612, output_1_1, output_0_612;
mixer gate_output_0_612(.a(output_1_612), .b(output_1_1), .y(output_0_612));
wire output_2_612, output_2_1, output_1_612;
mixer gate_output_1_612(.a(output_2_612), .b(output_2_1), .y(output_1_612));
wire output_3_612, output_3_1, output_2_612;
mixer gate_output_2_612(.a(output_3_612), .b(output_3_1), .y(output_2_612));
wire output_1_613, output_1_2, output_0_613;
mixer gate_output_0_613(.a(output_1_613), .b(output_1_2), .y(output_0_613));
wire output_2_613, output_2_2, output_1_613;
mixer gate_output_1_613(.a(output_2_613), .b(output_2_2), .y(output_1_613));
wire output_3_613, output_3_2, output_2_613;
mixer gate_output_2_613(.a(output_3_613), .b(output_3_2), .y(output_2_613));
wire output_1_614, output_1_0, output_0_614;
mixer gate_output_0_614(.a(output_1_614), .b(output_1_0), .y(output_0_614));
wire output_2_614, output_2_0, output_1_614;
mixer gate_output_1_614(.a(output_2_614), .b(output_2_0), .y(output_1_614));
wire output_3_614, output_3_0, output_2_614;
mixer gate_output_2_614(.a(output_3_614), .b(output_3_0), .y(output_2_614));
wire output_1_615, output_1_1, output_0_615;
mixer gate_output_0_615(.a(output_1_615), .b(output_1_1), .y(output_0_615));
wire output_2_615, output_2_1, output_1_615;
mixer gate_output_1_615(.a(output_2_615), .b(output_2_1), .y(output_1_615));
wire output_3_615, output_3_1, output_2_615;
mixer gate_output_2_615(.a(output_3_615), .b(output_3_1), .y(output_2_615));
wire output_1_616, output_1_2, output_0_616;
mixer gate_output_0_616(.a(output_1_616), .b(output_1_2), .y(output_0_616));
wire output_2_616, output_2_2, output_1_616;
mixer gate_output_1_616(.a(output_2_616), .b(output_2_2), .y(output_1_616));
wire output_3_616, output_3_2, output_2_616;
mixer gate_output_2_616(.a(output_3_616), .b(output_3_2), .y(output_2_616));
wire output_1_617, output_1_0, output_0_617;
mixer gate_output_0_617(.a(output_1_617), .b(output_1_0), .y(output_0_617));
wire output_2_617, output_2_0, output_1_617;
mixer gate_output_1_617(.a(output_2_617), .b(output_2_0), .y(output_1_617));
wire output_3_617, output_3_0, output_2_617;
mixer gate_output_2_617(.a(output_3_617), .b(output_3_0), .y(output_2_617));
wire output_1_618, output_1_1, output_0_618;
mixer gate_output_0_618(.a(output_1_618), .b(output_1_1), .y(output_0_618));
wire output_2_618, output_2_1, output_1_618;
mixer gate_output_1_618(.a(output_2_618), .b(output_2_1), .y(output_1_618));
wire output_3_618, output_3_1, output_2_618;
mixer gate_output_2_618(.a(output_3_618), .b(output_3_1), .y(output_2_618));
wire output_1_619, output_1_2, output_0_619;
mixer gate_output_0_619(.a(output_1_619), .b(output_1_2), .y(output_0_619));
wire output_2_619, output_2_2, output_1_619;
mixer gate_output_1_619(.a(output_2_619), .b(output_2_2), .y(output_1_619));
wire output_3_619, output_3_2, output_2_619;
mixer gate_output_2_619(.a(output_3_619), .b(output_3_2), .y(output_2_619));
wire output_1_620, output_1_0, output_0_620;
mixer gate_output_0_620(.a(output_1_620), .b(output_1_0), .y(output_0_620));
wire output_2_620, output_2_0, output_1_620;
mixer gate_output_1_620(.a(output_2_620), .b(output_2_0), .y(output_1_620));
wire output_3_620, output_3_0, output_2_620;
mixer gate_output_2_620(.a(output_3_620), .b(output_3_0), .y(output_2_620));
wire output_1_621, output_1_1, output_0_621;
mixer gate_output_0_621(.a(output_1_621), .b(output_1_1), .y(output_0_621));
wire output_2_621, output_2_1, output_1_621;
mixer gate_output_1_621(.a(output_2_621), .b(output_2_1), .y(output_1_621));
wire output_3_621, output_3_1, output_2_621;
mixer gate_output_2_621(.a(output_3_621), .b(output_3_1), .y(output_2_621));
wire output_1_622, output_1_2, output_0_622;
mixer gate_output_0_622(.a(output_1_622), .b(output_1_2), .y(output_0_622));
wire output_2_622, output_2_2, output_1_622;
mixer gate_output_1_622(.a(output_2_622), .b(output_2_2), .y(output_1_622));
wire output_3_622, output_3_2, output_2_622;
mixer gate_output_2_622(.a(output_3_622), .b(output_3_2), .y(output_2_622));
wire output_1_623, output_1_0, output_0_623;
mixer gate_output_0_623(.a(output_1_623), .b(output_1_0), .y(output_0_623));
wire output_2_623, output_2_0, output_1_623;
mixer gate_output_1_623(.a(output_2_623), .b(output_2_0), .y(output_1_623));
wire output_3_623, output_3_0, output_2_623;
mixer gate_output_2_623(.a(output_3_623), .b(output_3_0), .y(output_2_623));
wire output_1_624, output_1_1, output_0_624;
mixer gate_output_0_624(.a(output_1_624), .b(output_1_1), .y(output_0_624));
wire output_2_624, output_2_1, output_1_624;
mixer gate_output_1_624(.a(output_2_624), .b(output_2_1), .y(output_1_624));
wire output_3_624, output_3_1, output_2_624;
mixer gate_output_2_624(.a(output_3_624), .b(output_3_1), .y(output_2_624));
wire output_1_625, output_1_2, output_0_625;
mixer gate_output_0_625(.a(output_1_625), .b(output_1_2), .y(output_0_625));
wire output_2_625, output_2_2, output_1_625;
mixer gate_output_1_625(.a(output_2_625), .b(output_2_2), .y(output_1_625));
wire output_3_625, output_3_2, output_2_625;
mixer gate_output_2_625(.a(output_3_625), .b(output_3_2), .y(output_2_625));
wire output_1_626, output_1_0, output_0_626;
mixer gate_output_0_626(.a(output_1_626), .b(output_1_0), .y(output_0_626));
wire output_2_626, output_2_0, output_1_626;
mixer gate_output_1_626(.a(output_2_626), .b(output_2_0), .y(output_1_626));
wire output_3_626, output_3_0, output_2_626;
mixer gate_output_2_626(.a(output_3_626), .b(output_3_0), .y(output_2_626));
wire output_1_627, output_1_1, output_0_627;
mixer gate_output_0_627(.a(output_1_627), .b(output_1_1), .y(output_0_627));
wire output_2_627, output_2_1, output_1_627;
mixer gate_output_1_627(.a(output_2_627), .b(output_2_1), .y(output_1_627));
wire output_3_627, output_3_1, output_2_627;
mixer gate_output_2_627(.a(output_3_627), .b(output_3_1), .y(output_2_627));
wire output_1_628, output_1_2, output_0_628;
mixer gate_output_0_628(.a(output_1_628), .b(output_1_2), .y(output_0_628));
wire output_2_628, output_2_2, output_1_628;
mixer gate_output_1_628(.a(output_2_628), .b(output_2_2), .y(output_1_628));
wire output_3_628, output_3_2, output_2_628;
mixer gate_output_2_628(.a(output_3_628), .b(output_3_2), .y(output_2_628));
wire output_1_629, output_1_0, output_0_629;
mixer gate_output_0_629(.a(output_1_629), .b(output_1_0), .y(output_0_629));
wire output_2_629, output_2_0, output_1_629;
mixer gate_output_1_629(.a(output_2_629), .b(output_2_0), .y(output_1_629));
wire output_3_629, output_3_0, output_2_629;
mixer gate_output_2_629(.a(output_3_629), .b(output_3_0), .y(output_2_629));
wire output_1_630, output_1_1, output_0_630;
mixer gate_output_0_630(.a(output_1_630), .b(output_1_1), .y(output_0_630));
wire output_2_630, output_2_1, output_1_630;
mixer gate_output_1_630(.a(output_2_630), .b(output_2_1), .y(output_1_630));
wire output_3_630, output_3_1, output_2_630;
mixer gate_output_2_630(.a(output_3_630), .b(output_3_1), .y(output_2_630));
wire output_1_631, output_1_2, output_0_631;
mixer gate_output_0_631(.a(output_1_631), .b(output_1_2), .y(output_0_631));
wire output_2_631, output_2_2, output_1_631;
mixer gate_output_1_631(.a(output_2_631), .b(output_2_2), .y(output_1_631));
wire output_3_631, output_3_2, output_2_631;
mixer gate_output_2_631(.a(output_3_631), .b(output_3_2), .y(output_2_631));
wire output_1_632, output_1_0, output_0_632;
mixer gate_output_0_632(.a(output_1_632), .b(output_1_0), .y(output_0_632));
wire output_2_632, output_2_0, output_1_632;
mixer gate_output_1_632(.a(output_2_632), .b(output_2_0), .y(output_1_632));
wire output_3_632, output_3_0, output_2_632;
mixer gate_output_2_632(.a(output_3_632), .b(output_3_0), .y(output_2_632));
wire output_1_633, output_1_1, output_0_633;
mixer gate_output_0_633(.a(output_1_633), .b(output_1_1), .y(output_0_633));
wire output_2_633, output_2_1, output_1_633;
mixer gate_output_1_633(.a(output_2_633), .b(output_2_1), .y(output_1_633));
wire output_3_633, output_3_1, output_2_633;
mixer gate_output_2_633(.a(output_3_633), .b(output_3_1), .y(output_2_633));
wire output_1_634, output_1_2, output_0_634;
mixer gate_output_0_634(.a(output_1_634), .b(output_1_2), .y(output_0_634));
wire output_2_634, output_2_2, output_1_634;
mixer gate_output_1_634(.a(output_2_634), .b(output_2_2), .y(output_1_634));
wire output_3_634, output_3_2, output_2_634;
mixer gate_output_2_634(.a(output_3_634), .b(output_3_2), .y(output_2_634));
wire output_1_635, output_1_0, output_0_635;
mixer gate_output_0_635(.a(output_1_635), .b(output_1_0), .y(output_0_635));
wire output_2_635, output_2_0, output_1_635;
mixer gate_output_1_635(.a(output_2_635), .b(output_2_0), .y(output_1_635));
wire output_3_635, output_3_0, output_2_635;
mixer gate_output_2_635(.a(output_3_635), .b(output_3_0), .y(output_2_635));
wire output_1_636, output_1_1, output_0_636;
mixer gate_output_0_636(.a(output_1_636), .b(output_1_1), .y(output_0_636));
wire output_2_636, output_2_1, output_1_636;
mixer gate_output_1_636(.a(output_2_636), .b(output_2_1), .y(output_1_636));
wire output_3_636, output_3_1, output_2_636;
mixer gate_output_2_636(.a(output_3_636), .b(output_3_1), .y(output_2_636));
wire output_1_637, output_1_2, output_0_637;
mixer gate_output_0_637(.a(output_1_637), .b(output_1_2), .y(output_0_637));
wire output_2_637, output_2_2, output_1_637;
mixer gate_output_1_637(.a(output_2_637), .b(output_2_2), .y(output_1_637));
wire output_3_637, output_3_2, output_2_637;
mixer gate_output_2_637(.a(output_3_637), .b(output_3_2), .y(output_2_637));
wire output_1_638, output_1_0, output_0_638;
mixer gate_output_0_638(.a(output_1_638), .b(output_1_0), .y(output_0_638));
wire output_2_638, output_2_0, output_1_638;
mixer gate_output_1_638(.a(output_2_638), .b(output_2_0), .y(output_1_638));
wire output_3_638, output_3_0, output_2_638;
mixer gate_output_2_638(.a(output_3_638), .b(output_3_0), .y(output_2_638));
wire output_1_639, output_1_1, output_0_639;
mixer gate_output_0_639(.a(output_1_639), .b(output_1_1), .y(output_0_639));
wire output_2_639, output_2_1, output_1_639;
mixer gate_output_1_639(.a(output_2_639), .b(output_2_1), .y(output_1_639));
wire output_3_639, output_3_1, output_2_639;
mixer gate_output_2_639(.a(output_3_639), .b(output_3_1), .y(output_2_639));
wire output_1_640, output_1_2, output_0_640;
mixer gate_output_0_640(.a(output_1_640), .b(output_1_2), .y(output_0_640));
wire output_2_640, output_2_2, output_1_640;
mixer gate_output_1_640(.a(output_2_640), .b(output_2_2), .y(output_1_640));
wire output_3_640, output_3_2, output_2_640;
mixer gate_output_2_640(.a(output_3_640), .b(output_3_2), .y(output_2_640));
wire output_1_641, output_1_0, output_0_641;
mixer gate_output_0_641(.a(output_1_641), .b(output_1_0), .y(output_0_641));
wire output_2_641, output_2_0, output_1_641;
mixer gate_output_1_641(.a(output_2_641), .b(output_2_0), .y(output_1_641));
wire output_3_641, output_3_0, output_2_641;
mixer gate_output_2_641(.a(output_3_641), .b(output_3_0), .y(output_2_641));
wire output_1_642, output_1_1, output_0_642;
mixer gate_output_0_642(.a(output_1_642), .b(output_1_1), .y(output_0_642));
wire output_2_642, output_2_1, output_1_642;
mixer gate_output_1_642(.a(output_2_642), .b(output_2_1), .y(output_1_642));
wire output_3_642, output_3_1, output_2_642;
mixer gate_output_2_642(.a(output_3_642), .b(output_3_1), .y(output_2_642));
wire output_1_643, output_1_2, output_0_643;
mixer gate_output_0_643(.a(output_1_643), .b(output_1_2), .y(output_0_643));
wire output_2_643, output_2_2, output_1_643;
mixer gate_output_1_643(.a(output_2_643), .b(output_2_2), .y(output_1_643));
wire output_3_643, output_3_2, output_2_643;
mixer gate_output_2_643(.a(output_3_643), .b(output_3_2), .y(output_2_643));
wire output_1_644, output_1_0, output_0_644;
mixer gate_output_0_644(.a(output_1_644), .b(output_1_0), .y(output_0_644));
wire output_2_644, output_2_0, output_1_644;
mixer gate_output_1_644(.a(output_2_644), .b(output_2_0), .y(output_1_644));
wire output_3_644, output_3_0, output_2_644;
mixer gate_output_2_644(.a(output_3_644), .b(output_3_0), .y(output_2_644));
wire output_1_645, output_1_1, output_0_645;
mixer gate_output_0_645(.a(output_1_645), .b(output_1_1), .y(output_0_645));
wire output_2_645, output_2_1, output_1_645;
mixer gate_output_1_645(.a(output_2_645), .b(output_2_1), .y(output_1_645));
wire output_3_645, output_3_1, output_2_645;
mixer gate_output_2_645(.a(output_3_645), .b(output_3_1), .y(output_2_645));
wire output_1_646, output_1_2, output_0_646;
mixer gate_output_0_646(.a(output_1_646), .b(output_1_2), .y(output_0_646));
wire output_2_646, output_2_2, output_1_646;
mixer gate_output_1_646(.a(output_2_646), .b(output_2_2), .y(output_1_646));
wire output_3_646, output_3_2, output_2_646;
mixer gate_output_2_646(.a(output_3_646), .b(output_3_2), .y(output_2_646));
wire output_1_647, output_1_0, output_0_647;
mixer gate_output_0_647(.a(output_1_647), .b(output_1_0), .y(output_0_647));
wire output_2_647, output_2_0, output_1_647;
mixer gate_output_1_647(.a(output_2_647), .b(output_2_0), .y(output_1_647));
wire output_3_647, output_3_0, output_2_647;
mixer gate_output_2_647(.a(output_3_647), .b(output_3_0), .y(output_2_647));
wire output_1_648, output_1_1, output_0_648;
mixer gate_output_0_648(.a(output_1_648), .b(output_1_1), .y(output_0_648));
wire output_2_648, output_2_1, output_1_648;
mixer gate_output_1_648(.a(output_2_648), .b(output_2_1), .y(output_1_648));
wire output_3_648, output_3_1, output_2_648;
mixer gate_output_2_648(.a(output_3_648), .b(output_3_1), .y(output_2_648));
wire output_1_649, output_1_2, output_0_649;
mixer gate_output_0_649(.a(output_1_649), .b(output_1_2), .y(output_0_649));
wire output_2_649, output_2_2, output_1_649;
mixer gate_output_1_649(.a(output_2_649), .b(output_2_2), .y(output_1_649));
wire output_3_649, output_3_2, output_2_649;
mixer gate_output_2_649(.a(output_3_649), .b(output_3_2), .y(output_2_649));
wire output_1_650, output_1_0, output_0_650;
mixer gate_output_0_650(.a(output_1_650), .b(output_1_0), .y(output_0_650));
wire output_2_650, output_2_0, output_1_650;
mixer gate_output_1_650(.a(output_2_650), .b(output_2_0), .y(output_1_650));
wire output_3_650, output_3_0, output_2_650;
mixer gate_output_2_650(.a(output_3_650), .b(output_3_0), .y(output_2_650));
wire output_1_651, output_1_1, output_0_651;
mixer gate_output_0_651(.a(output_1_651), .b(output_1_1), .y(output_0_651));
wire output_2_651, output_2_1, output_1_651;
mixer gate_output_1_651(.a(output_2_651), .b(output_2_1), .y(output_1_651));
wire output_3_651, output_3_1, output_2_651;
mixer gate_output_2_651(.a(output_3_651), .b(output_3_1), .y(output_2_651));
wire output_1_652, output_1_2, output_0_652;
mixer gate_output_0_652(.a(output_1_652), .b(output_1_2), .y(output_0_652));
wire output_2_652, output_2_2, output_1_652;
mixer gate_output_1_652(.a(output_2_652), .b(output_2_2), .y(output_1_652));
wire output_3_652, output_3_2, output_2_652;
mixer gate_output_2_652(.a(output_3_652), .b(output_3_2), .y(output_2_652));
wire output_1_653, output_1_0, output_0_653;
mixer gate_output_0_653(.a(output_1_653), .b(output_1_0), .y(output_0_653));
wire output_2_653, output_2_0, output_1_653;
mixer gate_output_1_653(.a(output_2_653), .b(output_2_0), .y(output_1_653));
wire output_3_653, output_3_0, output_2_653;
mixer gate_output_2_653(.a(output_3_653), .b(output_3_0), .y(output_2_653));
wire output_1_654, output_1_1, output_0_654;
mixer gate_output_0_654(.a(output_1_654), .b(output_1_1), .y(output_0_654));
wire output_2_654, output_2_1, output_1_654;
mixer gate_output_1_654(.a(output_2_654), .b(output_2_1), .y(output_1_654));
wire output_3_654, output_3_1, output_2_654;
mixer gate_output_2_654(.a(output_3_654), .b(output_3_1), .y(output_2_654));
wire output_1_655, output_1_2, output_0_655;
mixer gate_output_0_655(.a(output_1_655), .b(output_1_2), .y(output_0_655));
wire output_2_655, output_2_2, output_1_655;
mixer gate_output_1_655(.a(output_2_655), .b(output_2_2), .y(output_1_655));
wire output_3_655, output_3_2, output_2_655;
mixer gate_output_2_655(.a(output_3_655), .b(output_3_2), .y(output_2_655));
wire output_1_656, output_1_0, output_0_656;
mixer gate_output_0_656(.a(output_1_656), .b(output_1_0), .y(output_0_656));
wire output_2_656, output_2_0, output_1_656;
mixer gate_output_1_656(.a(output_2_656), .b(output_2_0), .y(output_1_656));
wire output_3_656, output_3_0, output_2_656;
mixer gate_output_2_656(.a(output_3_656), .b(output_3_0), .y(output_2_656));
wire output_1_657, output_1_1, output_0_657;
mixer gate_output_0_657(.a(output_1_657), .b(output_1_1), .y(output_0_657));
wire output_2_657, output_2_1, output_1_657;
mixer gate_output_1_657(.a(output_2_657), .b(output_2_1), .y(output_1_657));
wire output_3_657, output_3_1, output_2_657;
mixer gate_output_2_657(.a(output_3_657), .b(output_3_1), .y(output_2_657));
wire output_1_658, output_1_2, output_0_658;
mixer gate_output_0_658(.a(output_1_658), .b(output_1_2), .y(output_0_658));
wire output_2_658, output_2_2, output_1_658;
mixer gate_output_1_658(.a(output_2_658), .b(output_2_2), .y(output_1_658));
wire output_3_658, output_3_2, output_2_658;
mixer gate_output_2_658(.a(output_3_658), .b(output_3_2), .y(output_2_658));
wire output_1_659, output_1_0, output_0_659;
mixer gate_output_0_659(.a(output_1_659), .b(output_1_0), .y(output_0_659));
wire output_2_659, output_2_0, output_1_659;
mixer gate_output_1_659(.a(output_2_659), .b(output_2_0), .y(output_1_659));
wire output_3_659, output_3_0, output_2_659;
mixer gate_output_2_659(.a(output_3_659), .b(output_3_0), .y(output_2_659));
wire output_1_660, output_1_1, output_0_660;
mixer gate_output_0_660(.a(output_1_660), .b(output_1_1), .y(output_0_660));
wire output_2_660, output_2_1, output_1_660;
mixer gate_output_1_660(.a(output_2_660), .b(output_2_1), .y(output_1_660));
wire output_3_660, output_3_1, output_2_660;
mixer gate_output_2_660(.a(output_3_660), .b(output_3_1), .y(output_2_660));
wire output_1_661, output_1_2, output_0_661;
mixer gate_output_0_661(.a(output_1_661), .b(output_1_2), .y(output_0_661));
wire output_2_661, output_2_2, output_1_661;
mixer gate_output_1_661(.a(output_2_661), .b(output_2_2), .y(output_1_661));
wire output_3_661, output_3_2, output_2_661;
mixer gate_output_2_661(.a(output_3_661), .b(output_3_2), .y(output_2_661));
wire output_1_662, output_1_0, output_0_662;
mixer gate_output_0_662(.a(output_1_662), .b(output_1_0), .y(output_0_662));
wire output_2_662, output_2_0, output_1_662;
mixer gate_output_1_662(.a(output_2_662), .b(output_2_0), .y(output_1_662));
wire output_3_662, output_3_0, output_2_662;
mixer gate_output_2_662(.a(output_3_662), .b(output_3_0), .y(output_2_662));
wire output_1_663, output_1_1, output_0_663;
mixer gate_output_0_663(.a(output_1_663), .b(output_1_1), .y(output_0_663));
wire output_2_663, output_2_1, output_1_663;
mixer gate_output_1_663(.a(output_2_663), .b(output_2_1), .y(output_1_663));
wire output_3_663, output_3_1, output_2_663;
mixer gate_output_2_663(.a(output_3_663), .b(output_3_1), .y(output_2_663));
wire output_1_664, output_1_2, output_0_664;
mixer gate_output_0_664(.a(output_1_664), .b(output_1_2), .y(output_0_664));
wire output_2_664, output_2_2, output_1_664;
mixer gate_output_1_664(.a(output_2_664), .b(output_2_2), .y(output_1_664));
wire output_3_664, output_3_2, output_2_664;
mixer gate_output_2_664(.a(output_3_664), .b(output_3_2), .y(output_2_664));
wire output_1_665, output_1_0, output_0_665;
mixer gate_output_0_665(.a(output_1_665), .b(output_1_0), .y(output_0_665));
wire output_2_665, output_2_0, output_1_665;
mixer gate_output_1_665(.a(output_2_665), .b(output_2_0), .y(output_1_665));
wire output_3_665, output_3_0, output_2_665;
mixer gate_output_2_665(.a(output_3_665), .b(output_3_0), .y(output_2_665));
wire output_1_666, output_1_1, output_0_666;
mixer gate_output_0_666(.a(output_1_666), .b(output_1_1), .y(output_0_666));
wire output_2_666, output_2_1, output_1_666;
mixer gate_output_1_666(.a(output_2_666), .b(output_2_1), .y(output_1_666));
wire output_3_666, output_3_1, output_2_666;
mixer gate_output_2_666(.a(output_3_666), .b(output_3_1), .y(output_2_666));
wire output_1_667, output_1_2, output_0_667;
mixer gate_output_0_667(.a(output_1_667), .b(output_1_2), .y(output_0_667));
wire output_2_667, output_2_2, output_1_667;
mixer gate_output_1_667(.a(output_2_667), .b(output_2_2), .y(output_1_667));
wire output_3_667, output_3_2, output_2_667;
mixer gate_output_2_667(.a(output_3_667), .b(output_3_2), .y(output_2_667));
wire output_1_668, output_1_0, output_0_668;
mixer gate_output_0_668(.a(output_1_668), .b(output_1_0), .y(output_0_668));
wire output_2_668, output_2_0, output_1_668;
mixer gate_output_1_668(.a(output_2_668), .b(output_2_0), .y(output_1_668));
wire output_3_668, output_3_0, output_2_668;
mixer gate_output_2_668(.a(output_3_668), .b(output_3_0), .y(output_2_668));
wire output_1_669, output_1_1, output_0_669;
mixer gate_output_0_669(.a(output_1_669), .b(output_1_1), .y(output_0_669));
wire output_2_669, output_2_1, output_1_669;
mixer gate_output_1_669(.a(output_2_669), .b(output_2_1), .y(output_1_669));
wire output_3_669, output_3_1, output_2_669;
mixer gate_output_2_669(.a(output_3_669), .b(output_3_1), .y(output_2_669));
wire output_1_670, output_1_2, output_0_670;
mixer gate_output_0_670(.a(output_1_670), .b(output_1_2), .y(output_0_670));
wire output_2_670, output_2_2, output_1_670;
mixer gate_output_1_670(.a(output_2_670), .b(output_2_2), .y(output_1_670));
wire output_3_670, output_3_2, output_2_670;
mixer gate_output_2_670(.a(output_3_670), .b(output_3_2), .y(output_2_670));
wire output_1_671, output_1_0, output_0_671;
mixer gate_output_0_671(.a(output_1_671), .b(output_1_0), .y(output_0_671));
wire output_2_671, output_2_0, output_1_671;
mixer gate_output_1_671(.a(output_2_671), .b(output_2_0), .y(output_1_671));
wire output_3_671, output_3_0, output_2_671;
mixer gate_output_2_671(.a(output_3_671), .b(output_3_0), .y(output_2_671));
wire output_1_672, output_1_1, output_0_672;
mixer gate_output_0_672(.a(output_1_672), .b(output_1_1), .y(output_0_672));
wire output_2_672, output_2_1, output_1_672;
mixer gate_output_1_672(.a(output_2_672), .b(output_2_1), .y(output_1_672));
wire output_3_672, output_3_1, output_2_672;
mixer gate_output_2_672(.a(output_3_672), .b(output_3_1), .y(output_2_672));
wire output_1_673, output_1_2, output_0_673;
mixer gate_output_0_673(.a(output_1_673), .b(output_1_2), .y(output_0_673));
wire output_2_673, output_2_2, output_1_673;
mixer gate_output_1_673(.a(output_2_673), .b(output_2_2), .y(output_1_673));
wire output_3_673, output_3_2, output_2_673;
mixer gate_output_2_673(.a(output_3_673), .b(output_3_2), .y(output_2_673));
wire output_1_674, output_1_0, output_0_674;
mixer gate_output_0_674(.a(output_1_674), .b(output_1_0), .y(output_0_674));
wire output_2_674, output_2_0, output_1_674;
mixer gate_output_1_674(.a(output_2_674), .b(output_2_0), .y(output_1_674));
wire output_3_674, output_3_0, output_2_674;
mixer gate_output_2_674(.a(output_3_674), .b(output_3_0), .y(output_2_674));
wire output_1_675, output_1_1, output_0_675;
mixer gate_output_0_675(.a(output_1_675), .b(output_1_1), .y(output_0_675));
wire output_2_675, output_2_1, output_1_675;
mixer gate_output_1_675(.a(output_2_675), .b(output_2_1), .y(output_1_675));
wire output_3_675, output_3_1, output_2_675;
mixer gate_output_2_675(.a(output_3_675), .b(output_3_1), .y(output_2_675));
wire output_1_676, output_1_2, output_0_676;
mixer gate_output_0_676(.a(output_1_676), .b(output_1_2), .y(output_0_676));
wire output_2_676, output_2_2, output_1_676;
mixer gate_output_1_676(.a(output_2_676), .b(output_2_2), .y(output_1_676));
wire output_3_676, output_3_2, output_2_676;
mixer gate_output_2_676(.a(output_3_676), .b(output_3_2), .y(output_2_676));
wire output_1_677, output_1_0, output_0_677;
mixer gate_output_0_677(.a(output_1_677), .b(output_1_0), .y(output_0_677));
wire output_2_677, output_2_0, output_1_677;
mixer gate_output_1_677(.a(output_2_677), .b(output_2_0), .y(output_1_677));
wire output_3_677, output_3_0, output_2_677;
mixer gate_output_2_677(.a(output_3_677), .b(output_3_0), .y(output_2_677));
wire output_1_678, output_1_1, output_0_678;
mixer gate_output_0_678(.a(output_1_678), .b(output_1_1), .y(output_0_678));
wire output_2_678, output_2_1, output_1_678;
mixer gate_output_1_678(.a(output_2_678), .b(output_2_1), .y(output_1_678));
wire output_3_678, output_3_1, output_2_678;
mixer gate_output_2_678(.a(output_3_678), .b(output_3_1), .y(output_2_678));
wire output_1_679, output_1_2, output_0_679;
mixer gate_output_0_679(.a(output_1_679), .b(output_1_2), .y(output_0_679));
wire output_2_679, output_2_2, output_1_679;
mixer gate_output_1_679(.a(output_2_679), .b(output_2_2), .y(output_1_679));
wire output_3_679, output_3_2, output_2_679;
mixer gate_output_2_679(.a(output_3_679), .b(output_3_2), .y(output_2_679));
wire output_1_680, output_1_0, output_0_680;
mixer gate_output_0_680(.a(output_1_680), .b(output_1_0), .y(output_0_680));
wire output_2_680, output_2_0, output_1_680;
mixer gate_output_1_680(.a(output_2_680), .b(output_2_0), .y(output_1_680));
wire output_3_680, output_3_0, output_2_680;
mixer gate_output_2_680(.a(output_3_680), .b(output_3_0), .y(output_2_680));
wire output_1_681, output_1_1, output_0_681;
mixer gate_output_0_681(.a(output_1_681), .b(output_1_1), .y(output_0_681));
wire output_2_681, output_2_1, output_1_681;
mixer gate_output_1_681(.a(output_2_681), .b(output_2_1), .y(output_1_681));
wire output_3_681, output_3_1, output_2_681;
mixer gate_output_2_681(.a(output_3_681), .b(output_3_1), .y(output_2_681));
wire output_1_682, output_1_2, output_0_682;
mixer gate_output_0_682(.a(output_1_682), .b(output_1_2), .y(output_0_682));
wire output_2_682, output_2_2, output_1_682;
mixer gate_output_1_682(.a(output_2_682), .b(output_2_2), .y(output_1_682));
wire output_3_682, output_3_2, output_2_682;
mixer gate_output_2_682(.a(output_3_682), .b(output_3_2), .y(output_2_682));
wire output_1_683, output_1_0, output_0_683;
mixer gate_output_0_683(.a(output_1_683), .b(output_1_0), .y(output_0_683));
wire output_2_683, output_2_0, output_1_683;
mixer gate_output_1_683(.a(output_2_683), .b(output_2_0), .y(output_1_683));
wire output_3_683, output_3_0, output_2_683;
mixer gate_output_2_683(.a(output_3_683), .b(output_3_0), .y(output_2_683));
wire output_1_684, output_1_1, output_0_684;
mixer gate_output_0_684(.a(output_1_684), .b(output_1_1), .y(output_0_684));
wire output_2_684, output_2_1, output_1_684;
mixer gate_output_1_684(.a(output_2_684), .b(output_2_1), .y(output_1_684));
wire output_3_684, output_3_1, output_2_684;
mixer gate_output_2_684(.a(output_3_684), .b(output_3_1), .y(output_2_684));
wire output_1_685, output_1_2, output_0_685;
mixer gate_output_0_685(.a(output_1_685), .b(output_1_2), .y(output_0_685));
wire output_2_685, output_2_2, output_1_685;
mixer gate_output_1_685(.a(output_2_685), .b(output_2_2), .y(output_1_685));
wire output_3_685, output_3_2, output_2_685;
mixer gate_output_2_685(.a(output_3_685), .b(output_3_2), .y(output_2_685));
wire output_1_686, output_1_0, output_0_686;
mixer gate_output_0_686(.a(output_1_686), .b(output_1_0), .y(output_0_686));
wire output_2_686, output_2_0, output_1_686;
mixer gate_output_1_686(.a(output_2_686), .b(output_2_0), .y(output_1_686));
wire output_3_686, output_3_0, output_2_686;
mixer gate_output_2_686(.a(output_3_686), .b(output_3_0), .y(output_2_686));
wire output_1_687, output_1_1, output_0_687;
mixer gate_output_0_687(.a(output_1_687), .b(output_1_1), .y(output_0_687));
wire output_2_687, output_2_1, output_1_687;
mixer gate_output_1_687(.a(output_2_687), .b(output_2_1), .y(output_1_687));
wire output_3_687, output_3_1, output_2_687;
mixer gate_output_2_687(.a(output_3_687), .b(output_3_1), .y(output_2_687));
wire output_1_688, output_1_2, output_0_688;
mixer gate_output_0_688(.a(output_1_688), .b(output_1_2), .y(output_0_688));
wire output_2_688, output_2_2, output_1_688;
mixer gate_output_1_688(.a(output_2_688), .b(output_2_2), .y(output_1_688));
wire output_3_688, output_3_2, output_2_688;
mixer gate_output_2_688(.a(output_3_688), .b(output_3_2), .y(output_2_688));
wire output_1_689, output_1_0, output_0_689;
mixer gate_output_0_689(.a(output_1_689), .b(output_1_0), .y(output_0_689));
wire output_2_689, output_2_0, output_1_689;
mixer gate_output_1_689(.a(output_2_689), .b(output_2_0), .y(output_1_689));
wire output_3_689, output_3_0, output_2_689;
mixer gate_output_2_689(.a(output_3_689), .b(output_3_0), .y(output_2_689));
wire output_1_690, output_1_1, output_0_690;
mixer gate_output_0_690(.a(output_1_690), .b(output_1_1), .y(output_0_690));
wire output_2_690, output_2_1, output_1_690;
mixer gate_output_1_690(.a(output_2_690), .b(output_2_1), .y(output_1_690));
wire output_3_690, output_3_1, output_2_690;
mixer gate_output_2_690(.a(output_3_690), .b(output_3_1), .y(output_2_690));
wire output_1_691, output_1_2, output_0_691;
mixer gate_output_0_691(.a(output_1_691), .b(output_1_2), .y(output_0_691));
wire output_2_691, output_2_2, output_1_691;
mixer gate_output_1_691(.a(output_2_691), .b(output_2_2), .y(output_1_691));
wire output_3_691, output_3_2, output_2_691;
mixer gate_output_2_691(.a(output_3_691), .b(output_3_2), .y(output_2_691));
wire output_1_692, output_1_0, output_0_692;
mixer gate_output_0_692(.a(output_1_692), .b(output_1_0), .y(output_0_692));
wire output_2_692, output_2_0, output_1_692;
mixer gate_output_1_692(.a(output_2_692), .b(output_2_0), .y(output_1_692));
wire output_3_692, output_3_0, output_2_692;
mixer gate_output_2_692(.a(output_3_692), .b(output_3_0), .y(output_2_692));
wire output_1_693, output_1_1, output_0_693;
mixer gate_output_0_693(.a(output_1_693), .b(output_1_1), .y(output_0_693));
wire output_2_693, output_2_1, output_1_693;
mixer gate_output_1_693(.a(output_2_693), .b(output_2_1), .y(output_1_693));
wire output_3_693, output_3_1, output_2_693;
mixer gate_output_2_693(.a(output_3_693), .b(output_3_1), .y(output_2_693));
wire output_1_694, output_1_2, output_0_694;
mixer gate_output_0_694(.a(output_1_694), .b(output_1_2), .y(output_0_694));
wire output_2_694, output_2_2, output_1_694;
mixer gate_output_1_694(.a(output_2_694), .b(output_2_2), .y(output_1_694));
wire output_3_694, output_3_2, output_2_694;
mixer gate_output_2_694(.a(output_3_694), .b(output_3_2), .y(output_2_694));
wire output_1_695, output_1_0, output_0_695;
mixer gate_output_0_695(.a(output_1_695), .b(output_1_0), .y(output_0_695));
wire output_2_695, output_2_0, output_1_695;
mixer gate_output_1_695(.a(output_2_695), .b(output_2_0), .y(output_1_695));
wire output_3_695, output_3_0, output_2_695;
mixer gate_output_2_695(.a(output_3_695), .b(output_3_0), .y(output_2_695));
wire output_1_696, output_1_1, output_0_696;
mixer gate_output_0_696(.a(output_1_696), .b(output_1_1), .y(output_0_696));
wire output_2_696, output_2_1, output_1_696;
mixer gate_output_1_696(.a(output_2_696), .b(output_2_1), .y(output_1_696));
wire output_3_696, output_3_1, output_2_696;
mixer gate_output_2_696(.a(output_3_696), .b(output_3_1), .y(output_2_696));
wire output_1_697, output_1_2, output_0_697;
mixer gate_output_0_697(.a(output_1_697), .b(output_1_2), .y(output_0_697));
wire output_2_697, output_2_2, output_1_697;
mixer gate_output_1_697(.a(output_2_697), .b(output_2_2), .y(output_1_697));
wire output_3_697, output_3_2, output_2_697;
mixer gate_output_2_697(.a(output_3_697), .b(output_3_2), .y(output_2_697));
wire output_1_698, output_1_0, output_0_698;
mixer gate_output_0_698(.a(output_1_698), .b(output_1_0), .y(output_0_698));
wire output_2_698, output_2_0, output_1_698;
mixer gate_output_1_698(.a(output_2_698), .b(output_2_0), .y(output_1_698));
wire output_3_698, output_3_0, output_2_698;
mixer gate_output_2_698(.a(output_3_698), .b(output_3_0), .y(output_2_698));
wire output_1_699, output_1_1, output_0_699;
mixer gate_output_0_699(.a(output_1_699), .b(output_1_1), .y(output_0_699));
wire output_2_699, output_2_1, output_1_699;
mixer gate_output_1_699(.a(output_2_699), .b(output_2_1), .y(output_1_699));
wire output_3_699, output_3_1, output_2_699;
mixer gate_output_2_699(.a(output_3_699), .b(output_3_1), .y(output_2_699));
wire output_1_700, output_1_2, output_0_700;
mixer gate_output_0_700(.a(output_1_700), .b(output_1_2), .y(output_0_700));
wire output_2_700, output_2_2, output_1_700;
mixer gate_output_1_700(.a(output_2_700), .b(output_2_2), .y(output_1_700));
wire output_3_700, output_3_2, output_2_700;
mixer gate_output_2_700(.a(output_3_700), .b(output_3_2), .y(output_2_700));
wire output_1_701, output_1_0, output_0_701;
mixer gate_output_0_701(.a(output_1_701), .b(output_1_0), .y(output_0_701));
wire output_2_701, output_2_0, output_1_701;
mixer gate_output_1_701(.a(output_2_701), .b(output_2_0), .y(output_1_701));
wire output_3_701, output_3_0, output_2_701;
mixer gate_output_2_701(.a(output_3_701), .b(output_3_0), .y(output_2_701));
wire output_1_702, output_1_1, output_0_702;
mixer gate_output_0_702(.a(output_1_702), .b(output_1_1), .y(output_0_702));
wire output_2_702, output_2_1, output_1_702;
mixer gate_output_1_702(.a(output_2_702), .b(output_2_1), .y(output_1_702));
wire output_3_702, output_3_1, output_2_702;
mixer gate_output_2_702(.a(output_3_702), .b(output_3_1), .y(output_2_702));
wire output_1_703, output_1_2, output_0_703;
mixer gate_output_0_703(.a(output_1_703), .b(output_1_2), .y(output_0_703));
wire output_2_703, output_2_2, output_1_703;
mixer gate_output_1_703(.a(output_2_703), .b(output_2_2), .y(output_1_703));
wire output_3_703, output_3_2, output_2_703;
mixer gate_output_2_703(.a(output_3_703), .b(output_3_2), .y(output_2_703));
wire output_1_704, output_1_0, output_0_704;
mixer gate_output_0_704(.a(output_1_704), .b(output_1_0), .y(output_0_704));
wire output_2_704, output_2_0, output_1_704;
mixer gate_output_1_704(.a(output_2_704), .b(output_2_0), .y(output_1_704));
wire output_3_704, output_3_0, output_2_704;
mixer gate_output_2_704(.a(output_3_704), .b(output_3_0), .y(output_2_704));
wire output_1_705, output_1_1, output_0_705;
mixer gate_output_0_705(.a(output_1_705), .b(output_1_1), .y(output_0_705));
wire output_2_705, output_2_1, output_1_705;
mixer gate_output_1_705(.a(output_2_705), .b(output_2_1), .y(output_1_705));
wire output_3_705, output_3_1, output_2_705;
mixer gate_output_2_705(.a(output_3_705), .b(output_3_1), .y(output_2_705));
wire output_1_706, output_1_2, output_0_706;
mixer gate_output_0_706(.a(output_1_706), .b(output_1_2), .y(output_0_706));
wire output_2_706, output_2_2, output_1_706;
mixer gate_output_1_706(.a(output_2_706), .b(output_2_2), .y(output_1_706));
wire output_3_706, output_3_2, output_2_706;
mixer gate_output_2_706(.a(output_3_706), .b(output_3_2), .y(output_2_706));
wire output_1_707, output_1_0, output_0_707;
mixer gate_output_0_707(.a(output_1_707), .b(output_1_0), .y(output_0_707));
wire output_2_707, output_2_0, output_1_707;
mixer gate_output_1_707(.a(output_2_707), .b(output_2_0), .y(output_1_707));
wire output_3_707, output_3_0, output_2_707;
mixer gate_output_2_707(.a(output_3_707), .b(output_3_0), .y(output_2_707));
wire output_1_708, output_1_1, output_0_708;
mixer gate_output_0_708(.a(output_1_708), .b(output_1_1), .y(output_0_708));
wire output_2_708, output_2_1, output_1_708;
mixer gate_output_1_708(.a(output_2_708), .b(output_2_1), .y(output_1_708));
wire output_3_708, output_3_1, output_2_708;
mixer gate_output_2_708(.a(output_3_708), .b(output_3_1), .y(output_2_708));
wire output_1_709, output_1_2, output_0_709;
mixer gate_output_0_709(.a(output_1_709), .b(output_1_2), .y(output_0_709));
wire output_2_709, output_2_2, output_1_709;
mixer gate_output_1_709(.a(output_2_709), .b(output_2_2), .y(output_1_709));
wire output_3_709, output_3_2, output_2_709;
mixer gate_output_2_709(.a(output_3_709), .b(output_3_2), .y(output_2_709));
wire output_1_710, output_1_0, output_0_710;
mixer gate_output_0_710(.a(output_1_710), .b(output_1_0), .y(output_0_710));
wire output_2_710, output_2_0, output_1_710;
mixer gate_output_1_710(.a(output_2_710), .b(output_2_0), .y(output_1_710));
wire output_3_710, output_3_0, output_2_710;
mixer gate_output_2_710(.a(output_3_710), .b(output_3_0), .y(output_2_710));
wire output_1_711, output_1_1, output_0_711;
mixer gate_output_0_711(.a(output_1_711), .b(output_1_1), .y(output_0_711));
wire output_2_711, output_2_1, output_1_711;
mixer gate_output_1_711(.a(output_2_711), .b(output_2_1), .y(output_1_711));
wire output_3_711, output_3_1, output_2_711;
mixer gate_output_2_711(.a(output_3_711), .b(output_3_1), .y(output_2_711));
wire output_1_712, output_1_2, output_0_712;
mixer gate_output_0_712(.a(output_1_712), .b(output_1_2), .y(output_0_712));
wire output_2_712, output_2_2, output_1_712;
mixer gate_output_1_712(.a(output_2_712), .b(output_2_2), .y(output_1_712));
wire output_3_712, output_3_2, output_2_712;
mixer gate_output_2_712(.a(output_3_712), .b(output_3_2), .y(output_2_712));
wire output_1_713, output_1_0, output_0_713;
mixer gate_output_0_713(.a(output_1_713), .b(output_1_0), .y(output_0_713));
wire output_2_713, output_2_0, output_1_713;
mixer gate_output_1_713(.a(output_2_713), .b(output_2_0), .y(output_1_713));
wire output_3_713, output_3_0, output_2_713;
mixer gate_output_2_713(.a(output_3_713), .b(output_3_0), .y(output_2_713));
wire output_1_714, output_1_1, output_0_714;
mixer gate_output_0_714(.a(output_1_714), .b(output_1_1), .y(output_0_714));
wire output_2_714, output_2_1, output_1_714;
mixer gate_output_1_714(.a(output_2_714), .b(output_2_1), .y(output_1_714));
wire output_3_714, output_3_1, output_2_714;
mixer gate_output_2_714(.a(output_3_714), .b(output_3_1), .y(output_2_714));
wire output_1_715, output_1_2, output_0_715;
mixer gate_output_0_715(.a(output_1_715), .b(output_1_2), .y(output_0_715));
wire output_2_715, output_2_2, output_1_715;
mixer gate_output_1_715(.a(output_2_715), .b(output_2_2), .y(output_1_715));
wire output_3_715, output_3_2, output_2_715;
mixer gate_output_2_715(.a(output_3_715), .b(output_3_2), .y(output_2_715));
wire output_1_716, output_1_0, output_0_716;
mixer gate_output_0_716(.a(output_1_716), .b(output_1_0), .y(output_0_716));
wire output_2_716, output_2_0, output_1_716;
mixer gate_output_1_716(.a(output_2_716), .b(output_2_0), .y(output_1_716));
wire output_3_716, output_3_0, output_2_716;
mixer gate_output_2_716(.a(output_3_716), .b(output_3_0), .y(output_2_716));
wire output_1_717, output_1_1, output_0_717;
mixer gate_output_0_717(.a(output_1_717), .b(output_1_1), .y(output_0_717));
wire output_2_717, output_2_1, output_1_717;
mixer gate_output_1_717(.a(output_2_717), .b(output_2_1), .y(output_1_717));
wire output_3_717, output_3_1, output_2_717;
mixer gate_output_2_717(.a(output_3_717), .b(output_3_1), .y(output_2_717));
wire output_1_718, output_1_2, output_0_718;
mixer gate_output_0_718(.a(output_1_718), .b(output_1_2), .y(output_0_718));
wire output_2_718, output_2_2, output_1_718;
mixer gate_output_1_718(.a(output_2_718), .b(output_2_2), .y(output_1_718));
wire output_3_718, output_3_2, output_2_718;
mixer gate_output_2_718(.a(output_3_718), .b(output_3_2), .y(output_2_718));
wire output_1_719, output_1_0, output_0_719;
mixer gate_output_0_719(.a(output_1_719), .b(output_1_0), .y(output_0_719));
wire output_2_719, output_2_0, output_1_719;
mixer gate_output_1_719(.a(output_2_719), .b(output_2_0), .y(output_1_719));
wire output_3_719, output_3_0, output_2_719;
mixer gate_output_2_719(.a(output_3_719), .b(output_3_0), .y(output_2_719));
wire output_1_720, output_1_1, output_0_720;
mixer gate_output_0_720(.a(output_1_720), .b(output_1_1), .y(output_0_720));
wire output_2_720, output_2_1, output_1_720;
mixer gate_output_1_720(.a(output_2_720), .b(output_2_1), .y(output_1_720));
wire output_3_720, output_3_1, output_2_720;
mixer gate_output_2_720(.a(output_3_720), .b(output_3_1), .y(output_2_720));
wire output_1_721, output_1_2, output_0_721;
mixer gate_output_0_721(.a(output_1_721), .b(output_1_2), .y(output_0_721));
wire output_2_721, output_2_2, output_1_721;
mixer gate_output_1_721(.a(output_2_721), .b(output_2_2), .y(output_1_721));
wire output_3_721, output_3_2, output_2_721;
mixer gate_output_2_721(.a(output_3_721), .b(output_3_2), .y(output_2_721));
wire output_1_722, output_1_0, output_0_722;
mixer gate_output_0_722(.a(output_1_722), .b(output_1_0), .y(output_0_722));
wire output_2_722, output_2_0, output_1_722;
mixer gate_output_1_722(.a(output_2_722), .b(output_2_0), .y(output_1_722));
wire output_3_722, output_3_0, output_2_722;
mixer gate_output_2_722(.a(output_3_722), .b(output_3_0), .y(output_2_722));
wire output_1_723, output_1_1, output_0_723;
mixer gate_output_0_723(.a(output_1_723), .b(output_1_1), .y(output_0_723));
wire output_2_723, output_2_1, output_1_723;
mixer gate_output_1_723(.a(output_2_723), .b(output_2_1), .y(output_1_723));
wire output_3_723, output_3_1, output_2_723;
mixer gate_output_2_723(.a(output_3_723), .b(output_3_1), .y(output_2_723));
wire output_1_724, output_1_2, output_0_724;
mixer gate_output_0_724(.a(output_1_724), .b(output_1_2), .y(output_0_724));
wire output_2_724, output_2_2, output_1_724;
mixer gate_output_1_724(.a(output_2_724), .b(output_2_2), .y(output_1_724));
wire output_3_724, output_3_2, output_2_724;
mixer gate_output_2_724(.a(output_3_724), .b(output_3_2), .y(output_2_724));
wire output_1_725, output_1_0, output_0_725;
mixer gate_output_0_725(.a(output_1_725), .b(output_1_0), .y(output_0_725));
wire output_2_725, output_2_0, output_1_725;
mixer gate_output_1_725(.a(output_2_725), .b(output_2_0), .y(output_1_725));
wire output_3_725, output_3_0, output_2_725;
mixer gate_output_2_725(.a(output_3_725), .b(output_3_0), .y(output_2_725));
wire output_1_726, output_1_1, output_0_726;
mixer gate_output_0_726(.a(output_1_726), .b(output_1_1), .y(output_0_726));
wire output_2_726, output_2_1, output_1_726;
mixer gate_output_1_726(.a(output_2_726), .b(output_2_1), .y(output_1_726));
wire output_3_726, output_3_1, output_2_726;
mixer gate_output_2_726(.a(output_3_726), .b(output_3_1), .y(output_2_726));
wire output_1_727, output_1_2, output_0_727;
mixer gate_output_0_727(.a(output_1_727), .b(output_1_2), .y(output_0_727));
wire output_2_727, output_2_2, output_1_727;
mixer gate_output_1_727(.a(output_2_727), .b(output_2_2), .y(output_1_727));
wire output_3_727, output_3_2, output_2_727;
mixer gate_output_2_727(.a(output_3_727), .b(output_3_2), .y(output_2_727));
wire output_1_728, output_1_0, output_0_728;
mixer gate_output_0_728(.a(output_1_728), .b(output_1_0), .y(output_0_728));
wire output_2_728, output_2_0, output_1_728;
mixer gate_output_1_728(.a(output_2_728), .b(output_2_0), .y(output_1_728));
wire output_3_728, output_3_0, output_2_728;
mixer gate_output_2_728(.a(output_3_728), .b(output_3_0), .y(output_2_728));
wire output_1_729, output_1_1, output_0_729;
mixer gate_output_0_729(.a(output_1_729), .b(output_1_1), .y(output_0_729));
wire output_2_729, output_2_1, output_1_729;
mixer gate_output_1_729(.a(output_2_729), .b(output_2_1), .y(output_1_729));
wire output_3_729, output_3_1, output_2_729;
mixer gate_output_2_729(.a(output_3_729), .b(output_3_1), .y(output_2_729));
wire output_1_730, output_1_2, output_0_730;
mixer gate_output_0_730(.a(output_1_730), .b(output_1_2), .y(output_0_730));
wire output_2_730, output_2_2, output_1_730;
mixer gate_output_1_730(.a(output_2_730), .b(output_2_2), .y(output_1_730));
wire output_3_730, output_3_2, output_2_730;
mixer gate_output_2_730(.a(output_3_730), .b(output_3_2), .y(output_2_730));
wire output_1_731, output_1_0, output_0_731;
mixer gate_output_0_731(.a(output_1_731), .b(output_1_0), .y(output_0_731));
wire output_2_731, output_2_0, output_1_731;
mixer gate_output_1_731(.a(output_2_731), .b(output_2_0), .y(output_1_731));
wire output_3_731, output_3_0, output_2_731;
mixer gate_output_2_731(.a(output_3_731), .b(output_3_0), .y(output_2_731));
wire output_1_732, output_1_1, output_0_732;
mixer gate_output_0_732(.a(output_1_732), .b(output_1_1), .y(output_0_732));
wire output_2_732, output_2_1, output_1_732;
mixer gate_output_1_732(.a(output_2_732), .b(output_2_1), .y(output_1_732));
wire output_3_732, output_3_1, output_2_732;
mixer gate_output_2_732(.a(output_3_732), .b(output_3_1), .y(output_2_732));
wire output_1_733, output_1_2, output_0_733;
mixer gate_output_0_733(.a(output_1_733), .b(output_1_2), .y(output_0_733));
wire output_2_733, output_2_2, output_1_733;
mixer gate_output_1_733(.a(output_2_733), .b(output_2_2), .y(output_1_733));
wire output_3_733, output_3_2, output_2_733;
mixer gate_output_2_733(.a(output_3_733), .b(output_3_2), .y(output_2_733));
wire output_1_734, output_1_0, output_0_734;
mixer gate_output_0_734(.a(output_1_734), .b(output_1_0), .y(output_0_734));
wire output_2_734, output_2_0, output_1_734;
mixer gate_output_1_734(.a(output_2_734), .b(output_2_0), .y(output_1_734));
wire output_3_734, output_3_0, output_2_734;
mixer gate_output_2_734(.a(output_3_734), .b(output_3_0), .y(output_2_734));
wire output_1_735, output_1_1, output_0_735;
mixer gate_output_0_735(.a(output_1_735), .b(output_1_1), .y(output_0_735));
wire output_2_735, output_2_1, output_1_735;
mixer gate_output_1_735(.a(output_2_735), .b(output_2_1), .y(output_1_735));
wire output_3_735, output_3_1, output_2_735;
mixer gate_output_2_735(.a(output_3_735), .b(output_3_1), .y(output_2_735));
wire output_1_736, output_1_2, output_0_736;
mixer gate_output_0_736(.a(output_1_736), .b(output_1_2), .y(output_0_736));
wire output_2_736, output_2_2, output_1_736;
mixer gate_output_1_736(.a(output_2_736), .b(output_2_2), .y(output_1_736));
wire output_3_736, output_3_2, output_2_736;
mixer gate_output_2_736(.a(output_3_736), .b(output_3_2), .y(output_2_736));
wire output_1_737, output_1_0, output_0_737;
mixer gate_output_0_737(.a(output_1_737), .b(output_1_0), .y(output_0_737));
wire output_2_737, output_2_0, output_1_737;
mixer gate_output_1_737(.a(output_2_737), .b(output_2_0), .y(output_1_737));
wire output_3_737, output_3_0, output_2_737;
mixer gate_output_2_737(.a(output_3_737), .b(output_3_0), .y(output_2_737));
wire output_1_738, output_1_1, output_0_738;
mixer gate_output_0_738(.a(output_1_738), .b(output_1_1), .y(output_0_738));
wire output_2_738, output_2_1, output_1_738;
mixer gate_output_1_738(.a(output_2_738), .b(output_2_1), .y(output_1_738));
wire output_3_738, output_3_1, output_2_738;
mixer gate_output_2_738(.a(output_3_738), .b(output_3_1), .y(output_2_738));
wire output_1_739, output_1_2, output_0_739;
mixer gate_output_0_739(.a(output_1_739), .b(output_1_2), .y(output_0_739));
wire output_2_739, output_2_2, output_1_739;
mixer gate_output_1_739(.a(output_2_739), .b(output_2_2), .y(output_1_739));
wire output_3_739, output_3_2, output_2_739;
mixer gate_output_2_739(.a(output_3_739), .b(output_3_2), .y(output_2_739));
wire output_1_740, output_1_0, output_0_740;
mixer gate_output_0_740(.a(output_1_740), .b(output_1_0), .y(output_0_740));
wire output_2_740, output_2_0, output_1_740;
mixer gate_output_1_740(.a(output_2_740), .b(output_2_0), .y(output_1_740));
wire output_3_740, output_3_0, output_2_740;
mixer gate_output_2_740(.a(output_3_740), .b(output_3_0), .y(output_2_740));
wire output_1_741, output_1_1, output_0_741;
mixer gate_output_0_741(.a(output_1_741), .b(output_1_1), .y(output_0_741));
wire output_2_741, output_2_1, output_1_741;
mixer gate_output_1_741(.a(output_2_741), .b(output_2_1), .y(output_1_741));
wire output_3_741, output_3_1, output_2_741;
mixer gate_output_2_741(.a(output_3_741), .b(output_3_1), .y(output_2_741));
wire output_1_742, output_1_2, output_0_742;
mixer gate_output_0_742(.a(output_1_742), .b(output_1_2), .y(output_0_742));
wire output_2_742, output_2_2, output_1_742;
mixer gate_output_1_742(.a(output_2_742), .b(output_2_2), .y(output_1_742));
wire output_3_742, output_3_2, output_2_742;
mixer gate_output_2_742(.a(output_3_742), .b(output_3_2), .y(output_2_742));
wire output_1_743, output_1_0, output_0_743;
mixer gate_output_0_743(.a(output_1_743), .b(output_1_0), .y(output_0_743));
wire output_2_743, output_2_0, output_1_743;
mixer gate_output_1_743(.a(output_2_743), .b(output_2_0), .y(output_1_743));
wire output_3_743, output_3_0, output_2_743;
mixer gate_output_2_743(.a(output_3_743), .b(output_3_0), .y(output_2_743));
wire output_1_744, output_1_1, output_0_744;
mixer gate_output_0_744(.a(output_1_744), .b(output_1_1), .y(output_0_744));
wire output_2_744, output_2_1, output_1_744;
mixer gate_output_1_744(.a(output_2_744), .b(output_2_1), .y(output_1_744));
wire output_3_744, output_3_1, output_2_744;
mixer gate_output_2_744(.a(output_3_744), .b(output_3_1), .y(output_2_744));
wire output_1_745, output_1_2, output_0_745;
mixer gate_output_0_745(.a(output_1_745), .b(output_1_2), .y(output_0_745));
wire output_2_745, output_2_2, output_1_745;
mixer gate_output_1_745(.a(output_2_745), .b(output_2_2), .y(output_1_745));
wire output_3_745, output_3_2, output_2_745;
mixer gate_output_2_745(.a(output_3_745), .b(output_3_2), .y(output_2_745));
wire output_1_746, output_1_0, output_0_746;
mixer gate_output_0_746(.a(output_1_746), .b(output_1_0), .y(output_0_746));
wire output_2_746, output_2_0, output_1_746;
mixer gate_output_1_746(.a(output_2_746), .b(output_2_0), .y(output_1_746));
wire output_3_746, output_3_0, output_2_746;
mixer gate_output_2_746(.a(output_3_746), .b(output_3_0), .y(output_2_746));
wire output_1_747, output_1_1, output_0_747;
mixer gate_output_0_747(.a(output_1_747), .b(output_1_1), .y(output_0_747));
wire output_2_747, output_2_1, output_1_747;
mixer gate_output_1_747(.a(output_2_747), .b(output_2_1), .y(output_1_747));
wire output_3_747, output_3_1, output_2_747;
mixer gate_output_2_747(.a(output_3_747), .b(output_3_1), .y(output_2_747));
wire output_1_748, output_1_2, output_0_748;
mixer gate_output_0_748(.a(output_1_748), .b(output_1_2), .y(output_0_748));
wire output_2_748, output_2_2, output_1_748;
mixer gate_output_1_748(.a(output_2_748), .b(output_2_2), .y(output_1_748));
wire output_3_748, output_3_2, output_2_748;
mixer gate_output_2_748(.a(output_3_748), .b(output_3_2), .y(output_2_748));
wire output_1_749, output_1_0, output_0_749;
mixer gate_output_0_749(.a(output_1_749), .b(output_1_0), .y(output_0_749));
wire output_2_749, output_2_0, output_1_749;
mixer gate_output_1_749(.a(output_2_749), .b(output_2_0), .y(output_1_749));
wire output_3_749, output_3_0, output_2_749;
mixer gate_output_2_749(.a(output_3_749), .b(output_3_0), .y(output_2_749));
wire output_1_750, output_1_1, output_0_750;
mixer gate_output_0_750(.a(output_1_750), .b(output_1_1), .y(output_0_750));
wire output_2_750, output_2_1, output_1_750;
mixer gate_output_1_750(.a(output_2_750), .b(output_2_1), .y(output_1_750));
wire output_3_750, output_3_1, output_2_750;
mixer gate_output_2_750(.a(output_3_750), .b(output_3_1), .y(output_2_750));
wire output_1_751, output_1_2, output_0_751;
mixer gate_output_0_751(.a(output_1_751), .b(output_1_2), .y(output_0_751));
wire output_2_751, output_2_2, output_1_751;
mixer gate_output_1_751(.a(output_2_751), .b(output_2_2), .y(output_1_751));
wire output_3_751, output_3_2, output_2_751;
mixer gate_output_2_751(.a(output_3_751), .b(output_3_2), .y(output_2_751));
wire output_1_752, output_1_0, output_0_752;
mixer gate_output_0_752(.a(output_1_752), .b(output_1_0), .y(output_0_752));
wire output_2_752, output_2_0, output_1_752;
mixer gate_output_1_752(.a(output_2_752), .b(output_2_0), .y(output_1_752));
wire output_3_752, output_3_0, output_2_752;
mixer gate_output_2_752(.a(output_3_752), .b(output_3_0), .y(output_2_752));
wire output_1_753, output_1_1, output_0_753;
mixer gate_output_0_753(.a(output_1_753), .b(output_1_1), .y(output_0_753));
wire output_2_753, output_2_1, output_1_753;
mixer gate_output_1_753(.a(output_2_753), .b(output_2_1), .y(output_1_753));
wire output_3_753, output_3_1, output_2_753;
mixer gate_output_2_753(.a(output_3_753), .b(output_3_1), .y(output_2_753));
wire output_1_754, output_1_2, output_0_754;
mixer gate_output_0_754(.a(output_1_754), .b(output_1_2), .y(output_0_754));
wire output_2_754, output_2_2, output_1_754;
mixer gate_output_1_754(.a(output_2_754), .b(output_2_2), .y(output_1_754));
wire output_3_754, output_3_2, output_2_754;
mixer gate_output_2_754(.a(output_3_754), .b(output_3_2), .y(output_2_754));
wire output_1_755, output_1_0, output_0_755;
mixer gate_output_0_755(.a(output_1_755), .b(output_1_0), .y(output_0_755));
wire output_2_755, output_2_0, output_1_755;
mixer gate_output_1_755(.a(output_2_755), .b(output_2_0), .y(output_1_755));
wire output_3_755, output_3_0, output_2_755;
mixer gate_output_2_755(.a(output_3_755), .b(output_3_0), .y(output_2_755));
wire output_1_756, output_1_1, output_0_756;
mixer gate_output_0_756(.a(output_1_756), .b(output_1_1), .y(output_0_756));
wire output_2_756, output_2_1, output_1_756;
mixer gate_output_1_756(.a(output_2_756), .b(output_2_1), .y(output_1_756));
wire output_3_756, output_3_1, output_2_756;
mixer gate_output_2_756(.a(output_3_756), .b(output_3_1), .y(output_2_756));
wire output_1_757, output_1_2, output_0_757;
mixer gate_output_0_757(.a(output_1_757), .b(output_1_2), .y(output_0_757));
wire output_2_757, output_2_2, output_1_757;
mixer gate_output_1_757(.a(output_2_757), .b(output_2_2), .y(output_1_757));
wire output_3_757, output_3_2, output_2_757;
mixer gate_output_2_757(.a(output_3_757), .b(output_3_2), .y(output_2_757));
wire output_1_758, output_1_0, output_0_758;
mixer gate_output_0_758(.a(output_1_758), .b(output_1_0), .y(output_0_758));
wire output_2_758, output_2_0, output_1_758;
mixer gate_output_1_758(.a(output_2_758), .b(output_2_0), .y(output_1_758));
wire output_3_758, output_3_0, output_2_758;
mixer gate_output_2_758(.a(output_3_758), .b(output_3_0), .y(output_2_758));
wire output_1_759, output_1_1, output_0_759;
mixer gate_output_0_759(.a(output_1_759), .b(output_1_1), .y(output_0_759));
wire output_2_759, output_2_1, output_1_759;
mixer gate_output_1_759(.a(output_2_759), .b(output_2_1), .y(output_1_759));
wire output_3_759, output_3_1, output_2_759;
mixer gate_output_2_759(.a(output_3_759), .b(output_3_1), .y(output_2_759));
wire output_1_760, output_1_2, output_0_760;
mixer gate_output_0_760(.a(output_1_760), .b(output_1_2), .y(output_0_760));
wire output_2_760, output_2_2, output_1_760;
mixer gate_output_1_760(.a(output_2_760), .b(output_2_2), .y(output_1_760));
wire output_3_760, output_3_2, output_2_760;
mixer gate_output_2_760(.a(output_3_760), .b(output_3_2), .y(output_2_760));
wire output_1_761, output_1_0, output_0_761;
mixer gate_output_0_761(.a(output_1_761), .b(output_1_0), .y(output_0_761));
wire output_2_761, output_2_0, output_1_761;
mixer gate_output_1_761(.a(output_2_761), .b(output_2_0), .y(output_1_761));
wire output_3_761, output_3_0, output_2_761;
mixer gate_output_2_761(.a(output_3_761), .b(output_3_0), .y(output_2_761));
wire output_1_762, output_1_1, output_0_762;
mixer gate_output_0_762(.a(output_1_762), .b(output_1_1), .y(output_0_762));
wire output_2_762, output_2_1, output_1_762;
mixer gate_output_1_762(.a(output_2_762), .b(output_2_1), .y(output_1_762));
wire output_3_762, output_3_1, output_2_762;
mixer gate_output_2_762(.a(output_3_762), .b(output_3_1), .y(output_2_762));
wire output_1_763, output_1_2, output_0_763;
mixer gate_output_0_763(.a(output_1_763), .b(output_1_2), .y(output_0_763));
wire output_2_763, output_2_2, output_1_763;
mixer gate_output_1_763(.a(output_2_763), .b(output_2_2), .y(output_1_763));
wire output_3_763, output_3_2, output_2_763;
mixer gate_output_2_763(.a(output_3_763), .b(output_3_2), .y(output_2_763));
wire output_1_764, output_1_0, output_0_764;
mixer gate_output_0_764(.a(output_1_764), .b(output_1_0), .y(output_0_764));
wire output_2_764, output_2_0, output_1_764;
mixer gate_output_1_764(.a(output_2_764), .b(output_2_0), .y(output_1_764));
wire output_3_764, output_3_0, output_2_764;
mixer gate_output_2_764(.a(output_3_764), .b(output_3_0), .y(output_2_764));
wire output_1_765, output_1_1, output_0_765;
mixer gate_output_0_765(.a(output_1_765), .b(output_1_1), .y(output_0_765));
wire output_2_765, output_2_1, output_1_765;
mixer gate_output_1_765(.a(output_2_765), .b(output_2_1), .y(output_1_765));
wire output_3_765, output_3_1, output_2_765;
mixer gate_output_2_765(.a(output_3_765), .b(output_3_1), .y(output_2_765));
wire output_1_766, output_1_2, output_0_766;
mixer gate_output_0_766(.a(output_1_766), .b(output_1_2), .y(output_0_766));
wire output_2_766, output_2_2, output_1_766;
mixer gate_output_1_766(.a(output_2_766), .b(output_2_2), .y(output_1_766));
wire output_3_766, output_3_2, output_2_766;
mixer gate_output_2_766(.a(output_3_766), .b(output_3_2), .y(output_2_766));
wire output_1_767, output_1_0, output_0_767;
mixer gate_output_0_767(.a(output_1_767), .b(output_1_0), .y(output_0_767));
wire output_2_767, output_2_0, output_1_767;
mixer gate_output_1_767(.a(output_2_767), .b(output_2_0), .y(output_1_767));
wire output_3_767, output_3_0, output_2_767;
mixer gate_output_2_767(.a(output_3_767), .b(output_3_0), .y(output_2_767));
wire output_1_768, output_1_1, output_0_768;
mixer gate_output_0_768(.a(output_1_768), .b(output_1_1), .y(output_0_768));
wire output_2_768, output_2_1, output_1_768;
mixer gate_output_1_768(.a(output_2_768), .b(output_2_1), .y(output_1_768));
wire output_3_768, output_3_1, output_2_768;
mixer gate_output_2_768(.a(output_3_768), .b(output_3_1), .y(output_2_768));
wire output_1_769, output_1_2, output_0_769;
mixer gate_output_0_769(.a(output_1_769), .b(output_1_2), .y(output_0_769));
wire output_2_769, output_2_2, output_1_769;
mixer gate_output_1_769(.a(output_2_769), .b(output_2_2), .y(output_1_769));
wire output_3_769, output_3_2, output_2_769;
mixer gate_output_2_769(.a(output_3_769), .b(output_3_2), .y(output_2_769));
wire output_1_770, output_1_0, output_0_770;
mixer gate_output_0_770(.a(output_1_770), .b(output_1_0), .y(output_0_770));
wire output_2_770, output_2_0, output_1_770;
mixer gate_output_1_770(.a(output_2_770), .b(output_2_0), .y(output_1_770));
wire output_3_770, output_3_0, output_2_770;
mixer gate_output_2_770(.a(output_3_770), .b(output_3_0), .y(output_2_770));
wire output_1_771, output_1_1, output_0_771;
mixer gate_output_0_771(.a(output_1_771), .b(output_1_1), .y(output_0_771));
wire output_2_771, output_2_1, output_1_771;
mixer gate_output_1_771(.a(output_2_771), .b(output_2_1), .y(output_1_771));
wire output_3_771, output_3_1, output_2_771;
mixer gate_output_2_771(.a(output_3_771), .b(output_3_1), .y(output_2_771));
wire output_1_772, output_1_2, output_0_772;
mixer gate_output_0_772(.a(output_1_772), .b(output_1_2), .y(output_0_772));
wire output_2_772, output_2_2, output_1_772;
mixer gate_output_1_772(.a(output_2_772), .b(output_2_2), .y(output_1_772));
wire output_3_772, output_3_2, output_2_772;
mixer gate_output_2_772(.a(output_3_772), .b(output_3_2), .y(output_2_772));
wire output_1_773, output_1_0, output_0_773;
mixer gate_output_0_773(.a(output_1_773), .b(output_1_0), .y(output_0_773));
wire output_2_773, output_2_0, output_1_773;
mixer gate_output_1_773(.a(output_2_773), .b(output_2_0), .y(output_1_773));
wire output_3_773, output_3_0, output_2_773;
mixer gate_output_2_773(.a(output_3_773), .b(output_3_0), .y(output_2_773));
wire output_1_774, output_1_1, output_0_774;
mixer gate_output_0_774(.a(output_1_774), .b(output_1_1), .y(output_0_774));
wire output_2_774, output_2_1, output_1_774;
mixer gate_output_1_774(.a(output_2_774), .b(output_2_1), .y(output_1_774));
wire output_3_774, output_3_1, output_2_774;
mixer gate_output_2_774(.a(output_3_774), .b(output_3_1), .y(output_2_774));
wire output_1_775, output_1_2, output_0_775;
mixer gate_output_0_775(.a(output_1_775), .b(output_1_2), .y(output_0_775));
wire output_2_775, output_2_2, output_1_775;
mixer gate_output_1_775(.a(output_2_775), .b(output_2_2), .y(output_1_775));
wire output_3_775, output_3_2, output_2_775;
mixer gate_output_2_775(.a(output_3_775), .b(output_3_2), .y(output_2_775));
wire output_1_776, output_1_0, output_0_776;
mixer gate_output_0_776(.a(output_1_776), .b(output_1_0), .y(output_0_776));
wire output_2_776, output_2_0, output_1_776;
mixer gate_output_1_776(.a(output_2_776), .b(output_2_0), .y(output_1_776));
wire output_3_776, output_3_0, output_2_776;
mixer gate_output_2_776(.a(output_3_776), .b(output_3_0), .y(output_2_776));
wire output_1_777, output_1_1, output_0_777;
mixer gate_output_0_777(.a(output_1_777), .b(output_1_1), .y(output_0_777));
wire output_2_777, output_2_1, output_1_777;
mixer gate_output_1_777(.a(output_2_777), .b(output_2_1), .y(output_1_777));
wire output_3_777, output_3_1, output_2_777;
mixer gate_output_2_777(.a(output_3_777), .b(output_3_1), .y(output_2_777));
wire output_1_778, output_1_2, output_0_778;
mixer gate_output_0_778(.a(output_1_778), .b(output_1_2), .y(output_0_778));
wire output_2_778, output_2_2, output_1_778;
mixer gate_output_1_778(.a(output_2_778), .b(output_2_2), .y(output_1_778));
wire output_3_778, output_3_2, output_2_778;
mixer gate_output_2_778(.a(output_3_778), .b(output_3_2), .y(output_2_778));
wire output_1_779, output_1_0, output_0_779;
mixer gate_output_0_779(.a(output_1_779), .b(output_1_0), .y(output_0_779));
wire output_2_779, output_2_0, output_1_779;
mixer gate_output_1_779(.a(output_2_779), .b(output_2_0), .y(output_1_779));
wire output_3_779, output_3_0, output_2_779;
mixer gate_output_2_779(.a(output_3_779), .b(output_3_0), .y(output_2_779));
wire output_1_780, output_1_1, output_0_780;
mixer gate_output_0_780(.a(output_1_780), .b(output_1_1), .y(output_0_780));
wire output_2_780, output_2_1, output_1_780;
mixer gate_output_1_780(.a(output_2_780), .b(output_2_1), .y(output_1_780));
wire output_3_780, output_3_1, output_2_780;
mixer gate_output_2_780(.a(output_3_780), .b(output_3_1), .y(output_2_780));
wire output_1_781, output_1_2, output_0_781;
mixer gate_output_0_781(.a(output_1_781), .b(output_1_2), .y(output_0_781));
wire output_2_781, output_2_2, output_1_781;
mixer gate_output_1_781(.a(output_2_781), .b(output_2_2), .y(output_1_781));
wire output_3_781, output_3_2, output_2_781;
mixer gate_output_2_781(.a(output_3_781), .b(output_3_2), .y(output_2_781));
wire output_1_782, output_1_0, output_0_782;
mixer gate_output_0_782(.a(output_1_782), .b(output_1_0), .y(output_0_782));
wire output_2_782, output_2_0, output_1_782;
mixer gate_output_1_782(.a(output_2_782), .b(output_2_0), .y(output_1_782));
wire output_3_782, output_3_0, output_2_782;
mixer gate_output_2_782(.a(output_3_782), .b(output_3_0), .y(output_2_782));
wire output_1_783, output_1_1, output_0_783;
mixer gate_output_0_783(.a(output_1_783), .b(output_1_1), .y(output_0_783));
wire output_2_783, output_2_1, output_1_783;
mixer gate_output_1_783(.a(output_2_783), .b(output_2_1), .y(output_1_783));
wire output_3_783, output_3_1, output_2_783;
mixer gate_output_2_783(.a(output_3_783), .b(output_3_1), .y(output_2_783));
wire output_1_784, output_1_2, output_0_784;
mixer gate_output_0_784(.a(output_1_784), .b(output_1_2), .y(output_0_784));
wire output_2_784, output_2_2, output_1_784;
mixer gate_output_1_784(.a(output_2_784), .b(output_2_2), .y(output_1_784));
wire output_3_784, output_3_2, output_2_784;
mixer gate_output_2_784(.a(output_3_784), .b(output_3_2), .y(output_2_784));
wire output_1_785, output_1_0, output_0_785;
mixer gate_output_0_785(.a(output_1_785), .b(output_1_0), .y(output_0_785));
wire output_2_785, output_2_0, output_1_785;
mixer gate_output_1_785(.a(output_2_785), .b(output_2_0), .y(output_1_785));
wire output_3_785, output_3_0, output_2_785;
mixer gate_output_2_785(.a(output_3_785), .b(output_3_0), .y(output_2_785));
wire output_1_786, output_1_1, output_0_786;
mixer gate_output_0_786(.a(output_1_786), .b(output_1_1), .y(output_0_786));
wire output_2_786, output_2_1, output_1_786;
mixer gate_output_1_786(.a(output_2_786), .b(output_2_1), .y(output_1_786));
wire output_3_786, output_3_1, output_2_786;
mixer gate_output_2_786(.a(output_3_786), .b(output_3_1), .y(output_2_786));
wire output_1_787, output_1_2, output_0_787;
mixer gate_output_0_787(.a(output_1_787), .b(output_1_2), .y(output_0_787));
wire output_2_787, output_2_2, output_1_787;
mixer gate_output_1_787(.a(output_2_787), .b(output_2_2), .y(output_1_787));
wire output_3_787, output_3_2, output_2_787;
mixer gate_output_2_787(.a(output_3_787), .b(output_3_2), .y(output_2_787));
wire output_1_788, output_1_0, output_0_788;
mixer gate_output_0_788(.a(output_1_788), .b(output_1_0), .y(output_0_788));
wire output_2_788, output_2_0, output_1_788;
mixer gate_output_1_788(.a(output_2_788), .b(output_2_0), .y(output_1_788));
wire output_3_788, output_3_0, output_2_788;
mixer gate_output_2_788(.a(output_3_788), .b(output_3_0), .y(output_2_788));
wire output_1_789, output_1_1, output_0_789;
mixer gate_output_0_789(.a(output_1_789), .b(output_1_1), .y(output_0_789));
wire output_2_789, output_2_1, output_1_789;
mixer gate_output_1_789(.a(output_2_789), .b(output_2_1), .y(output_1_789));
wire output_3_789, output_3_1, output_2_789;
mixer gate_output_2_789(.a(output_3_789), .b(output_3_1), .y(output_2_789));
wire output_1_790, output_1_2, output_0_790;
mixer gate_output_0_790(.a(output_1_790), .b(output_1_2), .y(output_0_790));
wire output_2_790, output_2_2, output_1_790;
mixer gate_output_1_790(.a(output_2_790), .b(output_2_2), .y(output_1_790));
wire output_3_790, output_3_2, output_2_790;
mixer gate_output_2_790(.a(output_3_790), .b(output_3_2), .y(output_2_790));
wire output_1_791, output_1_0, output_0_791;
mixer gate_output_0_791(.a(output_1_791), .b(output_1_0), .y(output_0_791));
wire output_2_791, output_2_0, output_1_791;
mixer gate_output_1_791(.a(output_2_791), .b(output_2_0), .y(output_1_791));
wire output_3_791, output_3_0, output_2_791;
mixer gate_output_2_791(.a(output_3_791), .b(output_3_0), .y(output_2_791));
wire output_1_792, output_1_1, output_0_792;
mixer gate_output_0_792(.a(output_1_792), .b(output_1_1), .y(output_0_792));
wire output_2_792, output_2_1, output_1_792;
mixer gate_output_1_792(.a(output_2_792), .b(output_2_1), .y(output_1_792));
wire output_3_792, output_3_1, output_2_792;
mixer gate_output_2_792(.a(output_3_792), .b(output_3_1), .y(output_2_792));
wire output_1_793, output_1_2, output_0_793;
mixer gate_output_0_793(.a(output_1_793), .b(output_1_2), .y(output_0_793));
wire output_2_793, output_2_2, output_1_793;
mixer gate_output_1_793(.a(output_2_793), .b(output_2_2), .y(output_1_793));
wire output_3_793, output_3_2, output_2_793;
mixer gate_output_2_793(.a(output_3_793), .b(output_3_2), .y(output_2_793));
wire output_1_794, output_1_0, output_0_794;
mixer gate_output_0_794(.a(output_1_794), .b(output_1_0), .y(output_0_794));
wire output_2_794, output_2_0, output_1_794;
mixer gate_output_1_794(.a(output_2_794), .b(output_2_0), .y(output_1_794));
wire output_3_794, output_3_0, output_2_794;
mixer gate_output_2_794(.a(output_3_794), .b(output_3_0), .y(output_2_794));
wire output_1_795, output_1_1, output_0_795;
mixer gate_output_0_795(.a(output_1_795), .b(output_1_1), .y(output_0_795));
wire output_2_795, output_2_1, output_1_795;
mixer gate_output_1_795(.a(output_2_795), .b(output_2_1), .y(output_1_795));
wire output_3_795, output_3_1, output_2_795;
mixer gate_output_2_795(.a(output_3_795), .b(output_3_1), .y(output_2_795));
wire output_1_796, output_1_2, output_0_796;
mixer gate_output_0_796(.a(output_1_796), .b(output_1_2), .y(output_0_796));
wire output_2_796, output_2_2, output_1_796;
mixer gate_output_1_796(.a(output_2_796), .b(output_2_2), .y(output_1_796));
wire output_3_796, output_3_2, output_2_796;
mixer gate_output_2_796(.a(output_3_796), .b(output_3_2), .y(output_2_796));
wire output_1_797, output_1_0, output_0_797;
mixer gate_output_0_797(.a(output_1_797), .b(output_1_0), .y(output_0_797));
wire output_2_797, output_2_0, output_1_797;
mixer gate_output_1_797(.a(output_2_797), .b(output_2_0), .y(output_1_797));
wire output_3_797, output_3_0, output_2_797;
mixer gate_output_2_797(.a(output_3_797), .b(output_3_0), .y(output_2_797));
wire output_1_798, output_1_1, output_0_798;
mixer gate_output_0_798(.a(output_1_798), .b(output_1_1), .y(output_0_798));
wire output_2_798, output_2_1, output_1_798;
mixer gate_output_1_798(.a(output_2_798), .b(output_2_1), .y(output_1_798));
wire output_3_798, output_3_1, output_2_798;
mixer gate_output_2_798(.a(output_3_798), .b(output_3_1), .y(output_2_798));
wire output_1_799, output_1_2, output_0_799;
mixer gate_output_0_799(.a(output_1_799), .b(output_1_2), .y(output_0_799));
wire output_2_799, output_2_2, output_1_799;
mixer gate_output_1_799(.a(output_2_799), .b(output_2_2), .y(output_1_799));
wire output_3_799, output_3_2, output_2_799;
mixer gate_output_2_799(.a(output_3_799), .b(output_3_2), .y(output_2_799));
wire output_1_800, output_1_0, output_0_800;
mixer gate_output_0_800(.a(output_1_800), .b(output_1_0), .y(output_0_800));
wire output_2_800, output_2_0, output_1_800;
mixer gate_output_1_800(.a(output_2_800), .b(output_2_0), .y(output_1_800));
wire output_3_800, output_3_0, output_2_800;
mixer gate_output_2_800(.a(output_3_800), .b(output_3_0), .y(output_2_800));
wire output_1_801, output_1_1, output_0_801;
mixer gate_output_0_801(.a(output_1_801), .b(output_1_1), .y(output_0_801));
wire output_2_801, output_2_1, output_1_801;
mixer gate_output_1_801(.a(output_2_801), .b(output_2_1), .y(output_1_801));
wire output_3_801, output_3_1, output_2_801;
mixer gate_output_2_801(.a(output_3_801), .b(output_3_1), .y(output_2_801));
wire output_1_802, output_1_2, output_0_802;
mixer gate_output_0_802(.a(output_1_802), .b(output_1_2), .y(output_0_802));
wire output_2_802, output_2_2, output_1_802;
mixer gate_output_1_802(.a(output_2_802), .b(output_2_2), .y(output_1_802));
wire output_3_802, output_3_2, output_2_802;
mixer gate_output_2_802(.a(output_3_802), .b(output_3_2), .y(output_2_802));
wire output_1_803, output_1_0, output_0_803;
mixer gate_output_0_803(.a(output_1_803), .b(output_1_0), .y(output_0_803));
wire output_2_803, output_2_0, output_1_803;
mixer gate_output_1_803(.a(output_2_803), .b(output_2_0), .y(output_1_803));
wire output_3_803, output_3_0, output_2_803;
mixer gate_output_2_803(.a(output_3_803), .b(output_3_0), .y(output_2_803));
wire output_1_804, output_1_1, output_0_804;
mixer gate_output_0_804(.a(output_1_804), .b(output_1_1), .y(output_0_804));
wire output_2_804, output_2_1, output_1_804;
mixer gate_output_1_804(.a(output_2_804), .b(output_2_1), .y(output_1_804));
wire output_3_804, output_3_1, output_2_804;
mixer gate_output_2_804(.a(output_3_804), .b(output_3_1), .y(output_2_804));
wire output_1_805, output_1_2, output_0_805;
mixer gate_output_0_805(.a(output_1_805), .b(output_1_2), .y(output_0_805));
wire output_2_805, output_2_2, output_1_805;
mixer gate_output_1_805(.a(output_2_805), .b(output_2_2), .y(output_1_805));
wire output_3_805, output_3_2, output_2_805;
mixer gate_output_2_805(.a(output_3_805), .b(output_3_2), .y(output_2_805));
wire output_1_806, output_1_0, output_0_806;
mixer gate_output_0_806(.a(output_1_806), .b(output_1_0), .y(output_0_806));
wire output_2_806, output_2_0, output_1_806;
mixer gate_output_1_806(.a(output_2_806), .b(output_2_0), .y(output_1_806));
wire output_3_806, output_3_0, output_2_806;
mixer gate_output_2_806(.a(output_3_806), .b(output_3_0), .y(output_2_806));
wire output_1_807, output_1_1, output_0_807;
mixer gate_output_0_807(.a(output_1_807), .b(output_1_1), .y(output_0_807));
wire output_2_807, output_2_1, output_1_807;
mixer gate_output_1_807(.a(output_2_807), .b(output_2_1), .y(output_1_807));
wire output_3_807, output_3_1, output_2_807;
mixer gate_output_2_807(.a(output_3_807), .b(output_3_1), .y(output_2_807));
wire output_1_808, output_1_2, output_0_808;
mixer gate_output_0_808(.a(output_1_808), .b(output_1_2), .y(output_0_808));
wire output_2_808, output_2_2, output_1_808;
mixer gate_output_1_808(.a(output_2_808), .b(output_2_2), .y(output_1_808));
wire output_3_808, output_3_2, output_2_808;
mixer gate_output_2_808(.a(output_3_808), .b(output_3_2), .y(output_2_808));
wire output_1_809, output_1_0, output_0_809;
mixer gate_output_0_809(.a(output_1_809), .b(output_1_0), .y(output_0_809));
wire output_2_809, output_2_0, output_1_809;
mixer gate_output_1_809(.a(output_2_809), .b(output_2_0), .y(output_1_809));
wire output_3_809, output_3_0, output_2_809;
mixer gate_output_2_809(.a(output_3_809), .b(output_3_0), .y(output_2_809));
wire output_1_810, output_1_1, output_0_810;
mixer gate_output_0_810(.a(output_1_810), .b(output_1_1), .y(output_0_810));
wire output_2_810, output_2_1, output_1_810;
mixer gate_output_1_810(.a(output_2_810), .b(output_2_1), .y(output_1_810));
wire output_3_810, output_3_1, output_2_810;
mixer gate_output_2_810(.a(output_3_810), .b(output_3_1), .y(output_2_810));
wire output_1_811, output_1_2, output_0_811;
mixer gate_output_0_811(.a(output_1_811), .b(output_1_2), .y(output_0_811));
wire output_2_811, output_2_2, output_1_811;
mixer gate_output_1_811(.a(output_2_811), .b(output_2_2), .y(output_1_811));
wire output_3_811, output_3_2, output_2_811;
mixer gate_output_2_811(.a(output_3_811), .b(output_3_2), .y(output_2_811));
wire output_1_812, output_1_0, output_0_812;
mixer gate_output_0_812(.a(output_1_812), .b(output_1_0), .y(output_0_812));
wire output_2_812, output_2_0, output_1_812;
mixer gate_output_1_812(.a(output_2_812), .b(output_2_0), .y(output_1_812));
wire output_3_812, output_3_0, output_2_812;
mixer gate_output_2_812(.a(output_3_812), .b(output_3_0), .y(output_2_812));
wire output_1_813, output_1_1, output_0_813;
mixer gate_output_0_813(.a(output_1_813), .b(output_1_1), .y(output_0_813));
wire output_2_813, output_2_1, output_1_813;
mixer gate_output_1_813(.a(output_2_813), .b(output_2_1), .y(output_1_813));
wire output_3_813, output_3_1, output_2_813;
mixer gate_output_2_813(.a(output_3_813), .b(output_3_1), .y(output_2_813));
wire output_1_814, output_1_2, output_0_814;
mixer gate_output_0_814(.a(output_1_814), .b(output_1_2), .y(output_0_814));
wire output_2_814, output_2_2, output_1_814;
mixer gate_output_1_814(.a(output_2_814), .b(output_2_2), .y(output_1_814));
wire output_3_814, output_3_2, output_2_814;
mixer gate_output_2_814(.a(output_3_814), .b(output_3_2), .y(output_2_814));
wire output_1_815, output_1_0, output_0_815;
mixer gate_output_0_815(.a(output_1_815), .b(output_1_0), .y(output_0_815));
wire output_2_815, output_2_0, output_1_815;
mixer gate_output_1_815(.a(output_2_815), .b(output_2_0), .y(output_1_815));
wire output_3_815, output_3_0, output_2_815;
mixer gate_output_2_815(.a(output_3_815), .b(output_3_0), .y(output_2_815));
wire output_1_816, output_1_1, output_0_816;
mixer gate_output_0_816(.a(output_1_816), .b(output_1_1), .y(output_0_816));
wire output_2_816, output_2_1, output_1_816;
mixer gate_output_1_816(.a(output_2_816), .b(output_2_1), .y(output_1_816));
wire output_3_816, output_3_1, output_2_816;
mixer gate_output_2_816(.a(output_3_816), .b(output_3_1), .y(output_2_816));
wire output_1_817, output_1_2, output_0_817;
mixer gate_output_0_817(.a(output_1_817), .b(output_1_2), .y(output_0_817));
wire output_2_817, output_2_2, output_1_817;
mixer gate_output_1_817(.a(output_2_817), .b(output_2_2), .y(output_1_817));
wire output_3_817, output_3_2, output_2_817;
mixer gate_output_2_817(.a(output_3_817), .b(output_3_2), .y(output_2_817));
wire output_1_818, output_1_0, output_0_818;
mixer gate_output_0_818(.a(output_1_818), .b(output_1_0), .y(output_0_818));
wire output_2_818, output_2_0, output_1_818;
mixer gate_output_1_818(.a(output_2_818), .b(output_2_0), .y(output_1_818));
wire output_3_818, output_3_0, output_2_818;
mixer gate_output_2_818(.a(output_3_818), .b(output_3_0), .y(output_2_818));
wire output_1_819, output_1_1, output_0_819;
mixer gate_output_0_819(.a(output_1_819), .b(output_1_1), .y(output_0_819));
wire output_2_819, output_2_1, output_1_819;
mixer gate_output_1_819(.a(output_2_819), .b(output_2_1), .y(output_1_819));
wire output_3_819, output_3_1, output_2_819;
mixer gate_output_2_819(.a(output_3_819), .b(output_3_1), .y(output_2_819));
wire output_1_820, output_1_2, output_0_820;
mixer gate_output_0_820(.a(output_1_820), .b(output_1_2), .y(output_0_820));
wire output_2_820, output_2_2, output_1_820;
mixer gate_output_1_820(.a(output_2_820), .b(output_2_2), .y(output_1_820));
wire output_3_820, output_3_2, output_2_820;
mixer gate_output_2_820(.a(output_3_820), .b(output_3_2), .y(output_2_820));
wire output_1_821, output_1_0, output_0_821;
mixer gate_output_0_821(.a(output_1_821), .b(output_1_0), .y(output_0_821));
wire output_2_821, output_2_0, output_1_821;
mixer gate_output_1_821(.a(output_2_821), .b(output_2_0), .y(output_1_821));
wire output_3_821, output_3_0, output_2_821;
mixer gate_output_2_821(.a(output_3_821), .b(output_3_0), .y(output_2_821));
wire output_1_822, output_1_1, output_0_822;
mixer gate_output_0_822(.a(output_1_822), .b(output_1_1), .y(output_0_822));
wire output_2_822, output_2_1, output_1_822;
mixer gate_output_1_822(.a(output_2_822), .b(output_2_1), .y(output_1_822));
wire output_3_822, output_3_1, output_2_822;
mixer gate_output_2_822(.a(output_3_822), .b(output_3_1), .y(output_2_822));
wire output_1_823, output_1_2, output_0_823;
mixer gate_output_0_823(.a(output_1_823), .b(output_1_2), .y(output_0_823));
wire output_2_823, output_2_2, output_1_823;
mixer gate_output_1_823(.a(output_2_823), .b(output_2_2), .y(output_1_823));
wire output_3_823, output_3_2, output_2_823;
mixer gate_output_2_823(.a(output_3_823), .b(output_3_2), .y(output_2_823));
wire output_1_824, output_1_0, output_0_824;
mixer gate_output_0_824(.a(output_1_824), .b(output_1_0), .y(output_0_824));
wire output_2_824, output_2_0, output_1_824;
mixer gate_output_1_824(.a(output_2_824), .b(output_2_0), .y(output_1_824));
wire output_3_824, output_3_0, output_2_824;
mixer gate_output_2_824(.a(output_3_824), .b(output_3_0), .y(output_2_824));
wire output_1_825, output_1_1, output_0_825;
mixer gate_output_0_825(.a(output_1_825), .b(output_1_1), .y(output_0_825));
wire output_2_825, output_2_1, output_1_825;
mixer gate_output_1_825(.a(output_2_825), .b(output_2_1), .y(output_1_825));
wire output_3_825, output_3_1, output_2_825;
mixer gate_output_2_825(.a(output_3_825), .b(output_3_1), .y(output_2_825));
wire output_1_826, output_1_2, output_0_826;
mixer gate_output_0_826(.a(output_1_826), .b(output_1_2), .y(output_0_826));
wire output_2_826, output_2_2, output_1_826;
mixer gate_output_1_826(.a(output_2_826), .b(output_2_2), .y(output_1_826));
wire output_3_826, output_3_2, output_2_826;
mixer gate_output_2_826(.a(output_3_826), .b(output_3_2), .y(output_2_826));
wire output_1_827, output_1_0, output_0_827;
mixer gate_output_0_827(.a(output_1_827), .b(output_1_0), .y(output_0_827));
wire output_2_827, output_2_0, output_1_827;
mixer gate_output_1_827(.a(output_2_827), .b(output_2_0), .y(output_1_827));
wire output_3_827, output_3_0, output_2_827;
mixer gate_output_2_827(.a(output_3_827), .b(output_3_0), .y(output_2_827));
wire output_1_828, output_1_1, output_0_828;
mixer gate_output_0_828(.a(output_1_828), .b(output_1_1), .y(output_0_828));
wire output_2_828, output_2_1, output_1_828;
mixer gate_output_1_828(.a(output_2_828), .b(output_2_1), .y(output_1_828));
wire output_3_828, output_3_1, output_2_828;
mixer gate_output_2_828(.a(output_3_828), .b(output_3_1), .y(output_2_828));
wire output_1_829, output_1_2, output_0_829;
mixer gate_output_0_829(.a(output_1_829), .b(output_1_2), .y(output_0_829));
wire output_2_829, output_2_2, output_1_829;
mixer gate_output_1_829(.a(output_2_829), .b(output_2_2), .y(output_1_829));
wire output_3_829, output_3_2, output_2_829;
mixer gate_output_2_829(.a(output_3_829), .b(output_3_2), .y(output_2_829));
wire output_1_830, output_1_0, output_0_830;
mixer gate_output_0_830(.a(output_1_830), .b(output_1_0), .y(output_0_830));
wire output_2_830, output_2_0, output_1_830;
mixer gate_output_1_830(.a(output_2_830), .b(output_2_0), .y(output_1_830));
wire output_3_830, output_3_0, output_2_830;
mixer gate_output_2_830(.a(output_3_830), .b(output_3_0), .y(output_2_830));
wire output_1_831, output_1_1, output_0_831;
mixer gate_output_0_831(.a(output_1_831), .b(output_1_1), .y(output_0_831));
wire output_2_831, output_2_1, output_1_831;
mixer gate_output_1_831(.a(output_2_831), .b(output_2_1), .y(output_1_831));
wire output_3_831, output_3_1, output_2_831;
mixer gate_output_2_831(.a(output_3_831), .b(output_3_1), .y(output_2_831));
wire output_1_832, output_1_2, output_0_832;
mixer gate_output_0_832(.a(output_1_832), .b(output_1_2), .y(output_0_832));
wire output_2_832, output_2_2, output_1_832;
mixer gate_output_1_832(.a(output_2_832), .b(output_2_2), .y(output_1_832));
wire output_3_832, output_3_2, output_2_832;
mixer gate_output_2_832(.a(output_3_832), .b(output_3_2), .y(output_2_832));
wire output_1_833, output_1_0, output_0_833;
mixer gate_output_0_833(.a(output_1_833), .b(output_1_0), .y(output_0_833));
wire output_2_833, output_2_0, output_1_833;
mixer gate_output_1_833(.a(output_2_833), .b(output_2_0), .y(output_1_833));
wire output_3_833, output_3_0, output_2_833;
mixer gate_output_2_833(.a(output_3_833), .b(output_3_0), .y(output_2_833));
wire output_1_834, output_1_1, output_0_834;
mixer gate_output_0_834(.a(output_1_834), .b(output_1_1), .y(output_0_834));
wire output_2_834, output_2_1, output_1_834;
mixer gate_output_1_834(.a(output_2_834), .b(output_2_1), .y(output_1_834));
wire output_3_834, output_3_1, output_2_834;
mixer gate_output_2_834(.a(output_3_834), .b(output_3_1), .y(output_2_834));
wire output_1_835, output_1_2, output_0_835;
mixer gate_output_0_835(.a(output_1_835), .b(output_1_2), .y(output_0_835));
wire output_2_835, output_2_2, output_1_835;
mixer gate_output_1_835(.a(output_2_835), .b(output_2_2), .y(output_1_835));
wire output_3_835, output_3_2, output_2_835;
mixer gate_output_2_835(.a(output_3_835), .b(output_3_2), .y(output_2_835));
wire output_1_836, output_1_0, output_0_836;
mixer gate_output_0_836(.a(output_1_836), .b(output_1_0), .y(output_0_836));
wire output_2_836, output_2_0, output_1_836;
mixer gate_output_1_836(.a(output_2_836), .b(output_2_0), .y(output_1_836));
wire output_3_836, output_3_0, output_2_836;
mixer gate_output_2_836(.a(output_3_836), .b(output_3_0), .y(output_2_836));
wire output_1_837, output_1_1, output_0_837;
mixer gate_output_0_837(.a(output_1_837), .b(output_1_1), .y(output_0_837));
wire output_2_837, output_2_1, output_1_837;
mixer gate_output_1_837(.a(output_2_837), .b(output_2_1), .y(output_1_837));
wire output_3_837, output_3_1, output_2_837;
mixer gate_output_2_837(.a(output_3_837), .b(output_3_1), .y(output_2_837));
wire output_1_838, output_1_2, output_0_838;
mixer gate_output_0_838(.a(output_1_838), .b(output_1_2), .y(output_0_838));
wire output_2_838, output_2_2, output_1_838;
mixer gate_output_1_838(.a(output_2_838), .b(output_2_2), .y(output_1_838));
wire output_3_838, output_3_2, output_2_838;
mixer gate_output_2_838(.a(output_3_838), .b(output_3_2), .y(output_2_838));
wire output_1_839, output_1_0, output_0_839;
mixer gate_output_0_839(.a(output_1_839), .b(output_1_0), .y(output_0_839));
wire output_2_839, output_2_0, output_1_839;
mixer gate_output_1_839(.a(output_2_839), .b(output_2_0), .y(output_1_839));
wire output_3_839, output_3_0, output_2_839;
mixer gate_output_2_839(.a(output_3_839), .b(output_3_0), .y(output_2_839));
wire output_1_840, output_1_1, output_0_840;
mixer gate_output_0_840(.a(output_1_840), .b(output_1_1), .y(output_0_840));
wire output_2_840, output_2_1, output_1_840;
mixer gate_output_1_840(.a(output_2_840), .b(output_2_1), .y(output_1_840));
wire output_3_840, output_3_1, output_2_840;
mixer gate_output_2_840(.a(output_3_840), .b(output_3_1), .y(output_2_840));
wire output_1_841, output_1_2, output_0_841;
mixer gate_output_0_841(.a(output_1_841), .b(output_1_2), .y(output_0_841));
wire output_2_841, output_2_2, output_1_841;
mixer gate_output_1_841(.a(output_2_841), .b(output_2_2), .y(output_1_841));
wire output_3_841, output_3_2, output_2_841;
mixer gate_output_2_841(.a(output_3_841), .b(output_3_2), .y(output_2_841));
wire output_1_842, output_1_0, output_0_842;
mixer gate_output_0_842(.a(output_1_842), .b(output_1_0), .y(output_0_842));
wire output_2_842, output_2_0, output_1_842;
mixer gate_output_1_842(.a(output_2_842), .b(output_2_0), .y(output_1_842));
wire output_3_842, output_3_0, output_2_842;
mixer gate_output_2_842(.a(output_3_842), .b(output_3_0), .y(output_2_842));
wire output_1_843, output_1_1, output_0_843;
mixer gate_output_0_843(.a(output_1_843), .b(output_1_1), .y(output_0_843));
wire output_2_843, output_2_1, output_1_843;
mixer gate_output_1_843(.a(output_2_843), .b(output_2_1), .y(output_1_843));
wire output_3_843, output_3_1, output_2_843;
mixer gate_output_2_843(.a(output_3_843), .b(output_3_1), .y(output_2_843));
wire output_1_844, output_1_2, output_0_844;
mixer gate_output_0_844(.a(output_1_844), .b(output_1_2), .y(output_0_844));
wire output_2_844, output_2_2, output_1_844;
mixer gate_output_1_844(.a(output_2_844), .b(output_2_2), .y(output_1_844));
wire output_3_844, output_3_2, output_2_844;
mixer gate_output_2_844(.a(output_3_844), .b(output_3_2), .y(output_2_844));
wire output_1_845, output_1_0, output_0_845;
mixer gate_output_0_845(.a(output_1_845), .b(output_1_0), .y(output_0_845));
wire output_2_845, output_2_0, output_1_845;
mixer gate_output_1_845(.a(output_2_845), .b(output_2_0), .y(output_1_845));
wire output_3_845, output_3_0, output_2_845;
mixer gate_output_2_845(.a(output_3_845), .b(output_3_0), .y(output_2_845));
wire output_1_846, output_1_1, output_0_846;
mixer gate_output_0_846(.a(output_1_846), .b(output_1_1), .y(output_0_846));
wire output_2_846, output_2_1, output_1_846;
mixer gate_output_1_846(.a(output_2_846), .b(output_2_1), .y(output_1_846));
wire output_3_846, output_3_1, output_2_846;
mixer gate_output_2_846(.a(output_3_846), .b(output_3_1), .y(output_2_846));
wire output_1_847, output_1_2, output_0_847;
mixer gate_output_0_847(.a(output_1_847), .b(output_1_2), .y(output_0_847));
wire output_2_847, output_2_2, output_1_847;
mixer gate_output_1_847(.a(output_2_847), .b(output_2_2), .y(output_1_847));
wire output_3_847, output_3_2, output_2_847;
mixer gate_output_2_847(.a(output_3_847), .b(output_3_2), .y(output_2_847));
wire output_1_848, output_1_0, output_0_848;
mixer gate_output_0_848(.a(output_1_848), .b(output_1_0), .y(output_0_848));
wire output_2_848, output_2_0, output_1_848;
mixer gate_output_1_848(.a(output_2_848), .b(output_2_0), .y(output_1_848));
wire output_3_848, output_3_0, output_2_848;
mixer gate_output_2_848(.a(output_3_848), .b(output_3_0), .y(output_2_848));
wire output_1_849, output_1_1, output_0_849;
mixer gate_output_0_849(.a(output_1_849), .b(output_1_1), .y(output_0_849));
wire output_2_849, output_2_1, output_1_849;
mixer gate_output_1_849(.a(output_2_849), .b(output_2_1), .y(output_1_849));
wire output_3_849, output_3_1, output_2_849;
mixer gate_output_2_849(.a(output_3_849), .b(output_3_1), .y(output_2_849));
wire output_1_850, output_1_2, output_0_850;
mixer gate_output_0_850(.a(output_1_850), .b(output_1_2), .y(output_0_850));
wire output_2_850, output_2_2, output_1_850;
mixer gate_output_1_850(.a(output_2_850), .b(output_2_2), .y(output_1_850));
wire output_3_850, output_3_2, output_2_850;
mixer gate_output_2_850(.a(output_3_850), .b(output_3_2), .y(output_2_850));
wire output_1_851, output_1_0, output_0_851;
mixer gate_output_0_851(.a(output_1_851), .b(output_1_0), .y(output_0_851));
wire output_2_851, output_2_0, output_1_851;
mixer gate_output_1_851(.a(output_2_851), .b(output_2_0), .y(output_1_851));
wire output_3_851, output_3_0, output_2_851;
mixer gate_output_2_851(.a(output_3_851), .b(output_3_0), .y(output_2_851));
wire output_1_852, output_1_1, output_0_852;
mixer gate_output_0_852(.a(output_1_852), .b(output_1_1), .y(output_0_852));
wire output_2_852, output_2_1, output_1_852;
mixer gate_output_1_852(.a(output_2_852), .b(output_2_1), .y(output_1_852));
wire output_3_852, output_3_1, output_2_852;
mixer gate_output_2_852(.a(output_3_852), .b(output_3_1), .y(output_2_852));
wire output_1_853, output_1_2, output_0_853;
mixer gate_output_0_853(.a(output_1_853), .b(output_1_2), .y(output_0_853));
wire output_2_853, output_2_2, output_1_853;
mixer gate_output_1_853(.a(output_2_853), .b(output_2_2), .y(output_1_853));
wire output_3_853, output_3_2, output_2_853;
mixer gate_output_2_853(.a(output_3_853), .b(output_3_2), .y(output_2_853));
wire output_1_854, output_1_0, output_0_854;
mixer gate_output_0_854(.a(output_1_854), .b(output_1_0), .y(output_0_854));
wire output_2_854, output_2_0, output_1_854;
mixer gate_output_1_854(.a(output_2_854), .b(output_2_0), .y(output_1_854));
wire output_3_854, output_3_0, output_2_854;
mixer gate_output_2_854(.a(output_3_854), .b(output_3_0), .y(output_2_854));
wire output_1_855, output_1_1, output_0_855;
mixer gate_output_0_855(.a(output_1_855), .b(output_1_1), .y(output_0_855));
wire output_2_855, output_2_1, output_1_855;
mixer gate_output_1_855(.a(output_2_855), .b(output_2_1), .y(output_1_855));
wire output_3_855, output_3_1, output_2_855;
mixer gate_output_2_855(.a(output_3_855), .b(output_3_1), .y(output_2_855));
wire output_1_856, output_1_2, output_0_856;
mixer gate_output_0_856(.a(output_1_856), .b(output_1_2), .y(output_0_856));
wire output_2_856, output_2_2, output_1_856;
mixer gate_output_1_856(.a(output_2_856), .b(output_2_2), .y(output_1_856));
wire output_3_856, output_3_2, output_2_856;
mixer gate_output_2_856(.a(output_3_856), .b(output_3_2), .y(output_2_856));
wire output_1_857, output_1_0, output_0_857;
mixer gate_output_0_857(.a(output_1_857), .b(output_1_0), .y(output_0_857));
wire output_2_857, output_2_0, output_1_857;
mixer gate_output_1_857(.a(output_2_857), .b(output_2_0), .y(output_1_857));
wire output_3_857, output_3_0, output_2_857;
mixer gate_output_2_857(.a(output_3_857), .b(output_3_0), .y(output_2_857));
wire output_1_858, output_1_1, output_0_858;
mixer gate_output_0_858(.a(output_1_858), .b(output_1_1), .y(output_0_858));
wire output_2_858, output_2_1, output_1_858;
mixer gate_output_1_858(.a(output_2_858), .b(output_2_1), .y(output_1_858));
wire output_3_858, output_3_1, output_2_858;
mixer gate_output_2_858(.a(output_3_858), .b(output_3_1), .y(output_2_858));
wire output_1_859, output_1_2, output_0_859;
mixer gate_output_0_859(.a(output_1_859), .b(output_1_2), .y(output_0_859));
wire output_2_859, output_2_2, output_1_859;
mixer gate_output_1_859(.a(output_2_859), .b(output_2_2), .y(output_1_859));
wire output_3_859, output_3_2, output_2_859;
mixer gate_output_2_859(.a(output_3_859), .b(output_3_2), .y(output_2_859));
wire output_1_860, output_1_0, output_0_860;
mixer gate_output_0_860(.a(output_1_860), .b(output_1_0), .y(output_0_860));
wire output_2_860, output_2_0, output_1_860;
mixer gate_output_1_860(.a(output_2_860), .b(output_2_0), .y(output_1_860));
wire output_3_860, output_3_0, output_2_860;
mixer gate_output_2_860(.a(output_3_860), .b(output_3_0), .y(output_2_860));
wire output_1_861, output_1_1, output_0_861;
mixer gate_output_0_861(.a(output_1_861), .b(output_1_1), .y(output_0_861));
wire output_2_861, output_2_1, output_1_861;
mixer gate_output_1_861(.a(output_2_861), .b(output_2_1), .y(output_1_861));
wire output_3_861, output_3_1, output_2_861;
mixer gate_output_2_861(.a(output_3_861), .b(output_3_1), .y(output_2_861));
wire output_1_862, output_1_2, output_0_862;
mixer gate_output_0_862(.a(output_1_862), .b(output_1_2), .y(output_0_862));
wire output_2_862, output_2_2, output_1_862;
mixer gate_output_1_862(.a(output_2_862), .b(output_2_2), .y(output_1_862));
wire output_3_862, output_3_2, output_2_862;
mixer gate_output_2_862(.a(output_3_862), .b(output_3_2), .y(output_2_862));
wire output_1_863, output_1_0, output_0_863;
mixer gate_output_0_863(.a(output_1_863), .b(output_1_0), .y(output_0_863));
wire output_2_863, output_2_0, output_1_863;
mixer gate_output_1_863(.a(output_2_863), .b(output_2_0), .y(output_1_863));
wire output_3_863, output_3_0, output_2_863;
mixer gate_output_2_863(.a(output_3_863), .b(output_3_0), .y(output_2_863));
wire output_1_864, output_1_1, output_0_864;
mixer gate_output_0_864(.a(output_1_864), .b(output_1_1), .y(output_0_864));
wire output_2_864, output_2_1, output_1_864;
mixer gate_output_1_864(.a(output_2_864), .b(output_2_1), .y(output_1_864));
wire output_3_864, output_3_1, output_2_864;
mixer gate_output_2_864(.a(output_3_864), .b(output_3_1), .y(output_2_864));
wire output_1_865, output_1_2, output_0_865;
mixer gate_output_0_865(.a(output_1_865), .b(output_1_2), .y(output_0_865));
wire output_2_865, output_2_2, output_1_865;
mixer gate_output_1_865(.a(output_2_865), .b(output_2_2), .y(output_1_865));
wire output_3_865, output_3_2, output_2_865;
mixer gate_output_2_865(.a(output_3_865), .b(output_3_2), .y(output_2_865));
wire output_1_866, output_1_0, output_0_866;
mixer gate_output_0_866(.a(output_1_866), .b(output_1_0), .y(output_0_866));
wire output_2_866, output_2_0, output_1_866;
mixer gate_output_1_866(.a(output_2_866), .b(output_2_0), .y(output_1_866));
wire output_3_866, output_3_0, output_2_866;
mixer gate_output_2_866(.a(output_3_866), .b(output_3_0), .y(output_2_866));
wire output_1_867, output_1_1, output_0_867;
mixer gate_output_0_867(.a(output_1_867), .b(output_1_1), .y(output_0_867));
wire output_2_867, output_2_1, output_1_867;
mixer gate_output_1_867(.a(output_2_867), .b(output_2_1), .y(output_1_867));
wire output_3_867, output_3_1, output_2_867;
mixer gate_output_2_867(.a(output_3_867), .b(output_3_1), .y(output_2_867));
wire output_1_868, output_1_2, output_0_868;
mixer gate_output_0_868(.a(output_1_868), .b(output_1_2), .y(output_0_868));
wire output_2_868, output_2_2, output_1_868;
mixer gate_output_1_868(.a(output_2_868), .b(output_2_2), .y(output_1_868));
wire output_3_868, output_3_2, output_2_868;
mixer gate_output_2_868(.a(output_3_868), .b(output_3_2), .y(output_2_868));
wire output_1_869, output_1_0, output_0_869;
mixer gate_output_0_869(.a(output_1_869), .b(output_1_0), .y(output_0_869));
wire output_2_869, output_2_0, output_1_869;
mixer gate_output_1_869(.a(output_2_869), .b(output_2_0), .y(output_1_869));
wire output_3_869, output_3_0, output_2_869;
mixer gate_output_2_869(.a(output_3_869), .b(output_3_0), .y(output_2_869));
wire output_1_870, output_1_1, output_0_870;
mixer gate_output_0_870(.a(output_1_870), .b(output_1_1), .y(output_0_870));
wire output_2_870, output_2_1, output_1_870;
mixer gate_output_1_870(.a(output_2_870), .b(output_2_1), .y(output_1_870));
wire output_3_870, output_3_1, output_2_870;
mixer gate_output_2_870(.a(output_3_870), .b(output_3_1), .y(output_2_870));
wire output_1_871, output_1_2, output_0_871;
mixer gate_output_0_871(.a(output_1_871), .b(output_1_2), .y(output_0_871));
wire output_2_871, output_2_2, output_1_871;
mixer gate_output_1_871(.a(output_2_871), .b(output_2_2), .y(output_1_871));
wire output_3_871, output_3_2, output_2_871;
mixer gate_output_2_871(.a(output_3_871), .b(output_3_2), .y(output_2_871));
wire output_1_872, output_1_0, output_0_872;
mixer gate_output_0_872(.a(output_1_872), .b(output_1_0), .y(output_0_872));
wire output_2_872, output_2_0, output_1_872;
mixer gate_output_1_872(.a(output_2_872), .b(output_2_0), .y(output_1_872));
wire output_3_872, output_3_0, output_2_872;
mixer gate_output_2_872(.a(output_3_872), .b(output_3_0), .y(output_2_872));
wire output_1_873, output_1_1, output_0_873;
mixer gate_output_0_873(.a(output_1_873), .b(output_1_1), .y(output_0_873));
wire output_2_873, output_2_1, output_1_873;
mixer gate_output_1_873(.a(output_2_873), .b(output_2_1), .y(output_1_873));
wire output_3_873, output_3_1, output_2_873;
mixer gate_output_2_873(.a(output_3_873), .b(output_3_1), .y(output_2_873));
wire output_1_874, output_1_2, output_0_874;
mixer gate_output_0_874(.a(output_1_874), .b(output_1_2), .y(output_0_874));
wire output_2_874, output_2_2, output_1_874;
mixer gate_output_1_874(.a(output_2_874), .b(output_2_2), .y(output_1_874));
wire output_3_874, output_3_2, output_2_874;
mixer gate_output_2_874(.a(output_3_874), .b(output_3_2), .y(output_2_874));
wire output_1_875, output_1_0, output_0_875;
mixer gate_output_0_875(.a(output_1_875), .b(output_1_0), .y(output_0_875));
wire output_2_875, output_2_0, output_1_875;
mixer gate_output_1_875(.a(output_2_875), .b(output_2_0), .y(output_1_875));
wire output_3_875, output_3_0, output_2_875;
mixer gate_output_2_875(.a(output_3_875), .b(output_3_0), .y(output_2_875));
wire output_1_876, output_1_1, output_0_876;
mixer gate_output_0_876(.a(output_1_876), .b(output_1_1), .y(output_0_876));
wire output_2_876, output_2_1, output_1_876;
mixer gate_output_1_876(.a(output_2_876), .b(output_2_1), .y(output_1_876));
wire output_3_876, output_3_1, output_2_876;
mixer gate_output_2_876(.a(output_3_876), .b(output_3_1), .y(output_2_876));
wire output_1_877, output_1_2, output_0_877;
mixer gate_output_0_877(.a(output_1_877), .b(output_1_2), .y(output_0_877));
wire output_2_877, output_2_2, output_1_877;
mixer gate_output_1_877(.a(output_2_877), .b(output_2_2), .y(output_1_877));
wire output_3_877, output_3_2, output_2_877;
mixer gate_output_2_877(.a(output_3_877), .b(output_3_2), .y(output_2_877));
wire output_1_878, output_1_0, output_0_878;
mixer gate_output_0_878(.a(output_1_878), .b(output_1_0), .y(output_0_878));
wire output_2_878, output_2_0, output_1_878;
mixer gate_output_1_878(.a(output_2_878), .b(output_2_0), .y(output_1_878));
wire output_3_878, output_3_0, output_2_878;
mixer gate_output_2_878(.a(output_3_878), .b(output_3_0), .y(output_2_878));
wire output_1_879, output_1_1, output_0_879;
mixer gate_output_0_879(.a(output_1_879), .b(output_1_1), .y(output_0_879));
wire output_2_879, output_2_1, output_1_879;
mixer gate_output_1_879(.a(output_2_879), .b(output_2_1), .y(output_1_879));
wire output_3_879, output_3_1, output_2_879;
mixer gate_output_2_879(.a(output_3_879), .b(output_3_1), .y(output_2_879));
wire output_1_880, output_1_2, output_0_880;
mixer gate_output_0_880(.a(output_1_880), .b(output_1_2), .y(output_0_880));
wire output_2_880, output_2_2, output_1_880;
mixer gate_output_1_880(.a(output_2_880), .b(output_2_2), .y(output_1_880));
wire output_3_880, output_3_2, output_2_880;
mixer gate_output_2_880(.a(output_3_880), .b(output_3_2), .y(output_2_880));
wire output_1_881, output_1_0, output_0_881;
mixer gate_output_0_881(.a(output_1_881), .b(output_1_0), .y(output_0_881));
wire output_2_881, output_2_0, output_1_881;
mixer gate_output_1_881(.a(output_2_881), .b(output_2_0), .y(output_1_881));
wire output_3_881, output_3_0, output_2_881;
mixer gate_output_2_881(.a(output_3_881), .b(output_3_0), .y(output_2_881));
wire output_1_882, output_1_1, output_0_882;
mixer gate_output_0_882(.a(output_1_882), .b(output_1_1), .y(output_0_882));
wire output_2_882, output_2_1, output_1_882;
mixer gate_output_1_882(.a(output_2_882), .b(output_2_1), .y(output_1_882));
wire output_3_882, output_3_1, output_2_882;
mixer gate_output_2_882(.a(output_3_882), .b(output_3_1), .y(output_2_882));
wire output_1_883, output_1_2, output_0_883;
mixer gate_output_0_883(.a(output_1_883), .b(output_1_2), .y(output_0_883));
wire output_2_883, output_2_2, output_1_883;
mixer gate_output_1_883(.a(output_2_883), .b(output_2_2), .y(output_1_883));
wire output_3_883, output_3_2, output_2_883;
mixer gate_output_2_883(.a(output_3_883), .b(output_3_2), .y(output_2_883));
wire output_1_884, output_1_0, output_0_884;
mixer gate_output_0_884(.a(output_1_884), .b(output_1_0), .y(output_0_884));
wire output_2_884, output_2_0, output_1_884;
mixer gate_output_1_884(.a(output_2_884), .b(output_2_0), .y(output_1_884));
wire output_3_884, output_3_0, output_2_884;
mixer gate_output_2_884(.a(output_3_884), .b(output_3_0), .y(output_2_884));
wire output_1_885, output_1_1, output_0_885;
mixer gate_output_0_885(.a(output_1_885), .b(output_1_1), .y(output_0_885));
wire output_2_885, output_2_1, output_1_885;
mixer gate_output_1_885(.a(output_2_885), .b(output_2_1), .y(output_1_885));
wire output_3_885, output_3_1, output_2_885;
mixer gate_output_2_885(.a(output_3_885), .b(output_3_1), .y(output_2_885));
wire output_1_886, output_1_2, output_0_886;
mixer gate_output_0_886(.a(output_1_886), .b(output_1_2), .y(output_0_886));
wire output_2_886, output_2_2, output_1_886;
mixer gate_output_1_886(.a(output_2_886), .b(output_2_2), .y(output_1_886));
wire output_3_886, output_3_2, output_2_886;
mixer gate_output_2_886(.a(output_3_886), .b(output_3_2), .y(output_2_886));
wire output_1_887, output_1_0, output_0_887;
mixer gate_output_0_887(.a(output_1_887), .b(output_1_0), .y(output_0_887));
wire output_2_887, output_2_0, output_1_887;
mixer gate_output_1_887(.a(output_2_887), .b(output_2_0), .y(output_1_887));
wire output_3_887, output_3_0, output_2_887;
mixer gate_output_2_887(.a(output_3_887), .b(output_3_0), .y(output_2_887));
wire output_1_888, output_1_1, output_0_888;
mixer gate_output_0_888(.a(output_1_888), .b(output_1_1), .y(output_0_888));
wire output_2_888, output_2_1, output_1_888;
mixer gate_output_1_888(.a(output_2_888), .b(output_2_1), .y(output_1_888));
wire output_3_888, output_3_1, output_2_888;
mixer gate_output_2_888(.a(output_3_888), .b(output_3_1), .y(output_2_888));
wire output_1_889, output_1_2, output_0_889;
mixer gate_output_0_889(.a(output_1_889), .b(output_1_2), .y(output_0_889));
wire output_2_889, output_2_2, output_1_889;
mixer gate_output_1_889(.a(output_2_889), .b(output_2_2), .y(output_1_889));
wire output_3_889, output_3_2, output_2_889;
mixer gate_output_2_889(.a(output_3_889), .b(output_3_2), .y(output_2_889));
wire output_1_890, output_1_0, output_0_890;
mixer gate_output_0_890(.a(output_1_890), .b(output_1_0), .y(output_0_890));
wire output_2_890, output_2_0, output_1_890;
mixer gate_output_1_890(.a(output_2_890), .b(output_2_0), .y(output_1_890));
wire output_3_890, output_3_0, output_2_890;
mixer gate_output_2_890(.a(output_3_890), .b(output_3_0), .y(output_2_890));
wire output_1_891, output_1_1, output_0_891;
mixer gate_output_0_891(.a(output_1_891), .b(output_1_1), .y(output_0_891));
wire output_2_891, output_2_1, output_1_891;
mixer gate_output_1_891(.a(output_2_891), .b(output_2_1), .y(output_1_891));
wire output_3_891, output_3_1, output_2_891;
mixer gate_output_2_891(.a(output_3_891), .b(output_3_1), .y(output_2_891));
wire output_1_892, output_1_2, output_0_892;
mixer gate_output_0_892(.a(output_1_892), .b(output_1_2), .y(output_0_892));
wire output_2_892, output_2_2, output_1_892;
mixer gate_output_1_892(.a(output_2_892), .b(output_2_2), .y(output_1_892));
wire output_3_892, output_3_2, output_2_892;
mixer gate_output_2_892(.a(output_3_892), .b(output_3_2), .y(output_2_892));
wire output_1_893, output_1_0, output_0_893;
mixer gate_output_0_893(.a(output_1_893), .b(output_1_0), .y(output_0_893));
wire output_2_893, output_2_0, output_1_893;
mixer gate_output_1_893(.a(output_2_893), .b(output_2_0), .y(output_1_893));
wire output_3_893, output_3_0, output_2_893;
mixer gate_output_2_893(.a(output_3_893), .b(output_3_0), .y(output_2_893));
wire output_1_894, output_1_1, output_0_894;
mixer gate_output_0_894(.a(output_1_894), .b(output_1_1), .y(output_0_894));
wire output_2_894, output_2_1, output_1_894;
mixer gate_output_1_894(.a(output_2_894), .b(output_2_1), .y(output_1_894));
wire output_3_894, output_3_1, output_2_894;
mixer gate_output_2_894(.a(output_3_894), .b(output_3_1), .y(output_2_894));
wire output_1_895, output_1_2, output_0_895;
mixer gate_output_0_895(.a(output_1_895), .b(output_1_2), .y(output_0_895));
wire output_2_895, output_2_2, output_1_895;
mixer gate_output_1_895(.a(output_2_895), .b(output_2_2), .y(output_1_895));
wire output_3_895, output_3_2, output_2_895;
mixer gate_output_2_895(.a(output_3_895), .b(output_3_2), .y(output_2_895));
wire output_1_896, output_1_0, output_0_896;
mixer gate_output_0_896(.a(output_1_896), .b(output_1_0), .y(output_0_896));
wire output_2_896, output_2_0, output_1_896;
mixer gate_output_1_896(.a(output_2_896), .b(output_2_0), .y(output_1_896));
wire output_3_896, output_3_0, output_2_896;
mixer gate_output_2_896(.a(output_3_896), .b(output_3_0), .y(output_2_896));
wire output_1_897, output_1_1, output_0_897;
mixer gate_output_0_897(.a(output_1_897), .b(output_1_1), .y(output_0_897));
wire output_2_897, output_2_1, output_1_897;
mixer gate_output_1_897(.a(output_2_897), .b(output_2_1), .y(output_1_897));
wire output_3_897, output_3_1, output_2_897;
mixer gate_output_2_897(.a(output_3_897), .b(output_3_1), .y(output_2_897));
wire output_1_898, output_1_2, output_0_898;
mixer gate_output_0_898(.a(output_1_898), .b(output_1_2), .y(output_0_898));
wire output_2_898, output_2_2, output_1_898;
mixer gate_output_1_898(.a(output_2_898), .b(output_2_2), .y(output_1_898));
wire output_3_898, output_3_2, output_2_898;
mixer gate_output_2_898(.a(output_3_898), .b(output_3_2), .y(output_2_898));
wire output_1_899, output_1_0, output_0_899;
mixer gate_output_0_899(.a(output_1_899), .b(output_1_0), .y(output_0_899));
wire output_2_899, output_2_0, output_1_899;
mixer gate_output_1_899(.a(output_2_899), .b(output_2_0), .y(output_1_899));
wire output_3_899, output_3_0, output_2_899;
mixer gate_output_2_899(.a(output_3_899), .b(output_3_0), .y(output_2_899));
wire output_1_900, output_1_1, output_0_900;
mixer gate_output_0_900(.a(output_1_900), .b(output_1_1), .y(output_0_900));
wire output_2_900, output_2_1, output_1_900;
mixer gate_output_1_900(.a(output_2_900), .b(output_2_1), .y(output_1_900));
wire output_3_900, output_3_1, output_2_900;
mixer gate_output_2_900(.a(output_3_900), .b(output_3_1), .y(output_2_900));
wire output_1_901, output_1_2, output_0_901;
mixer gate_output_0_901(.a(output_1_901), .b(output_1_2), .y(output_0_901));
wire output_2_901, output_2_2, output_1_901;
mixer gate_output_1_901(.a(output_2_901), .b(output_2_2), .y(output_1_901));
wire output_3_901, output_3_2, output_2_901;
mixer gate_output_2_901(.a(output_3_901), .b(output_3_2), .y(output_2_901));
wire output_1_902, output_1_0, output_0_902;
mixer gate_output_0_902(.a(output_1_902), .b(output_1_0), .y(output_0_902));
wire output_2_902, output_2_0, output_1_902;
mixer gate_output_1_902(.a(output_2_902), .b(output_2_0), .y(output_1_902));
wire output_3_902, output_3_0, output_2_902;
mixer gate_output_2_902(.a(output_3_902), .b(output_3_0), .y(output_2_902));
wire output_1_903, output_1_1, output_0_903;
mixer gate_output_0_903(.a(output_1_903), .b(output_1_1), .y(output_0_903));
wire output_2_903, output_2_1, output_1_903;
mixer gate_output_1_903(.a(output_2_903), .b(output_2_1), .y(output_1_903));
wire output_3_903, output_3_1, output_2_903;
mixer gate_output_2_903(.a(output_3_903), .b(output_3_1), .y(output_2_903));
wire output_1_904, output_1_2, output_0_904;
mixer gate_output_0_904(.a(output_1_904), .b(output_1_2), .y(output_0_904));
wire output_2_904, output_2_2, output_1_904;
mixer gate_output_1_904(.a(output_2_904), .b(output_2_2), .y(output_1_904));
wire output_3_904, output_3_2, output_2_904;
mixer gate_output_2_904(.a(output_3_904), .b(output_3_2), .y(output_2_904));
wire output_1_905, output_1_0, output_0_905;
mixer gate_output_0_905(.a(output_1_905), .b(output_1_0), .y(output_0_905));
wire output_2_905, output_2_0, output_1_905;
mixer gate_output_1_905(.a(output_2_905), .b(output_2_0), .y(output_1_905));
wire output_3_905, output_3_0, output_2_905;
mixer gate_output_2_905(.a(output_3_905), .b(output_3_0), .y(output_2_905));
wire output_1_906, output_1_1, output_0_906;
mixer gate_output_0_906(.a(output_1_906), .b(output_1_1), .y(output_0_906));
wire output_2_906, output_2_1, output_1_906;
mixer gate_output_1_906(.a(output_2_906), .b(output_2_1), .y(output_1_906));
wire output_3_906, output_3_1, output_2_906;
mixer gate_output_2_906(.a(output_3_906), .b(output_3_1), .y(output_2_906));
wire output_1_907, output_1_2, output_0_907;
mixer gate_output_0_907(.a(output_1_907), .b(output_1_2), .y(output_0_907));
wire output_2_907, output_2_2, output_1_907;
mixer gate_output_1_907(.a(output_2_907), .b(output_2_2), .y(output_1_907));
wire output_3_907, output_3_2, output_2_907;
mixer gate_output_2_907(.a(output_3_907), .b(output_3_2), .y(output_2_907));
wire output_1_908, output_1_0, output_0_908;
mixer gate_output_0_908(.a(output_1_908), .b(output_1_0), .y(output_0_908));
wire output_2_908, output_2_0, output_1_908;
mixer gate_output_1_908(.a(output_2_908), .b(output_2_0), .y(output_1_908));
wire output_3_908, output_3_0, output_2_908;
mixer gate_output_2_908(.a(output_3_908), .b(output_3_0), .y(output_2_908));
wire output_1_909, output_1_1, output_0_909;
mixer gate_output_0_909(.a(output_1_909), .b(output_1_1), .y(output_0_909));
wire output_2_909, output_2_1, output_1_909;
mixer gate_output_1_909(.a(output_2_909), .b(output_2_1), .y(output_1_909));
wire output_3_909, output_3_1, output_2_909;
mixer gate_output_2_909(.a(output_3_909), .b(output_3_1), .y(output_2_909));
wire output_1_910, output_1_2, output_0_910;
mixer gate_output_0_910(.a(output_1_910), .b(output_1_2), .y(output_0_910));
wire output_2_910, output_2_2, output_1_910;
mixer gate_output_1_910(.a(output_2_910), .b(output_2_2), .y(output_1_910));
wire output_3_910, output_3_2, output_2_910;
mixer gate_output_2_910(.a(output_3_910), .b(output_3_2), .y(output_2_910));
wire output_1_911, output_1_0, output_0_911;
mixer gate_output_0_911(.a(output_1_911), .b(output_1_0), .y(output_0_911));
wire output_2_911, output_2_0, output_1_911;
mixer gate_output_1_911(.a(output_2_911), .b(output_2_0), .y(output_1_911));
wire output_3_911, output_3_0, output_2_911;
mixer gate_output_2_911(.a(output_3_911), .b(output_3_0), .y(output_2_911));
wire output_1_912, output_1_1, output_0_912;
mixer gate_output_0_912(.a(output_1_912), .b(output_1_1), .y(output_0_912));
wire output_2_912, output_2_1, output_1_912;
mixer gate_output_1_912(.a(output_2_912), .b(output_2_1), .y(output_1_912));
wire output_3_912, output_3_1, output_2_912;
mixer gate_output_2_912(.a(output_3_912), .b(output_3_1), .y(output_2_912));
wire output_1_913, output_1_2, output_0_913;
mixer gate_output_0_913(.a(output_1_913), .b(output_1_2), .y(output_0_913));
wire output_2_913, output_2_2, output_1_913;
mixer gate_output_1_913(.a(output_2_913), .b(output_2_2), .y(output_1_913));
wire output_3_913, output_3_2, output_2_913;
mixer gate_output_2_913(.a(output_3_913), .b(output_3_2), .y(output_2_913));
wire output_1_914, output_1_0, output_0_914;
mixer gate_output_0_914(.a(output_1_914), .b(output_1_0), .y(output_0_914));
wire output_2_914, output_2_0, output_1_914;
mixer gate_output_1_914(.a(output_2_914), .b(output_2_0), .y(output_1_914));
wire output_3_914, output_3_0, output_2_914;
mixer gate_output_2_914(.a(output_3_914), .b(output_3_0), .y(output_2_914));
wire output_1_915, output_1_1, output_0_915;
mixer gate_output_0_915(.a(output_1_915), .b(output_1_1), .y(output_0_915));
wire output_2_915, output_2_1, output_1_915;
mixer gate_output_1_915(.a(output_2_915), .b(output_2_1), .y(output_1_915));
wire output_3_915, output_3_1, output_2_915;
mixer gate_output_2_915(.a(output_3_915), .b(output_3_1), .y(output_2_915));
wire output_1_916, output_1_2, output_0_916;
mixer gate_output_0_916(.a(output_1_916), .b(output_1_2), .y(output_0_916));
wire output_2_916, output_2_2, output_1_916;
mixer gate_output_1_916(.a(output_2_916), .b(output_2_2), .y(output_1_916));
wire output_3_916, output_3_2, output_2_916;
mixer gate_output_2_916(.a(output_3_916), .b(output_3_2), .y(output_2_916));
wire output_1_917, output_1_0, output_0_917;
mixer gate_output_0_917(.a(output_1_917), .b(output_1_0), .y(output_0_917));
wire output_2_917, output_2_0, output_1_917;
mixer gate_output_1_917(.a(output_2_917), .b(output_2_0), .y(output_1_917));
wire output_3_917, output_3_0, output_2_917;
mixer gate_output_2_917(.a(output_3_917), .b(output_3_0), .y(output_2_917));
wire output_1_918, output_1_1, output_0_918;
mixer gate_output_0_918(.a(output_1_918), .b(output_1_1), .y(output_0_918));
wire output_2_918, output_2_1, output_1_918;
mixer gate_output_1_918(.a(output_2_918), .b(output_2_1), .y(output_1_918));
wire output_3_918, output_3_1, output_2_918;
mixer gate_output_2_918(.a(output_3_918), .b(output_3_1), .y(output_2_918));
wire output_1_919, output_1_2, output_0_919;
mixer gate_output_0_919(.a(output_1_919), .b(output_1_2), .y(output_0_919));
wire output_2_919, output_2_2, output_1_919;
mixer gate_output_1_919(.a(output_2_919), .b(output_2_2), .y(output_1_919));
wire output_3_919, output_3_2, output_2_919;
mixer gate_output_2_919(.a(output_3_919), .b(output_3_2), .y(output_2_919));
wire output_1_920, output_1_0, output_0_920;
mixer gate_output_0_920(.a(output_1_920), .b(output_1_0), .y(output_0_920));
wire output_2_920, output_2_0, output_1_920;
mixer gate_output_1_920(.a(output_2_920), .b(output_2_0), .y(output_1_920));
wire output_3_920, output_3_0, output_2_920;
mixer gate_output_2_920(.a(output_3_920), .b(output_3_0), .y(output_2_920));
wire output_1_921, output_1_1, output_0_921;
mixer gate_output_0_921(.a(output_1_921), .b(output_1_1), .y(output_0_921));
wire output_2_921, output_2_1, output_1_921;
mixer gate_output_1_921(.a(output_2_921), .b(output_2_1), .y(output_1_921));
wire output_3_921, output_3_1, output_2_921;
mixer gate_output_2_921(.a(output_3_921), .b(output_3_1), .y(output_2_921));
wire output_1_922, output_1_2, output_0_922;
mixer gate_output_0_922(.a(output_1_922), .b(output_1_2), .y(output_0_922));
wire output_2_922, output_2_2, output_1_922;
mixer gate_output_1_922(.a(output_2_922), .b(output_2_2), .y(output_1_922));
wire output_3_922, output_3_2, output_2_922;
mixer gate_output_2_922(.a(output_3_922), .b(output_3_2), .y(output_2_922));
wire output_1_923, output_1_0, output_0_923;
mixer gate_output_0_923(.a(output_1_923), .b(output_1_0), .y(output_0_923));
wire output_2_923, output_2_0, output_1_923;
mixer gate_output_1_923(.a(output_2_923), .b(output_2_0), .y(output_1_923));
wire output_3_923, output_3_0, output_2_923;
mixer gate_output_2_923(.a(output_3_923), .b(output_3_0), .y(output_2_923));
wire output_1_924, output_1_1, output_0_924;
mixer gate_output_0_924(.a(output_1_924), .b(output_1_1), .y(output_0_924));
wire output_2_924, output_2_1, output_1_924;
mixer gate_output_1_924(.a(output_2_924), .b(output_2_1), .y(output_1_924));
wire output_3_924, output_3_1, output_2_924;
mixer gate_output_2_924(.a(output_3_924), .b(output_3_1), .y(output_2_924));
wire output_1_925, output_1_2, output_0_925;
mixer gate_output_0_925(.a(output_1_925), .b(output_1_2), .y(output_0_925));
wire output_2_925, output_2_2, output_1_925;
mixer gate_output_1_925(.a(output_2_925), .b(output_2_2), .y(output_1_925));
wire output_3_925, output_3_2, output_2_925;
mixer gate_output_2_925(.a(output_3_925), .b(output_3_2), .y(output_2_925));
wire output_1_926, output_1_0, output_0_926;
mixer gate_output_0_926(.a(output_1_926), .b(output_1_0), .y(output_0_926));
wire output_2_926, output_2_0, output_1_926;
mixer gate_output_1_926(.a(output_2_926), .b(output_2_0), .y(output_1_926));
wire output_3_926, output_3_0, output_2_926;
mixer gate_output_2_926(.a(output_3_926), .b(output_3_0), .y(output_2_926));
wire output_1_927, output_1_1, output_0_927;
mixer gate_output_0_927(.a(output_1_927), .b(output_1_1), .y(output_0_927));
wire output_2_927, output_2_1, output_1_927;
mixer gate_output_1_927(.a(output_2_927), .b(output_2_1), .y(output_1_927));
wire output_3_927, output_3_1, output_2_927;
mixer gate_output_2_927(.a(output_3_927), .b(output_3_1), .y(output_2_927));
wire output_1_928, output_1_2, output_0_928;
mixer gate_output_0_928(.a(output_1_928), .b(output_1_2), .y(output_0_928));
wire output_2_928, output_2_2, output_1_928;
mixer gate_output_1_928(.a(output_2_928), .b(output_2_2), .y(output_1_928));
wire output_3_928, output_3_2, output_2_928;
mixer gate_output_2_928(.a(output_3_928), .b(output_3_2), .y(output_2_928));
wire output_1_929, output_1_0, output_0_929;
mixer gate_output_0_929(.a(output_1_929), .b(output_1_0), .y(output_0_929));
wire output_2_929, output_2_0, output_1_929;
mixer gate_output_1_929(.a(output_2_929), .b(output_2_0), .y(output_1_929));
wire output_3_929, output_3_0, output_2_929;
mixer gate_output_2_929(.a(output_3_929), .b(output_3_0), .y(output_2_929));
wire output_1_930, output_1_1, output_0_930;
mixer gate_output_0_930(.a(output_1_930), .b(output_1_1), .y(output_0_930));
wire output_2_930, output_2_1, output_1_930;
mixer gate_output_1_930(.a(output_2_930), .b(output_2_1), .y(output_1_930));
wire output_3_930, output_3_1, output_2_930;
mixer gate_output_2_930(.a(output_3_930), .b(output_3_1), .y(output_2_930));
wire output_1_931, output_1_2, output_0_931;
mixer gate_output_0_931(.a(output_1_931), .b(output_1_2), .y(output_0_931));
wire output_2_931, output_2_2, output_1_931;
mixer gate_output_1_931(.a(output_2_931), .b(output_2_2), .y(output_1_931));
wire output_3_931, output_3_2, output_2_931;
mixer gate_output_2_931(.a(output_3_931), .b(output_3_2), .y(output_2_931));
wire output_1_932, output_1_0, output_0_932;
mixer gate_output_0_932(.a(output_1_932), .b(output_1_0), .y(output_0_932));
wire output_2_932, output_2_0, output_1_932;
mixer gate_output_1_932(.a(output_2_932), .b(output_2_0), .y(output_1_932));
wire output_3_932, output_3_0, output_2_932;
mixer gate_output_2_932(.a(output_3_932), .b(output_3_0), .y(output_2_932));
wire output_1_933, output_1_1, output_0_933;
mixer gate_output_0_933(.a(output_1_933), .b(output_1_1), .y(output_0_933));
wire output_2_933, output_2_1, output_1_933;
mixer gate_output_1_933(.a(output_2_933), .b(output_2_1), .y(output_1_933));
wire output_3_933, output_3_1, output_2_933;
mixer gate_output_2_933(.a(output_3_933), .b(output_3_1), .y(output_2_933));
wire output_1_934, output_1_2, output_0_934;
mixer gate_output_0_934(.a(output_1_934), .b(output_1_2), .y(output_0_934));
wire output_2_934, output_2_2, output_1_934;
mixer gate_output_1_934(.a(output_2_934), .b(output_2_2), .y(output_1_934));
wire output_3_934, output_3_2, output_2_934;
mixer gate_output_2_934(.a(output_3_934), .b(output_3_2), .y(output_2_934));
wire output_1_935, output_1_0, output_0_935;
mixer gate_output_0_935(.a(output_1_935), .b(output_1_0), .y(output_0_935));
wire output_2_935, output_2_0, output_1_935;
mixer gate_output_1_935(.a(output_2_935), .b(output_2_0), .y(output_1_935));
wire output_3_935, output_3_0, output_2_935;
mixer gate_output_2_935(.a(output_3_935), .b(output_3_0), .y(output_2_935));
wire output_1_936, output_1_1, output_0_936;
mixer gate_output_0_936(.a(output_1_936), .b(output_1_1), .y(output_0_936));
wire output_2_936, output_2_1, output_1_936;
mixer gate_output_1_936(.a(output_2_936), .b(output_2_1), .y(output_1_936));
wire output_3_936, output_3_1, output_2_936;
mixer gate_output_2_936(.a(output_3_936), .b(output_3_1), .y(output_2_936));
wire output_1_937, output_1_2, output_0_937;
mixer gate_output_0_937(.a(output_1_937), .b(output_1_2), .y(output_0_937));
wire output_2_937, output_2_2, output_1_937;
mixer gate_output_1_937(.a(output_2_937), .b(output_2_2), .y(output_1_937));
wire output_3_937, output_3_2, output_2_937;
mixer gate_output_2_937(.a(output_3_937), .b(output_3_2), .y(output_2_937));
wire output_1_938, output_1_0, output_0_938;
mixer gate_output_0_938(.a(output_1_938), .b(output_1_0), .y(output_0_938));
wire output_2_938, output_2_0, output_1_938;
mixer gate_output_1_938(.a(output_2_938), .b(output_2_0), .y(output_1_938));
wire output_3_938, output_3_0, output_2_938;
mixer gate_output_2_938(.a(output_3_938), .b(output_3_0), .y(output_2_938));
wire output_1_939, output_1_1, output_0_939;
mixer gate_output_0_939(.a(output_1_939), .b(output_1_1), .y(output_0_939));
wire output_2_939, output_2_1, output_1_939;
mixer gate_output_1_939(.a(output_2_939), .b(output_2_1), .y(output_1_939));
wire output_3_939, output_3_1, output_2_939;
mixer gate_output_2_939(.a(output_3_939), .b(output_3_1), .y(output_2_939));
wire output_1_940, output_1_2, output_0_940;
mixer gate_output_0_940(.a(output_1_940), .b(output_1_2), .y(output_0_940));
wire output_2_940, output_2_2, output_1_940;
mixer gate_output_1_940(.a(output_2_940), .b(output_2_2), .y(output_1_940));
wire output_3_940, output_3_2, output_2_940;
mixer gate_output_2_940(.a(output_3_940), .b(output_3_2), .y(output_2_940));
wire output_1_941, output_1_0, output_0_941;
mixer gate_output_0_941(.a(output_1_941), .b(output_1_0), .y(output_0_941));
wire output_2_941, output_2_0, output_1_941;
mixer gate_output_1_941(.a(output_2_941), .b(output_2_0), .y(output_1_941));
wire output_3_941, output_3_0, output_2_941;
mixer gate_output_2_941(.a(output_3_941), .b(output_3_0), .y(output_2_941));
wire output_1_942, output_1_1, output_0_942;
mixer gate_output_0_942(.a(output_1_942), .b(output_1_1), .y(output_0_942));
wire output_2_942, output_2_1, output_1_942;
mixer gate_output_1_942(.a(output_2_942), .b(output_2_1), .y(output_1_942));
wire output_3_942, output_3_1, output_2_942;
mixer gate_output_2_942(.a(output_3_942), .b(output_3_1), .y(output_2_942));
wire output_1_943, output_1_2, output_0_943;
mixer gate_output_0_943(.a(output_1_943), .b(output_1_2), .y(output_0_943));
wire output_2_943, output_2_2, output_1_943;
mixer gate_output_1_943(.a(output_2_943), .b(output_2_2), .y(output_1_943));
wire output_3_943, output_3_2, output_2_943;
mixer gate_output_2_943(.a(output_3_943), .b(output_3_2), .y(output_2_943));
wire output_1_944, output_1_0, output_0_944;
mixer gate_output_0_944(.a(output_1_944), .b(output_1_0), .y(output_0_944));
wire output_2_944, output_2_0, output_1_944;
mixer gate_output_1_944(.a(output_2_944), .b(output_2_0), .y(output_1_944));
wire output_3_944, output_3_0, output_2_944;
mixer gate_output_2_944(.a(output_3_944), .b(output_3_0), .y(output_2_944));
wire output_1_945, output_1_1, output_0_945;
mixer gate_output_0_945(.a(output_1_945), .b(output_1_1), .y(output_0_945));
wire output_2_945, output_2_1, output_1_945;
mixer gate_output_1_945(.a(output_2_945), .b(output_2_1), .y(output_1_945));
wire output_3_945, output_3_1, output_2_945;
mixer gate_output_2_945(.a(output_3_945), .b(output_3_1), .y(output_2_945));
wire output_1_946, output_1_2, output_0_946;
mixer gate_output_0_946(.a(output_1_946), .b(output_1_2), .y(output_0_946));
wire output_2_946, output_2_2, output_1_946;
mixer gate_output_1_946(.a(output_2_946), .b(output_2_2), .y(output_1_946));
wire output_3_946, output_3_2, output_2_946;
mixer gate_output_2_946(.a(output_3_946), .b(output_3_2), .y(output_2_946));
wire output_1_947, output_1_0, output_0_947;
mixer gate_output_0_947(.a(output_1_947), .b(output_1_0), .y(output_0_947));
wire output_2_947, output_2_0, output_1_947;
mixer gate_output_1_947(.a(output_2_947), .b(output_2_0), .y(output_1_947));
wire output_3_947, output_3_0, output_2_947;
mixer gate_output_2_947(.a(output_3_947), .b(output_3_0), .y(output_2_947));
wire output_1_948, output_1_1, output_0_948;
mixer gate_output_0_948(.a(output_1_948), .b(output_1_1), .y(output_0_948));
wire output_2_948, output_2_1, output_1_948;
mixer gate_output_1_948(.a(output_2_948), .b(output_2_1), .y(output_1_948));
wire output_3_948, output_3_1, output_2_948;
mixer gate_output_2_948(.a(output_3_948), .b(output_3_1), .y(output_2_948));
wire output_1_949, output_1_2, output_0_949;
mixer gate_output_0_949(.a(output_1_949), .b(output_1_2), .y(output_0_949));
wire output_2_949, output_2_2, output_1_949;
mixer gate_output_1_949(.a(output_2_949), .b(output_2_2), .y(output_1_949));
wire output_3_949, output_3_2, output_2_949;
mixer gate_output_2_949(.a(output_3_949), .b(output_3_2), .y(output_2_949));
wire output_1_950, output_1_0, output_0_950;
mixer gate_output_0_950(.a(output_1_950), .b(output_1_0), .y(output_0_950));
wire output_2_950, output_2_0, output_1_950;
mixer gate_output_1_950(.a(output_2_950), .b(output_2_0), .y(output_1_950));
wire output_3_950, output_3_0, output_2_950;
mixer gate_output_2_950(.a(output_3_950), .b(output_3_0), .y(output_2_950));
wire output_1_951, output_1_1, output_0_951;
mixer gate_output_0_951(.a(output_1_951), .b(output_1_1), .y(output_0_951));
wire output_2_951, output_2_1, output_1_951;
mixer gate_output_1_951(.a(output_2_951), .b(output_2_1), .y(output_1_951));
wire output_3_951, output_3_1, output_2_951;
mixer gate_output_2_951(.a(output_3_951), .b(output_3_1), .y(output_2_951));
wire output_1_952, output_1_2, output_0_952;
mixer gate_output_0_952(.a(output_1_952), .b(output_1_2), .y(output_0_952));
wire output_2_952, output_2_2, output_1_952;
mixer gate_output_1_952(.a(output_2_952), .b(output_2_2), .y(output_1_952));
wire output_3_952, output_3_2, output_2_952;
mixer gate_output_2_952(.a(output_3_952), .b(output_3_2), .y(output_2_952));
wire output_1_953, output_1_0, output_0_953;
mixer gate_output_0_953(.a(output_1_953), .b(output_1_0), .y(output_0_953));
wire output_2_953, output_2_0, output_1_953;
mixer gate_output_1_953(.a(output_2_953), .b(output_2_0), .y(output_1_953));
wire output_3_953, output_3_0, output_2_953;
mixer gate_output_2_953(.a(output_3_953), .b(output_3_0), .y(output_2_953));
wire output_1_954, output_1_1, output_0_954;
mixer gate_output_0_954(.a(output_1_954), .b(output_1_1), .y(output_0_954));
wire output_2_954, output_2_1, output_1_954;
mixer gate_output_1_954(.a(output_2_954), .b(output_2_1), .y(output_1_954));
wire output_3_954, output_3_1, output_2_954;
mixer gate_output_2_954(.a(output_3_954), .b(output_3_1), .y(output_2_954));
wire output_1_955, output_1_2, output_0_955;
mixer gate_output_0_955(.a(output_1_955), .b(output_1_2), .y(output_0_955));
wire output_2_955, output_2_2, output_1_955;
mixer gate_output_1_955(.a(output_2_955), .b(output_2_2), .y(output_1_955));
wire output_3_955, output_3_2, output_2_955;
mixer gate_output_2_955(.a(output_3_955), .b(output_3_2), .y(output_2_955));
wire output_1_956, output_1_0, output_0_956;
mixer gate_output_0_956(.a(output_1_956), .b(output_1_0), .y(output_0_956));
wire output_2_956, output_2_0, output_1_956;
mixer gate_output_1_956(.a(output_2_956), .b(output_2_0), .y(output_1_956));
wire output_3_956, output_3_0, output_2_956;
mixer gate_output_2_956(.a(output_3_956), .b(output_3_0), .y(output_2_956));
wire output_1_957, output_1_1, output_0_957;
mixer gate_output_0_957(.a(output_1_957), .b(output_1_1), .y(output_0_957));
wire output_2_957, output_2_1, output_1_957;
mixer gate_output_1_957(.a(output_2_957), .b(output_2_1), .y(output_1_957));
wire output_3_957, output_3_1, output_2_957;
mixer gate_output_2_957(.a(output_3_957), .b(output_3_1), .y(output_2_957));
wire output_1_958, output_1_2, output_0_958;
mixer gate_output_0_958(.a(output_1_958), .b(output_1_2), .y(output_0_958));
wire output_2_958, output_2_2, output_1_958;
mixer gate_output_1_958(.a(output_2_958), .b(output_2_2), .y(output_1_958));
wire output_3_958, output_3_2, output_2_958;
mixer gate_output_2_958(.a(output_3_958), .b(output_3_2), .y(output_2_958));
wire output_1_959, output_1_0, output_0_959;
mixer gate_output_0_959(.a(output_1_959), .b(output_1_0), .y(output_0_959));
wire output_2_959, output_2_0, output_1_959;
mixer gate_output_1_959(.a(output_2_959), .b(output_2_0), .y(output_1_959));
wire output_3_959, output_3_0, output_2_959;
mixer gate_output_2_959(.a(output_3_959), .b(output_3_0), .y(output_2_959));
wire output_1_960, output_1_1, output_0_960;
mixer gate_output_0_960(.a(output_1_960), .b(output_1_1), .y(output_0_960));
wire output_2_960, output_2_1, output_1_960;
mixer gate_output_1_960(.a(output_2_960), .b(output_2_1), .y(output_1_960));
wire output_3_960, output_3_1, output_2_960;
mixer gate_output_2_960(.a(output_3_960), .b(output_3_1), .y(output_2_960));
wire output_1_961, output_1_2, output_0_961;
mixer gate_output_0_961(.a(output_1_961), .b(output_1_2), .y(output_0_961));
wire output_2_961, output_2_2, output_1_961;
mixer gate_output_1_961(.a(output_2_961), .b(output_2_2), .y(output_1_961));
wire output_3_961, output_3_2, output_2_961;
mixer gate_output_2_961(.a(output_3_961), .b(output_3_2), .y(output_2_961));
wire output_1_962, output_1_0, output_0_962;
mixer gate_output_0_962(.a(output_1_962), .b(output_1_0), .y(output_0_962));
wire output_2_962, output_2_0, output_1_962;
mixer gate_output_1_962(.a(output_2_962), .b(output_2_0), .y(output_1_962));
wire output_3_962, output_3_0, output_2_962;
mixer gate_output_2_962(.a(output_3_962), .b(output_3_0), .y(output_2_962));
wire output_1_963, output_1_1, output_0_963;
mixer gate_output_0_963(.a(output_1_963), .b(output_1_1), .y(output_0_963));
wire output_2_963, output_2_1, output_1_963;
mixer gate_output_1_963(.a(output_2_963), .b(output_2_1), .y(output_1_963));
wire output_3_963, output_3_1, output_2_963;
mixer gate_output_2_963(.a(output_3_963), .b(output_3_1), .y(output_2_963));
wire output_1_964, output_1_2, output_0_964;
mixer gate_output_0_964(.a(output_1_964), .b(output_1_2), .y(output_0_964));
wire output_2_964, output_2_2, output_1_964;
mixer gate_output_1_964(.a(output_2_964), .b(output_2_2), .y(output_1_964));
wire output_3_964, output_3_2, output_2_964;
mixer gate_output_2_964(.a(output_3_964), .b(output_3_2), .y(output_2_964));
wire output_1_965, output_1_0, output_0_965;
mixer gate_output_0_965(.a(output_1_965), .b(output_1_0), .y(output_0_965));
wire output_2_965, output_2_0, output_1_965;
mixer gate_output_1_965(.a(output_2_965), .b(output_2_0), .y(output_1_965));
wire output_3_965, output_3_0, output_2_965;
mixer gate_output_2_965(.a(output_3_965), .b(output_3_0), .y(output_2_965));
wire output_1_966, output_1_1, output_0_966;
mixer gate_output_0_966(.a(output_1_966), .b(output_1_1), .y(output_0_966));
wire output_2_966, output_2_1, output_1_966;
mixer gate_output_1_966(.a(output_2_966), .b(output_2_1), .y(output_1_966));
wire output_3_966, output_3_1, output_2_966;
mixer gate_output_2_966(.a(output_3_966), .b(output_3_1), .y(output_2_966));
wire output_1_967, output_1_2, output_0_967;
mixer gate_output_0_967(.a(output_1_967), .b(output_1_2), .y(output_0_967));
wire output_2_967, output_2_2, output_1_967;
mixer gate_output_1_967(.a(output_2_967), .b(output_2_2), .y(output_1_967));
wire output_3_967, output_3_2, output_2_967;
mixer gate_output_2_967(.a(output_3_967), .b(output_3_2), .y(output_2_967));
wire output_1_968, output_1_0, output_0_968;
mixer gate_output_0_968(.a(output_1_968), .b(output_1_0), .y(output_0_968));
wire output_2_968, output_2_0, output_1_968;
mixer gate_output_1_968(.a(output_2_968), .b(output_2_0), .y(output_1_968));
wire output_3_968, output_3_0, output_2_968;
mixer gate_output_2_968(.a(output_3_968), .b(output_3_0), .y(output_2_968));
wire output_1_969, output_1_1, output_0_969;
mixer gate_output_0_969(.a(output_1_969), .b(output_1_1), .y(output_0_969));
wire output_2_969, output_2_1, output_1_969;
mixer gate_output_1_969(.a(output_2_969), .b(output_2_1), .y(output_1_969));
wire output_3_969, output_3_1, output_2_969;
mixer gate_output_2_969(.a(output_3_969), .b(output_3_1), .y(output_2_969));
wire output_1_970, output_1_2, output_0_970;
mixer gate_output_0_970(.a(output_1_970), .b(output_1_2), .y(output_0_970));
wire output_2_970, output_2_2, output_1_970;
mixer gate_output_1_970(.a(output_2_970), .b(output_2_2), .y(output_1_970));
wire output_3_970, output_3_2, output_2_970;
mixer gate_output_2_970(.a(output_3_970), .b(output_3_2), .y(output_2_970));
wire output_1_971, output_1_0, output_0_971;
mixer gate_output_0_971(.a(output_1_971), .b(output_1_0), .y(output_0_971));
wire output_2_971, output_2_0, output_1_971;
mixer gate_output_1_971(.a(output_2_971), .b(output_2_0), .y(output_1_971));
wire output_3_971, output_3_0, output_2_971;
mixer gate_output_2_971(.a(output_3_971), .b(output_3_0), .y(output_2_971));
wire output_1_972, output_1_1, output_0_972;
mixer gate_output_0_972(.a(output_1_972), .b(output_1_1), .y(output_0_972));
wire output_2_972, output_2_1, output_1_972;
mixer gate_output_1_972(.a(output_2_972), .b(output_2_1), .y(output_1_972));
wire output_3_972, output_3_1, output_2_972;
mixer gate_output_2_972(.a(output_3_972), .b(output_3_1), .y(output_2_972));
wire output_1_973, output_1_2, output_0_973;
mixer gate_output_0_973(.a(output_1_973), .b(output_1_2), .y(output_0_973));
wire output_2_973, output_2_2, output_1_973;
mixer gate_output_1_973(.a(output_2_973), .b(output_2_2), .y(output_1_973));
wire output_3_973, output_3_2, output_2_973;
mixer gate_output_2_973(.a(output_3_973), .b(output_3_2), .y(output_2_973));
wire output_1_974, output_1_0, output_0_974;
mixer gate_output_0_974(.a(output_1_974), .b(output_1_0), .y(output_0_974));
wire output_2_974, output_2_0, output_1_974;
mixer gate_output_1_974(.a(output_2_974), .b(output_2_0), .y(output_1_974));
wire output_3_974, output_3_0, output_2_974;
mixer gate_output_2_974(.a(output_3_974), .b(output_3_0), .y(output_2_974));
wire output_1_975, output_1_1, output_0_975;
mixer gate_output_0_975(.a(output_1_975), .b(output_1_1), .y(output_0_975));
wire output_2_975, output_2_1, output_1_975;
mixer gate_output_1_975(.a(output_2_975), .b(output_2_1), .y(output_1_975));
wire output_3_975, output_3_1, output_2_975;
mixer gate_output_2_975(.a(output_3_975), .b(output_3_1), .y(output_2_975));
wire output_1_976, output_1_2, output_0_976;
mixer gate_output_0_976(.a(output_1_976), .b(output_1_2), .y(output_0_976));
wire output_2_976, output_2_2, output_1_976;
mixer gate_output_1_976(.a(output_2_976), .b(output_2_2), .y(output_1_976));
wire output_3_976, output_3_2, output_2_976;
mixer gate_output_2_976(.a(output_3_976), .b(output_3_2), .y(output_2_976));
wire output_1_977, output_1_0, output_0_977;
mixer gate_output_0_977(.a(output_1_977), .b(output_1_0), .y(output_0_977));
wire output_2_977, output_2_0, output_1_977;
mixer gate_output_1_977(.a(output_2_977), .b(output_2_0), .y(output_1_977));
wire output_3_977, output_3_0, output_2_977;
mixer gate_output_2_977(.a(output_3_977), .b(output_3_0), .y(output_2_977));
wire output_1_978, output_1_1, output_0_978;
mixer gate_output_0_978(.a(output_1_978), .b(output_1_1), .y(output_0_978));
wire output_2_978, output_2_1, output_1_978;
mixer gate_output_1_978(.a(output_2_978), .b(output_2_1), .y(output_1_978));
wire output_3_978, output_3_1, output_2_978;
mixer gate_output_2_978(.a(output_3_978), .b(output_3_1), .y(output_2_978));
wire output_1_979, output_1_2, output_0_979;
mixer gate_output_0_979(.a(output_1_979), .b(output_1_2), .y(output_0_979));
wire output_2_979, output_2_2, output_1_979;
mixer gate_output_1_979(.a(output_2_979), .b(output_2_2), .y(output_1_979));
wire output_3_979, output_3_2, output_2_979;
mixer gate_output_2_979(.a(output_3_979), .b(output_3_2), .y(output_2_979));
wire output_1_980, output_1_0, output_0_980;
mixer gate_output_0_980(.a(output_1_980), .b(output_1_0), .y(output_0_980));
wire output_2_980, output_2_0, output_1_980;
mixer gate_output_1_980(.a(output_2_980), .b(output_2_0), .y(output_1_980));
wire output_3_980, output_3_0, output_2_980;
mixer gate_output_2_980(.a(output_3_980), .b(output_3_0), .y(output_2_980));
wire output_1_981, output_1_1, output_0_981;
mixer gate_output_0_981(.a(output_1_981), .b(output_1_1), .y(output_0_981));
wire output_2_981, output_2_1, output_1_981;
mixer gate_output_1_981(.a(output_2_981), .b(output_2_1), .y(output_1_981));
wire output_3_981, output_3_1, output_2_981;
mixer gate_output_2_981(.a(output_3_981), .b(output_3_1), .y(output_2_981));
wire output_1_982, output_1_2, output_0_982;
mixer gate_output_0_982(.a(output_1_982), .b(output_1_2), .y(output_0_982));
wire output_2_982, output_2_2, output_1_982;
mixer gate_output_1_982(.a(output_2_982), .b(output_2_2), .y(output_1_982));
wire output_3_982, output_3_2, output_2_982;
mixer gate_output_2_982(.a(output_3_982), .b(output_3_2), .y(output_2_982));
wire output_1_983, output_1_0, output_0_983;
mixer gate_output_0_983(.a(output_1_983), .b(output_1_0), .y(output_0_983));
wire output_2_983, output_2_0, output_1_983;
mixer gate_output_1_983(.a(output_2_983), .b(output_2_0), .y(output_1_983));
wire output_3_983, output_3_0, output_2_983;
mixer gate_output_2_983(.a(output_3_983), .b(output_3_0), .y(output_2_983));
wire output_1_984, output_1_1, output_0_984;
mixer gate_output_0_984(.a(output_1_984), .b(output_1_1), .y(output_0_984));
wire output_2_984, output_2_1, output_1_984;
mixer gate_output_1_984(.a(output_2_984), .b(output_2_1), .y(output_1_984));
wire output_3_984, output_3_1, output_2_984;
mixer gate_output_2_984(.a(output_3_984), .b(output_3_1), .y(output_2_984));
wire output_1_985, output_1_2, output_0_985;
mixer gate_output_0_985(.a(output_1_985), .b(output_1_2), .y(output_0_985));
wire output_2_985, output_2_2, output_1_985;
mixer gate_output_1_985(.a(output_2_985), .b(output_2_2), .y(output_1_985));
wire output_3_985, output_3_2, output_2_985;
mixer gate_output_2_985(.a(output_3_985), .b(output_3_2), .y(output_2_985));
wire output_1_986, output_1_0, output_0_986;
mixer gate_output_0_986(.a(output_1_986), .b(output_1_0), .y(output_0_986));
wire output_2_986, output_2_0, output_1_986;
mixer gate_output_1_986(.a(output_2_986), .b(output_2_0), .y(output_1_986));
wire output_3_986, output_3_0, output_2_986;
mixer gate_output_2_986(.a(output_3_986), .b(output_3_0), .y(output_2_986));
wire output_1_987, output_1_1, output_0_987;
mixer gate_output_0_987(.a(output_1_987), .b(output_1_1), .y(output_0_987));
wire output_2_987, output_2_1, output_1_987;
mixer gate_output_1_987(.a(output_2_987), .b(output_2_1), .y(output_1_987));
wire output_3_987, output_3_1, output_2_987;
mixer gate_output_2_987(.a(output_3_987), .b(output_3_1), .y(output_2_987));
wire output_1_988, output_1_2, output_0_988;
mixer gate_output_0_988(.a(output_1_988), .b(output_1_2), .y(output_0_988));
wire output_2_988, output_2_2, output_1_988;
mixer gate_output_1_988(.a(output_2_988), .b(output_2_2), .y(output_1_988));
wire output_3_988, output_3_2, output_2_988;
mixer gate_output_2_988(.a(output_3_988), .b(output_3_2), .y(output_2_988));
wire output_1_989, output_1_0, output_0_989;
mixer gate_output_0_989(.a(output_1_989), .b(output_1_0), .y(output_0_989));
wire output_2_989, output_2_0, output_1_989;
mixer gate_output_1_989(.a(output_2_989), .b(output_2_0), .y(output_1_989));
wire output_3_989, output_3_0, output_2_989;
mixer gate_output_2_989(.a(output_3_989), .b(output_3_0), .y(output_2_989));
wire output_1_990, output_1_1, output_0_990;
mixer gate_output_0_990(.a(output_1_990), .b(output_1_1), .y(output_0_990));
wire output_2_990, output_2_1, output_1_990;
mixer gate_output_1_990(.a(output_2_990), .b(output_2_1), .y(output_1_990));
wire output_3_990, output_3_1, output_2_990;
mixer gate_output_2_990(.a(output_3_990), .b(output_3_1), .y(output_2_990));
wire output_1_991, output_1_2, output_0_991;
mixer gate_output_0_991(.a(output_1_991), .b(output_1_2), .y(output_0_991));
wire output_2_991, output_2_2, output_1_991;
mixer gate_output_1_991(.a(output_2_991), .b(output_2_2), .y(output_1_991));
wire output_3_991, output_3_2, output_2_991;
mixer gate_output_2_991(.a(output_3_991), .b(output_3_2), .y(output_2_991));
wire output_1_992, output_1_0, output_0_992;
mixer gate_output_0_992(.a(output_1_992), .b(output_1_0), .y(output_0_992));
wire output_2_992, output_2_0, output_1_992;
mixer gate_output_1_992(.a(output_2_992), .b(output_2_0), .y(output_1_992));
wire output_3_992, output_3_0, output_2_992;
mixer gate_output_2_992(.a(output_3_992), .b(output_3_0), .y(output_2_992));
wire output_1_993, output_1_1, output_0_993;
mixer gate_output_0_993(.a(output_1_993), .b(output_1_1), .y(output_0_993));
wire output_2_993, output_2_1, output_1_993;
mixer gate_output_1_993(.a(output_2_993), .b(output_2_1), .y(output_1_993));
wire output_3_993, output_3_1, output_2_993;
mixer gate_output_2_993(.a(output_3_993), .b(output_3_1), .y(output_2_993));
wire output_1_994, output_1_2, output_0_994;
mixer gate_output_0_994(.a(output_1_994), .b(output_1_2), .y(output_0_994));
wire output_2_994, output_2_2, output_1_994;
mixer gate_output_1_994(.a(output_2_994), .b(output_2_2), .y(output_1_994));
wire output_3_994, output_3_2, output_2_994;
mixer gate_output_2_994(.a(output_3_994), .b(output_3_2), .y(output_2_994));
wire output_1_995, output_1_0, output_0_995;
mixer gate_output_0_995(.a(output_1_995), .b(output_1_0), .y(output_0_995));
wire output_2_995, output_2_0, output_1_995;
mixer gate_output_1_995(.a(output_2_995), .b(output_2_0), .y(output_1_995));
wire output_3_995, output_3_0, output_2_995;
mixer gate_output_2_995(.a(output_3_995), .b(output_3_0), .y(output_2_995));
wire output_1_996, output_1_1, output_0_996;
mixer gate_output_0_996(.a(output_1_996), .b(output_1_1), .y(output_0_996));
wire output_2_996, output_2_1, output_1_996;
mixer gate_output_1_996(.a(output_2_996), .b(output_2_1), .y(output_1_996));
wire output_3_996, output_3_1, output_2_996;
mixer gate_output_2_996(.a(output_3_996), .b(output_3_1), .y(output_2_996));
wire output_1_997, output_1_2, output_0_997;
mixer gate_output_0_997(.a(output_1_997), .b(output_1_2), .y(output_0_997));
wire output_2_997, output_2_2, output_1_997;
mixer gate_output_1_997(.a(output_2_997), .b(output_2_2), .y(output_1_997));
wire output_3_997, output_3_2, output_2_997;
mixer gate_output_2_997(.a(output_3_997), .b(output_3_2), .y(output_2_997));
wire output_1_998, output_1_0, output_0_998;
mixer gate_output_0_998(.a(output_1_998), .b(output_1_0), .y(output_0_998));
wire output_2_998, output_2_0, output_1_998;
mixer gate_output_1_998(.a(output_2_998), .b(output_2_0), .y(output_1_998));
wire output_3_998, output_3_0, output_2_998;
mixer gate_output_2_998(.a(output_3_998), .b(output_3_0), .y(output_2_998));
wire output_1_999, output_1_1, output_0_999;
mixer gate_output_0_999(.a(output_1_999), .b(output_1_1), .y(output_0_999));
wire output_2_999, output_2_1, output_1_999;
mixer gate_output_1_999(.a(output_2_999), .b(output_2_1), .y(output_1_999));
wire output_3_999, output_3_1, output_2_999;
mixer gate_output_2_999(.a(output_3_999), .b(output_3_1), .y(output_2_999));
wire output_1_1000, output_1_2, output_0_1000;
mixer gate_output_0_1000(.a(output_1_1000), .b(output_1_2), .y(output_0_1000));
wire output_2_1000, output_2_2, output_1_1000;
mixer gate_output_1_1000(.a(output_2_1000), .b(output_2_2), .y(output_1_1000));
wire output_3_1000, output_3_2, output_2_1000;
mixer gate_output_2_1000(.a(output_3_1000), .b(output_3_2), .y(output_2_1000));
wire output_1_1001, output_1_0, output_0_1001;
mixer gate_output_0_1001(.a(output_1_1001), .b(output_1_0), .y(output_0_1001));
wire output_2_1001, output_2_0, output_1_1001;
mixer gate_output_1_1001(.a(output_2_1001), .b(output_2_0), .y(output_1_1001));
wire output_3_1001, output_3_0, output_2_1001;
mixer gate_output_2_1001(.a(output_3_1001), .b(output_3_0), .y(output_2_1001));
wire output_1_1002, output_1_1, output_0_1002;
mixer gate_output_0_1002(.a(output_1_1002), .b(output_1_1), .y(output_0_1002));
wire output_2_1002, output_2_1, output_1_1002;
mixer gate_output_1_1002(.a(output_2_1002), .b(output_2_1), .y(output_1_1002));
wire output_3_1002, output_3_1, output_2_1002;
mixer gate_output_2_1002(.a(output_3_1002), .b(output_3_1), .y(output_2_1002));
wire output_1_1003, output_1_2, output_0_1003;
mixer gate_output_0_1003(.a(output_1_1003), .b(output_1_2), .y(output_0_1003));
wire output_2_1003, output_2_2, output_1_1003;
mixer gate_output_1_1003(.a(output_2_1003), .b(output_2_2), .y(output_1_1003));
wire output_3_1003, output_3_2, output_2_1003;
mixer gate_output_2_1003(.a(output_3_1003), .b(output_3_2), .y(output_2_1003));
wire output_1_1004, output_1_0, output_0_1004;
mixer gate_output_0_1004(.a(output_1_1004), .b(output_1_0), .y(output_0_1004));
wire output_2_1004, output_2_0, output_1_1004;
mixer gate_output_1_1004(.a(output_2_1004), .b(output_2_0), .y(output_1_1004));
wire output_3_1004, output_3_0, output_2_1004;
mixer gate_output_2_1004(.a(output_3_1004), .b(output_3_0), .y(output_2_1004));
wire output_1_1005, output_1_1, output_0_1005;
mixer gate_output_0_1005(.a(output_1_1005), .b(output_1_1), .y(output_0_1005));
wire output_2_1005, output_2_1, output_1_1005;
mixer gate_output_1_1005(.a(output_2_1005), .b(output_2_1), .y(output_1_1005));
wire output_3_1005, output_3_1, output_2_1005;
mixer gate_output_2_1005(.a(output_3_1005), .b(output_3_1), .y(output_2_1005));
wire output_1_1006, output_1_2, output_0_1006;
mixer gate_output_0_1006(.a(output_1_1006), .b(output_1_2), .y(output_0_1006));
wire output_2_1006, output_2_2, output_1_1006;
mixer gate_output_1_1006(.a(output_2_1006), .b(output_2_2), .y(output_1_1006));
wire output_3_1006, output_3_2, output_2_1006;
mixer gate_output_2_1006(.a(output_3_1006), .b(output_3_2), .y(output_2_1006));
wire output_1_1007, output_1_0, output_0_1007;
mixer gate_output_0_1007(.a(output_1_1007), .b(output_1_0), .y(output_0_1007));
wire output_2_1007, output_2_0, output_1_1007;
mixer gate_output_1_1007(.a(output_2_1007), .b(output_2_0), .y(output_1_1007));
wire output_3_1007, output_3_0, output_2_1007;
mixer gate_output_2_1007(.a(output_3_1007), .b(output_3_0), .y(output_2_1007));
wire output_1_1008, output_1_1, output_0_1008;
mixer gate_output_0_1008(.a(output_1_1008), .b(output_1_1), .y(output_0_1008));
wire output_2_1008, output_2_1, output_1_1008;
mixer gate_output_1_1008(.a(output_2_1008), .b(output_2_1), .y(output_1_1008));
wire output_3_1008, output_3_1, output_2_1008;
mixer gate_output_2_1008(.a(output_3_1008), .b(output_3_1), .y(output_2_1008));
wire output_1_1009, output_1_2, output_0_1009;
mixer gate_output_0_1009(.a(output_1_1009), .b(output_1_2), .y(output_0_1009));
wire output_2_1009, output_2_2, output_1_1009;
mixer gate_output_1_1009(.a(output_2_1009), .b(output_2_2), .y(output_1_1009));
wire output_3_1009, output_3_2, output_2_1009;
mixer gate_output_2_1009(.a(output_3_1009), .b(output_3_2), .y(output_2_1009));
wire output_1_1010, output_1_0, output_0_1010;
mixer gate_output_0_1010(.a(output_1_1010), .b(output_1_0), .y(output_0_1010));
wire output_2_1010, output_2_0, output_1_1010;
mixer gate_output_1_1010(.a(output_2_1010), .b(output_2_0), .y(output_1_1010));
wire output_3_1010, output_3_0, output_2_1010;
mixer gate_output_2_1010(.a(output_3_1010), .b(output_3_0), .y(output_2_1010));
wire output_1_1011, output_1_1, output_0_1011;
mixer gate_output_0_1011(.a(output_1_1011), .b(output_1_1), .y(output_0_1011));
wire output_2_1011, output_2_1, output_1_1011;
mixer gate_output_1_1011(.a(output_2_1011), .b(output_2_1), .y(output_1_1011));
wire output_3_1011, output_3_1, output_2_1011;
mixer gate_output_2_1011(.a(output_3_1011), .b(output_3_1), .y(output_2_1011));
wire output_1_1012, output_1_2, output_0_1012;
mixer gate_output_0_1012(.a(output_1_1012), .b(output_1_2), .y(output_0_1012));
wire output_2_1012, output_2_2, output_1_1012;
mixer gate_output_1_1012(.a(output_2_1012), .b(output_2_2), .y(output_1_1012));
wire output_3_1012, output_3_2, output_2_1012;
mixer gate_output_2_1012(.a(output_3_1012), .b(output_3_2), .y(output_2_1012));
wire output_1_1013, output_1_0, output_0_1013;
mixer gate_output_0_1013(.a(output_1_1013), .b(output_1_0), .y(output_0_1013));
wire output_2_1013, output_2_0, output_1_1013;
mixer gate_output_1_1013(.a(output_2_1013), .b(output_2_0), .y(output_1_1013));
wire output_3_1013, output_3_0, output_2_1013;
mixer gate_output_2_1013(.a(output_3_1013), .b(output_3_0), .y(output_2_1013));
wire output_1_1014, output_1_1, output_0_1014;
mixer gate_output_0_1014(.a(output_1_1014), .b(output_1_1), .y(output_0_1014));
wire output_2_1014, output_2_1, output_1_1014;
mixer gate_output_1_1014(.a(output_2_1014), .b(output_2_1), .y(output_1_1014));
wire output_3_1014, output_3_1, output_2_1014;
mixer gate_output_2_1014(.a(output_3_1014), .b(output_3_1), .y(output_2_1014));
wire output_1_1015, output_1_2, output_0_1015;
mixer gate_output_0_1015(.a(output_1_1015), .b(output_1_2), .y(output_0_1015));
wire output_2_1015, output_2_2, output_1_1015;
mixer gate_output_1_1015(.a(output_2_1015), .b(output_2_2), .y(output_1_1015));
wire output_3_1015, output_3_2, output_2_1015;
mixer gate_output_2_1015(.a(output_3_1015), .b(output_3_2), .y(output_2_1015));
wire output_1_1016, output_1_0, output_0_1016;
mixer gate_output_0_1016(.a(output_1_1016), .b(output_1_0), .y(output_0_1016));
wire output_2_1016, output_2_0, output_1_1016;
mixer gate_output_1_1016(.a(output_2_1016), .b(output_2_0), .y(output_1_1016));
wire output_3_1016, output_3_0, output_2_1016;
mixer gate_output_2_1016(.a(output_3_1016), .b(output_3_0), .y(output_2_1016));
wire output_1_1017, output_1_1, output_0_1017;
mixer gate_output_0_1017(.a(output_1_1017), .b(output_1_1), .y(output_0_1017));
wire output_2_1017, output_2_1, output_1_1017;
mixer gate_output_1_1017(.a(output_2_1017), .b(output_2_1), .y(output_1_1017));
wire output_3_1017, output_3_1, output_2_1017;
mixer gate_output_2_1017(.a(output_3_1017), .b(output_3_1), .y(output_2_1017));
wire output_1_1018, output_1_2, output_0_1018;
mixer gate_output_0_1018(.a(output_1_1018), .b(output_1_2), .y(output_0_1018));
wire output_2_1018, output_2_2, output_1_1018;
mixer gate_output_1_1018(.a(output_2_1018), .b(output_2_2), .y(output_1_1018));
wire output_3_1018, output_3_2, output_2_1018;
mixer gate_output_2_1018(.a(output_3_1018), .b(output_3_2), .y(output_2_1018));
wire output_1_1019, output_1_0, output_0_1019;
mixer gate_output_0_1019(.a(output_1_1019), .b(output_1_0), .y(output_0_1019));
wire output_2_1019, output_2_0, output_1_1019;
mixer gate_output_1_1019(.a(output_2_1019), .b(output_2_0), .y(output_1_1019));
wire output_3_1019, output_3_0, output_2_1019;
mixer gate_output_2_1019(.a(output_3_1019), .b(output_3_0), .y(output_2_1019));
wire output_1_1020, output_1_1, output_0_1020;
mixer gate_output_0_1020(.a(output_1_1020), .b(output_1_1), .y(output_0_1020));
wire output_2_1020, output_2_1, output_1_1020;
mixer gate_output_1_1020(.a(output_2_1020), .b(output_2_1), .y(output_1_1020));
wire output_3_1020, output_3_1, output_2_1020;
mixer gate_output_2_1020(.a(output_3_1020), .b(output_3_1), .y(output_2_1020));
wire output_1_1021, output_1_2, output_0_1021;
mixer gate_output_0_1021(.a(output_1_1021), .b(output_1_2), .y(output_0_1021));
wire output_2_1021, output_2_2, output_1_1021;
mixer gate_output_1_1021(.a(output_2_1021), .b(output_2_2), .y(output_1_1021));
wire output_3_1021, output_3_2, output_2_1021;
mixer gate_output_2_1021(.a(output_3_1021), .b(output_3_2), .y(output_2_1021));
wire output_1_1022, output_1_0, output_0_1022;
mixer gate_output_0_1022(.a(output_1_1022), .b(output_1_0), .y(output_0_1022));
wire output_2_1022, output_2_0, output_1_1022;
mixer gate_output_1_1022(.a(output_2_1022), .b(output_2_0), .y(output_1_1022));
wire output_3_1022, output_3_0, output_2_1022;
mixer gate_output_2_1022(.a(output_3_1022), .b(output_3_0), .y(output_2_1022));
wire output_1_1023, output_1_1, output_0_1023;
mixer gate_output_0_1023(.a(output_1_1023), .b(output_1_1), .y(output_0_1023));
wire output_2_1023, output_2_1, output_1_1023;
mixer gate_output_1_1023(.a(output_2_1023), .b(output_2_1), .y(output_1_1023));
wire output_3_1023, output_3_1, output_2_1023;
mixer gate_output_2_1023(.a(output_3_1023), .b(output_3_1), .y(output_2_1023));
assign output_0 = output_0_0;
wire output_0_1024;
assign output_0_1024 = input_0;
assign output_1 = output_1_0;
wire output_1_1024;
assign output_1_1024 = input_1;
assign output_2 = output_2_0;
wire output_2_1024;
assign output_2_1024 = input_2;
endmodule
