module rotary_cells (
inout pb1_1, pb1_2, pb1_3, pb1_4, p1, cb1_1, cb1_2, cb2_1, cb2_2, cb3_1, cb3_2, cb3_3, cb4_1, cb4_2, cb5_1, cb5_2, cb6_1, cb6_2
);
wire c1;
wire c2;
wire c3;
wire c4;
wire c5;
wire c6;
wire c7;
wire c8;
wire c9;
wire c10;
wire c11;
wire c12;
wire c13;
wire c14;
wire c15;
wire cc1;
wire cc2;
wire cc3;
wire cc4;
wire cc5;
wire cc6;
wire cc7;
wire cc8;
wire cc9;
wire cc10;
wire cc11;
wire cc12;
wire cc13;
MUX m1(.port5(c5),.port6(cc1),.port8(cc2),.port7(cc8),.port9(cc9),.port1(c1),.port2(c2),.port3(c3),.port4(c4));
MUX m2(.port2(c7),.port3(c8),.port4(c9),.port5(c10),.port7(cc6),.port9(cc7),.port6(cc12),.port8(cc13),.port1(c6));
assign c1 = pb1_1;
assign c2 = pb1_2;
assign c3 = pb1_3;
assign c4 = pb1_4;
ROTARY_MIXER rp(.port2(c6),.port3(cc3),.port6(cc4),.port7(cc5),.port4(cc10),.port5(cc11),.port1(c5));
LONG_CELL_TRAP b1_1(.port0(c11),.port0(c7));
LONG_CELL_TRAP b1_2(.port0(c12),.port0(c8));
LONG_CELL_TRAP b1_3(.port0(c13),.port0(c9));
LONG_CELL_TRAP b1_4(.port0(c14),.port0(c10));
TREE t1(.port1(c15),.port5(c11),.port4(c12),.port3(c13),.port2(c14));
assign c15 = p1;
assign cc1 = cb1_1;
assign cc2 = cb1_2;
assign cc8 = cb2_1;
assign cc9 = cb2_2;
assign cc3 = cb3_1;
assign cc4 = cb3_2;
assign cc5 = cb3_3;
assign cc10 = cb4_1;
assign cc11 = cb4_2;
assign cc6 = cb5_1;
assign cc7 = cb5_2;
assign cc12 = cb6_1;
assign cc13 = cb6_2;
endmodule
