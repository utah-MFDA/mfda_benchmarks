module fanout2_braid_16_256 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,output output_8,output output_9,output output_10,output output_11,output output_12,output output_13,output output_14,output output_15,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_9_0, output_9_1, output_8_0;
mixer gate_output_8_0(.a(output_9_0), .b(output_9_1), .y(output_8_0));
wire output_10_0, output_10_1, output_9_0;
mixer gate_output_9_0(.a(output_10_0), .b(output_10_1), .y(output_9_0));
wire output_11_0, output_11_1, output_10_0;
mixer gate_output_10_0(.a(output_11_0), .b(output_11_1), .y(output_10_0));
wire output_12_0, output_12_1, output_11_0;
mixer gate_output_11_0(.a(output_12_0), .b(output_12_1), .y(output_11_0));
wire output_13_0, output_13_1, output_12_0;
mixer gate_output_12_0(.a(output_13_0), .b(output_13_1), .y(output_12_0));
wire output_14_0, output_14_1, output_13_0;
mixer gate_output_13_0(.a(output_14_0), .b(output_14_1), .y(output_13_0));
wire output_15_0, output_15_1, output_14_0;
mixer gate_output_14_0(.a(output_15_0), .b(output_15_1), .y(output_14_0));
wire output_16_0, output_16_1, output_15_0;
mixer gate_output_15_0(.a(output_16_0), .b(output_16_1), .y(output_15_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_9_1, output_9_2, output_8_1;
mixer gate_output_8_1(.a(output_9_1), .b(output_9_2), .y(output_8_1));
wire output_10_1, output_10_2, output_9_1;
mixer gate_output_9_1(.a(output_10_1), .b(output_10_2), .y(output_9_1));
wire output_11_1, output_11_2, output_10_1;
mixer gate_output_10_1(.a(output_11_1), .b(output_11_2), .y(output_10_1));
wire output_12_1, output_12_2, output_11_1;
mixer gate_output_11_1(.a(output_12_1), .b(output_12_2), .y(output_11_1));
wire output_13_1, output_13_2, output_12_1;
mixer gate_output_12_1(.a(output_13_1), .b(output_13_2), .y(output_12_1));
wire output_14_1, output_14_2, output_13_1;
mixer gate_output_13_1(.a(output_14_1), .b(output_14_2), .y(output_13_1));
wire output_15_1, output_15_2, output_14_1;
mixer gate_output_14_1(.a(output_15_1), .b(output_15_2), .y(output_14_1));
wire output_16_1, output_16_2, output_15_1;
mixer gate_output_15_1(.a(output_16_1), .b(output_16_2), .y(output_15_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_9_2, output_9_3, output_8_2;
mixer gate_output_8_2(.a(output_9_2), .b(output_9_3), .y(output_8_2));
wire output_10_2, output_10_3, output_9_2;
mixer gate_output_9_2(.a(output_10_2), .b(output_10_3), .y(output_9_2));
wire output_11_2, output_11_3, output_10_2;
mixer gate_output_10_2(.a(output_11_2), .b(output_11_3), .y(output_10_2));
wire output_12_2, output_12_3, output_11_2;
mixer gate_output_11_2(.a(output_12_2), .b(output_12_3), .y(output_11_2));
wire output_13_2, output_13_3, output_12_2;
mixer gate_output_12_2(.a(output_13_2), .b(output_13_3), .y(output_12_2));
wire output_14_2, output_14_3, output_13_2;
mixer gate_output_13_2(.a(output_14_2), .b(output_14_3), .y(output_13_2));
wire output_15_2, output_15_3, output_14_2;
mixer gate_output_14_2(.a(output_15_2), .b(output_15_3), .y(output_14_2));
wire output_16_2, output_16_3, output_15_2;
mixer gate_output_15_2(.a(output_16_2), .b(output_16_3), .y(output_15_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_9_3, output_9_4, output_8_3;
mixer gate_output_8_3(.a(output_9_3), .b(output_9_4), .y(output_8_3));
wire output_10_3, output_10_4, output_9_3;
mixer gate_output_9_3(.a(output_10_3), .b(output_10_4), .y(output_9_3));
wire output_11_3, output_11_4, output_10_3;
mixer gate_output_10_3(.a(output_11_3), .b(output_11_4), .y(output_10_3));
wire output_12_3, output_12_4, output_11_3;
mixer gate_output_11_3(.a(output_12_3), .b(output_12_4), .y(output_11_3));
wire output_13_3, output_13_4, output_12_3;
mixer gate_output_12_3(.a(output_13_3), .b(output_13_4), .y(output_12_3));
wire output_14_3, output_14_4, output_13_3;
mixer gate_output_13_3(.a(output_14_3), .b(output_14_4), .y(output_13_3));
wire output_15_3, output_15_4, output_14_3;
mixer gate_output_14_3(.a(output_15_3), .b(output_15_4), .y(output_14_3));
wire output_16_3, output_16_4, output_15_3;
mixer gate_output_15_3(.a(output_16_3), .b(output_16_4), .y(output_15_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_9_4, output_9_5, output_8_4;
mixer gate_output_8_4(.a(output_9_4), .b(output_9_5), .y(output_8_4));
wire output_10_4, output_10_5, output_9_4;
mixer gate_output_9_4(.a(output_10_4), .b(output_10_5), .y(output_9_4));
wire output_11_4, output_11_5, output_10_4;
mixer gate_output_10_4(.a(output_11_4), .b(output_11_5), .y(output_10_4));
wire output_12_4, output_12_5, output_11_4;
mixer gate_output_11_4(.a(output_12_4), .b(output_12_5), .y(output_11_4));
wire output_13_4, output_13_5, output_12_4;
mixer gate_output_12_4(.a(output_13_4), .b(output_13_5), .y(output_12_4));
wire output_14_4, output_14_5, output_13_4;
mixer gate_output_13_4(.a(output_14_4), .b(output_14_5), .y(output_13_4));
wire output_15_4, output_15_5, output_14_4;
mixer gate_output_14_4(.a(output_15_4), .b(output_15_5), .y(output_14_4));
wire output_16_4, output_16_5, output_15_4;
mixer gate_output_15_4(.a(output_16_4), .b(output_16_5), .y(output_15_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_9_5, output_9_6, output_8_5;
mixer gate_output_8_5(.a(output_9_5), .b(output_9_6), .y(output_8_5));
wire output_10_5, output_10_6, output_9_5;
mixer gate_output_9_5(.a(output_10_5), .b(output_10_6), .y(output_9_5));
wire output_11_5, output_11_6, output_10_5;
mixer gate_output_10_5(.a(output_11_5), .b(output_11_6), .y(output_10_5));
wire output_12_5, output_12_6, output_11_5;
mixer gate_output_11_5(.a(output_12_5), .b(output_12_6), .y(output_11_5));
wire output_13_5, output_13_6, output_12_5;
mixer gate_output_12_5(.a(output_13_5), .b(output_13_6), .y(output_12_5));
wire output_14_5, output_14_6, output_13_5;
mixer gate_output_13_5(.a(output_14_5), .b(output_14_6), .y(output_13_5));
wire output_15_5, output_15_6, output_14_5;
mixer gate_output_14_5(.a(output_15_5), .b(output_15_6), .y(output_14_5));
wire output_16_5, output_16_6, output_15_5;
mixer gate_output_15_5(.a(output_16_5), .b(output_16_6), .y(output_15_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_9_6, output_9_7, output_8_6;
mixer gate_output_8_6(.a(output_9_6), .b(output_9_7), .y(output_8_6));
wire output_10_6, output_10_7, output_9_6;
mixer gate_output_9_6(.a(output_10_6), .b(output_10_7), .y(output_9_6));
wire output_11_6, output_11_7, output_10_6;
mixer gate_output_10_6(.a(output_11_6), .b(output_11_7), .y(output_10_6));
wire output_12_6, output_12_7, output_11_6;
mixer gate_output_11_6(.a(output_12_6), .b(output_12_7), .y(output_11_6));
wire output_13_6, output_13_7, output_12_6;
mixer gate_output_12_6(.a(output_13_6), .b(output_13_7), .y(output_12_6));
wire output_14_6, output_14_7, output_13_6;
mixer gate_output_13_6(.a(output_14_6), .b(output_14_7), .y(output_13_6));
wire output_15_6, output_15_7, output_14_6;
mixer gate_output_14_6(.a(output_15_6), .b(output_15_7), .y(output_14_6));
wire output_16_6, output_16_7, output_15_6;
mixer gate_output_15_6(.a(output_16_6), .b(output_16_7), .y(output_15_6));
wire output_1_7, output_1_8, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_8), .y(output_0_7));
wire output_2_7, output_2_8, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_8), .y(output_1_7));
wire output_3_7, output_3_8, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_8), .y(output_2_7));
wire output_4_7, output_4_8, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_8), .y(output_3_7));
wire output_5_7, output_5_8, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_8), .y(output_4_7));
wire output_6_7, output_6_8, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_8), .y(output_5_7));
wire output_7_7, output_7_8, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_8), .y(output_6_7));
wire output_8_7, output_8_8, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_8), .y(output_7_7));
wire output_9_7, output_9_8, output_8_7;
mixer gate_output_8_7(.a(output_9_7), .b(output_9_8), .y(output_8_7));
wire output_10_7, output_10_8, output_9_7;
mixer gate_output_9_7(.a(output_10_7), .b(output_10_8), .y(output_9_7));
wire output_11_7, output_11_8, output_10_7;
mixer gate_output_10_7(.a(output_11_7), .b(output_11_8), .y(output_10_7));
wire output_12_7, output_12_8, output_11_7;
mixer gate_output_11_7(.a(output_12_7), .b(output_12_8), .y(output_11_7));
wire output_13_7, output_13_8, output_12_7;
mixer gate_output_12_7(.a(output_13_7), .b(output_13_8), .y(output_12_7));
wire output_14_7, output_14_8, output_13_7;
mixer gate_output_13_7(.a(output_14_7), .b(output_14_8), .y(output_13_7));
wire output_15_7, output_15_8, output_14_7;
mixer gate_output_14_7(.a(output_15_7), .b(output_15_8), .y(output_14_7));
wire output_16_7, output_16_8, output_15_7;
mixer gate_output_15_7(.a(output_16_7), .b(output_16_8), .y(output_15_7));
wire output_1_8, output_1_9, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_9), .y(output_0_8));
wire output_2_8, output_2_9, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_9), .y(output_1_8));
wire output_3_8, output_3_9, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_9), .y(output_2_8));
wire output_4_8, output_4_9, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_9), .y(output_3_8));
wire output_5_8, output_5_9, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_9), .y(output_4_8));
wire output_6_8, output_6_9, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_9), .y(output_5_8));
wire output_7_8, output_7_9, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_9), .y(output_6_8));
wire output_8_8, output_8_9, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_9), .y(output_7_8));
wire output_9_8, output_9_9, output_8_8;
mixer gate_output_8_8(.a(output_9_8), .b(output_9_9), .y(output_8_8));
wire output_10_8, output_10_9, output_9_8;
mixer gate_output_9_8(.a(output_10_8), .b(output_10_9), .y(output_9_8));
wire output_11_8, output_11_9, output_10_8;
mixer gate_output_10_8(.a(output_11_8), .b(output_11_9), .y(output_10_8));
wire output_12_8, output_12_9, output_11_8;
mixer gate_output_11_8(.a(output_12_8), .b(output_12_9), .y(output_11_8));
wire output_13_8, output_13_9, output_12_8;
mixer gate_output_12_8(.a(output_13_8), .b(output_13_9), .y(output_12_8));
wire output_14_8, output_14_9, output_13_8;
mixer gate_output_13_8(.a(output_14_8), .b(output_14_9), .y(output_13_8));
wire output_15_8, output_15_9, output_14_8;
mixer gate_output_14_8(.a(output_15_8), .b(output_15_9), .y(output_14_8));
wire output_16_8, output_16_9, output_15_8;
mixer gate_output_15_8(.a(output_16_8), .b(output_16_9), .y(output_15_8));
wire output_1_9, output_1_10, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_10), .y(output_0_9));
wire output_2_9, output_2_10, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_10), .y(output_1_9));
wire output_3_9, output_3_10, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_10), .y(output_2_9));
wire output_4_9, output_4_10, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_10), .y(output_3_9));
wire output_5_9, output_5_10, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_10), .y(output_4_9));
wire output_6_9, output_6_10, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_10), .y(output_5_9));
wire output_7_9, output_7_10, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_10), .y(output_6_9));
wire output_8_9, output_8_10, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_10), .y(output_7_9));
wire output_9_9, output_9_10, output_8_9;
mixer gate_output_8_9(.a(output_9_9), .b(output_9_10), .y(output_8_9));
wire output_10_9, output_10_10, output_9_9;
mixer gate_output_9_9(.a(output_10_9), .b(output_10_10), .y(output_9_9));
wire output_11_9, output_11_10, output_10_9;
mixer gate_output_10_9(.a(output_11_9), .b(output_11_10), .y(output_10_9));
wire output_12_9, output_12_10, output_11_9;
mixer gate_output_11_9(.a(output_12_9), .b(output_12_10), .y(output_11_9));
wire output_13_9, output_13_10, output_12_9;
mixer gate_output_12_9(.a(output_13_9), .b(output_13_10), .y(output_12_9));
wire output_14_9, output_14_10, output_13_9;
mixer gate_output_13_9(.a(output_14_9), .b(output_14_10), .y(output_13_9));
wire output_15_9, output_15_10, output_14_9;
mixer gate_output_14_9(.a(output_15_9), .b(output_15_10), .y(output_14_9));
wire output_16_9, output_16_10, output_15_9;
mixer gate_output_15_9(.a(output_16_9), .b(output_16_10), .y(output_15_9));
wire output_1_10, output_1_11, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_11), .y(output_0_10));
wire output_2_10, output_2_11, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_11), .y(output_1_10));
wire output_3_10, output_3_11, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_11), .y(output_2_10));
wire output_4_10, output_4_11, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_11), .y(output_3_10));
wire output_5_10, output_5_11, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_11), .y(output_4_10));
wire output_6_10, output_6_11, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_11), .y(output_5_10));
wire output_7_10, output_7_11, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_11), .y(output_6_10));
wire output_8_10, output_8_11, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_11), .y(output_7_10));
wire output_9_10, output_9_11, output_8_10;
mixer gate_output_8_10(.a(output_9_10), .b(output_9_11), .y(output_8_10));
wire output_10_10, output_10_11, output_9_10;
mixer gate_output_9_10(.a(output_10_10), .b(output_10_11), .y(output_9_10));
wire output_11_10, output_11_11, output_10_10;
mixer gate_output_10_10(.a(output_11_10), .b(output_11_11), .y(output_10_10));
wire output_12_10, output_12_11, output_11_10;
mixer gate_output_11_10(.a(output_12_10), .b(output_12_11), .y(output_11_10));
wire output_13_10, output_13_11, output_12_10;
mixer gate_output_12_10(.a(output_13_10), .b(output_13_11), .y(output_12_10));
wire output_14_10, output_14_11, output_13_10;
mixer gate_output_13_10(.a(output_14_10), .b(output_14_11), .y(output_13_10));
wire output_15_10, output_15_11, output_14_10;
mixer gate_output_14_10(.a(output_15_10), .b(output_15_11), .y(output_14_10));
wire output_16_10, output_16_11, output_15_10;
mixer gate_output_15_10(.a(output_16_10), .b(output_16_11), .y(output_15_10));
wire output_1_11, output_1_12, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_12), .y(output_0_11));
wire output_2_11, output_2_12, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_12), .y(output_1_11));
wire output_3_11, output_3_12, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_12), .y(output_2_11));
wire output_4_11, output_4_12, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_12), .y(output_3_11));
wire output_5_11, output_5_12, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_12), .y(output_4_11));
wire output_6_11, output_6_12, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_12), .y(output_5_11));
wire output_7_11, output_7_12, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_12), .y(output_6_11));
wire output_8_11, output_8_12, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_12), .y(output_7_11));
wire output_9_11, output_9_12, output_8_11;
mixer gate_output_8_11(.a(output_9_11), .b(output_9_12), .y(output_8_11));
wire output_10_11, output_10_12, output_9_11;
mixer gate_output_9_11(.a(output_10_11), .b(output_10_12), .y(output_9_11));
wire output_11_11, output_11_12, output_10_11;
mixer gate_output_10_11(.a(output_11_11), .b(output_11_12), .y(output_10_11));
wire output_12_11, output_12_12, output_11_11;
mixer gate_output_11_11(.a(output_12_11), .b(output_12_12), .y(output_11_11));
wire output_13_11, output_13_12, output_12_11;
mixer gate_output_12_11(.a(output_13_11), .b(output_13_12), .y(output_12_11));
wire output_14_11, output_14_12, output_13_11;
mixer gate_output_13_11(.a(output_14_11), .b(output_14_12), .y(output_13_11));
wire output_15_11, output_15_12, output_14_11;
mixer gate_output_14_11(.a(output_15_11), .b(output_15_12), .y(output_14_11));
wire output_16_11, output_16_12, output_15_11;
mixer gate_output_15_11(.a(output_16_11), .b(output_16_12), .y(output_15_11));
wire output_1_12, output_1_13, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_13), .y(output_0_12));
wire output_2_12, output_2_13, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_13), .y(output_1_12));
wire output_3_12, output_3_13, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_13), .y(output_2_12));
wire output_4_12, output_4_13, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_13), .y(output_3_12));
wire output_5_12, output_5_13, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_13), .y(output_4_12));
wire output_6_12, output_6_13, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_13), .y(output_5_12));
wire output_7_12, output_7_13, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_13), .y(output_6_12));
wire output_8_12, output_8_13, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_13), .y(output_7_12));
wire output_9_12, output_9_13, output_8_12;
mixer gate_output_8_12(.a(output_9_12), .b(output_9_13), .y(output_8_12));
wire output_10_12, output_10_13, output_9_12;
mixer gate_output_9_12(.a(output_10_12), .b(output_10_13), .y(output_9_12));
wire output_11_12, output_11_13, output_10_12;
mixer gate_output_10_12(.a(output_11_12), .b(output_11_13), .y(output_10_12));
wire output_12_12, output_12_13, output_11_12;
mixer gate_output_11_12(.a(output_12_12), .b(output_12_13), .y(output_11_12));
wire output_13_12, output_13_13, output_12_12;
mixer gate_output_12_12(.a(output_13_12), .b(output_13_13), .y(output_12_12));
wire output_14_12, output_14_13, output_13_12;
mixer gate_output_13_12(.a(output_14_12), .b(output_14_13), .y(output_13_12));
wire output_15_12, output_15_13, output_14_12;
mixer gate_output_14_12(.a(output_15_12), .b(output_15_13), .y(output_14_12));
wire output_16_12, output_16_13, output_15_12;
mixer gate_output_15_12(.a(output_16_12), .b(output_16_13), .y(output_15_12));
wire output_1_13, output_1_14, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_14), .y(output_0_13));
wire output_2_13, output_2_14, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_14), .y(output_1_13));
wire output_3_13, output_3_14, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_14), .y(output_2_13));
wire output_4_13, output_4_14, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_14), .y(output_3_13));
wire output_5_13, output_5_14, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_14), .y(output_4_13));
wire output_6_13, output_6_14, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_14), .y(output_5_13));
wire output_7_13, output_7_14, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_14), .y(output_6_13));
wire output_8_13, output_8_14, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_14), .y(output_7_13));
wire output_9_13, output_9_14, output_8_13;
mixer gate_output_8_13(.a(output_9_13), .b(output_9_14), .y(output_8_13));
wire output_10_13, output_10_14, output_9_13;
mixer gate_output_9_13(.a(output_10_13), .b(output_10_14), .y(output_9_13));
wire output_11_13, output_11_14, output_10_13;
mixer gate_output_10_13(.a(output_11_13), .b(output_11_14), .y(output_10_13));
wire output_12_13, output_12_14, output_11_13;
mixer gate_output_11_13(.a(output_12_13), .b(output_12_14), .y(output_11_13));
wire output_13_13, output_13_14, output_12_13;
mixer gate_output_12_13(.a(output_13_13), .b(output_13_14), .y(output_12_13));
wire output_14_13, output_14_14, output_13_13;
mixer gate_output_13_13(.a(output_14_13), .b(output_14_14), .y(output_13_13));
wire output_15_13, output_15_14, output_14_13;
mixer gate_output_14_13(.a(output_15_13), .b(output_15_14), .y(output_14_13));
wire output_16_13, output_16_14, output_15_13;
mixer gate_output_15_13(.a(output_16_13), .b(output_16_14), .y(output_15_13));
wire output_1_14, output_1_15, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_15), .y(output_0_14));
wire output_2_14, output_2_15, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_15), .y(output_1_14));
wire output_3_14, output_3_15, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_15), .y(output_2_14));
wire output_4_14, output_4_15, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_15), .y(output_3_14));
wire output_5_14, output_5_15, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_15), .y(output_4_14));
wire output_6_14, output_6_15, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_15), .y(output_5_14));
wire output_7_14, output_7_15, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_15), .y(output_6_14));
wire output_8_14, output_8_15, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_15), .y(output_7_14));
wire output_9_14, output_9_15, output_8_14;
mixer gate_output_8_14(.a(output_9_14), .b(output_9_15), .y(output_8_14));
wire output_10_14, output_10_15, output_9_14;
mixer gate_output_9_14(.a(output_10_14), .b(output_10_15), .y(output_9_14));
wire output_11_14, output_11_15, output_10_14;
mixer gate_output_10_14(.a(output_11_14), .b(output_11_15), .y(output_10_14));
wire output_12_14, output_12_15, output_11_14;
mixer gate_output_11_14(.a(output_12_14), .b(output_12_15), .y(output_11_14));
wire output_13_14, output_13_15, output_12_14;
mixer gate_output_12_14(.a(output_13_14), .b(output_13_15), .y(output_12_14));
wire output_14_14, output_14_15, output_13_14;
mixer gate_output_13_14(.a(output_14_14), .b(output_14_15), .y(output_13_14));
wire output_15_14, output_15_15, output_14_14;
mixer gate_output_14_14(.a(output_15_14), .b(output_15_15), .y(output_14_14));
wire output_16_14, output_16_15, output_15_14;
mixer gate_output_15_14(.a(output_16_14), .b(output_16_15), .y(output_15_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
wire output_9_15, output_9_0, output_8_15;
mixer gate_output_8_15(.a(output_9_15), .b(output_9_0), .y(output_8_15));
wire output_10_15, output_10_0, output_9_15;
mixer gate_output_9_15(.a(output_10_15), .b(output_10_0), .y(output_9_15));
wire output_11_15, output_11_0, output_10_15;
mixer gate_output_10_15(.a(output_11_15), .b(output_11_0), .y(output_10_15));
wire output_12_15, output_12_0, output_11_15;
mixer gate_output_11_15(.a(output_12_15), .b(output_12_0), .y(output_11_15));
wire output_13_15, output_13_0, output_12_15;
mixer gate_output_12_15(.a(output_13_15), .b(output_13_0), .y(output_12_15));
wire output_14_15, output_14_0, output_13_15;
mixer gate_output_13_15(.a(output_14_15), .b(output_14_0), .y(output_13_15));
wire output_15_15, output_15_0, output_14_15;
mixer gate_output_14_15(.a(output_15_15), .b(output_15_0), .y(output_14_15));
wire output_16_15, output_16_0, output_15_15;
mixer gate_output_15_15(.a(output_16_15), .b(output_16_0), .y(output_15_15));
wire output_1_16, output_1_1, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_1), .y(output_0_16));
wire output_2_16, output_2_1, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_1), .y(output_1_16));
wire output_3_16, output_3_1, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_1), .y(output_2_16));
wire output_4_16, output_4_1, output_3_16;
mixer gate_output_3_16(.a(output_4_16), .b(output_4_1), .y(output_3_16));
wire output_5_16, output_5_1, output_4_16;
mixer gate_output_4_16(.a(output_5_16), .b(output_5_1), .y(output_4_16));
wire output_6_16, output_6_1, output_5_16;
mixer gate_output_5_16(.a(output_6_16), .b(output_6_1), .y(output_5_16));
wire output_7_16, output_7_1, output_6_16;
mixer gate_output_6_16(.a(output_7_16), .b(output_7_1), .y(output_6_16));
wire output_8_16, output_8_1, output_7_16;
mixer gate_output_7_16(.a(output_8_16), .b(output_8_1), .y(output_7_16));
wire output_9_16, output_9_1, output_8_16;
mixer gate_output_8_16(.a(output_9_16), .b(output_9_1), .y(output_8_16));
wire output_10_16, output_10_1, output_9_16;
mixer gate_output_9_16(.a(output_10_16), .b(output_10_1), .y(output_9_16));
wire output_11_16, output_11_1, output_10_16;
mixer gate_output_10_16(.a(output_11_16), .b(output_11_1), .y(output_10_16));
wire output_12_16, output_12_1, output_11_16;
mixer gate_output_11_16(.a(output_12_16), .b(output_12_1), .y(output_11_16));
wire output_13_16, output_13_1, output_12_16;
mixer gate_output_12_16(.a(output_13_16), .b(output_13_1), .y(output_12_16));
wire output_14_16, output_14_1, output_13_16;
mixer gate_output_13_16(.a(output_14_16), .b(output_14_1), .y(output_13_16));
wire output_15_16, output_15_1, output_14_16;
mixer gate_output_14_16(.a(output_15_16), .b(output_15_1), .y(output_14_16));
wire output_16_16, output_16_1, output_15_16;
mixer gate_output_15_16(.a(output_16_16), .b(output_16_1), .y(output_15_16));
wire output_1_17, output_1_2, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_2), .y(output_0_17));
wire output_2_17, output_2_2, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_2), .y(output_1_17));
wire output_3_17, output_3_2, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_2), .y(output_2_17));
wire output_4_17, output_4_2, output_3_17;
mixer gate_output_3_17(.a(output_4_17), .b(output_4_2), .y(output_3_17));
wire output_5_17, output_5_2, output_4_17;
mixer gate_output_4_17(.a(output_5_17), .b(output_5_2), .y(output_4_17));
wire output_6_17, output_6_2, output_5_17;
mixer gate_output_5_17(.a(output_6_17), .b(output_6_2), .y(output_5_17));
wire output_7_17, output_7_2, output_6_17;
mixer gate_output_6_17(.a(output_7_17), .b(output_7_2), .y(output_6_17));
wire output_8_17, output_8_2, output_7_17;
mixer gate_output_7_17(.a(output_8_17), .b(output_8_2), .y(output_7_17));
wire output_9_17, output_9_2, output_8_17;
mixer gate_output_8_17(.a(output_9_17), .b(output_9_2), .y(output_8_17));
wire output_10_17, output_10_2, output_9_17;
mixer gate_output_9_17(.a(output_10_17), .b(output_10_2), .y(output_9_17));
wire output_11_17, output_11_2, output_10_17;
mixer gate_output_10_17(.a(output_11_17), .b(output_11_2), .y(output_10_17));
wire output_12_17, output_12_2, output_11_17;
mixer gate_output_11_17(.a(output_12_17), .b(output_12_2), .y(output_11_17));
wire output_13_17, output_13_2, output_12_17;
mixer gate_output_12_17(.a(output_13_17), .b(output_13_2), .y(output_12_17));
wire output_14_17, output_14_2, output_13_17;
mixer gate_output_13_17(.a(output_14_17), .b(output_14_2), .y(output_13_17));
wire output_15_17, output_15_2, output_14_17;
mixer gate_output_14_17(.a(output_15_17), .b(output_15_2), .y(output_14_17));
wire output_16_17, output_16_2, output_15_17;
mixer gate_output_15_17(.a(output_16_17), .b(output_16_2), .y(output_15_17));
wire output_1_18, output_1_3, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_3), .y(output_0_18));
wire output_2_18, output_2_3, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_3), .y(output_1_18));
wire output_3_18, output_3_3, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_3), .y(output_2_18));
wire output_4_18, output_4_3, output_3_18;
mixer gate_output_3_18(.a(output_4_18), .b(output_4_3), .y(output_3_18));
wire output_5_18, output_5_3, output_4_18;
mixer gate_output_4_18(.a(output_5_18), .b(output_5_3), .y(output_4_18));
wire output_6_18, output_6_3, output_5_18;
mixer gate_output_5_18(.a(output_6_18), .b(output_6_3), .y(output_5_18));
wire output_7_18, output_7_3, output_6_18;
mixer gate_output_6_18(.a(output_7_18), .b(output_7_3), .y(output_6_18));
wire output_8_18, output_8_3, output_7_18;
mixer gate_output_7_18(.a(output_8_18), .b(output_8_3), .y(output_7_18));
wire output_9_18, output_9_3, output_8_18;
mixer gate_output_8_18(.a(output_9_18), .b(output_9_3), .y(output_8_18));
wire output_10_18, output_10_3, output_9_18;
mixer gate_output_9_18(.a(output_10_18), .b(output_10_3), .y(output_9_18));
wire output_11_18, output_11_3, output_10_18;
mixer gate_output_10_18(.a(output_11_18), .b(output_11_3), .y(output_10_18));
wire output_12_18, output_12_3, output_11_18;
mixer gate_output_11_18(.a(output_12_18), .b(output_12_3), .y(output_11_18));
wire output_13_18, output_13_3, output_12_18;
mixer gate_output_12_18(.a(output_13_18), .b(output_13_3), .y(output_12_18));
wire output_14_18, output_14_3, output_13_18;
mixer gate_output_13_18(.a(output_14_18), .b(output_14_3), .y(output_13_18));
wire output_15_18, output_15_3, output_14_18;
mixer gate_output_14_18(.a(output_15_18), .b(output_15_3), .y(output_14_18));
wire output_16_18, output_16_3, output_15_18;
mixer gate_output_15_18(.a(output_16_18), .b(output_16_3), .y(output_15_18));
wire output_1_19, output_1_4, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_4), .y(output_0_19));
wire output_2_19, output_2_4, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_4), .y(output_1_19));
wire output_3_19, output_3_4, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_4), .y(output_2_19));
wire output_4_19, output_4_4, output_3_19;
mixer gate_output_3_19(.a(output_4_19), .b(output_4_4), .y(output_3_19));
wire output_5_19, output_5_4, output_4_19;
mixer gate_output_4_19(.a(output_5_19), .b(output_5_4), .y(output_4_19));
wire output_6_19, output_6_4, output_5_19;
mixer gate_output_5_19(.a(output_6_19), .b(output_6_4), .y(output_5_19));
wire output_7_19, output_7_4, output_6_19;
mixer gate_output_6_19(.a(output_7_19), .b(output_7_4), .y(output_6_19));
wire output_8_19, output_8_4, output_7_19;
mixer gate_output_7_19(.a(output_8_19), .b(output_8_4), .y(output_7_19));
wire output_9_19, output_9_4, output_8_19;
mixer gate_output_8_19(.a(output_9_19), .b(output_9_4), .y(output_8_19));
wire output_10_19, output_10_4, output_9_19;
mixer gate_output_9_19(.a(output_10_19), .b(output_10_4), .y(output_9_19));
wire output_11_19, output_11_4, output_10_19;
mixer gate_output_10_19(.a(output_11_19), .b(output_11_4), .y(output_10_19));
wire output_12_19, output_12_4, output_11_19;
mixer gate_output_11_19(.a(output_12_19), .b(output_12_4), .y(output_11_19));
wire output_13_19, output_13_4, output_12_19;
mixer gate_output_12_19(.a(output_13_19), .b(output_13_4), .y(output_12_19));
wire output_14_19, output_14_4, output_13_19;
mixer gate_output_13_19(.a(output_14_19), .b(output_14_4), .y(output_13_19));
wire output_15_19, output_15_4, output_14_19;
mixer gate_output_14_19(.a(output_15_19), .b(output_15_4), .y(output_14_19));
wire output_16_19, output_16_4, output_15_19;
mixer gate_output_15_19(.a(output_16_19), .b(output_16_4), .y(output_15_19));
wire output_1_20, output_1_5, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_5), .y(output_0_20));
wire output_2_20, output_2_5, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_5), .y(output_1_20));
wire output_3_20, output_3_5, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_5), .y(output_2_20));
wire output_4_20, output_4_5, output_3_20;
mixer gate_output_3_20(.a(output_4_20), .b(output_4_5), .y(output_3_20));
wire output_5_20, output_5_5, output_4_20;
mixer gate_output_4_20(.a(output_5_20), .b(output_5_5), .y(output_4_20));
wire output_6_20, output_6_5, output_5_20;
mixer gate_output_5_20(.a(output_6_20), .b(output_6_5), .y(output_5_20));
wire output_7_20, output_7_5, output_6_20;
mixer gate_output_6_20(.a(output_7_20), .b(output_7_5), .y(output_6_20));
wire output_8_20, output_8_5, output_7_20;
mixer gate_output_7_20(.a(output_8_20), .b(output_8_5), .y(output_7_20));
wire output_9_20, output_9_5, output_8_20;
mixer gate_output_8_20(.a(output_9_20), .b(output_9_5), .y(output_8_20));
wire output_10_20, output_10_5, output_9_20;
mixer gate_output_9_20(.a(output_10_20), .b(output_10_5), .y(output_9_20));
wire output_11_20, output_11_5, output_10_20;
mixer gate_output_10_20(.a(output_11_20), .b(output_11_5), .y(output_10_20));
wire output_12_20, output_12_5, output_11_20;
mixer gate_output_11_20(.a(output_12_20), .b(output_12_5), .y(output_11_20));
wire output_13_20, output_13_5, output_12_20;
mixer gate_output_12_20(.a(output_13_20), .b(output_13_5), .y(output_12_20));
wire output_14_20, output_14_5, output_13_20;
mixer gate_output_13_20(.a(output_14_20), .b(output_14_5), .y(output_13_20));
wire output_15_20, output_15_5, output_14_20;
mixer gate_output_14_20(.a(output_15_20), .b(output_15_5), .y(output_14_20));
wire output_16_20, output_16_5, output_15_20;
mixer gate_output_15_20(.a(output_16_20), .b(output_16_5), .y(output_15_20));
wire output_1_21, output_1_6, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_6), .y(output_0_21));
wire output_2_21, output_2_6, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_6), .y(output_1_21));
wire output_3_21, output_3_6, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_6), .y(output_2_21));
wire output_4_21, output_4_6, output_3_21;
mixer gate_output_3_21(.a(output_4_21), .b(output_4_6), .y(output_3_21));
wire output_5_21, output_5_6, output_4_21;
mixer gate_output_4_21(.a(output_5_21), .b(output_5_6), .y(output_4_21));
wire output_6_21, output_6_6, output_5_21;
mixer gate_output_5_21(.a(output_6_21), .b(output_6_6), .y(output_5_21));
wire output_7_21, output_7_6, output_6_21;
mixer gate_output_6_21(.a(output_7_21), .b(output_7_6), .y(output_6_21));
wire output_8_21, output_8_6, output_7_21;
mixer gate_output_7_21(.a(output_8_21), .b(output_8_6), .y(output_7_21));
wire output_9_21, output_9_6, output_8_21;
mixer gate_output_8_21(.a(output_9_21), .b(output_9_6), .y(output_8_21));
wire output_10_21, output_10_6, output_9_21;
mixer gate_output_9_21(.a(output_10_21), .b(output_10_6), .y(output_9_21));
wire output_11_21, output_11_6, output_10_21;
mixer gate_output_10_21(.a(output_11_21), .b(output_11_6), .y(output_10_21));
wire output_12_21, output_12_6, output_11_21;
mixer gate_output_11_21(.a(output_12_21), .b(output_12_6), .y(output_11_21));
wire output_13_21, output_13_6, output_12_21;
mixer gate_output_12_21(.a(output_13_21), .b(output_13_6), .y(output_12_21));
wire output_14_21, output_14_6, output_13_21;
mixer gate_output_13_21(.a(output_14_21), .b(output_14_6), .y(output_13_21));
wire output_15_21, output_15_6, output_14_21;
mixer gate_output_14_21(.a(output_15_21), .b(output_15_6), .y(output_14_21));
wire output_16_21, output_16_6, output_15_21;
mixer gate_output_15_21(.a(output_16_21), .b(output_16_6), .y(output_15_21));
wire output_1_22, output_1_7, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_7), .y(output_0_22));
wire output_2_22, output_2_7, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_7), .y(output_1_22));
wire output_3_22, output_3_7, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_7), .y(output_2_22));
wire output_4_22, output_4_7, output_3_22;
mixer gate_output_3_22(.a(output_4_22), .b(output_4_7), .y(output_3_22));
wire output_5_22, output_5_7, output_4_22;
mixer gate_output_4_22(.a(output_5_22), .b(output_5_7), .y(output_4_22));
wire output_6_22, output_6_7, output_5_22;
mixer gate_output_5_22(.a(output_6_22), .b(output_6_7), .y(output_5_22));
wire output_7_22, output_7_7, output_6_22;
mixer gate_output_6_22(.a(output_7_22), .b(output_7_7), .y(output_6_22));
wire output_8_22, output_8_7, output_7_22;
mixer gate_output_7_22(.a(output_8_22), .b(output_8_7), .y(output_7_22));
wire output_9_22, output_9_7, output_8_22;
mixer gate_output_8_22(.a(output_9_22), .b(output_9_7), .y(output_8_22));
wire output_10_22, output_10_7, output_9_22;
mixer gate_output_9_22(.a(output_10_22), .b(output_10_7), .y(output_9_22));
wire output_11_22, output_11_7, output_10_22;
mixer gate_output_10_22(.a(output_11_22), .b(output_11_7), .y(output_10_22));
wire output_12_22, output_12_7, output_11_22;
mixer gate_output_11_22(.a(output_12_22), .b(output_12_7), .y(output_11_22));
wire output_13_22, output_13_7, output_12_22;
mixer gate_output_12_22(.a(output_13_22), .b(output_13_7), .y(output_12_22));
wire output_14_22, output_14_7, output_13_22;
mixer gate_output_13_22(.a(output_14_22), .b(output_14_7), .y(output_13_22));
wire output_15_22, output_15_7, output_14_22;
mixer gate_output_14_22(.a(output_15_22), .b(output_15_7), .y(output_14_22));
wire output_16_22, output_16_7, output_15_22;
mixer gate_output_15_22(.a(output_16_22), .b(output_16_7), .y(output_15_22));
wire output_1_23, output_1_8, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_8), .y(output_0_23));
wire output_2_23, output_2_8, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_8), .y(output_1_23));
wire output_3_23, output_3_8, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_8), .y(output_2_23));
wire output_4_23, output_4_8, output_3_23;
mixer gate_output_3_23(.a(output_4_23), .b(output_4_8), .y(output_3_23));
wire output_5_23, output_5_8, output_4_23;
mixer gate_output_4_23(.a(output_5_23), .b(output_5_8), .y(output_4_23));
wire output_6_23, output_6_8, output_5_23;
mixer gate_output_5_23(.a(output_6_23), .b(output_6_8), .y(output_5_23));
wire output_7_23, output_7_8, output_6_23;
mixer gate_output_6_23(.a(output_7_23), .b(output_7_8), .y(output_6_23));
wire output_8_23, output_8_8, output_7_23;
mixer gate_output_7_23(.a(output_8_23), .b(output_8_8), .y(output_7_23));
wire output_9_23, output_9_8, output_8_23;
mixer gate_output_8_23(.a(output_9_23), .b(output_9_8), .y(output_8_23));
wire output_10_23, output_10_8, output_9_23;
mixer gate_output_9_23(.a(output_10_23), .b(output_10_8), .y(output_9_23));
wire output_11_23, output_11_8, output_10_23;
mixer gate_output_10_23(.a(output_11_23), .b(output_11_8), .y(output_10_23));
wire output_12_23, output_12_8, output_11_23;
mixer gate_output_11_23(.a(output_12_23), .b(output_12_8), .y(output_11_23));
wire output_13_23, output_13_8, output_12_23;
mixer gate_output_12_23(.a(output_13_23), .b(output_13_8), .y(output_12_23));
wire output_14_23, output_14_8, output_13_23;
mixer gate_output_13_23(.a(output_14_23), .b(output_14_8), .y(output_13_23));
wire output_15_23, output_15_8, output_14_23;
mixer gate_output_14_23(.a(output_15_23), .b(output_15_8), .y(output_14_23));
wire output_16_23, output_16_8, output_15_23;
mixer gate_output_15_23(.a(output_16_23), .b(output_16_8), .y(output_15_23));
wire output_1_24, output_1_9, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_9), .y(output_0_24));
wire output_2_24, output_2_9, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_9), .y(output_1_24));
wire output_3_24, output_3_9, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_9), .y(output_2_24));
wire output_4_24, output_4_9, output_3_24;
mixer gate_output_3_24(.a(output_4_24), .b(output_4_9), .y(output_3_24));
wire output_5_24, output_5_9, output_4_24;
mixer gate_output_4_24(.a(output_5_24), .b(output_5_9), .y(output_4_24));
wire output_6_24, output_6_9, output_5_24;
mixer gate_output_5_24(.a(output_6_24), .b(output_6_9), .y(output_5_24));
wire output_7_24, output_7_9, output_6_24;
mixer gate_output_6_24(.a(output_7_24), .b(output_7_9), .y(output_6_24));
wire output_8_24, output_8_9, output_7_24;
mixer gate_output_7_24(.a(output_8_24), .b(output_8_9), .y(output_7_24));
wire output_9_24, output_9_9, output_8_24;
mixer gate_output_8_24(.a(output_9_24), .b(output_9_9), .y(output_8_24));
wire output_10_24, output_10_9, output_9_24;
mixer gate_output_9_24(.a(output_10_24), .b(output_10_9), .y(output_9_24));
wire output_11_24, output_11_9, output_10_24;
mixer gate_output_10_24(.a(output_11_24), .b(output_11_9), .y(output_10_24));
wire output_12_24, output_12_9, output_11_24;
mixer gate_output_11_24(.a(output_12_24), .b(output_12_9), .y(output_11_24));
wire output_13_24, output_13_9, output_12_24;
mixer gate_output_12_24(.a(output_13_24), .b(output_13_9), .y(output_12_24));
wire output_14_24, output_14_9, output_13_24;
mixer gate_output_13_24(.a(output_14_24), .b(output_14_9), .y(output_13_24));
wire output_15_24, output_15_9, output_14_24;
mixer gate_output_14_24(.a(output_15_24), .b(output_15_9), .y(output_14_24));
wire output_16_24, output_16_9, output_15_24;
mixer gate_output_15_24(.a(output_16_24), .b(output_16_9), .y(output_15_24));
wire output_1_25, output_1_10, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_10), .y(output_0_25));
wire output_2_25, output_2_10, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_10), .y(output_1_25));
wire output_3_25, output_3_10, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_10), .y(output_2_25));
wire output_4_25, output_4_10, output_3_25;
mixer gate_output_3_25(.a(output_4_25), .b(output_4_10), .y(output_3_25));
wire output_5_25, output_5_10, output_4_25;
mixer gate_output_4_25(.a(output_5_25), .b(output_5_10), .y(output_4_25));
wire output_6_25, output_6_10, output_5_25;
mixer gate_output_5_25(.a(output_6_25), .b(output_6_10), .y(output_5_25));
wire output_7_25, output_7_10, output_6_25;
mixer gate_output_6_25(.a(output_7_25), .b(output_7_10), .y(output_6_25));
wire output_8_25, output_8_10, output_7_25;
mixer gate_output_7_25(.a(output_8_25), .b(output_8_10), .y(output_7_25));
wire output_9_25, output_9_10, output_8_25;
mixer gate_output_8_25(.a(output_9_25), .b(output_9_10), .y(output_8_25));
wire output_10_25, output_10_10, output_9_25;
mixer gate_output_9_25(.a(output_10_25), .b(output_10_10), .y(output_9_25));
wire output_11_25, output_11_10, output_10_25;
mixer gate_output_10_25(.a(output_11_25), .b(output_11_10), .y(output_10_25));
wire output_12_25, output_12_10, output_11_25;
mixer gate_output_11_25(.a(output_12_25), .b(output_12_10), .y(output_11_25));
wire output_13_25, output_13_10, output_12_25;
mixer gate_output_12_25(.a(output_13_25), .b(output_13_10), .y(output_12_25));
wire output_14_25, output_14_10, output_13_25;
mixer gate_output_13_25(.a(output_14_25), .b(output_14_10), .y(output_13_25));
wire output_15_25, output_15_10, output_14_25;
mixer gate_output_14_25(.a(output_15_25), .b(output_15_10), .y(output_14_25));
wire output_16_25, output_16_10, output_15_25;
mixer gate_output_15_25(.a(output_16_25), .b(output_16_10), .y(output_15_25));
wire output_1_26, output_1_11, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_11), .y(output_0_26));
wire output_2_26, output_2_11, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_11), .y(output_1_26));
wire output_3_26, output_3_11, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_11), .y(output_2_26));
wire output_4_26, output_4_11, output_3_26;
mixer gate_output_3_26(.a(output_4_26), .b(output_4_11), .y(output_3_26));
wire output_5_26, output_5_11, output_4_26;
mixer gate_output_4_26(.a(output_5_26), .b(output_5_11), .y(output_4_26));
wire output_6_26, output_6_11, output_5_26;
mixer gate_output_5_26(.a(output_6_26), .b(output_6_11), .y(output_5_26));
wire output_7_26, output_7_11, output_6_26;
mixer gate_output_6_26(.a(output_7_26), .b(output_7_11), .y(output_6_26));
wire output_8_26, output_8_11, output_7_26;
mixer gate_output_7_26(.a(output_8_26), .b(output_8_11), .y(output_7_26));
wire output_9_26, output_9_11, output_8_26;
mixer gate_output_8_26(.a(output_9_26), .b(output_9_11), .y(output_8_26));
wire output_10_26, output_10_11, output_9_26;
mixer gate_output_9_26(.a(output_10_26), .b(output_10_11), .y(output_9_26));
wire output_11_26, output_11_11, output_10_26;
mixer gate_output_10_26(.a(output_11_26), .b(output_11_11), .y(output_10_26));
wire output_12_26, output_12_11, output_11_26;
mixer gate_output_11_26(.a(output_12_26), .b(output_12_11), .y(output_11_26));
wire output_13_26, output_13_11, output_12_26;
mixer gate_output_12_26(.a(output_13_26), .b(output_13_11), .y(output_12_26));
wire output_14_26, output_14_11, output_13_26;
mixer gate_output_13_26(.a(output_14_26), .b(output_14_11), .y(output_13_26));
wire output_15_26, output_15_11, output_14_26;
mixer gate_output_14_26(.a(output_15_26), .b(output_15_11), .y(output_14_26));
wire output_16_26, output_16_11, output_15_26;
mixer gate_output_15_26(.a(output_16_26), .b(output_16_11), .y(output_15_26));
wire output_1_27, output_1_12, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_12), .y(output_0_27));
wire output_2_27, output_2_12, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_12), .y(output_1_27));
wire output_3_27, output_3_12, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_12), .y(output_2_27));
wire output_4_27, output_4_12, output_3_27;
mixer gate_output_3_27(.a(output_4_27), .b(output_4_12), .y(output_3_27));
wire output_5_27, output_5_12, output_4_27;
mixer gate_output_4_27(.a(output_5_27), .b(output_5_12), .y(output_4_27));
wire output_6_27, output_6_12, output_5_27;
mixer gate_output_5_27(.a(output_6_27), .b(output_6_12), .y(output_5_27));
wire output_7_27, output_7_12, output_6_27;
mixer gate_output_6_27(.a(output_7_27), .b(output_7_12), .y(output_6_27));
wire output_8_27, output_8_12, output_7_27;
mixer gate_output_7_27(.a(output_8_27), .b(output_8_12), .y(output_7_27));
wire output_9_27, output_9_12, output_8_27;
mixer gate_output_8_27(.a(output_9_27), .b(output_9_12), .y(output_8_27));
wire output_10_27, output_10_12, output_9_27;
mixer gate_output_9_27(.a(output_10_27), .b(output_10_12), .y(output_9_27));
wire output_11_27, output_11_12, output_10_27;
mixer gate_output_10_27(.a(output_11_27), .b(output_11_12), .y(output_10_27));
wire output_12_27, output_12_12, output_11_27;
mixer gate_output_11_27(.a(output_12_27), .b(output_12_12), .y(output_11_27));
wire output_13_27, output_13_12, output_12_27;
mixer gate_output_12_27(.a(output_13_27), .b(output_13_12), .y(output_12_27));
wire output_14_27, output_14_12, output_13_27;
mixer gate_output_13_27(.a(output_14_27), .b(output_14_12), .y(output_13_27));
wire output_15_27, output_15_12, output_14_27;
mixer gate_output_14_27(.a(output_15_27), .b(output_15_12), .y(output_14_27));
wire output_16_27, output_16_12, output_15_27;
mixer gate_output_15_27(.a(output_16_27), .b(output_16_12), .y(output_15_27));
wire output_1_28, output_1_13, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_13), .y(output_0_28));
wire output_2_28, output_2_13, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_13), .y(output_1_28));
wire output_3_28, output_3_13, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_13), .y(output_2_28));
wire output_4_28, output_4_13, output_3_28;
mixer gate_output_3_28(.a(output_4_28), .b(output_4_13), .y(output_3_28));
wire output_5_28, output_5_13, output_4_28;
mixer gate_output_4_28(.a(output_5_28), .b(output_5_13), .y(output_4_28));
wire output_6_28, output_6_13, output_5_28;
mixer gate_output_5_28(.a(output_6_28), .b(output_6_13), .y(output_5_28));
wire output_7_28, output_7_13, output_6_28;
mixer gate_output_6_28(.a(output_7_28), .b(output_7_13), .y(output_6_28));
wire output_8_28, output_8_13, output_7_28;
mixer gate_output_7_28(.a(output_8_28), .b(output_8_13), .y(output_7_28));
wire output_9_28, output_9_13, output_8_28;
mixer gate_output_8_28(.a(output_9_28), .b(output_9_13), .y(output_8_28));
wire output_10_28, output_10_13, output_9_28;
mixer gate_output_9_28(.a(output_10_28), .b(output_10_13), .y(output_9_28));
wire output_11_28, output_11_13, output_10_28;
mixer gate_output_10_28(.a(output_11_28), .b(output_11_13), .y(output_10_28));
wire output_12_28, output_12_13, output_11_28;
mixer gate_output_11_28(.a(output_12_28), .b(output_12_13), .y(output_11_28));
wire output_13_28, output_13_13, output_12_28;
mixer gate_output_12_28(.a(output_13_28), .b(output_13_13), .y(output_12_28));
wire output_14_28, output_14_13, output_13_28;
mixer gate_output_13_28(.a(output_14_28), .b(output_14_13), .y(output_13_28));
wire output_15_28, output_15_13, output_14_28;
mixer gate_output_14_28(.a(output_15_28), .b(output_15_13), .y(output_14_28));
wire output_16_28, output_16_13, output_15_28;
mixer gate_output_15_28(.a(output_16_28), .b(output_16_13), .y(output_15_28));
wire output_1_29, output_1_14, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_14), .y(output_0_29));
wire output_2_29, output_2_14, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_14), .y(output_1_29));
wire output_3_29, output_3_14, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_14), .y(output_2_29));
wire output_4_29, output_4_14, output_3_29;
mixer gate_output_3_29(.a(output_4_29), .b(output_4_14), .y(output_3_29));
wire output_5_29, output_5_14, output_4_29;
mixer gate_output_4_29(.a(output_5_29), .b(output_5_14), .y(output_4_29));
wire output_6_29, output_6_14, output_5_29;
mixer gate_output_5_29(.a(output_6_29), .b(output_6_14), .y(output_5_29));
wire output_7_29, output_7_14, output_6_29;
mixer gate_output_6_29(.a(output_7_29), .b(output_7_14), .y(output_6_29));
wire output_8_29, output_8_14, output_7_29;
mixer gate_output_7_29(.a(output_8_29), .b(output_8_14), .y(output_7_29));
wire output_9_29, output_9_14, output_8_29;
mixer gate_output_8_29(.a(output_9_29), .b(output_9_14), .y(output_8_29));
wire output_10_29, output_10_14, output_9_29;
mixer gate_output_9_29(.a(output_10_29), .b(output_10_14), .y(output_9_29));
wire output_11_29, output_11_14, output_10_29;
mixer gate_output_10_29(.a(output_11_29), .b(output_11_14), .y(output_10_29));
wire output_12_29, output_12_14, output_11_29;
mixer gate_output_11_29(.a(output_12_29), .b(output_12_14), .y(output_11_29));
wire output_13_29, output_13_14, output_12_29;
mixer gate_output_12_29(.a(output_13_29), .b(output_13_14), .y(output_12_29));
wire output_14_29, output_14_14, output_13_29;
mixer gate_output_13_29(.a(output_14_29), .b(output_14_14), .y(output_13_29));
wire output_15_29, output_15_14, output_14_29;
mixer gate_output_14_29(.a(output_15_29), .b(output_15_14), .y(output_14_29));
wire output_16_29, output_16_14, output_15_29;
mixer gate_output_15_29(.a(output_16_29), .b(output_16_14), .y(output_15_29));
wire output_1_30, output_1_15, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_15), .y(output_0_30));
wire output_2_30, output_2_15, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_15), .y(output_1_30));
wire output_3_30, output_3_15, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_15), .y(output_2_30));
wire output_4_30, output_4_15, output_3_30;
mixer gate_output_3_30(.a(output_4_30), .b(output_4_15), .y(output_3_30));
wire output_5_30, output_5_15, output_4_30;
mixer gate_output_4_30(.a(output_5_30), .b(output_5_15), .y(output_4_30));
wire output_6_30, output_6_15, output_5_30;
mixer gate_output_5_30(.a(output_6_30), .b(output_6_15), .y(output_5_30));
wire output_7_30, output_7_15, output_6_30;
mixer gate_output_6_30(.a(output_7_30), .b(output_7_15), .y(output_6_30));
wire output_8_30, output_8_15, output_7_30;
mixer gate_output_7_30(.a(output_8_30), .b(output_8_15), .y(output_7_30));
wire output_9_30, output_9_15, output_8_30;
mixer gate_output_8_30(.a(output_9_30), .b(output_9_15), .y(output_8_30));
wire output_10_30, output_10_15, output_9_30;
mixer gate_output_9_30(.a(output_10_30), .b(output_10_15), .y(output_9_30));
wire output_11_30, output_11_15, output_10_30;
mixer gate_output_10_30(.a(output_11_30), .b(output_11_15), .y(output_10_30));
wire output_12_30, output_12_15, output_11_30;
mixer gate_output_11_30(.a(output_12_30), .b(output_12_15), .y(output_11_30));
wire output_13_30, output_13_15, output_12_30;
mixer gate_output_12_30(.a(output_13_30), .b(output_13_15), .y(output_12_30));
wire output_14_30, output_14_15, output_13_30;
mixer gate_output_13_30(.a(output_14_30), .b(output_14_15), .y(output_13_30));
wire output_15_30, output_15_15, output_14_30;
mixer gate_output_14_30(.a(output_15_30), .b(output_15_15), .y(output_14_30));
wire output_16_30, output_16_15, output_15_30;
mixer gate_output_15_30(.a(output_16_30), .b(output_16_15), .y(output_15_30));
wire output_1_31, output_1_0, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_0), .y(output_0_31));
wire output_2_31, output_2_0, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_0), .y(output_1_31));
wire output_3_31, output_3_0, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_0), .y(output_2_31));
wire output_4_31, output_4_0, output_3_31;
mixer gate_output_3_31(.a(output_4_31), .b(output_4_0), .y(output_3_31));
wire output_5_31, output_5_0, output_4_31;
mixer gate_output_4_31(.a(output_5_31), .b(output_5_0), .y(output_4_31));
wire output_6_31, output_6_0, output_5_31;
mixer gate_output_5_31(.a(output_6_31), .b(output_6_0), .y(output_5_31));
wire output_7_31, output_7_0, output_6_31;
mixer gate_output_6_31(.a(output_7_31), .b(output_7_0), .y(output_6_31));
wire output_8_31, output_8_0, output_7_31;
mixer gate_output_7_31(.a(output_8_31), .b(output_8_0), .y(output_7_31));
wire output_9_31, output_9_0, output_8_31;
mixer gate_output_8_31(.a(output_9_31), .b(output_9_0), .y(output_8_31));
wire output_10_31, output_10_0, output_9_31;
mixer gate_output_9_31(.a(output_10_31), .b(output_10_0), .y(output_9_31));
wire output_11_31, output_11_0, output_10_31;
mixer gate_output_10_31(.a(output_11_31), .b(output_11_0), .y(output_10_31));
wire output_12_31, output_12_0, output_11_31;
mixer gate_output_11_31(.a(output_12_31), .b(output_12_0), .y(output_11_31));
wire output_13_31, output_13_0, output_12_31;
mixer gate_output_12_31(.a(output_13_31), .b(output_13_0), .y(output_12_31));
wire output_14_31, output_14_0, output_13_31;
mixer gate_output_13_31(.a(output_14_31), .b(output_14_0), .y(output_13_31));
wire output_15_31, output_15_0, output_14_31;
mixer gate_output_14_31(.a(output_15_31), .b(output_15_0), .y(output_14_31));
wire output_16_31, output_16_0, output_15_31;
mixer gate_output_15_31(.a(output_16_31), .b(output_16_0), .y(output_15_31));
wire output_1_32, output_1_1, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_1), .y(output_0_32));
wire output_2_32, output_2_1, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_1), .y(output_1_32));
wire output_3_32, output_3_1, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_1), .y(output_2_32));
wire output_4_32, output_4_1, output_3_32;
mixer gate_output_3_32(.a(output_4_32), .b(output_4_1), .y(output_3_32));
wire output_5_32, output_5_1, output_4_32;
mixer gate_output_4_32(.a(output_5_32), .b(output_5_1), .y(output_4_32));
wire output_6_32, output_6_1, output_5_32;
mixer gate_output_5_32(.a(output_6_32), .b(output_6_1), .y(output_5_32));
wire output_7_32, output_7_1, output_6_32;
mixer gate_output_6_32(.a(output_7_32), .b(output_7_1), .y(output_6_32));
wire output_8_32, output_8_1, output_7_32;
mixer gate_output_7_32(.a(output_8_32), .b(output_8_1), .y(output_7_32));
wire output_9_32, output_9_1, output_8_32;
mixer gate_output_8_32(.a(output_9_32), .b(output_9_1), .y(output_8_32));
wire output_10_32, output_10_1, output_9_32;
mixer gate_output_9_32(.a(output_10_32), .b(output_10_1), .y(output_9_32));
wire output_11_32, output_11_1, output_10_32;
mixer gate_output_10_32(.a(output_11_32), .b(output_11_1), .y(output_10_32));
wire output_12_32, output_12_1, output_11_32;
mixer gate_output_11_32(.a(output_12_32), .b(output_12_1), .y(output_11_32));
wire output_13_32, output_13_1, output_12_32;
mixer gate_output_12_32(.a(output_13_32), .b(output_13_1), .y(output_12_32));
wire output_14_32, output_14_1, output_13_32;
mixer gate_output_13_32(.a(output_14_32), .b(output_14_1), .y(output_13_32));
wire output_15_32, output_15_1, output_14_32;
mixer gate_output_14_32(.a(output_15_32), .b(output_15_1), .y(output_14_32));
wire output_16_32, output_16_1, output_15_32;
mixer gate_output_15_32(.a(output_16_32), .b(output_16_1), .y(output_15_32));
wire output_1_33, output_1_2, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_2), .y(output_0_33));
wire output_2_33, output_2_2, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_2), .y(output_1_33));
wire output_3_33, output_3_2, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_2), .y(output_2_33));
wire output_4_33, output_4_2, output_3_33;
mixer gate_output_3_33(.a(output_4_33), .b(output_4_2), .y(output_3_33));
wire output_5_33, output_5_2, output_4_33;
mixer gate_output_4_33(.a(output_5_33), .b(output_5_2), .y(output_4_33));
wire output_6_33, output_6_2, output_5_33;
mixer gate_output_5_33(.a(output_6_33), .b(output_6_2), .y(output_5_33));
wire output_7_33, output_7_2, output_6_33;
mixer gate_output_6_33(.a(output_7_33), .b(output_7_2), .y(output_6_33));
wire output_8_33, output_8_2, output_7_33;
mixer gate_output_7_33(.a(output_8_33), .b(output_8_2), .y(output_7_33));
wire output_9_33, output_9_2, output_8_33;
mixer gate_output_8_33(.a(output_9_33), .b(output_9_2), .y(output_8_33));
wire output_10_33, output_10_2, output_9_33;
mixer gate_output_9_33(.a(output_10_33), .b(output_10_2), .y(output_9_33));
wire output_11_33, output_11_2, output_10_33;
mixer gate_output_10_33(.a(output_11_33), .b(output_11_2), .y(output_10_33));
wire output_12_33, output_12_2, output_11_33;
mixer gate_output_11_33(.a(output_12_33), .b(output_12_2), .y(output_11_33));
wire output_13_33, output_13_2, output_12_33;
mixer gate_output_12_33(.a(output_13_33), .b(output_13_2), .y(output_12_33));
wire output_14_33, output_14_2, output_13_33;
mixer gate_output_13_33(.a(output_14_33), .b(output_14_2), .y(output_13_33));
wire output_15_33, output_15_2, output_14_33;
mixer gate_output_14_33(.a(output_15_33), .b(output_15_2), .y(output_14_33));
wire output_16_33, output_16_2, output_15_33;
mixer gate_output_15_33(.a(output_16_33), .b(output_16_2), .y(output_15_33));
wire output_1_34, output_1_3, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_3), .y(output_0_34));
wire output_2_34, output_2_3, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_3), .y(output_1_34));
wire output_3_34, output_3_3, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_3), .y(output_2_34));
wire output_4_34, output_4_3, output_3_34;
mixer gate_output_3_34(.a(output_4_34), .b(output_4_3), .y(output_3_34));
wire output_5_34, output_5_3, output_4_34;
mixer gate_output_4_34(.a(output_5_34), .b(output_5_3), .y(output_4_34));
wire output_6_34, output_6_3, output_5_34;
mixer gate_output_5_34(.a(output_6_34), .b(output_6_3), .y(output_5_34));
wire output_7_34, output_7_3, output_6_34;
mixer gate_output_6_34(.a(output_7_34), .b(output_7_3), .y(output_6_34));
wire output_8_34, output_8_3, output_7_34;
mixer gate_output_7_34(.a(output_8_34), .b(output_8_3), .y(output_7_34));
wire output_9_34, output_9_3, output_8_34;
mixer gate_output_8_34(.a(output_9_34), .b(output_9_3), .y(output_8_34));
wire output_10_34, output_10_3, output_9_34;
mixer gate_output_9_34(.a(output_10_34), .b(output_10_3), .y(output_9_34));
wire output_11_34, output_11_3, output_10_34;
mixer gate_output_10_34(.a(output_11_34), .b(output_11_3), .y(output_10_34));
wire output_12_34, output_12_3, output_11_34;
mixer gate_output_11_34(.a(output_12_34), .b(output_12_3), .y(output_11_34));
wire output_13_34, output_13_3, output_12_34;
mixer gate_output_12_34(.a(output_13_34), .b(output_13_3), .y(output_12_34));
wire output_14_34, output_14_3, output_13_34;
mixer gate_output_13_34(.a(output_14_34), .b(output_14_3), .y(output_13_34));
wire output_15_34, output_15_3, output_14_34;
mixer gate_output_14_34(.a(output_15_34), .b(output_15_3), .y(output_14_34));
wire output_16_34, output_16_3, output_15_34;
mixer gate_output_15_34(.a(output_16_34), .b(output_16_3), .y(output_15_34));
wire output_1_35, output_1_4, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_4), .y(output_0_35));
wire output_2_35, output_2_4, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_4), .y(output_1_35));
wire output_3_35, output_3_4, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_4), .y(output_2_35));
wire output_4_35, output_4_4, output_3_35;
mixer gate_output_3_35(.a(output_4_35), .b(output_4_4), .y(output_3_35));
wire output_5_35, output_5_4, output_4_35;
mixer gate_output_4_35(.a(output_5_35), .b(output_5_4), .y(output_4_35));
wire output_6_35, output_6_4, output_5_35;
mixer gate_output_5_35(.a(output_6_35), .b(output_6_4), .y(output_5_35));
wire output_7_35, output_7_4, output_6_35;
mixer gate_output_6_35(.a(output_7_35), .b(output_7_4), .y(output_6_35));
wire output_8_35, output_8_4, output_7_35;
mixer gate_output_7_35(.a(output_8_35), .b(output_8_4), .y(output_7_35));
wire output_9_35, output_9_4, output_8_35;
mixer gate_output_8_35(.a(output_9_35), .b(output_9_4), .y(output_8_35));
wire output_10_35, output_10_4, output_9_35;
mixer gate_output_9_35(.a(output_10_35), .b(output_10_4), .y(output_9_35));
wire output_11_35, output_11_4, output_10_35;
mixer gate_output_10_35(.a(output_11_35), .b(output_11_4), .y(output_10_35));
wire output_12_35, output_12_4, output_11_35;
mixer gate_output_11_35(.a(output_12_35), .b(output_12_4), .y(output_11_35));
wire output_13_35, output_13_4, output_12_35;
mixer gate_output_12_35(.a(output_13_35), .b(output_13_4), .y(output_12_35));
wire output_14_35, output_14_4, output_13_35;
mixer gate_output_13_35(.a(output_14_35), .b(output_14_4), .y(output_13_35));
wire output_15_35, output_15_4, output_14_35;
mixer gate_output_14_35(.a(output_15_35), .b(output_15_4), .y(output_14_35));
wire output_16_35, output_16_4, output_15_35;
mixer gate_output_15_35(.a(output_16_35), .b(output_16_4), .y(output_15_35));
wire output_1_36, output_1_5, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_5), .y(output_0_36));
wire output_2_36, output_2_5, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_5), .y(output_1_36));
wire output_3_36, output_3_5, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_5), .y(output_2_36));
wire output_4_36, output_4_5, output_3_36;
mixer gate_output_3_36(.a(output_4_36), .b(output_4_5), .y(output_3_36));
wire output_5_36, output_5_5, output_4_36;
mixer gate_output_4_36(.a(output_5_36), .b(output_5_5), .y(output_4_36));
wire output_6_36, output_6_5, output_5_36;
mixer gate_output_5_36(.a(output_6_36), .b(output_6_5), .y(output_5_36));
wire output_7_36, output_7_5, output_6_36;
mixer gate_output_6_36(.a(output_7_36), .b(output_7_5), .y(output_6_36));
wire output_8_36, output_8_5, output_7_36;
mixer gate_output_7_36(.a(output_8_36), .b(output_8_5), .y(output_7_36));
wire output_9_36, output_9_5, output_8_36;
mixer gate_output_8_36(.a(output_9_36), .b(output_9_5), .y(output_8_36));
wire output_10_36, output_10_5, output_9_36;
mixer gate_output_9_36(.a(output_10_36), .b(output_10_5), .y(output_9_36));
wire output_11_36, output_11_5, output_10_36;
mixer gate_output_10_36(.a(output_11_36), .b(output_11_5), .y(output_10_36));
wire output_12_36, output_12_5, output_11_36;
mixer gate_output_11_36(.a(output_12_36), .b(output_12_5), .y(output_11_36));
wire output_13_36, output_13_5, output_12_36;
mixer gate_output_12_36(.a(output_13_36), .b(output_13_5), .y(output_12_36));
wire output_14_36, output_14_5, output_13_36;
mixer gate_output_13_36(.a(output_14_36), .b(output_14_5), .y(output_13_36));
wire output_15_36, output_15_5, output_14_36;
mixer gate_output_14_36(.a(output_15_36), .b(output_15_5), .y(output_14_36));
wire output_16_36, output_16_5, output_15_36;
mixer gate_output_15_36(.a(output_16_36), .b(output_16_5), .y(output_15_36));
wire output_1_37, output_1_6, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_6), .y(output_0_37));
wire output_2_37, output_2_6, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_6), .y(output_1_37));
wire output_3_37, output_3_6, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_6), .y(output_2_37));
wire output_4_37, output_4_6, output_3_37;
mixer gate_output_3_37(.a(output_4_37), .b(output_4_6), .y(output_3_37));
wire output_5_37, output_5_6, output_4_37;
mixer gate_output_4_37(.a(output_5_37), .b(output_5_6), .y(output_4_37));
wire output_6_37, output_6_6, output_5_37;
mixer gate_output_5_37(.a(output_6_37), .b(output_6_6), .y(output_5_37));
wire output_7_37, output_7_6, output_6_37;
mixer gate_output_6_37(.a(output_7_37), .b(output_7_6), .y(output_6_37));
wire output_8_37, output_8_6, output_7_37;
mixer gate_output_7_37(.a(output_8_37), .b(output_8_6), .y(output_7_37));
wire output_9_37, output_9_6, output_8_37;
mixer gate_output_8_37(.a(output_9_37), .b(output_9_6), .y(output_8_37));
wire output_10_37, output_10_6, output_9_37;
mixer gate_output_9_37(.a(output_10_37), .b(output_10_6), .y(output_9_37));
wire output_11_37, output_11_6, output_10_37;
mixer gate_output_10_37(.a(output_11_37), .b(output_11_6), .y(output_10_37));
wire output_12_37, output_12_6, output_11_37;
mixer gate_output_11_37(.a(output_12_37), .b(output_12_6), .y(output_11_37));
wire output_13_37, output_13_6, output_12_37;
mixer gate_output_12_37(.a(output_13_37), .b(output_13_6), .y(output_12_37));
wire output_14_37, output_14_6, output_13_37;
mixer gate_output_13_37(.a(output_14_37), .b(output_14_6), .y(output_13_37));
wire output_15_37, output_15_6, output_14_37;
mixer gate_output_14_37(.a(output_15_37), .b(output_15_6), .y(output_14_37));
wire output_16_37, output_16_6, output_15_37;
mixer gate_output_15_37(.a(output_16_37), .b(output_16_6), .y(output_15_37));
wire output_1_38, output_1_7, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_7), .y(output_0_38));
wire output_2_38, output_2_7, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_7), .y(output_1_38));
wire output_3_38, output_3_7, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_7), .y(output_2_38));
wire output_4_38, output_4_7, output_3_38;
mixer gate_output_3_38(.a(output_4_38), .b(output_4_7), .y(output_3_38));
wire output_5_38, output_5_7, output_4_38;
mixer gate_output_4_38(.a(output_5_38), .b(output_5_7), .y(output_4_38));
wire output_6_38, output_6_7, output_5_38;
mixer gate_output_5_38(.a(output_6_38), .b(output_6_7), .y(output_5_38));
wire output_7_38, output_7_7, output_6_38;
mixer gate_output_6_38(.a(output_7_38), .b(output_7_7), .y(output_6_38));
wire output_8_38, output_8_7, output_7_38;
mixer gate_output_7_38(.a(output_8_38), .b(output_8_7), .y(output_7_38));
wire output_9_38, output_9_7, output_8_38;
mixer gate_output_8_38(.a(output_9_38), .b(output_9_7), .y(output_8_38));
wire output_10_38, output_10_7, output_9_38;
mixer gate_output_9_38(.a(output_10_38), .b(output_10_7), .y(output_9_38));
wire output_11_38, output_11_7, output_10_38;
mixer gate_output_10_38(.a(output_11_38), .b(output_11_7), .y(output_10_38));
wire output_12_38, output_12_7, output_11_38;
mixer gate_output_11_38(.a(output_12_38), .b(output_12_7), .y(output_11_38));
wire output_13_38, output_13_7, output_12_38;
mixer gate_output_12_38(.a(output_13_38), .b(output_13_7), .y(output_12_38));
wire output_14_38, output_14_7, output_13_38;
mixer gate_output_13_38(.a(output_14_38), .b(output_14_7), .y(output_13_38));
wire output_15_38, output_15_7, output_14_38;
mixer gate_output_14_38(.a(output_15_38), .b(output_15_7), .y(output_14_38));
wire output_16_38, output_16_7, output_15_38;
mixer gate_output_15_38(.a(output_16_38), .b(output_16_7), .y(output_15_38));
wire output_1_39, output_1_8, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_8), .y(output_0_39));
wire output_2_39, output_2_8, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_8), .y(output_1_39));
wire output_3_39, output_3_8, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_8), .y(output_2_39));
wire output_4_39, output_4_8, output_3_39;
mixer gate_output_3_39(.a(output_4_39), .b(output_4_8), .y(output_3_39));
wire output_5_39, output_5_8, output_4_39;
mixer gate_output_4_39(.a(output_5_39), .b(output_5_8), .y(output_4_39));
wire output_6_39, output_6_8, output_5_39;
mixer gate_output_5_39(.a(output_6_39), .b(output_6_8), .y(output_5_39));
wire output_7_39, output_7_8, output_6_39;
mixer gate_output_6_39(.a(output_7_39), .b(output_7_8), .y(output_6_39));
wire output_8_39, output_8_8, output_7_39;
mixer gate_output_7_39(.a(output_8_39), .b(output_8_8), .y(output_7_39));
wire output_9_39, output_9_8, output_8_39;
mixer gate_output_8_39(.a(output_9_39), .b(output_9_8), .y(output_8_39));
wire output_10_39, output_10_8, output_9_39;
mixer gate_output_9_39(.a(output_10_39), .b(output_10_8), .y(output_9_39));
wire output_11_39, output_11_8, output_10_39;
mixer gate_output_10_39(.a(output_11_39), .b(output_11_8), .y(output_10_39));
wire output_12_39, output_12_8, output_11_39;
mixer gate_output_11_39(.a(output_12_39), .b(output_12_8), .y(output_11_39));
wire output_13_39, output_13_8, output_12_39;
mixer gate_output_12_39(.a(output_13_39), .b(output_13_8), .y(output_12_39));
wire output_14_39, output_14_8, output_13_39;
mixer gate_output_13_39(.a(output_14_39), .b(output_14_8), .y(output_13_39));
wire output_15_39, output_15_8, output_14_39;
mixer gate_output_14_39(.a(output_15_39), .b(output_15_8), .y(output_14_39));
wire output_16_39, output_16_8, output_15_39;
mixer gate_output_15_39(.a(output_16_39), .b(output_16_8), .y(output_15_39));
wire output_1_40, output_1_9, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_9), .y(output_0_40));
wire output_2_40, output_2_9, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_9), .y(output_1_40));
wire output_3_40, output_3_9, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_9), .y(output_2_40));
wire output_4_40, output_4_9, output_3_40;
mixer gate_output_3_40(.a(output_4_40), .b(output_4_9), .y(output_3_40));
wire output_5_40, output_5_9, output_4_40;
mixer gate_output_4_40(.a(output_5_40), .b(output_5_9), .y(output_4_40));
wire output_6_40, output_6_9, output_5_40;
mixer gate_output_5_40(.a(output_6_40), .b(output_6_9), .y(output_5_40));
wire output_7_40, output_7_9, output_6_40;
mixer gate_output_6_40(.a(output_7_40), .b(output_7_9), .y(output_6_40));
wire output_8_40, output_8_9, output_7_40;
mixer gate_output_7_40(.a(output_8_40), .b(output_8_9), .y(output_7_40));
wire output_9_40, output_9_9, output_8_40;
mixer gate_output_8_40(.a(output_9_40), .b(output_9_9), .y(output_8_40));
wire output_10_40, output_10_9, output_9_40;
mixer gate_output_9_40(.a(output_10_40), .b(output_10_9), .y(output_9_40));
wire output_11_40, output_11_9, output_10_40;
mixer gate_output_10_40(.a(output_11_40), .b(output_11_9), .y(output_10_40));
wire output_12_40, output_12_9, output_11_40;
mixer gate_output_11_40(.a(output_12_40), .b(output_12_9), .y(output_11_40));
wire output_13_40, output_13_9, output_12_40;
mixer gate_output_12_40(.a(output_13_40), .b(output_13_9), .y(output_12_40));
wire output_14_40, output_14_9, output_13_40;
mixer gate_output_13_40(.a(output_14_40), .b(output_14_9), .y(output_13_40));
wire output_15_40, output_15_9, output_14_40;
mixer gate_output_14_40(.a(output_15_40), .b(output_15_9), .y(output_14_40));
wire output_16_40, output_16_9, output_15_40;
mixer gate_output_15_40(.a(output_16_40), .b(output_16_9), .y(output_15_40));
wire output_1_41, output_1_10, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_10), .y(output_0_41));
wire output_2_41, output_2_10, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_10), .y(output_1_41));
wire output_3_41, output_3_10, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_10), .y(output_2_41));
wire output_4_41, output_4_10, output_3_41;
mixer gate_output_3_41(.a(output_4_41), .b(output_4_10), .y(output_3_41));
wire output_5_41, output_5_10, output_4_41;
mixer gate_output_4_41(.a(output_5_41), .b(output_5_10), .y(output_4_41));
wire output_6_41, output_6_10, output_5_41;
mixer gate_output_5_41(.a(output_6_41), .b(output_6_10), .y(output_5_41));
wire output_7_41, output_7_10, output_6_41;
mixer gate_output_6_41(.a(output_7_41), .b(output_7_10), .y(output_6_41));
wire output_8_41, output_8_10, output_7_41;
mixer gate_output_7_41(.a(output_8_41), .b(output_8_10), .y(output_7_41));
wire output_9_41, output_9_10, output_8_41;
mixer gate_output_8_41(.a(output_9_41), .b(output_9_10), .y(output_8_41));
wire output_10_41, output_10_10, output_9_41;
mixer gate_output_9_41(.a(output_10_41), .b(output_10_10), .y(output_9_41));
wire output_11_41, output_11_10, output_10_41;
mixer gate_output_10_41(.a(output_11_41), .b(output_11_10), .y(output_10_41));
wire output_12_41, output_12_10, output_11_41;
mixer gate_output_11_41(.a(output_12_41), .b(output_12_10), .y(output_11_41));
wire output_13_41, output_13_10, output_12_41;
mixer gate_output_12_41(.a(output_13_41), .b(output_13_10), .y(output_12_41));
wire output_14_41, output_14_10, output_13_41;
mixer gate_output_13_41(.a(output_14_41), .b(output_14_10), .y(output_13_41));
wire output_15_41, output_15_10, output_14_41;
mixer gate_output_14_41(.a(output_15_41), .b(output_15_10), .y(output_14_41));
wire output_16_41, output_16_10, output_15_41;
mixer gate_output_15_41(.a(output_16_41), .b(output_16_10), .y(output_15_41));
wire output_1_42, output_1_11, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_11), .y(output_0_42));
wire output_2_42, output_2_11, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_11), .y(output_1_42));
wire output_3_42, output_3_11, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_11), .y(output_2_42));
wire output_4_42, output_4_11, output_3_42;
mixer gate_output_3_42(.a(output_4_42), .b(output_4_11), .y(output_3_42));
wire output_5_42, output_5_11, output_4_42;
mixer gate_output_4_42(.a(output_5_42), .b(output_5_11), .y(output_4_42));
wire output_6_42, output_6_11, output_5_42;
mixer gate_output_5_42(.a(output_6_42), .b(output_6_11), .y(output_5_42));
wire output_7_42, output_7_11, output_6_42;
mixer gate_output_6_42(.a(output_7_42), .b(output_7_11), .y(output_6_42));
wire output_8_42, output_8_11, output_7_42;
mixer gate_output_7_42(.a(output_8_42), .b(output_8_11), .y(output_7_42));
wire output_9_42, output_9_11, output_8_42;
mixer gate_output_8_42(.a(output_9_42), .b(output_9_11), .y(output_8_42));
wire output_10_42, output_10_11, output_9_42;
mixer gate_output_9_42(.a(output_10_42), .b(output_10_11), .y(output_9_42));
wire output_11_42, output_11_11, output_10_42;
mixer gate_output_10_42(.a(output_11_42), .b(output_11_11), .y(output_10_42));
wire output_12_42, output_12_11, output_11_42;
mixer gate_output_11_42(.a(output_12_42), .b(output_12_11), .y(output_11_42));
wire output_13_42, output_13_11, output_12_42;
mixer gate_output_12_42(.a(output_13_42), .b(output_13_11), .y(output_12_42));
wire output_14_42, output_14_11, output_13_42;
mixer gate_output_13_42(.a(output_14_42), .b(output_14_11), .y(output_13_42));
wire output_15_42, output_15_11, output_14_42;
mixer gate_output_14_42(.a(output_15_42), .b(output_15_11), .y(output_14_42));
wire output_16_42, output_16_11, output_15_42;
mixer gate_output_15_42(.a(output_16_42), .b(output_16_11), .y(output_15_42));
wire output_1_43, output_1_12, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_12), .y(output_0_43));
wire output_2_43, output_2_12, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_12), .y(output_1_43));
wire output_3_43, output_3_12, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_12), .y(output_2_43));
wire output_4_43, output_4_12, output_3_43;
mixer gate_output_3_43(.a(output_4_43), .b(output_4_12), .y(output_3_43));
wire output_5_43, output_5_12, output_4_43;
mixer gate_output_4_43(.a(output_5_43), .b(output_5_12), .y(output_4_43));
wire output_6_43, output_6_12, output_5_43;
mixer gate_output_5_43(.a(output_6_43), .b(output_6_12), .y(output_5_43));
wire output_7_43, output_7_12, output_6_43;
mixer gate_output_6_43(.a(output_7_43), .b(output_7_12), .y(output_6_43));
wire output_8_43, output_8_12, output_7_43;
mixer gate_output_7_43(.a(output_8_43), .b(output_8_12), .y(output_7_43));
wire output_9_43, output_9_12, output_8_43;
mixer gate_output_8_43(.a(output_9_43), .b(output_9_12), .y(output_8_43));
wire output_10_43, output_10_12, output_9_43;
mixer gate_output_9_43(.a(output_10_43), .b(output_10_12), .y(output_9_43));
wire output_11_43, output_11_12, output_10_43;
mixer gate_output_10_43(.a(output_11_43), .b(output_11_12), .y(output_10_43));
wire output_12_43, output_12_12, output_11_43;
mixer gate_output_11_43(.a(output_12_43), .b(output_12_12), .y(output_11_43));
wire output_13_43, output_13_12, output_12_43;
mixer gate_output_12_43(.a(output_13_43), .b(output_13_12), .y(output_12_43));
wire output_14_43, output_14_12, output_13_43;
mixer gate_output_13_43(.a(output_14_43), .b(output_14_12), .y(output_13_43));
wire output_15_43, output_15_12, output_14_43;
mixer gate_output_14_43(.a(output_15_43), .b(output_15_12), .y(output_14_43));
wire output_16_43, output_16_12, output_15_43;
mixer gate_output_15_43(.a(output_16_43), .b(output_16_12), .y(output_15_43));
wire output_1_44, output_1_13, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_13), .y(output_0_44));
wire output_2_44, output_2_13, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_13), .y(output_1_44));
wire output_3_44, output_3_13, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_13), .y(output_2_44));
wire output_4_44, output_4_13, output_3_44;
mixer gate_output_3_44(.a(output_4_44), .b(output_4_13), .y(output_3_44));
wire output_5_44, output_5_13, output_4_44;
mixer gate_output_4_44(.a(output_5_44), .b(output_5_13), .y(output_4_44));
wire output_6_44, output_6_13, output_5_44;
mixer gate_output_5_44(.a(output_6_44), .b(output_6_13), .y(output_5_44));
wire output_7_44, output_7_13, output_6_44;
mixer gate_output_6_44(.a(output_7_44), .b(output_7_13), .y(output_6_44));
wire output_8_44, output_8_13, output_7_44;
mixer gate_output_7_44(.a(output_8_44), .b(output_8_13), .y(output_7_44));
wire output_9_44, output_9_13, output_8_44;
mixer gate_output_8_44(.a(output_9_44), .b(output_9_13), .y(output_8_44));
wire output_10_44, output_10_13, output_9_44;
mixer gate_output_9_44(.a(output_10_44), .b(output_10_13), .y(output_9_44));
wire output_11_44, output_11_13, output_10_44;
mixer gate_output_10_44(.a(output_11_44), .b(output_11_13), .y(output_10_44));
wire output_12_44, output_12_13, output_11_44;
mixer gate_output_11_44(.a(output_12_44), .b(output_12_13), .y(output_11_44));
wire output_13_44, output_13_13, output_12_44;
mixer gate_output_12_44(.a(output_13_44), .b(output_13_13), .y(output_12_44));
wire output_14_44, output_14_13, output_13_44;
mixer gate_output_13_44(.a(output_14_44), .b(output_14_13), .y(output_13_44));
wire output_15_44, output_15_13, output_14_44;
mixer gate_output_14_44(.a(output_15_44), .b(output_15_13), .y(output_14_44));
wire output_16_44, output_16_13, output_15_44;
mixer gate_output_15_44(.a(output_16_44), .b(output_16_13), .y(output_15_44));
wire output_1_45, output_1_14, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_14), .y(output_0_45));
wire output_2_45, output_2_14, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_14), .y(output_1_45));
wire output_3_45, output_3_14, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_14), .y(output_2_45));
wire output_4_45, output_4_14, output_3_45;
mixer gate_output_3_45(.a(output_4_45), .b(output_4_14), .y(output_3_45));
wire output_5_45, output_5_14, output_4_45;
mixer gate_output_4_45(.a(output_5_45), .b(output_5_14), .y(output_4_45));
wire output_6_45, output_6_14, output_5_45;
mixer gate_output_5_45(.a(output_6_45), .b(output_6_14), .y(output_5_45));
wire output_7_45, output_7_14, output_6_45;
mixer gate_output_6_45(.a(output_7_45), .b(output_7_14), .y(output_6_45));
wire output_8_45, output_8_14, output_7_45;
mixer gate_output_7_45(.a(output_8_45), .b(output_8_14), .y(output_7_45));
wire output_9_45, output_9_14, output_8_45;
mixer gate_output_8_45(.a(output_9_45), .b(output_9_14), .y(output_8_45));
wire output_10_45, output_10_14, output_9_45;
mixer gate_output_9_45(.a(output_10_45), .b(output_10_14), .y(output_9_45));
wire output_11_45, output_11_14, output_10_45;
mixer gate_output_10_45(.a(output_11_45), .b(output_11_14), .y(output_10_45));
wire output_12_45, output_12_14, output_11_45;
mixer gate_output_11_45(.a(output_12_45), .b(output_12_14), .y(output_11_45));
wire output_13_45, output_13_14, output_12_45;
mixer gate_output_12_45(.a(output_13_45), .b(output_13_14), .y(output_12_45));
wire output_14_45, output_14_14, output_13_45;
mixer gate_output_13_45(.a(output_14_45), .b(output_14_14), .y(output_13_45));
wire output_15_45, output_15_14, output_14_45;
mixer gate_output_14_45(.a(output_15_45), .b(output_15_14), .y(output_14_45));
wire output_16_45, output_16_14, output_15_45;
mixer gate_output_15_45(.a(output_16_45), .b(output_16_14), .y(output_15_45));
wire output_1_46, output_1_15, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_15), .y(output_0_46));
wire output_2_46, output_2_15, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_15), .y(output_1_46));
wire output_3_46, output_3_15, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_15), .y(output_2_46));
wire output_4_46, output_4_15, output_3_46;
mixer gate_output_3_46(.a(output_4_46), .b(output_4_15), .y(output_3_46));
wire output_5_46, output_5_15, output_4_46;
mixer gate_output_4_46(.a(output_5_46), .b(output_5_15), .y(output_4_46));
wire output_6_46, output_6_15, output_5_46;
mixer gate_output_5_46(.a(output_6_46), .b(output_6_15), .y(output_5_46));
wire output_7_46, output_7_15, output_6_46;
mixer gate_output_6_46(.a(output_7_46), .b(output_7_15), .y(output_6_46));
wire output_8_46, output_8_15, output_7_46;
mixer gate_output_7_46(.a(output_8_46), .b(output_8_15), .y(output_7_46));
wire output_9_46, output_9_15, output_8_46;
mixer gate_output_8_46(.a(output_9_46), .b(output_9_15), .y(output_8_46));
wire output_10_46, output_10_15, output_9_46;
mixer gate_output_9_46(.a(output_10_46), .b(output_10_15), .y(output_9_46));
wire output_11_46, output_11_15, output_10_46;
mixer gate_output_10_46(.a(output_11_46), .b(output_11_15), .y(output_10_46));
wire output_12_46, output_12_15, output_11_46;
mixer gate_output_11_46(.a(output_12_46), .b(output_12_15), .y(output_11_46));
wire output_13_46, output_13_15, output_12_46;
mixer gate_output_12_46(.a(output_13_46), .b(output_13_15), .y(output_12_46));
wire output_14_46, output_14_15, output_13_46;
mixer gate_output_13_46(.a(output_14_46), .b(output_14_15), .y(output_13_46));
wire output_15_46, output_15_15, output_14_46;
mixer gate_output_14_46(.a(output_15_46), .b(output_15_15), .y(output_14_46));
wire output_16_46, output_16_15, output_15_46;
mixer gate_output_15_46(.a(output_16_46), .b(output_16_15), .y(output_15_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_4_47, output_4_0, output_3_47;
mixer gate_output_3_47(.a(output_4_47), .b(output_4_0), .y(output_3_47));
wire output_5_47, output_5_0, output_4_47;
mixer gate_output_4_47(.a(output_5_47), .b(output_5_0), .y(output_4_47));
wire output_6_47, output_6_0, output_5_47;
mixer gate_output_5_47(.a(output_6_47), .b(output_6_0), .y(output_5_47));
wire output_7_47, output_7_0, output_6_47;
mixer gate_output_6_47(.a(output_7_47), .b(output_7_0), .y(output_6_47));
wire output_8_47, output_8_0, output_7_47;
mixer gate_output_7_47(.a(output_8_47), .b(output_8_0), .y(output_7_47));
wire output_9_47, output_9_0, output_8_47;
mixer gate_output_8_47(.a(output_9_47), .b(output_9_0), .y(output_8_47));
wire output_10_47, output_10_0, output_9_47;
mixer gate_output_9_47(.a(output_10_47), .b(output_10_0), .y(output_9_47));
wire output_11_47, output_11_0, output_10_47;
mixer gate_output_10_47(.a(output_11_47), .b(output_11_0), .y(output_10_47));
wire output_12_47, output_12_0, output_11_47;
mixer gate_output_11_47(.a(output_12_47), .b(output_12_0), .y(output_11_47));
wire output_13_47, output_13_0, output_12_47;
mixer gate_output_12_47(.a(output_13_47), .b(output_13_0), .y(output_12_47));
wire output_14_47, output_14_0, output_13_47;
mixer gate_output_13_47(.a(output_14_47), .b(output_14_0), .y(output_13_47));
wire output_15_47, output_15_0, output_14_47;
mixer gate_output_14_47(.a(output_15_47), .b(output_15_0), .y(output_14_47));
wire output_16_47, output_16_0, output_15_47;
mixer gate_output_15_47(.a(output_16_47), .b(output_16_0), .y(output_15_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_4_48, output_4_1, output_3_48;
mixer gate_output_3_48(.a(output_4_48), .b(output_4_1), .y(output_3_48));
wire output_5_48, output_5_1, output_4_48;
mixer gate_output_4_48(.a(output_5_48), .b(output_5_1), .y(output_4_48));
wire output_6_48, output_6_1, output_5_48;
mixer gate_output_5_48(.a(output_6_48), .b(output_6_1), .y(output_5_48));
wire output_7_48, output_7_1, output_6_48;
mixer gate_output_6_48(.a(output_7_48), .b(output_7_1), .y(output_6_48));
wire output_8_48, output_8_1, output_7_48;
mixer gate_output_7_48(.a(output_8_48), .b(output_8_1), .y(output_7_48));
wire output_9_48, output_9_1, output_8_48;
mixer gate_output_8_48(.a(output_9_48), .b(output_9_1), .y(output_8_48));
wire output_10_48, output_10_1, output_9_48;
mixer gate_output_9_48(.a(output_10_48), .b(output_10_1), .y(output_9_48));
wire output_11_48, output_11_1, output_10_48;
mixer gate_output_10_48(.a(output_11_48), .b(output_11_1), .y(output_10_48));
wire output_12_48, output_12_1, output_11_48;
mixer gate_output_11_48(.a(output_12_48), .b(output_12_1), .y(output_11_48));
wire output_13_48, output_13_1, output_12_48;
mixer gate_output_12_48(.a(output_13_48), .b(output_13_1), .y(output_12_48));
wire output_14_48, output_14_1, output_13_48;
mixer gate_output_13_48(.a(output_14_48), .b(output_14_1), .y(output_13_48));
wire output_15_48, output_15_1, output_14_48;
mixer gate_output_14_48(.a(output_15_48), .b(output_15_1), .y(output_14_48));
wire output_16_48, output_16_1, output_15_48;
mixer gate_output_15_48(.a(output_16_48), .b(output_16_1), .y(output_15_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_4_49, output_4_2, output_3_49;
mixer gate_output_3_49(.a(output_4_49), .b(output_4_2), .y(output_3_49));
wire output_5_49, output_5_2, output_4_49;
mixer gate_output_4_49(.a(output_5_49), .b(output_5_2), .y(output_4_49));
wire output_6_49, output_6_2, output_5_49;
mixer gate_output_5_49(.a(output_6_49), .b(output_6_2), .y(output_5_49));
wire output_7_49, output_7_2, output_6_49;
mixer gate_output_6_49(.a(output_7_49), .b(output_7_2), .y(output_6_49));
wire output_8_49, output_8_2, output_7_49;
mixer gate_output_7_49(.a(output_8_49), .b(output_8_2), .y(output_7_49));
wire output_9_49, output_9_2, output_8_49;
mixer gate_output_8_49(.a(output_9_49), .b(output_9_2), .y(output_8_49));
wire output_10_49, output_10_2, output_9_49;
mixer gate_output_9_49(.a(output_10_49), .b(output_10_2), .y(output_9_49));
wire output_11_49, output_11_2, output_10_49;
mixer gate_output_10_49(.a(output_11_49), .b(output_11_2), .y(output_10_49));
wire output_12_49, output_12_2, output_11_49;
mixer gate_output_11_49(.a(output_12_49), .b(output_12_2), .y(output_11_49));
wire output_13_49, output_13_2, output_12_49;
mixer gate_output_12_49(.a(output_13_49), .b(output_13_2), .y(output_12_49));
wire output_14_49, output_14_2, output_13_49;
mixer gate_output_13_49(.a(output_14_49), .b(output_14_2), .y(output_13_49));
wire output_15_49, output_15_2, output_14_49;
mixer gate_output_14_49(.a(output_15_49), .b(output_15_2), .y(output_14_49));
wire output_16_49, output_16_2, output_15_49;
mixer gate_output_15_49(.a(output_16_49), .b(output_16_2), .y(output_15_49));
wire output_1_50, output_1_3, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_3), .y(output_0_50));
wire output_2_50, output_2_3, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_3), .y(output_1_50));
wire output_3_50, output_3_3, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_3), .y(output_2_50));
wire output_4_50, output_4_3, output_3_50;
mixer gate_output_3_50(.a(output_4_50), .b(output_4_3), .y(output_3_50));
wire output_5_50, output_5_3, output_4_50;
mixer gate_output_4_50(.a(output_5_50), .b(output_5_3), .y(output_4_50));
wire output_6_50, output_6_3, output_5_50;
mixer gate_output_5_50(.a(output_6_50), .b(output_6_3), .y(output_5_50));
wire output_7_50, output_7_3, output_6_50;
mixer gate_output_6_50(.a(output_7_50), .b(output_7_3), .y(output_6_50));
wire output_8_50, output_8_3, output_7_50;
mixer gate_output_7_50(.a(output_8_50), .b(output_8_3), .y(output_7_50));
wire output_9_50, output_9_3, output_8_50;
mixer gate_output_8_50(.a(output_9_50), .b(output_9_3), .y(output_8_50));
wire output_10_50, output_10_3, output_9_50;
mixer gate_output_9_50(.a(output_10_50), .b(output_10_3), .y(output_9_50));
wire output_11_50, output_11_3, output_10_50;
mixer gate_output_10_50(.a(output_11_50), .b(output_11_3), .y(output_10_50));
wire output_12_50, output_12_3, output_11_50;
mixer gate_output_11_50(.a(output_12_50), .b(output_12_3), .y(output_11_50));
wire output_13_50, output_13_3, output_12_50;
mixer gate_output_12_50(.a(output_13_50), .b(output_13_3), .y(output_12_50));
wire output_14_50, output_14_3, output_13_50;
mixer gate_output_13_50(.a(output_14_50), .b(output_14_3), .y(output_13_50));
wire output_15_50, output_15_3, output_14_50;
mixer gate_output_14_50(.a(output_15_50), .b(output_15_3), .y(output_14_50));
wire output_16_50, output_16_3, output_15_50;
mixer gate_output_15_50(.a(output_16_50), .b(output_16_3), .y(output_15_50));
wire output_1_51, output_1_4, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_4), .y(output_0_51));
wire output_2_51, output_2_4, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_4), .y(output_1_51));
wire output_3_51, output_3_4, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_4), .y(output_2_51));
wire output_4_51, output_4_4, output_3_51;
mixer gate_output_3_51(.a(output_4_51), .b(output_4_4), .y(output_3_51));
wire output_5_51, output_5_4, output_4_51;
mixer gate_output_4_51(.a(output_5_51), .b(output_5_4), .y(output_4_51));
wire output_6_51, output_6_4, output_5_51;
mixer gate_output_5_51(.a(output_6_51), .b(output_6_4), .y(output_5_51));
wire output_7_51, output_7_4, output_6_51;
mixer gate_output_6_51(.a(output_7_51), .b(output_7_4), .y(output_6_51));
wire output_8_51, output_8_4, output_7_51;
mixer gate_output_7_51(.a(output_8_51), .b(output_8_4), .y(output_7_51));
wire output_9_51, output_9_4, output_8_51;
mixer gate_output_8_51(.a(output_9_51), .b(output_9_4), .y(output_8_51));
wire output_10_51, output_10_4, output_9_51;
mixer gate_output_9_51(.a(output_10_51), .b(output_10_4), .y(output_9_51));
wire output_11_51, output_11_4, output_10_51;
mixer gate_output_10_51(.a(output_11_51), .b(output_11_4), .y(output_10_51));
wire output_12_51, output_12_4, output_11_51;
mixer gate_output_11_51(.a(output_12_51), .b(output_12_4), .y(output_11_51));
wire output_13_51, output_13_4, output_12_51;
mixer gate_output_12_51(.a(output_13_51), .b(output_13_4), .y(output_12_51));
wire output_14_51, output_14_4, output_13_51;
mixer gate_output_13_51(.a(output_14_51), .b(output_14_4), .y(output_13_51));
wire output_15_51, output_15_4, output_14_51;
mixer gate_output_14_51(.a(output_15_51), .b(output_15_4), .y(output_14_51));
wire output_16_51, output_16_4, output_15_51;
mixer gate_output_15_51(.a(output_16_51), .b(output_16_4), .y(output_15_51));
wire output_1_52, output_1_5, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_5), .y(output_0_52));
wire output_2_52, output_2_5, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_5), .y(output_1_52));
wire output_3_52, output_3_5, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_5), .y(output_2_52));
wire output_4_52, output_4_5, output_3_52;
mixer gate_output_3_52(.a(output_4_52), .b(output_4_5), .y(output_3_52));
wire output_5_52, output_5_5, output_4_52;
mixer gate_output_4_52(.a(output_5_52), .b(output_5_5), .y(output_4_52));
wire output_6_52, output_6_5, output_5_52;
mixer gate_output_5_52(.a(output_6_52), .b(output_6_5), .y(output_5_52));
wire output_7_52, output_7_5, output_6_52;
mixer gate_output_6_52(.a(output_7_52), .b(output_7_5), .y(output_6_52));
wire output_8_52, output_8_5, output_7_52;
mixer gate_output_7_52(.a(output_8_52), .b(output_8_5), .y(output_7_52));
wire output_9_52, output_9_5, output_8_52;
mixer gate_output_8_52(.a(output_9_52), .b(output_9_5), .y(output_8_52));
wire output_10_52, output_10_5, output_9_52;
mixer gate_output_9_52(.a(output_10_52), .b(output_10_5), .y(output_9_52));
wire output_11_52, output_11_5, output_10_52;
mixer gate_output_10_52(.a(output_11_52), .b(output_11_5), .y(output_10_52));
wire output_12_52, output_12_5, output_11_52;
mixer gate_output_11_52(.a(output_12_52), .b(output_12_5), .y(output_11_52));
wire output_13_52, output_13_5, output_12_52;
mixer gate_output_12_52(.a(output_13_52), .b(output_13_5), .y(output_12_52));
wire output_14_52, output_14_5, output_13_52;
mixer gate_output_13_52(.a(output_14_52), .b(output_14_5), .y(output_13_52));
wire output_15_52, output_15_5, output_14_52;
mixer gate_output_14_52(.a(output_15_52), .b(output_15_5), .y(output_14_52));
wire output_16_52, output_16_5, output_15_52;
mixer gate_output_15_52(.a(output_16_52), .b(output_16_5), .y(output_15_52));
wire output_1_53, output_1_6, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_6), .y(output_0_53));
wire output_2_53, output_2_6, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_6), .y(output_1_53));
wire output_3_53, output_3_6, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_6), .y(output_2_53));
wire output_4_53, output_4_6, output_3_53;
mixer gate_output_3_53(.a(output_4_53), .b(output_4_6), .y(output_3_53));
wire output_5_53, output_5_6, output_4_53;
mixer gate_output_4_53(.a(output_5_53), .b(output_5_6), .y(output_4_53));
wire output_6_53, output_6_6, output_5_53;
mixer gate_output_5_53(.a(output_6_53), .b(output_6_6), .y(output_5_53));
wire output_7_53, output_7_6, output_6_53;
mixer gate_output_6_53(.a(output_7_53), .b(output_7_6), .y(output_6_53));
wire output_8_53, output_8_6, output_7_53;
mixer gate_output_7_53(.a(output_8_53), .b(output_8_6), .y(output_7_53));
wire output_9_53, output_9_6, output_8_53;
mixer gate_output_8_53(.a(output_9_53), .b(output_9_6), .y(output_8_53));
wire output_10_53, output_10_6, output_9_53;
mixer gate_output_9_53(.a(output_10_53), .b(output_10_6), .y(output_9_53));
wire output_11_53, output_11_6, output_10_53;
mixer gate_output_10_53(.a(output_11_53), .b(output_11_6), .y(output_10_53));
wire output_12_53, output_12_6, output_11_53;
mixer gate_output_11_53(.a(output_12_53), .b(output_12_6), .y(output_11_53));
wire output_13_53, output_13_6, output_12_53;
mixer gate_output_12_53(.a(output_13_53), .b(output_13_6), .y(output_12_53));
wire output_14_53, output_14_6, output_13_53;
mixer gate_output_13_53(.a(output_14_53), .b(output_14_6), .y(output_13_53));
wire output_15_53, output_15_6, output_14_53;
mixer gate_output_14_53(.a(output_15_53), .b(output_15_6), .y(output_14_53));
wire output_16_53, output_16_6, output_15_53;
mixer gate_output_15_53(.a(output_16_53), .b(output_16_6), .y(output_15_53));
wire output_1_54, output_1_7, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_7), .y(output_0_54));
wire output_2_54, output_2_7, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_7), .y(output_1_54));
wire output_3_54, output_3_7, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_7), .y(output_2_54));
wire output_4_54, output_4_7, output_3_54;
mixer gate_output_3_54(.a(output_4_54), .b(output_4_7), .y(output_3_54));
wire output_5_54, output_5_7, output_4_54;
mixer gate_output_4_54(.a(output_5_54), .b(output_5_7), .y(output_4_54));
wire output_6_54, output_6_7, output_5_54;
mixer gate_output_5_54(.a(output_6_54), .b(output_6_7), .y(output_5_54));
wire output_7_54, output_7_7, output_6_54;
mixer gate_output_6_54(.a(output_7_54), .b(output_7_7), .y(output_6_54));
wire output_8_54, output_8_7, output_7_54;
mixer gate_output_7_54(.a(output_8_54), .b(output_8_7), .y(output_7_54));
wire output_9_54, output_9_7, output_8_54;
mixer gate_output_8_54(.a(output_9_54), .b(output_9_7), .y(output_8_54));
wire output_10_54, output_10_7, output_9_54;
mixer gate_output_9_54(.a(output_10_54), .b(output_10_7), .y(output_9_54));
wire output_11_54, output_11_7, output_10_54;
mixer gate_output_10_54(.a(output_11_54), .b(output_11_7), .y(output_10_54));
wire output_12_54, output_12_7, output_11_54;
mixer gate_output_11_54(.a(output_12_54), .b(output_12_7), .y(output_11_54));
wire output_13_54, output_13_7, output_12_54;
mixer gate_output_12_54(.a(output_13_54), .b(output_13_7), .y(output_12_54));
wire output_14_54, output_14_7, output_13_54;
mixer gate_output_13_54(.a(output_14_54), .b(output_14_7), .y(output_13_54));
wire output_15_54, output_15_7, output_14_54;
mixer gate_output_14_54(.a(output_15_54), .b(output_15_7), .y(output_14_54));
wire output_16_54, output_16_7, output_15_54;
mixer gate_output_15_54(.a(output_16_54), .b(output_16_7), .y(output_15_54));
wire output_1_55, output_1_8, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_8), .y(output_0_55));
wire output_2_55, output_2_8, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_8), .y(output_1_55));
wire output_3_55, output_3_8, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_8), .y(output_2_55));
wire output_4_55, output_4_8, output_3_55;
mixer gate_output_3_55(.a(output_4_55), .b(output_4_8), .y(output_3_55));
wire output_5_55, output_5_8, output_4_55;
mixer gate_output_4_55(.a(output_5_55), .b(output_5_8), .y(output_4_55));
wire output_6_55, output_6_8, output_5_55;
mixer gate_output_5_55(.a(output_6_55), .b(output_6_8), .y(output_5_55));
wire output_7_55, output_7_8, output_6_55;
mixer gate_output_6_55(.a(output_7_55), .b(output_7_8), .y(output_6_55));
wire output_8_55, output_8_8, output_7_55;
mixer gate_output_7_55(.a(output_8_55), .b(output_8_8), .y(output_7_55));
wire output_9_55, output_9_8, output_8_55;
mixer gate_output_8_55(.a(output_9_55), .b(output_9_8), .y(output_8_55));
wire output_10_55, output_10_8, output_9_55;
mixer gate_output_9_55(.a(output_10_55), .b(output_10_8), .y(output_9_55));
wire output_11_55, output_11_8, output_10_55;
mixer gate_output_10_55(.a(output_11_55), .b(output_11_8), .y(output_10_55));
wire output_12_55, output_12_8, output_11_55;
mixer gate_output_11_55(.a(output_12_55), .b(output_12_8), .y(output_11_55));
wire output_13_55, output_13_8, output_12_55;
mixer gate_output_12_55(.a(output_13_55), .b(output_13_8), .y(output_12_55));
wire output_14_55, output_14_8, output_13_55;
mixer gate_output_13_55(.a(output_14_55), .b(output_14_8), .y(output_13_55));
wire output_15_55, output_15_8, output_14_55;
mixer gate_output_14_55(.a(output_15_55), .b(output_15_8), .y(output_14_55));
wire output_16_55, output_16_8, output_15_55;
mixer gate_output_15_55(.a(output_16_55), .b(output_16_8), .y(output_15_55));
wire output_1_56, output_1_9, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_9), .y(output_0_56));
wire output_2_56, output_2_9, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_9), .y(output_1_56));
wire output_3_56, output_3_9, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_9), .y(output_2_56));
wire output_4_56, output_4_9, output_3_56;
mixer gate_output_3_56(.a(output_4_56), .b(output_4_9), .y(output_3_56));
wire output_5_56, output_5_9, output_4_56;
mixer gate_output_4_56(.a(output_5_56), .b(output_5_9), .y(output_4_56));
wire output_6_56, output_6_9, output_5_56;
mixer gate_output_5_56(.a(output_6_56), .b(output_6_9), .y(output_5_56));
wire output_7_56, output_7_9, output_6_56;
mixer gate_output_6_56(.a(output_7_56), .b(output_7_9), .y(output_6_56));
wire output_8_56, output_8_9, output_7_56;
mixer gate_output_7_56(.a(output_8_56), .b(output_8_9), .y(output_7_56));
wire output_9_56, output_9_9, output_8_56;
mixer gate_output_8_56(.a(output_9_56), .b(output_9_9), .y(output_8_56));
wire output_10_56, output_10_9, output_9_56;
mixer gate_output_9_56(.a(output_10_56), .b(output_10_9), .y(output_9_56));
wire output_11_56, output_11_9, output_10_56;
mixer gate_output_10_56(.a(output_11_56), .b(output_11_9), .y(output_10_56));
wire output_12_56, output_12_9, output_11_56;
mixer gate_output_11_56(.a(output_12_56), .b(output_12_9), .y(output_11_56));
wire output_13_56, output_13_9, output_12_56;
mixer gate_output_12_56(.a(output_13_56), .b(output_13_9), .y(output_12_56));
wire output_14_56, output_14_9, output_13_56;
mixer gate_output_13_56(.a(output_14_56), .b(output_14_9), .y(output_13_56));
wire output_15_56, output_15_9, output_14_56;
mixer gate_output_14_56(.a(output_15_56), .b(output_15_9), .y(output_14_56));
wire output_16_56, output_16_9, output_15_56;
mixer gate_output_15_56(.a(output_16_56), .b(output_16_9), .y(output_15_56));
wire output_1_57, output_1_10, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_10), .y(output_0_57));
wire output_2_57, output_2_10, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_10), .y(output_1_57));
wire output_3_57, output_3_10, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_10), .y(output_2_57));
wire output_4_57, output_4_10, output_3_57;
mixer gate_output_3_57(.a(output_4_57), .b(output_4_10), .y(output_3_57));
wire output_5_57, output_5_10, output_4_57;
mixer gate_output_4_57(.a(output_5_57), .b(output_5_10), .y(output_4_57));
wire output_6_57, output_6_10, output_5_57;
mixer gate_output_5_57(.a(output_6_57), .b(output_6_10), .y(output_5_57));
wire output_7_57, output_7_10, output_6_57;
mixer gate_output_6_57(.a(output_7_57), .b(output_7_10), .y(output_6_57));
wire output_8_57, output_8_10, output_7_57;
mixer gate_output_7_57(.a(output_8_57), .b(output_8_10), .y(output_7_57));
wire output_9_57, output_9_10, output_8_57;
mixer gate_output_8_57(.a(output_9_57), .b(output_9_10), .y(output_8_57));
wire output_10_57, output_10_10, output_9_57;
mixer gate_output_9_57(.a(output_10_57), .b(output_10_10), .y(output_9_57));
wire output_11_57, output_11_10, output_10_57;
mixer gate_output_10_57(.a(output_11_57), .b(output_11_10), .y(output_10_57));
wire output_12_57, output_12_10, output_11_57;
mixer gate_output_11_57(.a(output_12_57), .b(output_12_10), .y(output_11_57));
wire output_13_57, output_13_10, output_12_57;
mixer gate_output_12_57(.a(output_13_57), .b(output_13_10), .y(output_12_57));
wire output_14_57, output_14_10, output_13_57;
mixer gate_output_13_57(.a(output_14_57), .b(output_14_10), .y(output_13_57));
wire output_15_57, output_15_10, output_14_57;
mixer gate_output_14_57(.a(output_15_57), .b(output_15_10), .y(output_14_57));
wire output_16_57, output_16_10, output_15_57;
mixer gate_output_15_57(.a(output_16_57), .b(output_16_10), .y(output_15_57));
wire output_1_58, output_1_11, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_11), .y(output_0_58));
wire output_2_58, output_2_11, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_11), .y(output_1_58));
wire output_3_58, output_3_11, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_11), .y(output_2_58));
wire output_4_58, output_4_11, output_3_58;
mixer gate_output_3_58(.a(output_4_58), .b(output_4_11), .y(output_3_58));
wire output_5_58, output_5_11, output_4_58;
mixer gate_output_4_58(.a(output_5_58), .b(output_5_11), .y(output_4_58));
wire output_6_58, output_6_11, output_5_58;
mixer gate_output_5_58(.a(output_6_58), .b(output_6_11), .y(output_5_58));
wire output_7_58, output_7_11, output_6_58;
mixer gate_output_6_58(.a(output_7_58), .b(output_7_11), .y(output_6_58));
wire output_8_58, output_8_11, output_7_58;
mixer gate_output_7_58(.a(output_8_58), .b(output_8_11), .y(output_7_58));
wire output_9_58, output_9_11, output_8_58;
mixer gate_output_8_58(.a(output_9_58), .b(output_9_11), .y(output_8_58));
wire output_10_58, output_10_11, output_9_58;
mixer gate_output_9_58(.a(output_10_58), .b(output_10_11), .y(output_9_58));
wire output_11_58, output_11_11, output_10_58;
mixer gate_output_10_58(.a(output_11_58), .b(output_11_11), .y(output_10_58));
wire output_12_58, output_12_11, output_11_58;
mixer gate_output_11_58(.a(output_12_58), .b(output_12_11), .y(output_11_58));
wire output_13_58, output_13_11, output_12_58;
mixer gate_output_12_58(.a(output_13_58), .b(output_13_11), .y(output_12_58));
wire output_14_58, output_14_11, output_13_58;
mixer gate_output_13_58(.a(output_14_58), .b(output_14_11), .y(output_13_58));
wire output_15_58, output_15_11, output_14_58;
mixer gate_output_14_58(.a(output_15_58), .b(output_15_11), .y(output_14_58));
wire output_16_58, output_16_11, output_15_58;
mixer gate_output_15_58(.a(output_16_58), .b(output_16_11), .y(output_15_58));
wire output_1_59, output_1_12, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_12), .y(output_0_59));
wire output_2_59, output_2_12, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_12), .y(output_1_59));
wire output_3_59, output_3_12, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_12), .y(output_2_59));
wire output_4_59, output_4_12, output_3_59;
mixer gate_output_3_59(.a(output_4_59), .b(output_4_12), .y(output_3_59));
wire output_5_59, output_5_12, output_4_59;
mixer gate_output_4_59(.a(output_5_59), .b(output_5_12), .y(output_4_59));
wire output_6_59, output_6_12, output_5_59;
mixer gate_output_5_59(.a(output_6_59), .b(output_6_12), .y(output_5_59));
wire output_7_59, output_7_12, output_6_59;
mixer gate_output_6_59(.a(output_7_59), .b(output_7_12), .y(output_6_59));
wire output_8_59, output_8_12, output_7_59;
mixer gate_output_7_59(.a(output_8_59), .b(output_8_12), .y(output_7_59));
wire output_9_59, output_9_12, output_8_59;
mixer gate_output_8_59(.a(output_9_59), .b(output_9_12), .y(output_8_59));
wire output_10_59, output_10_12, output_9_59;
mixer gate_output_9_59(.a(output_10_59), .b(output_10_12), .y(output_9_59));
wire output_11_59, output_11_12, output_10_59;
mixer gate_output_10_59(.a(output_11_59), .b(output_11_12), .y(output_10_59));
wire output_12_59, output_12_12, output_11_59;
mixer gate_output_11_59(.a(output_12_59), .b(output_12_12), .y(output_11_59));
wire output_13_59, output_13_12, output_12_59;
mixer gate_output_12_59(.a(output_13_59), .b(output_13_12), .y(output_12_59));
wire output_14_59, output_14_12, output_13_59;
mixer gate_output_13_59(.a(output_14_59), .b(output_14_12), .y(output_13_59));
wire output_15_59, output_15_12, output_14_59;
mixer gate_output_14_59(.a(output_15_59), .b(output_15_12), .y(output_14_59));
wire output_16_59, output_16_12, output_15_59;
mixer gate_output_15_59(.a(output_16_59), .b(output_16_12), .y(output_15_59));
wire output_1_60, output_1_13, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_13), .y(output_0_60));
wire output_2_60, output_2_13, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_13), .y(output_1_60));
wire output_3_60, output_3_13, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_13), .y(output_2_60));
wire output_4_60, output_4_13, output_3_60;
mixer gate_output_3_60(.a(output_4_60), .b(output_4_13), .y(output_3_60));
wire output_5_60, output_5_13, output_4_60;
mixer gate_output_4_60(.a(output_5_60), .b(output_5_13), .y(output_4_60));
wire output_6_60, output_6_13, output_5_60;
mixer gate_output_5_60(.a(output_6_60), .b(output_6_13), .y(output_5_60));
wire output_7_60, output_7_13, output_6_60;
mixer gate_output_6_60(.a(output_7_60), .b(output_7_13), .y(output_6_60));
wire output_8_60, output_8_13, output_7_60;
mixer gate_output_7_60(.a(output_8_60), .b(output_8_13), .y(output_7_60));
wire output_9_60, output_9_13, output_8_60;
mixer gate_output_8_60(.a(output_9_60), .b(output_9_13), .y(output_8_60));
wire output_10_60, output_10_13, output_9_60;
mixer gate_output_9_60(.a(output_10_60), .b(output_10_13), .y(output_9_60));
wire output_11_60, output_11_13, output_10_60;
mixer gate_output_10_60(.a(output_11_60), .b(output_11_13), .y(output_10_60));
wire output_12_60, output_12_13, output_11_60;
mixer gate_output_11_60(.a(output_12_60), .b(output_12_13), .y(output_11_60));
wire output_13_60, output_13_13, output_12_60;
mixer gate_output_12_60(.a(output_13_60), .b(output_13_13), .y(output_12_60));
wire output_14_60, output_14_13, output_13_60;
mixer gate_output_13_60(.a(output_14_60), .b(output_14_13), .y(output_13_60));
wire output_15_60, output_15_13, output_14_60;
mixer gate_output_14_60(.a(output_15_60), .b(output_15_13), .y(output_14_60));
wire output_16_60, output_16_13, output_15_60;
mixer gate_output_15_60(.a(output_16_60), .b(output_16_13), .y(output_15_60));
wire output_1_61, output_1_14, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_14), .y(output_0_61));
wire output_2_61, output_2_14, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_14), .y(output_1_61));
wire output_3_61, output_3_14, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_14), .y(output_2_61));
wire output_4_61, output_4_14, output_3_61;
mixer gate_output_3_61(.a(output_4_61), .b(output_4_14), .y(output_3_61));
wire output_5_61, output_5_14, output_4_61;
mixer gate_output_4_61(.a(output_5_61), .b(output_5_14), .y(output_4_61));
wire output_6_61, output_6_14, output_5_61;
mixer gate_output_5_61(.a(output_6_61), .b(output_6_14), .y(output_5_61));
wire output_7_61, output_7_14, output_6_61;
mixer gate_output_6_61(.a(output_7_61), .b(output_7_14), .y(output_6_61));
wire output_8_61, output_8_14, output_7_61;
mixer gate_output_7_61(.a(output_8_61), .b(output_8_14), .y(output_7_61));
wire output_9_61, output_9_14, output_8_61;
mixer gate_output_8_61(.a(output_9_61), .b(output_9_14), .y(output_8_61));
wire output_10_61, output_10_14, output_9_61;
mixer gate_output_9_61(.a(output_10_61), .b(output_10_14), .y(output_9_61));
wire output_11_61, output_11_14, output_10_61;
mixer gate_output_10_61(.a(output_11_61), .b(output_11_14), .y(output_10_61));
wire output_12_61, output_12_14, output_11_61;
mixer gate_output_11_61(.a(output_12_61), .b(output_12_14), .y(output_11_61));
wire output_13_61, output_13_14, output_12_61;
mixer gate_output_12_61(.a(output_13_61), .b(output_13_14), .y(output_12_61));
wire output_14_61, output_14_14, output_13_61;
mixer gate_output_13_61(.a(output_14_61), .b(output_14_14), .y(output_13_61));
wire output_15_61, output_15_14, output_14_61;
mixer gate_output_14_61(.a(output_15_61), .b(output_15_14), .y(output_14_61));
wire output_16_61, output_16_14, output_15_61;
mixer gate_output_15_61(.a(output_16_61), .b(output_16_14), .y(output_15_61));
wire output_1_62, output_1_15, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_15), .y(output_0_62));
wire output_2_62, output_2_15, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_15), .y(output_1_62));
wire output_3_62, output_3_15, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_15), .y(output_2_62));
wire output_4_62, output_4_15, output_3_62;
mixer gate_output_3_62(.a(output_4_62), .b(output_4_15), .y(output_3_62));
wire output_5_62, output_5_15, output_4_62;
mixer gate_output_4_62(.a(output_5_62), .b(output_5_15), .y(output_4_62));
wire output_6_62, output_6_15, output_5_62;
mixer gate_output_5_62(.a(output_6_62), .b(output_6_15), .y(output_5_62));
wire output_7_62, output_7_15, output_6_62;
mixer gate_output_6_62(.a(output_7_62), .b(output_7_15), .y(output_6_62));
wire output_8_62, output_8_15, output_7_62;
mixer gate_output_7_62(.a(output_8_62), .b(output_8_15), .y(output_7_62));
wire output_9_62, output_9_15, output_8_62;
mixer gate_output_8_62(.a(output_9_62), .b(output_9_15), .y(output_8_62));
wire output_10_62, output_10_15, output_9_62;
mixer gate_output_9_62(.a(output_10_62), .b(output_10_15), .y(output_9_62));
wire output_11_62, output_11_15, output_10_62;
mixer gate_output_10_62(.a(output_11_62), .b(output_11_15), .y(output_10_62));
wire output_12_62, output_12_15, output_11_62;
mixer gate_output_11_62(.a(output_12_62), .b(output_12_15), .y(output_11_62));
wire output_13_62, output_13_15, output_12_62;
mixer gate_output_12_62(.a(output_13_62), .b(output_13_15), .y(output_12_62));
wire output_14_62, output_14_15, output_13_62;
mixer gate_output_13_62(.a(output_14_62), .b(output_14_15), .y(output_13_62));
wire output_15_62, output_15_15, output_14_62;
mixer gate_output_14_62(.a(output_15_62), .b(output_15_15), .y(output_14_62));
wire output_16_62, output_16_15, output_15_62;
mixer gate_output_15_62(.a(output_16_62), .b(output_16_15), .y(output_15_62));
wire output_1_63, output_1_0, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_0), .y(output_0_63));
wire output_2_63, output_2_0, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_0), .y(output_1_63));
wire output_3_63, output_3_0, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_0), .y(output_2_63));
wire output_4_63, output_4_0, output_3_63;
mixer gate_output_3_63(.a(output_4_63), .b(output_4_0), .y(output_3_63));
wire output_5_63, output_5_0, output_4_63;
mixer gate_output_4_63(.a(output_5_63), .b(output_5_0), .y(output_4_63));
wire output_6_63, output_6_0, output_5_63;
mixer gate_output_5_63(.a(output_6_63), .b(output_6_0), .y(output_5_63));
wire output_7_63, output_7_0, output_6_63;
mixer gate_output_6_63(.a(output_7_63), .b(output_7_0), .y(output_6_63));
wire output_8_63, output_8_0, output_7_63;
mixer gate_output_7_63(.a(output_8_63), .b(output_8_0), .y(output_7_63));
wire output_9_63, output_9_0, output_8_63;
mixer gate_output_8_63(.a(output_9_63), .b(output_9_0), .y(output_8_63));
wire output_10_63, output_10_0, output_9_63;
mixer gate_output_9_63(.a(output_10_63), .b(output_10_0), .y(output_9_63));
wire output_11_63, output_11_0, output_10_63;
mixer gate_output_10_63(.a(output_11_63), .b(output_11_0), .y(output_10_63));
wire output_12_63, output_12_0, output_11_63;
mixer gate_output_11_63(.a(output_12_63), .b(output_12_0), .y(output_11_63));
wire output_13_63, output_13_0, output_12_63;
mixer gate_output_12_63(.a(output_13_63), .b(output_13_0), .y(output_12_63));
wire output_14_63, output_14_0, output_13_63;
mixer gate_output_13_63(.a(output_14_63), .b(output_14_0), .y(output_13_63));
wire output_15_63, output_15_0, output_14_63;
mixer gate_output_14_63(.a(output_15_63), .b(output_15_0), .y(output_14_63));
wire output_16_63, output_16_0, output_15_63;
mixer gate_output_15_63(.a(output_16_63), .b(output_16_0), .y(output_15_63));
wire output_1_64, output_1_1, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_1), .y(output_0_64));
wire output_2_64, output_2_1, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_1), .y(output_1_64));
wire output_3_64, output_3_1, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_1), .y(output_2_64));
wire output_4_64, output_4_1, output_3_64;
mixer gate_output_3_64(.a(output_4_64), .b(output_4_1), .y(output_3_64));
wire output_5_64, output_5_1, output_4_64;
mixer gate_output_4_64(.a(output_5_64), .b(output_5_1), .y(output_4_64));
wire output_6_64, output_6_1, output_5_64;
mixer gate_output_5_64(.a(output_6_64), .b(output_6_1), .y(output_5_64));
wire output_7_64, output_7_1, output_6_64;
mixer gate_output_6_64(.a(output_7_64), .b(output_7_1), .y(output_6_64));
wire output_8_64, output_8_1, output_7_64;
mixer gate_output_7_64(.a(output_8_64), .b(output_8_1), .y(output_7_64));
wire output_9_64, output_9_1, output_8_64;
mixer gate_output_8_64(.a(output_9_64), .b(output_9_1), .y(output_8_64));
wire output_10_64, output_10_1, output_9_64;
mixer gate_output_9_64(.a(output_10_64), .b(output_10_1), .y(output_9_64));
wire output_11_64, output_11_1, output_10_64;
mixer gate_output_10_64(.a(output_11_64), .b(output_11_1), .y(output_10_64));
wire output_12_64, output_12_1, output_11_64;
mixer gate_output_11_64(.a(output_12_64), .b(output_12_1), .y(output_11_64));
wire output_13_64, output_13_1, output_12_64;
mixer gate_output_12_64(.a(output_13_64), .b(output_13_1), .y(output_12_64));
wire output_14_64, output_14_1, output_13_64;
mixer gate_output_13_64(.a(output_14_64), .b(output_14_1), .y(output_13_64));
wire output_15_64, output_15_1, output_14_64;
mixer gate_output_14_64(.a(output_15_64), .b(output_15_1), .y(output_14_64));
wire output_16_64, output_16_1, output_15_64;
mixer gate_output_15_64(.a(output_16_64), .b(output_16_1), .y(output_15_64));
wire output_1_65, output_1_2, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_2), .y(output_0_65));
wire output_2_65, output_2_2, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_2), .y(output_1_65));
wire output_3_65, output_3_2, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_2), .y(output_2_65));
wire output_4_65, output_4_2, output_3_65;
mixer gate_output_3_65(.a(output_4_65), .b(output_4_2), .y(output_3_65));
wire output_5_65, output_5_2, output_4_65;
mixer gate_output_4_65(.a(output_5_65), .b(output_5_2), .y(output_4_65));
wire output_6_65, output_6_2, output_5_65;
mixer gate_output_5_65(.a(output_6_65), .b(output_6_2), .y(output_5_65));
wire output_7_65, output_7_2, output_6_65;
mixer gate_output_6_65(.a(output_7_65), .b(output_7_2), .y(output_6_65));
wire output_8_65, output_8_2, output_7_65;
mixer gate_output_7_65(.a(output_8_65), .b(output_8_2), .y(output_7_65));
wire output_9_65, output_9_2, output_8_65;
mixer gate_output_8_65(.a(output_9_65), .b(output_9_2), .y(output_8_65));
wire output_10_65, output_10_2, output_9_65;
mixer gate_output_9_65(.a(output_10_65), .b(output_10_2), .y(output_9_65));
wire output_11_65, output_11_2, output_10_65;
mixer gate_output_10_65(.a(output_11_65), .b(output_11_2), .y(output_10_65));
wire output_12_65, output_12_2, output_11_65;
mixer gate_output_11_65(.a(output_12_65), .b(output_12_2), .y(output_11_65));
wire output_13_65, output_13_2, output_12_65;
mixer gate_output_12_65(.a(output_13_65), .b(output_13_2), .y(output_12_65));
wire output_14_65, output_14_2, output_13_65;
mixer gate_output_13_65(.a(output_14_65), .b(output_14_2), .y(output_13_65));
wire output_15_65, output_15_2, output_14_65;
mixer gate_output_14_65(.a(output_15_65), .b(output_15_2), .y(output_14_65));
wire output_16_65, output_16_2, output_15_65;
mixer gate_output_15_65(.a(output_16_65), .b(output_16_2), .y(output_15_65));
wire output_1_66, output_1_3, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_3), .y(output_0_66));
wire output_2_66, output_2_3, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_3), .y(output_1_66));
wire output_3_66, output_3_3, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_3), .y(output_2_66));
wire output_4_66, output_4_3, output_3_66;
mixer gate_output_3_66(.a(output_4_66), .b(output_4_3), .y(output_3_66));
wire output_5_66, output_5_3, output_4_66;
mixer gate_output_4_66(.a(output_5_66), .b(output_5_3), .y(output_4_66));
wire output_6_66, output_6_3, output_5_66;
mixer gate_output_5_66(.a(output_6_66), .b(output_6_3), .y(output_5_66));
wire output_7_66, output_7_3, output_6_66;
mixer gate_output_6_66(.a(output_7_66), .b(output_7_3), .y(output_6_66));
wire output_8_66, output_8_3, output_7_66;
mixer gate_output_7_66(.a(output_8_66), .b(output_8_3), .y(output_7_66));
wire output_9_66, output_9_3, output_8_66;
mixer gate_output_8_66(.a(output_9_66), .b(output_9_3), .y(output_8_66));
wire output_10_66, output_10_3, output_9_66;
mixer gate_output_9_66(.a(output_10_66), .b(output_10_3), .y(output_9_66));
wire output_11_66, output_11_3, output_10_66;
mixer gate_output_10_66(.a(output_11_66), .b(output_11_3), .y(output_10_66));
wire output_12_66, output_12_3, output_11_66;
mixer gate_output_11_66(.a(output_12_66), .b(output_12_3), .y(output_11_66));
wire output_13_66, output_13_3, output_12_66;
mixer gate_output_12_66(.a(output_13_66), .b(output_13_3), .y(output_12_66));
wire output_14_66, output_14_3, output_13_66;
mixer gate_output_13_66(.a(output_14_66), .b(output_14_3), .y(output_13_66));
wire output_15_66, output_15_3, output_14_66;
mixer gate_output_14_66(.a(output_15_66), .b(output_15_3), .y(output_14_66));
wire output_16_66, output_16_3, output_15_66;
mixer gate_output_15_66(.a(output_16_66), .b(output_16_3), .y(output_15_66));
wire output_1_67, output_1_4, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_4), .y(output_0_67));
wire output_2_67, output_2_4, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_4), .y(output_1_67));
wire output_3_67, output_3_4, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_4), .y(output_2_67));
wire output_4_67, output_4_4, output_3_67;
mixer gate_output_3_67(.a(output_4_67), .b(output_4_4), .y(output_3_67));
wire output_5_67, output_5_4, output_4_67;
mixer gate_output_4_67(.a(output_5_67), .b(output_5_4), .y(output_4_67));
wire output_6_67, output_6_4, output_5_67;
mixer gate_output_5_67(.a(output_6_67), .b(output_6_4), .y(output_5_67));
wire output_7_67, output_7_4, output_6_67;
mixer gate_output_6_67(.a(output_7_67), .b(output_7_4), .y(output_6_67));
wire output_8_67, output_8_4, output_7_67;
mixer gate_output_7_67(.a(output_8_67), .b(output_8_4), .y(output_7_67));
wire output_9_67, output_9_4, output_8_67;
mixer gate_output_8_67(.a(output_9_67), .b(output_9_4), .y(output_8_67));
wire output_10_67, output_10_4, output_9_67;
mixer gate_output_9_67(.a(output_10_67), .b(output_10_4), .y(output_9_67));
wire output_11_67, output_11_4, output_10_67;
mixer gate_output_10_67(.a(output_11_67), .b(output_11_4), .y(output_10_67));
wire output_12_67, output_12_4, output_11_67;
mixer gate_output_11_67(.a(output_12_67), .b(output_12_4), .y(output_11_67));
wire output_13_67, output_13_4, output_12_67;
mixer gate_output_12_67(.a(output_13_67), .b(output_13_4), .y(output_12_67));
wire output_14_67, output_14_4, output_13_67;
mixer gate_output_13_67(.a(output_14_67), .b(output_14_4), .y(output_13_67));
wire output_15_67, output_15_4, output_14_67;
mixer gate_output_14_67(.a(output_15_67), .b(output_15_4), .y(output_14_67));
wire output_16_67, output_16_4, output_15_67;
mixer gate_output_15_67(.a(output_16_67), .b(output_16_4), .y(output_15_67));
wire output_1_68, output_1_5, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_5), .y(output_0_68));
wire output_2_68, output_2_5, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_5), .y(output_1_68));
wire output_3_68, output_3_5, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_5), .y(output_2_68));
wire output_4_68, output_4_5, output_3_68;
mixer gate_output_3_68(.a(output_4_68), .b(output_4_5), .y(output_3_68));
wire output_5_68, output_5_5, output_4_68;
mixer gate_output_4_68(.a(output_5_68), .b(output_5_5), .y(output_4_68));
wire output_6_68, output_6_5, output_5_68;
mixer gate_output_5_68(.a(output_6_68), .b(output_6_5), .y(output_5_68));
wire output_7_68, output_7_5, output_6_68;
mixer gate_output_6_68(.a(output_7_68), .b(output_7_5), .y(output_6_68));
wire output_8_68, output_8_5, output_7_68;
mixer gate_output_7_68(.a(output_8_68), .b(output_8_5), .y(output_7_68));
wire output_9_68, output_9_5, output_8_68;
mixer gate_output_8_68(.a(output_9_68), .b(output_9_5), .y(output_8_68));
wire output_10_68, output_10_5, output_9_68;
mixer gate_output_9_68(.a(output_10_68), .b(output_10_5), .y(output_9_68));
wire output_11_68, output_11_5, output_10_68;
mixer gate_output_10_68(.a(output_11_68), .b(output_11_5), .y(output_10_68));
wire output_12_68, output_12_5, output_11_68;
mixer gate_output_11_68(.a(output_12_68), .b(output_12_5), .y(output_11_68));
wire output_13_68, output_13_5, output_12_68;
mixer gate_output_12_68(.a(output_13_68), .b(output_13_5), .y(output_12_68));
wire output_14_68, output_14_5, output_13_68;
mixer gate_output_13_68(.a(output_14_68), .b(output_14_5), .y(output_13_68));
wire output_15_68, output_15_5, output_14_68;
mixer gate_output_14_68(.a(output_15_68), .b(output_15_5), .y(output_14_68));
wire output_16_68, output_16_5, output_15_68;
mixer gate_output_15_68(.a(output_16_68), .b(output_16_5), .y(output_15_68));
wire output_1_69, output_1_6, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_6), .y(output_0_69));
wire output_2_69, output_2_6, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_6), .y(output_1_69));
wire output_3_69, output_3_6, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_6), .y(output_2_69));
wire output_4_69, output_4_6, output_3_69;
mixer gate_output_3_69(.a(output_4_69), .b(output_4_6), .y(output_3_69));
wire output_5_69, output_5_6, output_4_69;
mixer gate_output_4_69(.a(output_5_69), .b(output_5_6), .y(output_4_69));
wire output_6_69, output_6_6, output_5_69;
mixer gate_output_5_69(.a(output_6_69), .b(output_6_6), .y(output_5_69));
wire output_7_69, output_7_6, output_6_69;
mixer gate_output_6_69(.a(output_7_69), .b(output_7_6), .y(output_6_69));
wire output_8_69, output_8_6, output_7_69;
mixer gate_output_7_69(.a(output_8_69), .b(output_8_6), .y(output_7_69));
wire output_9_69, output_9_6, output_8_69;
mixer gate_output_8_69(.a(output_9_69), .b(output_9_6), .y(output_8_69));
wire output_10_69, output_10_6, output_9_69;
mixer gate_output_9_69(.a(output_10_69), .b(output_10_6), .y(output_9_69));
wire output_11_69, output_11_6, output_10_69;
mixer gate_output_10_69(.a(output_11_69), .b(output_11_6), .y(output_10_69));
wire output_12_69, output_12_6, output_11_69;
mixer gate_output_11_69(.a(output_12_69), .b(output_12_6), .y(output_11_69));
wire output_13_69, output_13_6, output_12_69;
mixer gate_output_12_69(.a(output_13_69), .b(output_13_6), .y(output_12_69));
wire output_14_69, output_14_6, output_13_69;
mixer gate_output_13_69(.a(output_14_69), .b(output_14_6), .y(output_13_69));
wire output_15_69, output_15_6, output_14_69;
mixer gate_output_14_69(.a(output_15_69), .b(output_15_6), .y(output_14_69));
wire output_16_69, output_16_6, output_15_69;
mixer gate_output_15_69(.a(output_16_69), .b(output_16_6), .y(output_15_69));
wire output_1_70, output_1_7, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_7), .y(output_0_70));
wire output_2_70, output_2_7, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_7), .y(output_1_70));
wire output_3_70, output_3_7, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_7), .y(output_2_70));
wire output_4_70, output_4_7, output_3_70;
mixer gate_output_3_70(.a(output_4_70), .b(output_4_7), .y(output_3_70));
wire output_5_70, output_5_7, output_4_70;
mixer gate_output_4_70(.a(output_5_70), .b(output_5_7), .y(output_4_70));
wire output_6_70, output_6_7, output_5_70;
mixer gate_output_5_70(.a(output_6_70), .b(output_6_7), .y(output_5_70));
wire output_7_70, output_7_7, output_6_70;
mixer gate_output_6_70(.a(output_7_70), .b(output_7_7), .y(output_6_70));
wire output_8_70, output_8_7, output_7_70;
mixer gate_output_7_70(.a(output_8_70), .b(output_8_7), .y(output_7_70));
wire output_9_70, output_9_7, output_8_70;
mixer gate_output_8_70(.a(output_9_70), .b(output_9_7), .y(output_8_70));
wire output_10_70, output_10_7, output_9_70;
mixer gate_output_9_70(.a(output_10_70), .b(output_10_7), .y(output_9_70));
wire output_11_70, output_11_7, output_10_70;
mixer gate_output_10_70(.a(output_11_70), .b(output_11_7), .y(output_10_70));
wire output_12_70, output_12_7, output_11_70;
mixer gate_output_11_70(.a(output_12_70), .b(output_12_7), .y(output_11_70));
wire output_13_70, output_13_7, output_12_70;
mixer gate_output_12_70(.a(output_13_70), .b(output_13_7), .y(output_12_70));
wire output_14_70, output_14_7, output_13_70;
mixer gate_output_13_70(.a(output_14_70), .b(output_14_7), .y(output_13_70));
wire output_15_70, output_15_7, output_14_70;
mixer gate_output_14_70(.a(output_15_70), .b(output_15_7), .y(output_14_70));
wire output_16_70, output_16_7, output_15_70;
mixer gate_output_15_70(.a(output_16_70), .b(output_16_7), .y(output_15_70));
wire output_1_71, output_1_8, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_8), .y(output_0_71));
wire output_2_71, output_2_8, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_8), .y(output_1_71));
wire output_3_71, output_3_8, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_8), .y(output_2_71));
wire output_4_71, output_4_8, output_3_71;
mixer gate_output_3_71(.a(output_4_71), .b(output_4_8), .y(output_3_71));
wire output_5_71, output_5_8, output_4_71;
mixer gate_output_4_71(.a(output_5_71), .b(output_5_8), .y(output_4_71));
wire output_6_71, output_6_8, output_5_71;
mixer gate_output_5_71(.a(output_6_71), .b(output_6_8), .y(output_5_71));
wire output_7_71, output_7_8, output_6_71;
mixer gate_output_6_71(.a(output_7_71), .b(output_7_8), .y(output_6_71));
wire output_8_71, output_8_8, output_7_71;
mixer gate_output_7_71(.a(output_8_71), .b(output_8_8), .y(output_7_71));
wire output_9_71, output_9_8, output_8_71;
mixer gate_output_8_71(.a(output_9_71), .b(output_9_8), .y(output_8_71));
wire output_10_71, output_10_8, output_9_71;
mixer gate_output_9_71(.a(output_10_71), .b(output_10_8), .y(output_9_71));
wire output_11_71, output_11_8, output_10_71;
mixer gate_output_10_71(.a(output_11_71), .b(output_11_8), .y(output_10_71));
wire output_12_71, output_12_8, output_11_71;
mixer gate_output_11_71(.a(output_12_71), .b(output_12_8), .y(output_11_71));
wire output_13_71, output_13_8, output_12_71;
mixer gate_output_12_71(.a(output_13_71), .b(output_13_8), .y(output_12_71));
wire output_14_71, output_14_8, output_13_71;
mixer gate_output_13_71(.a(output_14_71), .b(output_14_8), .y(output_13_71));
wire output_15_71, output_15_8, output_14_71;
mixer gate_output_14_71(.a(output_15_71), .b(output_15_8), .y(output_14_71));
wire output_16_71, output_16_8, output_15_71;
mixer gate_output_15_71(.a(output_16_71), .b(output_16_8), .y(output_15_71));
wire output_1_72, output_1_9, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_9), .y(output_0_72));
wire output_2_72, output_2_9, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_9), .y(output_1_72));
wire output_3_72, output_3_9, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_9), .y(output_2_72));
wire output_4_72, output_4_9, output_3_72;
mixer gate_output_3_72(.a(output_4_72), .b(output_4_9), .y(output_3_72));
wire output_5_72, output_5_9, output_4_72;
mixer gate_output_4_72(.a(output_5_72), .b(output_5_9), .y(output_4_72));
wire output_6_72, output_6_9, output_5_72;
mixer gate_output_5_72(.a(output_6_72), .b(output_6_9), .y(output_5_72));
wire output_7_72, output_7_9, output_6_72;
mixer gate_output_6_72(.a(output_7_72), .b(output_7_9), .y(output_6_72));
wire output_8_72, output_8_9, output_7_72;
mixer gate_output_7_72(.a(output_8_72), .b(output_8_9), .y(output_7_72));
wire output_9_72, output_9_9, output_8_72;
mixer gate_output_8_72(.a(output_9_72), .b(output_9_9), .y(output_8_72));
wire output_10_72, output_10_9, output_9_72;
mixer gate_output_9_72(.a(output_10_72), .b(output_10_9), .y(output_9_72));
wire output_11_72, output_11_9, output_10_72;
mixer gate_output_10_72(.a(output_11_72), .b(output_11_9), .y(output_10_72));
wire output_12_72, output_12_9, output_11_72;
mixer gate_output_11_72(.a(output_12_72), .b(output_12_9), .y(output_11_72));
wire output_13_72, output_13_9, output_12_72;
mixer gate_output_12_72(.a(output_13_72), .b(output_13_9), .y(output_12_72));
wire output_14_72, output_14_9, output_13_72;
mixer gate_output_13_72(.a(output_14_72), .b(output_14_9), .y(output_13_72));
wire output_15_72, output_15_9, output_14_72;
mixer gate_output_14_72(.a(output_15_72), .b(output_15_9), .y(output_14_72));
wire output_16_72, output_16_9, output_15_72;
mixer gate_output_15_72(.a(output_16_72), .b(output_16_9), .y(output_15_72));
wire output_1_73, output_1_10, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_10), .y(output_0_73));
wire output_2_73, output_2_10, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_10), .y(output_1_73));
wire output_3_73, output_3_10, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_10), .y(output_2_73));
wire output_4_73, output_4_10, output_3_73;
mixer gate_output_3_73(.a(output_4_73), .b(output_4_10), .y(output_3_73));
wire output_5_73, output_5_10, output_4_73;
mixer gate_output_4_73(.a(output_5_73), .b(output_5_10), .y(output_4_73));
wire output_6_73, output_6_10, output_5_73;
mixer gate_output_5_73(.a(output_6_73), .b(output_6_10), .y(output_5_73));
wire output_7_73, output_7_10, output_6_73;
mixer gate_output_6_73(.a(output_7_73), .b(output_7_10), .y(output_6_73));
wire output_8_73, output_8_10, output_7_73;
mixer gate_output_7_73(.a(output_8_73), .b(output_8_10), .y(output_7_73));
wire output_9_73, output_9_10, output_8_73;
mixer gate_output_8_73(.a(output_9_73), .b(output_9_10), .y(output_8_73));
wire output_10_73, output_10_10, output_9_73;
mixer gate_output_9_73(.a(output_10_73), .b(output_10_10), .y(output_9_73));
wire output_11_73, output_11_10, output_10_73;
mixer gate_output_10_73(.a(output_11_73), .b(output_11_10), .y(output_10_73));
wire output_12_73, output_12_10, output_11_73;
mixer gate_output_11_73(.a(output_12_73), .b(output_12_10), .y(output_11_73));
wire output_13_73, output_13_10, output_12_73;
mixer gate_output_12_73(.a(output_13_73), .b(output_13_10), .y(output_12_73));
wire output_14_73, output_14_10, output_13_73;
mixer gate_output_13_73(.a(output_14_73), .b(output_14_10), .y(output_13_73));
wire output_15_73, output_15_10, output_14_73;
mixer gate_output_14_73(.a(output_15_73), .b(output_15_10), .y(output_14_73));
wire output_16_73, output_16_10, output_15_73;
mixer gate_output_15_73(.a(output_16_73), .b(output_16_10), .y(output_15_73));
wire output_1_74, output_1_11, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_11), .y(output_0_74));
wire output_2_74, output_2_11, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_11), .y(output_1_74));
wire output_3_74, output_3_11, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_11), .y(output_2_74));
wire output_4_74, output_4_11, output_3_74;
mixer gate_output_3_74(.a(output_4_74), .b(output_4_11), .y(output_3_74));
wire output_5_74, output_5_11, output_4_74;
mixer gate_output_4_74(.a(output_5_74), .b(output_5_11), .y(output_4_74));
wire output_6_74, output_6_11, output_5_74;
mixer gate_output_5_74(.a(output_6_74), .b(output_6_11), .y(output_5_74));
wire output_7_74, output_7_11, output_6_74;
mixer gate_output_6_74(.a(output_7_74), .b(output_7_11), .y(output_6_74));
wire output_8_74, output_8_11, output_7_74;
mixer gate_output_7_74(.a(output_8_74), .b(output_8_11), .y(output_7_74));
wire output_9_74, output_9_11, output_8_74;
mixer gate_output_8_74(.a(output_9_74), .b(output_9_11), .y(output_8_74));
wire output_10_74, output_10_11, output_9_74;
mixer gate_output_9_74(.a(output_10_74), .b(output_10_11), .y(output_9_74));
wire output_11_74, output_11_11, output_10_74;
mixer gate_output_10_74(.a(output_11_74), .b(output_11_11), .y(output_10_74));
wire output_12_74, output_12_11, output_11_74;
mixer gate_output_11_74(.a(output_12_74), .b(output_12_11), .y(output_11_74));
wire output_13_74, output_13_11, output_12_74;
mixer gate_output_12_74(.a(output_13_74), .b(output_13_11), .y(output_12_74));
wire output_14_74, output_14_11, output_13_74;
mixer gate_output_13_74(.a(output_14_74), .b(output_14_11), .y(output_13_74));
wire output_15_74, output_15_11, output_14_74;
mixer gate_output_14_74(.a(output_15_74), .b(output_15_11), .y(output_14_74));
wire output_16_74, output_16_11, output_15_74;
mixer gate_output_15_74(.a(output_16_74), .b(output_16_11), .y(output_15_74));
wire output_1_75, output_1_12, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_12), .y(output_0_75));
wire output_2_75, output_2_12, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_12), .y(output_1_75));
wire output_3_75, output_3_12, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_12), .y(output_2_75));
wire output_4_75, output_4_12, output_3_75;
mixer gate_output_3_75(.a(output_4_75), .b(output_4_12), .y(output_3_75));
wire output_5_75, output_5_12, output_4_75;
mixer gate_output_4_75(.a(output_5_75), .b(output_5_12), .y(output_4_75));
wire output_6_75, output_6_12, output_5_75;
mixer gate_output_5_75(.a(output_6_75), .b(output_6_12), .y(output_5_75));
wire output_7_75, output_7_12, output_6_75;
mixer gate_output_6_75(.a(output_7_75), .b(output_7_12), .y(output_6_75));
wire output_8_75, output_8_12, output_7_75;
mixer gate_output_7_75(.a(output_8_75), .b(output_8_12), .y(output_7_75));
wire output_9_75, output_9_12, output_8_75;
mixer gate_output_8_75(.a(output_9_75), .b(output_9_12), .y(output_8_75));
wire output_10_75, output_10_12, output_9_75;
mixer gate_output_9_75(.a(output_10_75), .b(output_10_12), .y(output_9_75));
wire output_11_75, output_11_12, output_10_75;
mixer gate_output_10_75(.a(output_11_75), .b(output_11_12), .y(output_10_75));
wire output_12_75, output_12_12, output_11_75;
mixer gate_output_11_75(.a(output_12_75), .b(output_12_12), .y(output_11_75));
wire output_13_75, output_13_12, output_12_75;
mixer gate_output_12_75(.a(output_13_75), .b(output_13_12), .y(output_12_75));
wire output_14_75, output_14_12, output_13_75;
mixer gate_output_13_75(.a(output_14_75), .b(output_14_12), .y(output_13_75));
wire output_15_75, output_15_12, output_14_75;
mixer gate_output_14_75(.a(output_15_75), .b(output_15_12), .y(output_14_75));
wire output_16_75, output_16_12, output_15_75;
mixer gate_output_15_75(.a(output_16_75), .b(output_16_12), .y(output_15_75));
wire output_1_76, output_1_13, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_13), .y(output_0_76));
wire output_2_76, output_2_13, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_13), .y(output_1_76));
wire output_3_76, output_3_13, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_13), .y(output_2_76));
wire output_4_76, output_4_13, output_3_76;
mixer gate_output_3_76(.a(output_4_76), .b(output_4_13), .y(output_3_76));
wire output_5_76, output_5_13, output_4_76;
mixer gate_output_4_76(.a(output_5_76), .b(output_5_13), .y(output_4_76));
wire output_6_76, output_6_13, output_5_76;
mixer gate_output_5_76(.a(output_6_76), .b(output_6_13), .y(output_5_76));
wire output_7_76, output_7_13, output_6_76;
mixer gate_output_6_76(.a(output_7_76), .b(output_7_13), .y(output_6_76));
wire output_8_76, output_8_13, output_7_76;
mixer gate_output_7_76(.a(output_8_76), .b(output_8_13), .y(output_7_76));
wire output_9_76, output_9_13, output_8_76;
mixer gate_output_8_76(.a(output_9_76), .b(output_9_13), .y(output_8_76));
wire output_10_76, output_10_13, output_9_76;
mixer gate_output_9_76(.a(output_10_76), .b(output_10_13), .y(output_9_76));
wire output_11_76, output_11_13, output_10_76;
mixer gate_output_10_76(.a(output_11_76), .b(output_11_13), .y(output_10_76));
wire output_12_76, output_12_13, output_11_76;
mixer gate_output_11_76(.a(output_12_76), .b(output_12_13), .y(output_11_76));
wire output_13_76, output_13_13, output_12_76;
mixer gate_output_12_76(.a(output_13_76), .b(output_13_13), .y(output_12_76));
wire output_14_76, output_14_13, output_13_76;
mixer gate_output_13_76(.a(output_14_76), .b(output_14_13), .y(output_13_76));
wire output_15_76, output_15_13, output_14_76;
mixer gate_output_14_76(.a(output_15_76), .b(output_15_13), .y(output_14_76));
wire output_16_76, output_16_13, output_15_76;
mixer gate_output_15_76(.a(output_16_76), .b(output_16_13), .y(output_15_76));
wire output_1_77, output_1_14, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_14), .y(output_0_77));
wire output_2_77, output_2_14, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_14), .y(output_1_77));
wire output_3_77, output_3_14, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_14), .y(output_2_77));
wire output_4_77, output_4_14, output_3_77;
mixer gate_output_3_77(.a(output_4_77), .b(output_4_14), .y(output_3_77));
wire output_5_77, output_5_14, output_4_77;
mixer gate_output_4_77(.a(output_5_77), .b(output_5_14), .y(output_4_77));
wire output_6_77, output_6_14, output_5_77;
mixer gate_output_5_77(.a(output_6_77), .b(output_6_14), .y(output_5_77));
wire output_7_77, output_7_14, output_6_77;
mixer gate_output_6_77(.a(output_7_77), .b(output_7_14), .y(output_6_77));
wire output_8_77, output_8_14, output_7_77;
mixer gate_output_7_77(.a(output_8_77), .b(output_8_14), .y(output_7_77));
wire output_9_77, output_9_14, output_8_77;
mixer gate_output_8_77(.a(output_9_77), .b(output_9_14), .y(output_8_77));
wire output_10_77, output_10_14, output_9_77;
mixer gate_output_9_77(.a(output_10_77), .b(output_10_14), .y(output_9_77));
wire output_11_77, output_11_14, output_10_77;
mixer gate_output_10_77(.a(output_11_77), .b(output_11_14), .y(output_10_77));
wire output_12_77, output_12_14, output_11_77;
mixer gate_output_11_77(.a(output_12_77), .b(output_12_14), .y(output_11_77));
wire output_13_77, output_13_14, output_12_77;
mixer gate_output_12_77(.a(output_13_77), .b(output_13_14), .y(output_12_77));
wire output_14_77, output_14_14, output_13_77;
mixer gate_output_13_77(.a(output_14_77), .b(output_14_14), .y(output_13_77));
wire output_15_77, output_15_14, output_14_77;
mixer gate_output_14_77(.a(output_15_77), .b(output_15_14), .y(output_14_77));
wire output_16_77, output_16_14, output_15_77;
mixer gate_output_15_77(.a(output_16_77), .b(output_16_14), .y(output_15_77));
wire output_1_78, output_1_15, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_15), .y(output_0_78));
wire output_2_78, output_2_15, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_15), .y(output_1_78));
wire output_3_78, output_3_15, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_15), .y(output_2_78));
wire output_4_78, output_4_15, output_3_78;
mixer gate_output_3_78(.a(output_4_78), .b(output_4_15), .y(output_3_78));
wire output_5_78, output_5_15, output_4_78;
mixer gate_output_4_78(.a(output_5_78), .b(output_5_15), .y(output_4_78));
wire output_6_78, output_6_15, output_5_78;
mixer gate_output_5_78(.a(output_6_78), .b(output_6_15), .y(output_5_78));
wire output_7_78, output_7_15, output_6_78;
mixer gate_output_6_78(.a(output_7_78), .b(output_7_15), .y(output_6_78));
wire output_8_78, output_8_15, output_7_78;
mixer gate_output_7_78(.a(output_8_78), .b(output_8_15), .y(output_7_78));
wire output_9_78, output_9_15, output_8_78;
mixer gate_output_8_78(.a(output_9_78), .b(output_9_15), .y(output_8_78));
wire output_10_78, output_10_15, output_9_78;
mixer gate_output_9_78(.a(output_10_78), .b(output_10_15), .y(output_9_78));
wire output_11_78, output_11_15, output_10_78;
mixer gate_output_10_78(.a(output_11_78), .b(output_11_15), .y(output_10_78));
wire output_12_78, output_12_15, output_11_78;
mixer gate_output_11_78(.a(output_12_78), .b(output_12_15), .y(output_11_78));
wire output_13_78, output_13_15, output_12_78;
mixer gate_output_12_78(.a(output_13_78), .b(output_13_15), .y(output_12_78));
wire output_14_78, output_14_15, output_13_78;
mixer gate_output_13_78(.a(output_14_78), .b(output_14_15), .y(output_13_78));
wire output_15_78, output_15_15, output_14_78;
mixer gate_output_14_78(.a(output_15_78), .b(output_15_15), .y(output_14_78));
wire output_16_78, output_16_15, output_15_78;
mixer gate_output_15_78(.a(output_16_78), .b(output_16_15), .y(output_15_78));
wire output_1_79, output_1_0, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_0), .y(output_0_79));
wire output_2_79, output_2_0, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_0), .y(output_1_79));
wire output_3_79, output_3_0, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_0), .y(output_2_79));
wire output_4_79, output_4_0, output_3_79;
mixer gate_output_3_79(.a(output_4_79), .b(output_4_0), .y(output_3_79));
wire output_5_79, output_5_0, output_4_79;
mixer gate_output_4_79(.a(output_5_79), .b(output_5_0), .y(output_4_79));
wire output_6_79, output_6_0, output_5_79;
mixer gate_output_5_79(.a(output_6_79), .b(output_6_0), .y(output_5_79));
wire output_7_79, output_7_0, output_6_79;
mixer gate_output_6_79(.a(output_7_79), .b(output_7_0), .y(output_6_79));
wire output_8_79, output_8_0, output_7_79;
mixer gate_output_7_79(.a(output_8_79), .b(output_8_0), .y(output_7_79));
wire output_9_79, output_9_0, output_8_79;
mixer gate_output_8_79(.a(output_9_79), .b(output_9_0), .y(output_8_79));
wire output_10_79, output_10_0, output_9_79;
mixer gate_output_9_79(.a(output_10_79), .b(output_10_0), .y(output_9_79));
wire output_11_79, output_11_0, output_10_79;
mixer gate_output_10_79(.a(output_11_79), .b(output_11_0), .y(output_10_79));
wire output_12_79, output_12_0, output_11_79;
mixer gate_output_11_79(.a(output_12_79), .b(output_12_0), .y(output_11_79));
wire output_13_79, output_13_0, output_12_79;
mixer gate_output_12_79(.a(output_13_79), .b(output_13_0), .y(output_12_79));
wire output_14_79, output_14_0, output_13_79;
mixer gate_output_13_79(.a(output_14_79), .b(output_14_0), .y(output_13_79));
wire output_15_79, output_15_0, output_14_79;
mixer gate_output_14_79(.a(output_15_79), .b(output_15_0), .y(output_14_79));
wire output_16_79, output_16_0, output_15_79;
mixer gate_output_15_79(.a(output_16_79), .b(output_16_0), .y(output_15_79));
wire output_1_80, output_1_1, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_1), .y(output_0_80));
wire output_2_80, output_2_1, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_1), .y(output_1_80));
wire output_3_80, output_3_1, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_1), .y(output_2_80));
wire output_4_80, output_4_1, output_3_80;
mixer gate_output_3_80(.a(output_4_80), .b(output_4_1), .y(output_3_80));
wire output_5_80, output_5_1, output_4_80;
mixer gate_output_4_80(.a(output_5_80), .b(output_5_1), .y(output_4_80));
wire output_6_80, output_6_1, output_5_80;
mixer gate_output_5_80(.a(output_6_80), .b(output_6_1), .y(output_5_80));
wire output_7_80, output_7_1, output_6_80;
mixer gate_output_6_80(.a(output_7_80), .b(output_7_1), .y(output_6_80));
wire output_8_80, output_8_1, output_7_80;
mixer gate_output_7_80(.a(output_8_80), .b(output_8_1), .y(output_7_80));
wire output_9_80, output_9_1, output_8_80;
mixer gate_output_8_80(.a(output_9_80), .b(output_9_1), .y(output_8_80));
wire output_10_80, output_10_1, output_9_80;
mixer gate_output_9_80(.a(output_10_80), .b(output_10_1), .y(output_9_80));
wire output_11_80, output_11_1, output_10_80;
mixer gate_output_10_80(.a(output_11_80), .b(output_11_1), .y(output_10_80));
wire output_12_80, output_12_1, output_11_80;
mixer gate_output_11_80(.a(output_12_80), .b(output_12_1), .y(output_11_80));
wire output_13_80, output_13_1, output_12_80;
mixer gate_output_12_80(.a(output_13_80), .b(output_13_1), .y(output_12_80));
wire output_14_80, output_14_1, output_13_80;
mixer gate_output_13_80(.a(output_14_80), .b(output_14_1), .y(output_13_80));
wire output_15_80, output_15_1, output_14_80;
mixer gate_output_14_80(.a(output_15_80), .b(output_15_1), .y(output_14_80));
wire output_16_80, output_16_1, output_15_80;
mixer gate_output_15_80(.a(output_16_80), .b(output_16_1), .y(output_15_80));
wire output_1_81, output_1_2, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_2), .y(output_0_81));
wire output_2_81, output_2_2, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_2), .y(output_1_81));
wire output_3_81, output_3_2, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_2), .y(output_2_81));
wire output_4_81, output_4_2, output_3_81;
mixer gate_output_3_81(.a(output_4_81), .b(output_4_2), .y(output_3_81));
wire output_5_81, output_5_2, output_4_81;
mixer gate_output_4_81(.a(output_5_81), .b(output_5_2), .y(output_4_81));
wire output_6_81, output_6_2, output_5_81;
mixer gate_output_5_81(.a(output_6_81), .b(output_6_2), .y(output_5_81));
wire output_7_81, output_7_2, output_6_81;
mixer gate_output_6_81(.a(output_7_81), .b(output_7_2), .y(output_6_81));
wire output_8_81, output_8_2, output_7_81;
mixer gate_output_7_81(.a(output_8_81), .b(output_8_2), .y(output_7_81));
wire output_9_81, output_9_2, output_8_81;
mixer gate_output_8_81(.a(output_9_81), .b(output_9_2), .y(output_8_81));
wire output_10_81, output_10_2, output_9_81;
mixer gate_output_9_81(.a(output_10_81), .b(output_10_2), .y(output_9_81));
wire output_11_81, output_11_2, output_10_81;
mixer gate_output_10_81(.a(output_11_81), .b(output_11_2), .y(output_10_81));
wire output_12_81, output_12_2, output_11_81;
mixer gate_output_11_81(.a(output_12_81), .b(output_12_2), .y(output_11_81));
wire output_13_81, output_13_2, output_12_81;
mixer gate_output_12_81(.a(output_13_81), .b(output_13_2), .y(output_12_81));
wire output_14_81, output_14_2, output_13_81;
mixer gate_output_13_81(.a(output_14_81), .b(output_14_2), .y(output_13_81));
wire output_15_81, output_15_2, output_14_81;
mixer gate_output_14_81(.a(output_15_81), .b(output_15_2), .y(output_14_81));
wire output_16_81, output_16_2, output_15_81;
mixer gate_output_15_81(.a(output_16_81), .b(output_16_2), .y(output_15_81));
wire output_1_82, output_1_3, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_3), .y(output_0_82));
wire output_2_82, output_2_3, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_3), .y(output_1_82));
wire output_3_82, output_3_3, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_3), .y(output_2_82));
wire output_4_82, output_4_3, output_3_82;
mixer gate_output_3_82(.a(output_4_82), .b(output_4_3), .y(output_3_82));
wire output_5_82, output_5_3, output_4_82;
mixer gate_output_4_82(.a(output_5_82), .b(output_5_3), .y(output_4_82));
wire output_6_82, output_6_3, output_5_82;
mixer gate_output_5_82(.a(output_6_82), .b(output_6_3), .y(output_5_82));
wire output_7_82, output_7_3, output_6_82;
mixer gate_output_6_82(.a(output_7_82), .b(output_7_3), .y(output_6_82));
wire output_8_82, output_8_3, output_7_82;
mixer gate_output_7_82(.a(output_8_82), .b(output_8_3), .y(output_7_82));
wire output_9_82, output_9_3, output_8_82;
mixer gate_output_8_82(.a(output_9_82), .b(output_9_3), .y(output_8_82));
wire output_10_82, output_10_3, output_9_82;
mixer gate_output_9_82(.a(output_10_82), .b(output_10_3), .y(output_9_82));
wire output_11_82, output_11_3, output_10_82;
mixer gate_output_10_82(.a(output_11_82), .b(output_11_3), .y(output_10_82));
wire output_12_82, output_12_3, output_11_82;
mixer gate_output_11_82(.a(output_12_82), .b(output_12_3), .y(output_11_82));
wire output_13_82, output_13_3, output_12_82;
mixer gate_output_12_82(.a(output_13_82), .b(output_13_3), .y(output_12_82));
wire output_14_82, output_14_3, output_13_82;
mixer gate_output_13_82(.a(output_14_82), .b(output_14_3), .y(output_13_82));
wire output_15_82, output_15_3, output_14_82;
mixer gate_output_14_82(.a(output_15_82), .b(output_15_3), .y(output_14_82));
wire output_16_82, output_16_3, output_15_82;
mixer gate_output_15_82(.a(output_16_82), .b(output_16_3), .y(output_15_82));
wire output_1_83, output_1_4, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_4), .y(output_0_83));
wire output_2_83, output_2_4, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_4), .y(output_1_83));
wire output_3_83, output_3_4, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_4), .y(output_2_83));
wire output_4_83, output_4_4, output_3_83;
mixer gate_output_3_83(.a(output_4_83), .b(output_4_4), .y(output_3_83));
wire output_5_83, output_5_4, output_4_83;
mixer gate_output_4_83(.a(output_5_83), .b(output_5_4), .y(output_4_83));
wire output_6_83, output_6_4, output_5_83;
mixer gate_output_5_83(.a(output_6_83), .b(output_6_4), .y(output_5_83));
wire output_7_83, output_7_4, output_6_83;
mixer gate_output_6_83(.a(output_7_83), .b(output_7_4), .y(output_6_83));
wire output_8_83, output_8_4, output_7_83;
mixer gate_output_7_83(.a(output_8_83), .b(output_8_4), .y(output_7_83));
wire output_9_83, output_9_4, output_8_83;
mixer gate_output_8_83(.a(output_9_83), .b(output_9_4), .y(output_8_83));
wire output_10_83, output_10_4, output_9_83;
mixer gate_output_9_83(.a(output_10_83), .b(output_10_4), .y(output_9_83));
wire output_11_83, output_11_4, output_10_83;
mixer gate_output_10_83(.a(output_11_83), .b(output_11_4), .y(output_10_83));
wire output_12_83, output_12_4, output_11_83;
mixer gate_output_11_83(.a(output_12_83), .b(output_12_4), .y(output_11_83));
wire output_13_83, output_13_4, output_12_83;
mixer gate_output_12_83(.a(output_13_83), .b(output_13_4), .y(output_12_83));
wire output_14_83, output_14_4, output_13_83;
mixer gate_output_13_83(.a(output_14_83), .b(output_14_4), .y(output_13_83));
wire output_15_83, output_15_4, output_14_83;
mixer gate_output_14_83(.a(output_15_83), .b(output_15_4), .y(output_14_83));
wire output_16_83, output_16_4, output_15_83;
mixer gate_output_15_83(.a(output_16_83), .b(output_16_4), .y(output_15_83));
wire output_1_84, output_1_5, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_5), .y(output_0_84));
wire output_2_84, output_2_5, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_5), .y(output_1_84));
wire output_3_84, output_3_5, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_5), .y(output_2_84));
wire output_4_84, output_4_5, output_3_84;
mixer gate_output_3_84(.a(output_4_84), .b(output_4_5), .y(output_3_84));
wire output_5_84, output_5_5, output_4_84;
mixer gate_output_4_84(.a(output_5_84), .b(output_5_5), .y(output_4_84));
wire output_6_84, output_6_5, output_5_84;
mixer gate_output_5_84(.a(output_6_84), .b(output_6_5), .y(output_5_84));
wire output_7_84, output_7_5, output_6_84;
mixer gate_output_6_84(.a(output_7_84), .b(output_7_5), .y(output_6_84));
wire output_8_84, output_8_5, output_7_84;
mixer gate_output_7_84(.a(output_8_84), .b(output_8_5), .y(output_7_84));
wire output_9_84, output_9_5, output_8_84;
mixer gate_output_8_84(.a(output_9_84), .b(output_9_5), .y(output_8_84));
wire output_10_84, output_10_5, output_9_84;
mixer gate_output_9_84(.a(output_10_84), .b(output_10_5), .y(output_9_84));
wire output_11_84, output_11_5, output_10_84;
mixer gate_output_10_84(.a(output_11_84), .b(output_11_5), .y(output_10_84));
wire output_12_84, output_12_5, output_11_84;
mixer gate_output_11_84(.a(output_12_84), .b(output_12_5), .y(output_11_84));
wire output_13_84, output_13_5, output_12_84;
mixer gate_output_12_84(.a(output_13_84), .b(output_13_5), .y(output_12_84));
wire output_14_84, output_14_5, output_13_84;
mixer gate_output_13_84(.a(output_14_84), .b(output_14_5), .y(output_13_84));
wire output_15_84, output_15_5, output_14_84;
mixer gate_output_14_84(.a(output_15_84), .b(output_15_5), .y(output_14_84));
wire output_16_84, output_16_5, output_15_84;
mixer gate_output_15_84(.a(output_16_84), .b(output_16_5), .y(output_15_84));
wire output_1_85, output_1_6, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_6), .y(output_0_85));
wire output_2_85, output_2_6, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_6), .y(output_1_85));
wire output_3_85, output_3_6, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_6), .y(output_2_85));
wire output_4_85, output_4_6, output_3_85;
mixer gate_output_3_85(.a(output_4_85), .b(output_4_6), .y(output_3_85));
wire output_5_85, output_5_6, output_4_85;
mixer gate_output_4_85(.a(output_5_85), .b(output_5_6), .y(output_4_85));
wire output_6_85, output_6_6, output_5_85;
mixer gate_output_5_85(.a(output_6_85), .b(output_6_6), .y(output_5_85));
wire output_7_85, output_7_6, output_6_85;
mixer gate_output_6_85(.a(output_7_85), .b(output_7_6), .y(output_6_85));
wire output_8_85, output_8_6, output_7_85;
mixer gate_output_7_85(.a(output_8_85), .b(output_8_6), .y(output_7_85));
wire output_9_85, output_9_6, output_8_85;
mixer gate_output_8_85(.a(output_9_85), .b(output_9_6), .y(output_8_85));
wire output_10_85, output_10_6, output_9_85;
mixer gate_output_9_85(.a(output_10_85), .b(output_10_6), .y(output_9_85));
wire output_11_85, output_11_6, output_10_85;
mixer gate_output_10_85(.a(output_11_85), .b(output_11_6), .y(output_10_85));
wire output_12_85, output_12_6, output_11_85;
mixer gate_output_11_85(.a(output_12_85), .b(output_12_6), .y(output_11_85));
wire output_13_85, output_13_6, output_12_85;
mixer gate_output_12_85(.a(output_13_85), .b(output_13_6), .y(output_12_85));
wire output_14_85, output_14_6, output_13_85;
mixer gate_output_13_85(.a(output_14_85), .b(output_14_6), .y(output_13_85));
wire output_15_85, output_15_6, output_14_85;
mixer gate_output_14_85(.a(output_15_85), .b(output_15_6), .y(output_14_85));
wire output_16_85, output_16_6, output_15_85;
mixer gate_output_15_85(.a(output_16_85), .b(output_16_6), .y(output_15_85));
wire output_1_86, output_1_7, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_7), .y(output_0_86));
wire output_2_86, output_2_7, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_7), .y(output_1_86));
wire output_3_86, output_3_7, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_7), .y(output_2_86));
wire output_4_86, output_4_7, output_3_86;
mixer gate_output_3_86(.a(output_4_86), .b(output_4_7), .y(output_3_86));
wire output_5_86, output_5_7, output_4_86;
mixer gate_output_4_86(.a(output_5_86), .b(output_5_7), .y(output_4_86));
wire output_6_86, output_6_7, output_5_86;
mixer gate_output_5_86(.a(output_6_86), .b(output_6_7), .y(output_5_86));
wire output_7_86, output_7_7, output_6_86;
mixer gate_output_6_86(.a(output_7_86), .b(output_7_7), .y(output_6_86));
wire output_8_86, output_8_7, output_7_86;
mixer gate_output_7_86(.a(output_8_86), .b(output_8_7), .y(output_7_86));
wire output_9_86, output_9_7, output_8_86;
mixer gate_output_8_86(.a(output_9_86), .b(output_9_7), .y(output_8_86));
wire output_10_86, output_10_7, output_9_86;
mixer gate_output_9_86(.a(output_10_86), .b(output_10_7), .y(output_9_86));
wire output_11_86, output_11_7, output_10_86;
mixer gate_output_10_86(.a(output_11_86), .b(output_11_7), .y(output_10_86));
wire output_12_86, output_12_7, output_11_86;
mixer gate_output_11_86(.a(output_12_86), .b(output_12_7), .y(output_11_86));
wire output_13_86, output_13_7, output_12_86;
mixer gate_output_12_86(.a(output_13_86), .b(output_13_7), .y(output_12_86));
wire output_14_86, output_14_7, output_13_86;
mixer gate_output_13_86(.a(output_14_86), .b(output_14_7), .y(output_13_86));
wire output_15_86, output_15_7, output_14_86;
mixer gate_output_14_86(.a(output_15_86), .b(output_15_7), .y(output_14_86));
wire output_16_86, output_16_7, output_15_86;
mixer gate_output_15_86(.a(output_16_86), .b(output_16_7), .y(output_15_86));
wire output_1_87, output_1_8, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_8), .y(output_0_87));
wire output_2_87, output_2_8, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_8), .y(output_1_87));
wire output_3_87, output_3_8, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_8), .y(output_2_87));
wire output_4_87, output_4_8, output_3_87;
mixer gate_output_3_87(.a(output_4_87), .b(output_4_8), .y(output_3_87));
wire output_5_87, output_5_8, output_4_87;
mixer gate_output_4_87(.a(output_5_87), .b(output_5_8), .y(output_4_87));
wire output_6_87, output_6_8, output_5_87;
mixer gate_output_5_87(.a(output_6_87), .b(output_6_8), .y(output_5_87));
wire output_7_87, output_7_8, output_6_87;
mixer gate_output_6_87(.a(output_7_87), .b(output_7_8), .y(output_6_87));
wire output_8_87, output_8_8, output_7_87;
mixer gate_output_7_87(.a(output_8_87), .b(output_8_8), .y(output_7_87));
wire output_9_87, output_9_8, output_8_87;
mixer gate_output_8_87(.a(output_9_87), .b(output_9_8), .y(output_8_87));
wire output_10_87, output_10_8, output_9_87;
mixer gate_output_9_87(.a(output_10_87), .b(output_10_8), .y(output_9_87));
wire output_11_87, output_11_8, output_10_87;
mixer gate_output_10_87(.a(output_11_87), .b(output_11_8), .y(output_10_87));
wire output_12_87, output_12_8, output_11_87;
mixer gate_output_11_87(.a(output_12_87), .b(output_12_8), .y(output_11_87));
wire output_13_87, output_13_8, output_12_87;
mixer gate_output_12_87(.a(output_13_87), .b(output_13_8), .y(output_12_87));
wire output_14_87, output_14_8, output_13_87;
mixer gate_output_13_87(.a(output_14_87), .b(output_14_8), .y(output_13_87));
wire output_15_87, output_15_8, output_14_87;
mixer gate_output_14_87(.a(output_15_87), .b(output_15_8), .y(output_14_87));
wire output_16_87, output_16_8, output_15_87;
mixer gate_output_15_87(.a(output_16_87), .b(output_16_8), .y(output_15_87));
wire output_1_88, output_1_9, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_9), .y(output_0_88));
wire output_2_88, output_2_9, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_9), .y(output_1_88));
wire output_3_88, output_3_9, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_9), .y(output_2_88));
wire output_4_88, output_4_9, output_3_88;
mixer gate_output_3_88(.a(output_4_88), .b(output_4_9), .y(output_3_88));
wire output_5_88, output_5_9, output_4_88;
mixer gate_output_4_88(.a(output_5_88), .b(output_5_9), .y(output_4_88));
wire output_6_88, output_6_9, output_5_88;
mixer gate_output_5_88(.a(output_6_88), .b(output_6_9), .y(output_5_88));
wire output_7_88, output_7_9, output_6_88;
mixer gate_output_6_88(.a(output_7_88), .b(output_7_9), .y(output_6_88));
wire output_8_88, output_8_9, output_7_88;
mixer gate_output_7_88(.a(output_8_88), .b(output_8_9), .y(output_7_88));
wire output_9_88, output_9_9, output_8_88;
mixer gate_output_8_88(.a(output_9_88), .b(output_9_9), .y(output_8_88));
wire output_10_88, output_10_9, output_9_88;
mixer gate_output_9_88(.a(output_10_88), .b(output_10_9), .y(output_9_88));
wire output_11_88, output_11_9, output_10_88;
mixer gate_output_10_88(.a(output_11_88), .b(output_11_9), .y(output_10_88));
wire output_12_88, output_12_9, output_11_88;
mixer gate_output_11_88(.a(output_12_88), .b(output_12_9), .y(output_11_88));
wire output_13_88, output_13_9, output_12_88;
mixer gate_output_12_88(.a(output_13_88), .b(output_13_9), .y(output_12_88));
wire output_14_88, output_14_9, output_13_88;
mixer gate_output_13_88(.a(output_14_88), .b(output_14_9), .y(output_13_88));
wire output_15_88, output_15_9, output_14_88;
mixer gate_output_14_88(.a(output_15_88), .b(output_15_9), .y(output_14_88));
wire output_16_88, output_16_9, output_15_88;
mixer gate_output_15_88(.a(output_16_88), .b(output_16_9), .y(output_15_88));
wire output_1_89, output_1_10, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_10), .y(output_0_89));
wire output_2_89, output_2_10, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_10), .y(output_1_89));
wire output_3_89, output_3_10, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_10), .y(output_2_89));
wire output_4_89, output_4_10, output_3_89;
mixer gate_output_3_89(.a(output_4_89), .b(output_4_10), .y(output_3_89));
wire output_5_89, output_5_10, output_4_89;
mixer gate_output_4_89(.a(output_5_89), .b(output_5_10), .y(output_4_89));
wire output_6_89, output_6_10, output_5_89;
mixer gate_output_5_89(.a(output_6_89), .b(output_6_10), .y(output_5_89));
wire output_7_89, output_7_10, output_6_89;
mixer gate_output_6_89(.a(output_7_89), .b(output_7_10), .y(output_6_89));
wire output_8_89, output_8_10, output_7_89;
mixer gate_output_7_89(.a(output_8_89), .b(output_8_10), .y(output_7_89));
wire output_9_89, output_9_10, output_8_89;
mixer gate_output_8_89(.a(output_9_89), .b(output_9_10), .y(output_8_89));
wire output_10_89, output_10_10, output_9_89;
mixer gate_output_9_89(.a(output_10_89), .b(output_10_10), .y(output_9_89));
wire output_11_89, output_11_10, output_10_89;
mixer gate_output_10_89(.a(output_11_89), .b(output_11_10), .y(output_10_89));
wire output_12_89, output_12_10, output_11_89;
mixer gate_output_11_89(.a(output_12_89), .b(output_12_10), .y(output_11_89));
wire output_13_89, output_13_10, output_12_89;
mixer gate_output_12_89(.a(output_13_89), .b(output_13_10), .y(output_12_89));
wire output_14_89, output_14_10, output_13_89;
mixer gate_output_13_89(.a(output_14_89), .b(output_14_10), .y(output_13_89));
wire output_15_89, output_15_10, output_14_89;
mixer gate_output_14_89(.a(output_15_89), .b(output_15_10), .y(output_14_89));
wire output_16_89, output_16_10, output_15_89;
mixer gate_output_15_89(.a(output_16_89), .b(output_16_10), .y(output_15_89));
wire output_1_90, output_1_11, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_11), .y(output_0_90));
wire output_2_90, output_2_11, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_11), .y(output_1_90));
wire output_3_90, output_3_11, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_11), .y(output_2_90));
wire output_4_90, output_4_11, output_3_90;
mixer gate_output_3_90(.a(output_4_90), .b(output_4_11), .y(output_3_90));
wire output_5_90, output_5_11, output_4_90;
mixer gate_output_4_90(.a(output_5_90), .b(output_5_11), .y(output_4_90));
wire output_6_90, output_6_11, output_5_90;
mixer gate_output_5_90(.a(output_6_90), .b(output_6_11), .y(output_5_90));
wire output_7_90, output_7_11, output_6_90;
mixer gate_output_6_90(.a(output_7_90), .b(output_7_11), .y(output_6_90));
wire output_8_90, output_8_11, output_7_90;
mixer gate_output_7_90(.a(output_8_90), .b(output_8_11), .y(output_7_90));
wire output_9_90, output_9_11, output_8_90;
mixer gate_output_8_90(.a(output_9_90), .b(output_9_11), .y(output_8_90));
wire output_10_90, output_10_11, output_9_90;
mixer gate_output_9_90(.a(output_10_90), .b(output_10_11), .y(output_9_90));
wire output_11_90, output_11_11, output_10_90;
mixer gate_output_10_90(.a(output_11_90), .b(output_11_11), .y(output_10_90));
wire output_12_90, output_12_11, output_11_90;
mixer gate_output_11_90(.a(output_12_90), .b(output_12_11), .y(output_11_90));
wire output_13_90, output_13_11, output_12_90;
mixer gate_output_12_90(.a(output_13_90), .b(output_13_11), .y(output_12_90));
wire output_14_90, output_14_11, output_13_90;
mixer gate_output_13_90(.a(output_14_90), .b(output_14_11), .y(output_13_90));
wire output_15_90, output_15_11, output_14_90;
mixer gate_output_14_90(.a(output_15_90), .b(output_15_11), .y(output_14_90));
wire output_16_90, output_16_11, output_15_90;
mixer gate_output_15_90(.a(output_16_90), .b(output_16_11), .y(output_15_90));
wire output_1_91, output_1_12, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_12), .y(output_0_91));
wire output_2_91, output_2_12, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_12), .y(output_1_91));
wire output_3_91, output_3_12, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_12), .y(output_2_91));
wire output_4_91, output_4_12, output_3_91;
mixer gate_output_3_91(.a(output_4_91), .b(output_4_12), .y(output_3_91));
wire output_5_91, output_5_12, output_4_91;
mixer gate_output_4_91(.a(output_5_91), .b(output_5_12), .y(output_4_91));
wire output_6_91, output_6_12, output_5_91;
mixer gate_output_5_91(.a(output_6_91), .b(output_6_12), .y(output_5_91));
wire output_7_91, output_7_12, output_6_91;
mixer gate_output_6_91(.a(output_7_91), .b(output_7_12), .y(output_6_91));
wire output_8_91, output_8_12, output_7_91;
mixer gate_output_7_91(.a(output_8_91), .b(output_8_12), .y(output_7_91));
wire output_9_91, output_9_12, output_8_91;
mixer gate_output_8_91(.a(output_9_91), .b(output_9_12), .y(output_8_91));
wire output_10_91, output_10_12, output_9_91;
mixer gate_output_9_91(.a(output_10_91), .b(output_10_12), .y(output_9_91));
wire output_11_91, output_11_12, output_10_91;
mixer gate_output_10_91(.a(output_11_91), .b(output_11_12), .y(output_10_91));
wire output_12_91, output_12_12, output_11_91;
mixer gate_output_11_91(.a(output_12_91), .b(output_12_12), .y(output_11_91));
wire output_13_91, output_13_12, output_12_91;
mixer gate_output_12_91(.a(output_13_91), .b(output_13_12), .y(output_12_91));
wire output_14_91, output_14_12, output_13_91;
mixer gate_output_13_91(.a(output_14_91), .b(output_14_12), .y(output_13_91));
wire output_15_91, output_15_12, output_14_91;
mixer gate_output_14_91(.a(output_15_91), .b(output_15_12), .y(output_14_91));
wire output_16_91, output_16_12, output_15_91;
mixer gate_output_15_91(.a(output_16_91), .b(output_16_12), .y(output_15_91));
wire output_1_92, output_1_13, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_13), .y(output_0_92));
wire output_2_92, output_2_13, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_13), .y(output_1_92));
wire output_3_92, output_3_13, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_13), .y(output_2_92));
wire output_4_92, output_4_13, output_3_92;
mixer gate_output_3_92(.a(output_4_92), .b(output_4_13), .y(output_3_92));
wire output_5_92, output_5_13, output_4_92;
mixer gate_output_4_92(.a(output_5_92), .b(output_5_13), .y(output_4_92));
wire output_6_92, output_6_13, output_5_92;
mixer gate_output_5_92(.a(output_6_92), .b(output_6_13), .y(output_5_92));
wire output_7_92, output_7_13, output_6_92;
mixer gate_output_6_92(.a(output_7_92), .b(output_7_13), .y(output_6_92));
wire output_8_92, output_8_13, output_7_92;
mixer gate_output_7_92(.a(output_8_92), .b(output_8_13), .y(output_7_92));
wire output_9_92, output_9_13, output_8_92;
mixer gate_output_8_92(.a(output_9_92), .b(output_9_13), .y(output_8_92));
wire output_10_92, output_10_13, output_9_92;
mixer gate_output_9_92(.a(output_10_92), .b(output_10_13), .y(output_9_92));
wire output_11_92, output_11_13, output_10_92;
mixer gate_output_10_92(.a(output_11_92), .b(output_11_13), .y(output_10_92));
wire output_12_92, output_12_13, output_11_92;
mixer gate_output_11_92(.a(output_12_92), .b(output_12_13), .y(output_11_92));
wire output_13_92, output_13_13, output_12_92;
mixer gate_output_12_92(.a(output_13_92), .b(output_13_13), .y(output_12_92));
wire output_14_92, output_14_13, output_13_92;
mixer gate_output_13_92(.a(output_14_92), .b(output_14_13), .y(output_13_92));
wire output_15_92, output_15_13, output_14_92;
mixer gate_output_14_92(.a(output_15_92), .b(output_15_13), .y(output_14_92));
wire output_16_92, output_16_13, output_15_92;
mixer gate_output_15_92(.a(output_16_92), .b(output_16_13), .y(output_15_92));
wire output_1_93, output_1_14, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_14), .y(output_0_93));
wire output_2_93, output_2_14, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_14), .y(output_1_93));
wire output_3_93, output_3_14, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_14), .y(output_2_93));
wire output_4_93, output_4_14, output_3_93;
mixer gate_output_3_93(.a(output_4_93), .b(output_4_14), .y(output_3_93));
wire output_5_93, output_5_14, output_4_93;
mixer gate_output_4_93(.a(output_5_93), .b(output_5_14), .y(output_4_93));
wire output_6_93, output_6_14, output_5_93;
mixer gate_output_5_93(.a(output_6_93), .b(output_6_14), .y(output_5_93));
wire output_7_93, output_7_14, output_6_93;
mixer gate_output_6_93(.a(output_7_93), .b(output_7_14), .y(output_6_93));
wire output_8_93, output_8_14, output_7_93;
mixer gate_output_7_93(.a(output_8_93), .b(output_8_14), .y(output_7_93));
wire output_9_93, output_9_14, output_8_93;
mixer gate_output_8_93(.a(output_9_93), .b(output_9_14), .y(output_8_93));
wire output_10_93, output_10_14, output_9_93;
mixer gate_output_9_93(.a(output_10_93), .b(output_10_14), .y(output_9_93));
wire output_11_93, output_11_14, output_10_93;
mixer gate_output_10_93(.a(output_11_93), .b(output_11_14), .y(output_10_93));
wire output_12_93, output_12_14, output_11_93;
mixer gate_output_11_93(.a(output_12_93), .b(output_12_14), .y(output_11_93));
wire output_13_93, output_13_14, output_12_93;
mixer gate_output_12_93(.a(output_13_93), .b(output_13_14), .y(output_12_93));
wire output_14_93, output_14_14, output_13_93;
mixer gate_output_13_93(.a(output_14_93), .b(output_14_14), .y(output_13_93));
wire output_15_93, output_15_14, output_14_93;
mixer gate_output_14_93(.a(output_15_93), .b(output_15_14), .y(output_14_93));
wire output_16_93, output_16_14, output_15_93;
mixer gate_output_15_93(.a(output_16_93), .b(output_16_14), .y(output_15_93));
wire output_1_94, output_1_15, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_15), .y(output_0_94));
wire output_2_94, output_2_15, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_15), .y(output_1_94));
wire output_3_94, output_3_15, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_15), .y(output_2_94));
wire output_4_94, output_4_15, output_3_94;
mixer gate_output_3_94(.a(output_4_94), .b(output_4_15), .y(output_3_94));
wire output_5_94, output_5_15, output_4_94;
mixer gate_output_4_94(.a(output_5_94), .b(output_5_15), .y(output_4_94));
wire output_6_94, output_6_15, output_5_94;
mixer gate_output_5_94(.a(output_6_94), .b(output_6_15), .y(output_5_94));
wire output_7_94, output_7_15, output_6_94;
mixer gate_output_6_94(.a(output_7_94), .b(output_7_15), .y(output_6_94));
wire output_8_94, output_8_15, output_7_94;
mixer gate_output_7_94(.a(output_8_94), .b(output_8_15), .y(output_7_94));
wire output_9_94, output_9_15, output_8_94;
mixer gate_output_8_94(.a(output_9_94), .b(output_9_15), .y(output_8_94));
wire output_10_94, output_10_15, output_9_94;
mixer gate_output_9_94(.a(output_10_94), .b(output_10_15), .y(output_9_94));
wire output_11_94, output_11_15, output_10_94;
mixer gate_output_10_94(.a(output_11_94), .b(output_11_15), .y(output_10_94));
wire output_12_94, output_12_15, output_11_94;
mixer gate_output_11_94(.a(output_12_94), .b(output_12_15), .y(output_11_94));
wire output_13_94, output_13_15, output_12_94;
mixer gate_output_12_94(.a(output_13_94), .b(output_13_15), .y(output_12_94));
wire output_14_94, output_14_15, output_13_94;
mixer gate_output_13_94(.a(output_14_94), .b(output_14_15), .y(output_13_94));
wire output_15_94, output_15_15, output_14_94;
mixer gate_output_14_94(.a(output_15_94), .b(output_15_15), .y(output_14_94));
wire output_16_94, output_16_15, output_15_94;
mixer gate_output_15_94(.a(output_16_94), .b(output_16_15), .y(output_15_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_4_95, output_4_0, output_3_95;
mixer gate_output_3_95(.a(output_4_95), .b(output_4_0), .y(output_3_95));
wire output_5_95, output_5_0, output_4_95;
mixer gate_output_4_95(.a(output_5_95), .b(output_5_0), .y(output_4_95));
wire output_6_95, output_6_0, output_5_95;
mixer gate_output_5_95(.a(output_6_95), .b(output_6_0), .y(output_5_95));
wire output_7_95, output_7_0, output_6_95;
mixer gate_output_6_95(.a(output_7_95), .b(output_7_0), .y(output_6_95));
wire output_8_95, output_8_0, output_7_95;
mixer gate_output_7_95(.a(output_8_95), .b(output_8_0), .y(output_7_95));
wire output_9_95, output_9_0, output_8_95;
mixer gate_output_8_95(.a(output_9_95), .b(output_9_0), .y(output_8_95));
wire output_10_95, output_10_0, output_9_95;
mixer gate_output_9_95(.a(output_10_95), .b(output_10_0), .y(output_9_95));
wire output_11_95, output_11_0, output_10_95;
mixer gate_output_10_95(.a(output_11_95), .b(output_11_0), .y(output_10_95));
wire output_12_95, output_12_0, output_11_95;
mixer gate_output_11_95(.a(output_12_95), .b(output_12_0), .y(output_11_95));
wire output_13_95, output_13_0, output_12_95;
mixer gate_output_12_95(.a(output_13_95), .b(output_13_0), .y(output_12_95));
wire output_14_95, output_14_0, output_13_95;
mixer gate_output_13_95(.a(output_14_95), .b(output_14_0), .y(output_13_95));
wire output_15_95, output_15_0, output_14_95;
mixer gate_output_14_95(.a(output_15_95), .b(output_15_0), .y(output_14_95));
wire output_16_95, output_16_0, output_15_95;
mixer gate_output_15_95(.a(output_16_95), .b(output_16_0), .y(output_15_95));
wire output_1_96, output_1_1, output_0_96;
mixer gate_output_0_96(.a(output_1_96), .b(output_1_1), .y(output_0_96));
wire output_2_96, output_2_1, output_1_96;
mixer gate_output_1_96(.a(output_2_96), .b(output_2_1), .y(output_1_96));
wire output_3_96, output_3_1, output_2_96;
mixer gate_output_2_96(.a(output_3_96), .b(output_3_1), .y(output_2_96));
wire output_4_96, output_4_1, output_3_96;
mixer gate_output_3_96(.a(output_4_96), .b(output_4_1), .y(output_3_96));
wire output_5_96, output_5_1, output_4_96;
mixer gate_output_4_96(.a(output_5_96), .b(output_5_1), .y(output_4_96));
wire output_6_96, output_6_1, output_5_96;
mixer gate_output_5_96(.a(output_6_96), .b(output_6_1), .y(output_5_96));
wire output_7_96, output_7_1, output_6_96;
mixer gate_output_6_96(.a(output_7_96), .b(output_7_1), .y(output_6_96));
wire output_8_96, output_8_1, output_7_96;
mixer gate_output_7_96(.a(output_8_96), .b(output_8_1), .y(output_7_96));
wire output_9_96, output_9_1, output_8_96;
mixer gate_output_8_96(.a(output_9_96), .b(output_9_1), .y(output_8_96));
wire output_10_96, output_10_1, output_9_96;
mixer gate_output_9_96(.a(output_10_96), .b(output_10_1), .y(output_9_96));
wire output_11_96, output_11_1, output_10_96;
mixer gate_output_10_96(.a(output_11_96), .b(output_11_1), .y(output_10_96));
wire output_12_96, output_12_1, output_11_96;
mixer gate_output_11_96(.a(output_12_96), .b(output_12_1), .y(output_11_96));
wire output_13_96, output_13_1, output_12_96;
mixer gate_output_12_96(.a(output_13_96), .b(output_13_1), .y(output_12_96));
wire output_14_96, output_14_1, output_13_96;
mixer gate_output_13_96(.a(output_14_96), .b(output_14_1), .y(output_13_96));
wire output_15_96, output_15_1, output_14_96;
mixer gate_output_14_96(.a(output_15_96), .b(output_15_1), .y(output_14_96));
wire output_16_96, output_16_1, output_15_96;
mixer gate_output_15_96(.a(output_16_96), .b(output_16_1), .y(output_15_96));
wire output_1_97, output_1_2, output_0_97;
mixer gate_output_0_97(.a(output_1_97), .b(output_1_2), .y(output_0_97));
wire output_2_97, output_2_2, output_1_97;
mixer gate_output_1_97(.a(output_2_97), .b(output_2_2), .y(output_1_97));
wire output_3_97, output_3_2, output_2_97;
mixer gate_output_2_97(.a(output_3_97), .b(output_3_2), .y(output_2_97));
wire output_4_97, output_4_2, output_3_97;
mixer gate_output_3_97(.a(output_4_97), .b(output_4_2), .y(output_3_97));
wire output_5_97, output_5_2, output_4_97;
mixer gate_output_4_97(.a(output_5_97), .b(output_5_2), .y(output_4_97));
wire output_6_97, output_6_2, output_5_97;
mixer gate_output_5_97(.a(output_6_97), .b(output_6_2), .y(output_5_97));
wire output_7_97, output_7_2, output_6_97;
mixer gate_output_6_97(.a(output_7_97), .b(output_7_2), .y(output_6_97));
wire output_8_97, output_8_2, output_7_97;
mixer gate_output_7_97(.a(output_8_97), .b(output_8_2), .y(output_7_97));
wire output_9_97, output_9_2, output_8_97;
mixer gate_output_8_97(.a(output_9_97), .b(output_9_2), .y(output_8_97));
wire output_10_97, output_10_2, output_9_97;
mixer gate_output_9_97(.a(output_10_97), .b(output_10_2), .y(output_9_97));
wire output_11_97, output_11_2, output_10_97;
mixer gate_output_10_97(.a(output_11_97), .b(output_11_2), .y(output_10_97));
wire output_12_97, output_12_2, output_11_97;
mixer gate_output_11_97(.a(output_12_97), .b(output_12_2), .y(output_11_97));
wire output_13_97, output_13_2, output_12_97;
mixer gate_output_12_97(.a(output_13_97), .b(output_13_2), .y(output_12_97));
wire output_14_97, output_14_2, output_13_97;
mixer gate_output_13_97(.a(output_14_97), .b(output_14_2), .y(output_13_97));
wire output_15_97, output_15_2, output_14_97;
mixer gate_output_14_97(.a(output_15_97), .b(output_15_2), .y(output_14_97));
wire output_16_97, output_16_2, output_15_97;
mixer gate_output_15_97(.a(output_16_97), .b(output_16_2), .y(output_15_97));
wire output_1_98, output_1_3, output_0_98;
mixer gate_output_0_98(.a(output_1_98), .b(output_1_3), .y(output_0_98));
wire output_2_98, output_2_3, output_1_98;
mixer gate_output_1_98(.a(output_2_98), .b(output_2_3), .y(output_1_98));
wire output_3_98, output_3_3, output_2_98;
mixer gate_output_2_98(.a(output_3_98), .b(output_3_3), .y(output_2_98));
wire output_4_98, output_4_3, output_3_98;
mixer gate_output_3_98(.a(output_4_98), .b(output_4_3), .y(output_3_98));
wire output_5_98, output_5_3, output_4_98;
mixer gate_output_4_98(.a(output_5_98), .b(output_5_3), .y(output_4_98));
wire output_6_98, output_6_3, output_5_98;
mixer gate_output_5_98(.a(output_6_98), .b(output_6_3), .y(output_5_98));
wire output_7_98, output_7_3, output_6_98;
mixer gate_output_6_98(.a(output_7_98), .b(output_7_3), .y(output_6_98));
wire output_8_98, output_8_3, output_7_98;
mixer gate_output_7_98(.a(output_8_98), .b(output_8_3), .y(output_7_98));
wire output_9_98, output_9_3, output_8_98;
mixer gate_output_8_98(.a(output_9_98), .b(output_9_3), .y(output_8_98));
wire output_10_98, output_10_3, output_9_98;
mixer gate_output_9_98(.a(output_10_98), .b(output_10_3), .y(output_9_98));
wire output_11_98, output_11_3, output_10_98;
mixer gate_output_10_98(.a(output_11_98), .b(output_11_3), .y(output_10_98));
wire output_12_98, output_12_3, output_11_98;
mixer gate_output_11_98(.a(output_12_98), .b(output_12_3), .y(output_11_98));
wire output_13_98, output_13_3, output_12_98;
mixer gate_output_12_98(.a(output_13_98), .b(output_13_3), .y(output_12_98));
wire output_14_98, output_14_3, output_13_98;
mixer gate_output_13_98(.a(output_14_98), .b(output_14_3), .y(output_13_98));
wire output_15_98, output_15_3, output_14_98;
mixer gate_output_14_98(.a(output_15_98), .b(output_15_3), .y(output_14_98));
wire output_16_98, output_16_3, output_15_98;
mixer gate_output_15_98(.a(output_16_98), .b(output_16_3), .y(output_15_98));
wire output_1_99, output_1_4, output_0_99;
mixer gate_output_0_99(.a(output_1_99), .b(output_1_4), .y(output_0_99));
wire output_2_99, output_2_4, output_1_99;
mixer gate_output_1_99(.a(output_2_99), .b(output_2_4), .y(output_1_99));
wire output_3_99, output_3_4, output_2_99;
mixer gate_output_2_99(.a(output_3_99), .b(output_3_4), .y(output_2_99));
wire output_4_99, output_4_4, output_3_99;
mixer gate_output_3_99(.a(output_4_99), .b(output_4_4), .y(output_3_99));
wire output_5_99, output_5_4, output_4_99;
mixer gate_output_4_99(.a(output_5_99), .b(output_5_4), .y(output_4_99));
wire output_6_99, output_6_4, output_5_99;
mixer gate_output_5_99(.a(output_6_99), .b(output_6_4), .y(output_5_99));
wire output_7_99, output_7_4, output_6_99;
mixer gate_output_6_99(.a(output_7_99), .b(output_7_4), .y(output_6_99));
wire output_8_99, output_8_4, output_7_99;
mixer gate_output_7_99(.a(output_8_99), .b(output_8_4), .y(output_7_99));
wire output_9_99, output_9_4, output_8_99;
mixer gate_output_8_99(.a(output_9_99), .b(output_9_4), .y(output_8_99));
wire output_10_99, output_10_4, output_9_99;
mixer gate_output_9_99(.a(output_10_99), .b(output_10_4), .y(output_9_99));
wire output_11_99, output_11_4, output_10_99;
mixer gate_output_10_99(.a(output_11_99), .b(output_11_4), .y(output_10_99));
wire output_12_99, output_12_4, output_11_99;
mixer gate_output_11_99(.a(output_12_99), .b(output_12_4), .y(output_11_99));
wire output_13_99, output_13_4, output_12_99;
mixer gate_output_12_99(.a(output_13_99), .b(output_13_4), .y(output_12_99));
wire output_14_99, output_14_4, output_13_99;
mixer gate_output_13_99(.a(output_14_99), .b(output_14_4), .y(output_13_99));
wire output_15_99, output_15_4, output_14_99;
mixer gate_output_14_99(.a(output_15_99), .b(output_15_4), .y(output_14_99));
wire output_16_99, output_16_4, output_15_99;
mixer gate_output_15_99(.a(output_16_99), .b(output_16_4), .y(output_15_99));
wire output_1_100, output_1_5, output_0_100;
mixer gate_output_0_100(.a(output_1_100), .b(output_1_5), .y(output_0_100));
wire output_2_100, output_2_5, output_1_100;
mixer gate_output_1_100(.a(output_2_100), .b(output_2_5), .y(output_1_100));
wire output_3_100, output_3_5, output_2_100;
mixer gate_output_2_100(.a(output_3_100), .b(output_3_5), .y(output_2_100));
wire output_4_100, output_4_5, output_3_100;
mixer gate_output_3_100(.a(output_4_100), .b(output_4_5), .y(output_3_100));
wire output_5_100, output_5_5, output_4_100;
mixer gate_output_4_100(.a(output_5_100), .b(output_5_5), .y(output_4_100));
wire output_6_100, output_6_5, output_5_100;
mixer gate_output_5_100(.a(output_6_100), .b(output_6_5), .y(output_5_100));
wire output_7_100, output_7_5, output_6_100;
mixer gate_output_6_100(.a(output_7_100), .b(output_7_5), .y(output_6_100));
wire output_8_100, output_8_5, output_7_100;
mixer gate_output_7_100(.a(output_8_100), .b(output_8_5), .y(output_7_100));
wire output_9_100, output_9_5, output_8_100;
mixer gate_output_8_100(.a(output_9_100), .b(output_9_5), .y(output_8_100));
wire output_10_100, output_10_5, output_9_100;
mixer gate_output_9_100(.a(output_10_100), .b(output_10_5), .y(output_9_100));
wire output_11_100, output_11_5, output_10_100;
mixer gate_output_10_100(.a(output_11_100), .b(output_11_5), .y(output_10_100));
wire output_12_100, output_12_5, output_11_100;
mixer gate_output_11_100(.a(output_12_100), .b(output_12_5), .y(output_11_100));
wire output_13_100, output_13_5, output_12_100;
mixer gate_output_12_100(.a(output_13_100), .b(output_13_5), .y(output_12_100));
wire output_14_100, output_14_5, output_13_100;
mixer gate_output_13_100(.a(output_14_100), .b(output_14_5), .y(output_13_100));
wire output_15_100, output_15_5, output_14_100;
mixer gate_output_14_100(.a(output_15_100), .b(output_15_5), .y(output_14_100));
wire output_16_100, output_16_5, output_15_100;
mixer gate_output_15_100(.a(output_16_100), .b(output_16_5), .y(output_15_100));
wire output_1_101, output_1_6, output_0_101;
mixer gate_output_0_101(.a(output_1_101), .b(output_1_6), .y(output_0_101));
wire output_2_101, output_2_6, output_1_101;
mixer gate_output_1_101(.a(output_2_101), .b(output_2_6), .y(output_1_101));
wire output_3_101, output_3_6, output_2_101;
mixer gate_output_2_101(.a(output_3_101), .b(output_3_6), .y(output_2_101));
wire output_4_101, output_4_6, output_3_101;
mixer gate_output_3_101(.a(output_4_101), .b(output_4_6), .y(output_3_101));
wire output_5_101, output_5_6, output_4_101;
mixer gate_output_4_101(.a(output_5_101), .b(output_5_6), .y(output_4_101));
wire output_6_101, output_6_6, output_5_101;
mixer gate_output_5_101(.a(output_6_101), .b(output_6_6), .y(output_5_101));
wire output_7_101, output_7_6, output_6_101;
mixer gate_output_6_101(.a(output_7_101), .b(output_7_6), .y(output_6_101));
wire output_8_101, output_8_6, output_7_101;
mixer gate_output_7_101(.a(output_8_101), .b(output_8_6), .y(output_7_101));
wire output_9_101, output_9_6, output_8_101;
mixer gate_output_8_101(.a(output_9_101), .b(output_9_6), .y(output_8_101));
wire output_10_101, output_10_6, output_9_101;
mixer gate_output_9_101(.a(output_10_101), .b(output_10_6), .y(output_9_101));
wire output_11_101, output_11_6, output_10_101;
mixer gate_output_10_101(.a(output_11_101), .b(output_11_6), .y(output_10_101));
wire output_12_101, output_12_6, output_11_101;
mixer gate_output_11_101(.a(output_12_101), .b(output_12_6), .y(output_11_101));
wire output_13_101, output_13_6, output_12_101;
mixer gate_output_12_101(.a(output_13_101), .b(output_13_6), .y(output_12_101));
wire output_14_101, output_14_6, output_13_101;
mixer gate_output_13_101(.a(output_14_101), .b(output_14_6), .y(output_13_101));
wire output_15_101, output_15_6, output_14_101;
mixer gate_output_14_101(.a(output_15_101), .b(output_15_6), .y(output_14_101));
wire output_16_101, output_16_6, output_15_101;
mixer gate_output_15_101(.a(output_16_101), .b(output_16_6), .y(output_15_101));
wire output_1_102, output_1_7, output_0_102;
mixer gate_output_0_102(.a(output_1_102), .b(output_1_7), .y(output_0_102));
wire output_2_102, output_2_7, output_1_102;
mixer gate_output_1_102(.a(output_2_102), .b(output_2_7), .y(output_1_102));
wire output_3_102, output_3_7, output_2_102;
mixer gate_output_2_102(.a(output_3_102), .b(output_3_7), .y(output_2_102));
wire output_4_102, output_4_7, output_3_102;
mixer gate_output_3_102(.a(output_4_102), .b(output_4_7), .y(output_3_102));
wire output_5_102, output_5_7, output_4_102;
mixer gate_output_4_102(.a(output_5_102), .b(output_5_7), .y(output_4_102));
wire output_6_102, output_6_7, output_5_102;
mixer gate_output_5_102(.a(output_6_102), .b(output_6_7), .y(output_5_102));
wire output_7_102, output_7_7, output_6_102;
mixer gate_output_6_102(.a(output_7_102), .b(output_7_7), .y(output_6_102));
wire output_8_102, output_8_7, output_7_102;
mixer gate_output_7_102(.a(output_8_102), .b(output_8_7), .y(output_7_102));
wire output_9_102, output_9_7, output_8_102;
mixer gate_output_8_102(.a(output_9_102), .b(output_9_7), .y(output_8_102));
wire output_10_102, output_10_7, output_9_102;
mixer gate_output_9_102(.a(output_10_102), .b(output_10_7), .y(output_9_102));
wire output_11_102, output_11_7, output_10_102;
mixer gate_output_10_102(.a(output_11_102), .b(output_11_7), .y(output_10_102));
wire output_12_102, output_12_7, output_11_102;
mixer gate_output_11_102(.a(output_12_102), .b(output_12_7), .y(output_11_102));
wire output_13_102, output_13_7, output_12_102;
mixer gate_output_12_102(.a(output_13_102), .b(output_13_7), .y(output_12_102));
wire output_14_102, output_14_7, output_13_102;
mixer gate_output_13_102(.a(output_14_102), .b(output_14_7), .y(output_13_102));
wire output_15_102, output_15_7, output_14_102;
mixer gate_output_14_102(.a(output_15_102), .b(output_15_7), .y(output_14_102));
wire output_16_102, output_16_7, output_15_102;
mixer gate_output_15_102(.a(output_16_102), .b(output_16_7), .y(output_15_102));
wire output_1_103, output_1_8, output_0_103;
mixer gate_output_0_103(.a(output_1_103), .b(output_1_8), .y(output_0_103));
wire output_2_103, output_2_8, output_1_103;
mixer gate_output_1_103(.a(output_2_103), .b(output_2_8), .y(output_1_103));
wire output_3_103, output_3_8, output_2_103;
mixer gate_output_2_103(.a(output_3_103), .b(output_3_8), .y(output_2_103));
wire output_4_103, output_4_8, output_3_103;
mixer gate_output_3_103(.a(output_4_103), .b(output_4_8), .y(output_3_103));
wire output_5_103, output_5_8, output_4_103;
mixer gate_output_4_103(.a(output_5_103), .b(output_5_8), .y(output_4_103));
wire output_6_103, output_6_8, output_5_103;
mixer gate_output_5_103(.a(output_6_103), .b(output_6_8), .y(output_5_103));
wire output_7_103, output_7_8, output_6_103;
mixer gate_output_6_103(.a(output_7_103), .b(output_7_8), .y(output_6_103));
wire output_8_103, output_8_8, output_7_103;
mixer gate_output_7_103(.a(output_8_103), .b(output_8_8), .y(output_7_103));
wire output_9_103, output_9_8, output_8_103;
mixer gate_output_8_103(.a(output_9_103), .b(output_9_8), .y(output_8_103));
wire output_10_103, output_10_8, output_9_103;
mixer gate_output_9_103(.a(output_10_103), .b(output_10_8), .y(output_9_103));
wire output_11_103, output_11_8, output_10_103;
mixer gate_output_10_103(.a(output_11_103), .b(output_11_8), .y(output_10_103));
wire output_12_103, output_12_8, output_11_103;
mixer gate_output_11_103(.a(output_12_103), .b(output_12_8), .y(output_11_103));
wire output_13_103, output_13_8, output_12_103;
mixer gate_output_12_103(.a(output_13_103), .b(output_13_8), .y(output_12_103));
wire output_14_103, output_14_8, output_13_103;
mixer gate_output_13_103(.a(output_14_103), .b(output_14_8), .y(output_13_103));
wire output_15_103, output_15_8, output_14_103;
mixer gate_output_14_103(.a(output_15_103), .b(output_15_8), .y(output_14_103));
wire output_16_103, output_16_8, output_15_103;
mixer gate_output_15_103(.a(output_16_103), .b(output_16_8), .y(output_15_103));
wire output_1_104, output_1_9, output_0_104;
mixer gate_output_0_104(.a(output_1_104), .b(output_1_9), .y(output_0_104));
wire output_2_104, output_2_9, output_1_104;
mixer gate_output_1_104(.a(output_2_104), .b(output_2_9), .y(output_1_104));
wire output_3_104, output_3_9, output_2_104;
mixer gate_output_2_104(.a(output_3_104), .b(output_3_9), .y(output_2_104));
wire output_4_104, output_4_9, output_3_104;
mixer gate_output_3_104(.a(output_4_104), .b(output_4_9), .y(output_3_104));
wire output_5_104, output_5_9, output_4_104;
mixer gate_output_4_104(.a(output_5_104), .b(output_5_9), .y(output_4_104));
wire output_6_104, output_6_9, output_5_104;
mixer gate_output_5_104(.a(output_6_104), .b(output_6_9), .y(output_5_104));
wire output_7_104, output_7_9, output_6_104;
mixer gate_output_6_104(.a(output_7_104), .b(output_7_9), .y(output_6_104));
wire output_8_104, output_8_9, output_7_104;
mixer gate_output_7_104(.a(output_8_104), .b(output_8_9), .y(output_7_104));
wire output_9_104, output_9_9, output_8_104;
mixer gate_output_8_104(.a(output_9_104), .b(output_9_9), .y(output_8_104));
wire output_10_104, output_10_9, output_9_104;
mixer gate_output_9_104(.a(output_10_104), .b(output_10_9), .y(output_9_104));
wire output_11_104, output_11_9, output_10_104;
mixer gate_output_10_104(.a(output_11_104), .b(output_11_9), .y(output_10_104));
wire output_12_104, output_12_9, output_11_104;
mixer gate_output_11_104(.a(output_12_104), .b(output_12_9), .y(output_11_104));
wire output_13_104, output_13_9, output_12_104;
mixer gate_output_12_104(.a(output_13_104), .b(output_13_9), .y(output_12_104));
wire output_14_104, output_14_9, output_13_104;
mixer gate_output_13_104(.a(output_14_104), .b(output_14_9), .y(output_13_104));
wire output_15_104, output_15_9, output_14_104;
mixer gate_output_14_104(.a(output_15_104), .b(output_15_9), .y(output_14_104));
wire output_16_104, output_16_9, output_15_104;
mixer gate_output_15_104(.a(output_16_104), .b(output_16_9), .y(output_15_104));
wire output_1_105, output_1_10, output_0_105;
mixer gate_output_0_105(.a(output_1_105), .b(output_1_10), .y(output_0_105));
wire output_2_105, output_2_10, output_1_105;
mixer gate_output_1_105(.a(output_2_105), .b(output_2_10), .y(output_1_105));
wire output_3_105, output_3_10, output_2_105;
mixer gate_output_2_105(.a(output_3_105), .b(output_3_10), .y(output_2_105));
wire output_4_105, output_4_10, output_3_105;
mixer gate_output_3_105(.a(output_4_105), .b(output_4_10), .y(output_3_105));
wire output_5_105, output_5_10, output_4_105;
mixer gate_output_4_105(.a(output_5_105), .b(output_5_10), .y(output_4_105));
wire output_6_105, output_6_10, output_5_105;
mixer gate_output_5_105(.a(output_6_105), .b(output_6_10), .y(output_5_105));
wire output_7_105, output_7_10, output_6_105;
mixer gate_output_6_105(.a(output_7_105), .b(output_7_10), .y(output_6_105));
wire output_8_105, output_8_10, output_7_105;
mixer gate_output_7_105(.a(output_8_105), .b(output_8_10), .y(output_7_105));
wire output_9_105, output_9_10, output_8_105;
mixer gate_output_8_105(.a(output_9_105), .b(output_9_10), .y(output_8_105));
wire output_10_105, output_10_10, output_9_105;
mixer gate_output_9_105(.a(output_10_105), .b(output_10_10), .y(output_9_105));
wire output_11_105, output_11_10, output_10_105;
mixer gate_output_10_105(.a(output_11_105), .b(output_11_10), .y(output_10_105));
wire output_12_105, output_12_10, output_11_105;
mixer gate_output_11_105(.a(output_12_105), .b(output_12_10), .y(output_11_105));
wire output_13_105, output_13_10, output_12_105;
mixer gate_output_12_105(.a(output_13_105), .b(output_13_10), .y(output_12_105));
wire output_14_105, output_14_10, output_13_105;
mixer gate_output_13_105(.a(output_14_105), .b(output_14_10), .y(output_13_105));
wire output_15_105, output_15_10, output_14_105;
mixer gate_output_14_105(.a(output_15_105), .b(output_15_10), .y(output_14_105));
wire output_16_105, output_16_10, output_15_105;
mixer gate_output_15_105(.a(output_16_105), .b(output_16_10), .y(output_15_105));
wire output_1_106, output_1_11, output_0_106;
mixer gate_output_0_106(.a(output_1_106), .b(output_1_11), .y(output_0_106));
wire output_2_106, output_2_11, output_1_106;
mixer gate_output_1_106(.a(output_2_106), .b(output_2_11), .y(output_1_106));
wire output_3_106, output_3_11, output_2_106;
mixer gate_output_2_106(.a(output_3_106), .b(output_3_11), .y(output_2_106));
wire output_4_106, output_4_11, output_3_106;
mixer gate_output_3_106(.a(output_4_106), .b(output_4_11), .y(output_3_106));
wire output_5_106, output_5_11, output_4_106;
mixer gate_output_4_106(.a(output_5_106), .b(output_5_11), .y(output_4_106));
wire output_6_106, output_6_11, output_5_106;
mixer gate_output_5_106(.a(output_6_106), .b(output_6_11), .y(output_5_106));
wire output_7_106, output_7_11, output_6_106;
mixer gate_output_6_106(.a(output_7_106), .b(output_7_11), .y(output_6_106));
wire output_8_106, output_8_11, output_7_106;
mixer gate_output_7_106(.a(output_8_106), .b(output_8_11), .y(output_7_106));
wire output_9_106, output_9_11, output_8_106;
mixer gate_output_8_106(.a(output_9_106), .b(output_9_11), .y(output_8_106));
wire output_10_106, output_10_11, output_9_106;
mixer gate_output_9_106(.a(output_10_106), .b(output_10_11), .y(output_9_106));
wire output_11_106, output_11_11, output_10_106;
mixer gate_output_10_106(.a(output_11_106), .b(output_11_11), .y(output_10_106));
wire output_12_106, output_12_11, output_11_106;
mixer gate_output_11_106(.a(output_12_106), .b(output_12_11), .y(output_11_106));
wire output_13_106, output_13_11, output_12_106;
mixer gate_output_12_106(.a(output_13_106), .b(output_13_11), .y(output_12_106));
wire output_14_106, output_14_11, output_13_106;
mixer gate_output_13_106(.a(output_14_106), .b(output_14_11), .y(output_13_106));
wire output_15_106, output_15_11, output_14_106;
mixer gate_output_14_106(.a(output_15_106), .b(output_15_11), .y(output_14_106));
wire output_16_106, output_16_11, output_15_106;
mixer gate_output_15_106(.a(output_16_106), .b(output_16_11), .y(output_15_106));
wire output_1_107, output_1_12, output_0_107;
mixer gate_output_0_107(.a(output_1_107), .b(output_1_12), .y(output_0_107));
wire output_2_107, output_2_12, output_1_107;
mixer gate_output_1_107(.a(output_2_107), .b(output_2_12), .y(output_1_107));
wire output_3_107, output_3_12, output_2_107;
mixer gate_output_2_107(.a(output_3_107), .b(output_3_12), .y(output_2_107));
wire output_4_107, output_4_12, output_3_107;
mixer gate_output_3_107(.a(output_4_107), .b(output_4_12), .y(output_3_107));
wire output_5_107, output_5_12, output_4_107;
mixer gate_output_4_107(.a(output_5_107), .b(output_5_12), .y(output_4_107));
wire output_6_107, output_6_12, output_5_107;
mixer gate_output_5_107(.a(output_6_107), .b(output_6_12), .y(output_5_107));
wire output_7_107, output_7_12, output_6_107;
mixer gate_output_6_107(.a(output_7_107), .b(output_7_12), .y(output_6_107));
wire output_8_107, output_8_12, output_7_107;
mixer gate_output_7_107(.a(output_8_107), .b(output_8_12), .y(output_7_107));
wire output_9_107, output_9_12, output_8_107;
mixer gate_output_8_107(.a(output_9_107), .b(output_9_12), .y(output_8_107));
wire output_10_107, output_10_12, output_9_107;
mixer gate_output_9_107(.a(output_10_107), .b(output_10_12), .y(output_9_107));
wire output_11_107, output_11_12, output_10_107;
mixer gate_output_10_107(.a(output_11_107), .b(output_11_12), .y(output_10_107));
wire output_12_107, output_12_12, output_11_107;
mixer gate_output_11_107(.a(output_12_107), .b(output_12_12), .y(output_11_107));
wire output_13_107, output_13_12, output_12_107;
mixer gate_output_12_107(.a(output_13_107), .b(output_13_12), .y(output_12_107));
wire output_14_107, output_14_12, output_13_107;
mixer gate_output_13_107(.a(output_14_107), .b(output_14_12), .y(output_13_107));
wire output_15_107, output_15_12, output_14_107;
mixer gate_output_14_107(.a(output_15_107), .b(output_15_12), .y(output_14_107));
wire output_16_107, output_16_12, output_15_107;
mixer gate_output_15_107(.a(output_16_107), .b(output_16_12), .y(output_15_107));
wire output_1_108, output_1_13, output_0_108;
mixer gate_output_0_108(.a(output_1_108), .b(output_1_13), .y(output_0_108));
wire output_2_108, output_2_13, output_1_108;
mixer gate_output_1_108(.a(output_2_108), .b(output_2_13), .y(output_1_108));
wire output_3_108, output_3_13, output_2_108;
mixer gate_output_2_108(.a(output_3_108), .b(output_3_13), .y(output_2_108));
wire output_4_108, output_4_13, output_3_108;
mixer gate_output_3_108(.a(output_4_108), .b(output_4_13), .y(output_3_108));
wire output_5_108, output_5_13, output_4_108;
mixer gate_output_4_108(.a(output_5_108), .b(output_5_13), .y(output_4_108));
wire output_6_108, output_6_13, output_5_108;
mixer gate_output_5_108(.a(output_6_108), .b(output_6_13), .y(output_5_108));
wire output_7_108, output_7_13, output_6_108;
mixer gate_output_6_108(.a(output_7_108), .b(output_7_13), .y(output_6_108));
wire output_8_108, output_8_13, output_7_108;
mixer gate_output_7_108(.a(output_8_108), .b(output_8_13), .y(output_7_108));
wire output_9_108, output_9_13, output_8_108;
mixer gate_output_8_108(.a(output_9_108), .b(output_9_13), .y(output_8_108));
wire output_10_108, output_10_13, output_9_108;
mixer gate_output_9_108(.a(output_10_108), .b(output_10_13), .y(output_9_108));
wire output_11_108, output_11_13, output_10_108;
mixer gate_output_10_108(.a(output_11_108), .b(output_11_13), .y(output_10_108));
wire output_12_108, output_12_13, output_11_108;
mixer gate_output_11_108(.a(output_12_108), .b(output_12_13), .y(output_11_108));
wire output_13_108, output_13_13, output_12_108;
mixer gate_output_12_108(.a(output_13_108), .b(output_13_13), .y(output_12_108));
wire output_14_108, output_14_13, output_13_108;
mixer gate_output_13_108(.a(output_14_108), .b(output_14_13), .y(output_13_108));
wire output_15_108, output_15_13, output_14_108;
mixer gate_output_14_108(.a(output_15_108), .b(output_15_13), .y(output_14_108));
wire output_16_108, output_16_13, output_15_108;
mixer gate_output_15_108(.a(output_16_108), .b(output_16_13), .y(output_15_108));
wire output_1_109, output_1_14, output_0_109;
mixer gate_output_0_109(.a(output_1_109), .b(output_1_14), .y(output_0_109));
wire output_2_109, output_2_14, output_1_109;
mixer gate_output_1_109(.a(output_2_109), .b(output_2_14), .y(output_1_109));
wire output_3_109, output_3_14, output_2_109;
mixer gate_output_2_109(.a(output_3_109), .b(output_3_14), .y(output_2_109));
wire output_4_109, output_4_14, output_3_109;
mixer gate_output_3_109(.a(output_4_109), .b(output_4_14), .y(output_3_109));
wire output_5_109, output_5_14, output_4_109;
mixer gate_output_4_109(.a(output_5_109), .b(output_5_14), .y(output_4_109));
wire output_6_109, output_6_14, output_5_109;
mixer gate_output_5_109(.a(output_6_109), .b(output_6_14), .y(output_5_109));
wire output_7_109, output_7_14, output_6_109;
mixer gate_output_6_109(.a(output_7_109), .b(output_7_14), .y(output_6_109));
wire output_8_109, output_8_14, output_7_109;
mixer gate_output_7_109(.a(output_8_109), .b(output_8_14), .y(output_7_109));
wire output_9_109, output_9_14, output_8_109;
mixer gate_output_8_109(.a(output_9_109), .b(output_9_14), .y(output_8_109));
wire output_10_109, output_10_14, output_9_109;
mixer gate_output_9_109(.a(output_10_109), .b(output_10_14), .y(output_9_109));
wire output_11_109, output_11_14, output_10_109;
mixer gate_output_10_109(.a(output_11_109), .b(output_11_14), .y(output_10_109));
wire output_12_109, output_12_14, output_11_109;
mixer gate_output_11_109(.a(output_12_109), .b(output_12_14), .y(output_11_109));
wire output_13_109, output_13_14, output_12_109;
mixer gate_output_12_109(.a(output_13_109), .b(output_13_14), .y(output_12_109));
wire output_14_109, output_14_14, output_13_109;
mixer gate_output_13_109(.a(output_14_109), .b(output_14_14), .y(output_13_109));
wire output_15_109, output_15_14, output_14_109;
mixer gate_output_14_109(.a(output_15_109), .b(output_15_14), .y(output_14_109));
wire output_16_109, output_16_14, output_15_109;
mixer gate_output_15_109(.a(output_16_109), .b(output_16_14), .y(output_15_109));
wire output_1_110, output_1_15, output_0_110;
mixer gate_output_0_110(.a(output_1_110), .b(output_1_15), .y(output_0_110));
wire output_2_110, output_2_15, output_1_110;
mixer gate_output_1_110(.a(output_2_110), .b(output_2_15), .y(output_1_110));
wire output_3_110, output_3_15, output_2_110;
mixer gate_output_2_110(.a(output_3_110), .b(output_3_15), .y(output_2_110));
wire output_4_110, output_4_15, output_3_110;
mixer gate_output_3_110(.a(output_4_110), .b(output_4_15), .y(output_3_110));
wire output_5_110, output_5_15, output_4_110;
mixer gate_output_4_110(.a(output_5_110), .b(output_5_15), .y(output_4_110));
wire output_6_110, output_6_15, output_5_110;
mixer gate_output_5_110(.a(output_6_110), .b(output_6_15), .y(output_5_110));
wire output_7_110, output_7_15, output_6_110;
mixer gate_output_6_110(.a(output_7_110), .b(output_7_15), .y(output_6_110));
wire output_8_110, output_8_15, output_7_110;
mixer gate_output_7_110(.a(output_8_110), .b(output_8_15), .y(output_7_110));
wire output_9_110, output_9_15, output_8_110;
mixer gate_output_8_110(.a(output_9_110), .b(output_9_15), .y(output_8_110));
wire output_10_110, output_10_15, output_9_110;
mixer gate_output_9_110(.a(output_10_110), .b(output_10_15), .y(output_9_110));
wire output_11_110, output_11_15, output_10_110;
mixer gate_output_10_110(.a(output_11_110), .b(output_11_15), .y(output_10_110));
wire output_12_110, output_12_15, output_11_110;
mixer gate_output_11_110(.a(output_12_110), .b(output_12_15), .y(output_11_110));
wire output_13_110, output_13_15, output_12_110;
mixer gate_output_12_110(.a(output_13_110), .b(output_13_15), .y(output_12_110));
wire output_14_110, output_14_15, output_13_110;
mixer gate_output_13_110(.a(output_14_110), .b(output_14_15), .y(output_13_110));
wire output_15_110, output_15_15, output_14_110;
mixer gate_output_14_110(.a(output_15_110), .b(output_15_15), .y(output_14_110));
wire output_16_110, output_16_15, output_15_110;
mixer gate_output_15_110(.a(output_16_110), .b(output_16_15), .y(output_15_110));
wire output_1_111, output_1_0, output_0_111;
mixer gate_output_0_111(.a(output_1_111), .b(output_1_0), .y(output_0_111));
wire output_2_111, output_2_0, output_1_111;
mixer gate_output_1_111(.a(output_2_111), .b(output_2_0), .y(output_1_111));
wire output_3_111, output_3_0, output_2_111;
mixer gate_output_2_111(.a(output_3_111), .b(output_3_0), .y(output_2_111));
wire output_4_111, output_4_0, output_3_111;
mixer gate_output_3_111(.a(output_4_111), .b(output_4_0), .y(output_3_111));
wire output_5_111, output_5_0, output_4_111;
mixer gate_output_4_111(.a(output_5_111), .b(output_5_0), .y(output_4_111));
wire output_6_111, output_6_0, output_5_111;
mixer gate_output_5_111(.a(output_6_111), .b(output_6_0), .y(output_5_111));
wire output_7_111, output_7_0, output_6_111;
mixer gate_output_6_111(.a(output_7_111), .b(output_7_0), .y(output_6_111));
wire output_8_111, output_8_0, output_7_111;
mixer gate_output_7_111(.a(output_8_111), .b(output_8_0), .y(output_7_111));
wire output_9_111, output_9_0, output_8_111;
mixer gate_output_8_111(.a(output_9_111), .b(output_9_0), .y(output_8_111));
wire output_10_111, output_10_0, output_9_111;
mixer gate_output_9_111(.a(output_10_111), .b(output_10_0), .y(output_9_111));
wire output_11_111, output_11_0, output_10_111;
mixer gate_output_10_111(.a(output_11_111), .b(output_11_0), .y(output_10_111));
wire output_12_111, output_12_0, output_11_111;
mixer gate_output_11_111(.a(output_12_111), .b(output_12_0), .y(output_11_111));
wire output_13_111, output_13_0, output_12_111;
mixer gate_output_12_111(.a(output_13_111), .b(output_13_0), .y(output_12_111));
wire output_14_111, output_14_0, output_13_111;
mixer gate_output_13_111(.a(output_14_111), .b(output_14_0), .y(output_13_111));
wire output_15_111, output_15_0, output_14_111;
mixer gate_output_14_111(.a(output_15_111), .b(output_15_0), .y(output_14_111));
wire output_16_111, output_16_0, output_15_111;
mixer gate_output_15_111(.a(output_16_111), .b(output_16_0), .y(output_15_111));
wire output_1_112, output_1_1, output_0_112;
mixer gate_output_0_112(.a(output_1_112), .b(output_1_1), .y(output_0_112));
wire output_2_112, output_2_1, output_1_112;
mixer gate_output_1_112(.a(output_2_112), .b(output_2_1), .y(output_1_112));
wire output_3_112, output_3_1, output_2_112;
mixer gate_output_2_112(.a(output_3_112), .b(output_3_1), .y(output_2_112));
wire output_4_112, output_4_1, output_3_112;
mixer gate_output_3_112(.a(output_4_112), .b(output_4_1), .y(output_3_112));
wire output_5_112, output_5_1, output_4_112;
mixer gate_output_4_112(.a(output_5_112), .b(output_5_1), .y(output_4_112));
wire output_6_112, output_6_1, output_5_112;
mixer gate_output_5_112(.a(output_6_112), .b(output_6_1), .y(output_5_112));
wire output_7_112, output_7_1, output_6_112;
mixer gate_output_6_112(.a(output_7_112), .b(output_7_1), .y(output_6_112));
wire output_8_112, output_8_1, output_7_112;
mixer gate_output_7_112(.a(output_8_112), .b(output_8_1), .y(output_7_112));
wire output_9_112, output_9_1, output_8_112;
mixer gate_output_8_112(.a(output_9_112), .b(output_9_1), .y(output_8_112));
wire output_10_112, output_10_1, output_9_112;
mixer gate_output_9_112(.a(output_10_112), .b(output_10_1), .y(output_9_112));
wire output_11_112, output_11_1, output_10_112;
mixer gate_output_10_112(.a(output_11_112), .b(output_11_1), .y(output_10_112));
wire output_12_112, output_12_1, output_11_112;
mixer gate_output_11_112(.a(output_12_112), .b(output_12_1), .y(output_11_112));
wire output_13_112, output_13_1, output_12_112;
mixer gate_output_12_112(.a(output_13_112), .b(output_13_1), .y(output_12_112));
wire output_14_112, output_14_1, output_13_112;
mixer gate_output_13_112(.a(output_14_112), .b(output_14_1), .y(output_13_112));
wire output_15_112, output_15_1, output_14_112;
mixer gate_output_14_112(.a(output_15_112), .b(output_15_1), .y(output_14_112));
wire output_16_112, output_16_1, output_15_112;
mixer gate_output_15_112(.a(output_16_112), .b(output_16_1), .y(output_15_112));
wire output_1_113, output_1_2, output_0_113;
mixer gate_output_0_113(.a(output_1_113), .b(output_1_2), .y(output_0_113));
wire output_2_113, output_2_2, output_1_113;
mixer gate_output_1_113(.a(output_2_113), .b(output_2_2), .y(output_1_113));
wire output_3_113, output_3_2, output_2_113;
mixer gate_output_2_113(.a(output_3_113), .b(output_3_2), .y(output_2_113));
wire output_4_113, output_4_2, output_3_113;
mixer gate_output_3_113(.a(output_4_113), .b(output_4_2), .y(output_3_113));
wire output_5_113, output_5_2, output_4_113;
mixer gate_output_4_113(.a(output_5_113), .b(output_5_2), .y(output_4_113));
wire output_6_113, output_6_2, output_5_113;
mixer gate_output_5_113(.a(output_6_113), .b(output_6_2), .y(output_5_113));
wire output_7_113, output_7_2, output_6_113;
mixer gate_output_6_113(.a(output_7_113), .b(output_7_2), .y(output_6_113));
wire output_8_113, output_8_2, output_7_113;
mixer gate_output_7_113(.a(output_8_113), .b(output_8_2), .y(output_7_113));
wire output_9_113, output_9_2, output_8_113;
mixer gate_output_8_113(.a(output_9_113), .b(output_9_2), .y(output_8_113));
wire output_10_113, output_10_2, output_9_113;
mixer gate_output_9_113(.a(output_10_113), .b(output_10_2), .y(output_9_113));
wire output_11_113, output_11_2, output_10_113;
mixer gate_output_10_113(.a(output_11_113), .b(output_11_2), .y(output_10_113));
wire output_12_113, output_12_2, output_11_113;
mixer gate_output_11_113(.a(output_12_113), .b(output_12_2), .y(output_11_113));
wire output_13_113, output_13_2, output_12_113;
mixer gate_output_12_113(.a(output_13_113), .b(output_13_2), .y(output_12_113));
wire output_14_113, output_14_2, output_13_113;
mixer gate_output_13_113(.a(output_14_113), .b(output_14_2), .y(output_13_113));
wire output_15_113, output_15_2, output_14_113;
mixer gate_output_14_113(.a(output_15_113), .b(output_15_2), .y(output_14_113));
wire output_16_113, output_16_2, output_15_113;
mixer gate_output_15_113(.a(output_16_113), .b(output_16_2), .y(output_15_113));
wire output_1_114, output_1_3, output_0_114;
mixer gate_output_0_114(.a(output_1_114), .b(output_1_3), .y(output_0_114));
wire output_2_114, output_2_3, output_1_114;
mixer gate_output_1_114(.a(output_2_114), .b(output_2_3), .y(output_1_114));
wire output_3_114, output_3_3, output_2_114;
mixer gate_output_2_114(.a(output_3_114), .b(output_3_3), .y(output_2_114));
wire output_4_114, output_4_3, output_3_114;
mixer gate_output_3_114(.a(output_4_114), .b(output_4_3), .y(output_3_114));
wire output_5_114, output_5_3, output_4_114;
mixer gate_output_4_114(.a(output_5_114), .b(output_5_3), .y(output_4_114));
wire output_6_114, output_6_3, output_5_114;
mixer gate_output_5_114(.a(output_6_114), .b(output_6_3), .y(output_5_114));
wire output_7_114, output_7_3, output_6_114;
mixer gate_output_6_114(.a(output_7_114), .b(output_7_3), .y(output_6_114));
wire output_8_114, output_8_3, output_7_114;
mixer gate_output_7_114(.a(output_8_114), .b(output_8_3), .y(output_7_114));
wire output_9_114, output_9_3, output_8_114;
mixer gate_output_8_114(.a(output_9_114), .b(output_9_3), .y(output_8_114));
wire output_10_114, output_10_3, output_9_114;
mixer gate_output_9_114(.a(output_10_114), .b(output_10_3), .y(output_9_114));
wire output_11_114, output_11_3, output_10_114;
mixer gate_output_10_114(.a(output_11_114), .b(output_11_3), .y(output_10_114));
wire output_12_114, output_12_3, output_11_114;
mixer gate_output_11_114(.a(output_12_114), .b(output_12_3), .y(output_11_114));
wire output_13_114, output_13_3, output_12_114;
mixer gate_output_12_114(.a(output_13_114), .b(output_13_3), .y(output_12_114));
wire output_14_114, output_14_3, output_13_114;
mixer gate_output_13_114(.a(output_14_114), .b(output_14_3), .y(output_13_114));
wire output_15_114, output_15_3, output_14_114;
mixer gate_output_14_114(.a(output_15_114), .b(output_15_3), .y(output_14_114));
wire output_16_114, output_16_3, output_15_114;
mixer gate_output_15_114(.a(output_16_114), .b(output_16_3), .y(output_15_114));
wire output_1_115, output_1_4, output_0_115;
mixer gate_output_0_115(.a(output_1_115), .b(output_1_4), .y(output_0_115));
wire output_2_115, output_2_4, output_1_115;
mixer gate_output_1_115(.a(output_2_115), .b(output_2_4), .y(output_1_115));
wire output_3_115, output_3_4, output_2_115;
mixer gate_output_2_115(.a(output_3_115), .b(output_3_4), .y(output_2_115));
wire output_4_115, output_4_4, output_3_115;
mixer gate_output_3_115(.a(output_4_115), .b(output_4_4), .y(output_3_115));
wire output_5_115, output_5_4, output_4_115;
mixer gate_output_4_115(.a(output_5_115), .b(output_5_4), .y(output_4_115));
wire output_6_115, output_6_4, output_5_115;
mixer gate_output_5_115(.a(output_6_115), .b(output_6_4), .y(output_5_115));
wire output_7_115, output_7_4, output_6_115;
mixer gate_output_6_115(.a(output_7_115), .b(output_7_4), .y(output_6_115));
wire output_8_115, output_8_4, output_7_115;
mixer gate_output_7_115(.a(output_8_115), .b(output_8_4), .y(output_7_115));
wire output_9_115, output_9_4, output_8_115;
mixer gate_output_8_115(.a(output_9_115), .b(output_9_4), .y(output_8_115));
wire output_10_115, output_10_4, output_9_115;
mixer gate_output_9_115(.a(output_10_115), .b(output_10_4), .y(output_9_115));
wire output_11_115, output_11_4, output_10_115;
mixer gate_output_10_115(.a(output_11_115), .b(output_11_4), .y(output_10_115));
wire output_12_115, output_12_4, output_11_115;
mixer gate_output_11_115(.a(output_12_115), .b(output_12_4), .y(output_11_115));
wire output_13_115, output_13_4, output_12_115;
mixer gate_output_12_115(.a(output_13_115), .b(output_13_4), .y(output_12_115));
wire output_14_115, output_14_4, output_13_115;
mixer gate_output_13_115(.a(output_14_115), .b(output_14_4), .y(output_13_115));
wire output_15_115, output_15_4, output_14_115;
mixer gate_output_14_115(.a(output_15_115), .b(output_15_4), .y(output_14_115));
wire output_16_115, output_16_4, output_15_115;
mixer gate_output_15_115(.a(output_16_115), .b(output_16_4), .y(output_15_115));
wire output_1_116, output_1_5, output_0_116;
mixer gate_output_0_116(.a(output_1_116), .b(output_1_5), .y(output_0_116));
wire output_2_116, output_2_5, output_1_116;
mixer gate_output_1_116(.a(output_2_116), .b(output_2_5), .y(output_1_116));
wire output_3_116, output_3_5, output_2_116;
mixer gate_output_2_116(.a(output_3_116), .b(output_3_5), .y(output_2_116));
wire output_4_116, output_4_5, output_3_116;
mixer gate_output_3_116(.a(output_4_116), .b(output_4_5), .y(output_3_116));
wire output_5_116, output_5_5, output_4_116;
mixer gate_output_4_116(.a(output_5_116), .b(output_5_5), .y(output_4_116));
wire output_6_116, output_6_5, output_5_116;
mixer gate_output_5_116(.a(output_6_116), .b(output_6_5), .y(output_5_116));
wire output_7_116, output_7_5, output_6_116;
mixer gate_output_6_116(.a(output_7_116), .b(output_7_5), .y(output_6_116));
wire output_8_116, output_8_5, output_7_116;
mixer gate_output_7_116(.a(output_8_116), .b(output_8_5), .y(output_7_116));
wire output_9_116, output_9_5, output_8_116;
mixer gate_output_8_116(.a(output_9_116), .b(output_9_5), .y(output_8_116));
wire output_10_116, output_10_5, output_9_116;
mixer gate_output_9_116(.a(output_10_116), .b(output_10_5), .y(output_9_116));
wire output_11_116, output_11_5, output_10_116;
mixer gate_output_10_116(.a(output_11_116), .b(output_11_5), .y(output_10_116));
wire output_12_116, output_12_5, output_11_116;
mixer gate_output_11_116(.a(output_12_116), .b(output_12_5), .y(output_11_116));
wire output_13_116, output_13_5, output_12_116;
mixer gate_output_12_116(.a(output_13_116), .b(output_13_5), .y(output_12_116));
wire output_14_116, output_14_5, output_13_116;
mixer gate_output_13_116(.a(output_14_116), .b(output_14_5), .y(output_13_116));
wire output_15_116, output_15_5, output_14_116;
mixer gate_output_14_116(.a(output_15_116), .b(output_15_5), .y(output_14_116));
wire output_16_116, output_16_5, output_15_116;
mixer gate_output_15_116(.a(output_16_116), .b(output_16_5), .y(output_15_116));
wire output_1_117, output_1_6, output_0_117;
mixer gate_output_0_117(.a(output_1_117), .b(output_1_6), .y(output_0_117));
wire output_2_117, output_2_6, output_1_117;
mixer gate_output_1_117(.a(output_2_117), .b(output_2_6), .y(output_1_117));
wire output_3_117, output_3_6, output_2_117;
mixer gate_output_2_117(.a(output_3_117), .b(output_3_6), .y(output_2_117));
wire output_4_117, output_4_6, output_3_117;
mixer gate_output_3_117(.a(output_4_117), .b(output_4_6), .y(output_3_117));
wire output_5_117, output_5_6, output_4_117;
mixer gate_output_4_117(.a(output_5_117), .b(output_5_6), .y(output_4_117));
wire output_6_117, output_6_6, output_5_117;
mixer gate_output_5_117(.a(output_6_117), .b(output_6_6), .y(output_5_117));
wire output_7_117, output_7_6, output_6_117;
mixer gate_output_6_117(.a(output_7_117), .b(output_7_6), .y(output_6_117));
wire output_8_117, output_8_6, output_7_117;
mixer gate_output_7_117(.a(output_8_117), .b(output_8_6), .y(output_7_117));
wire output_9_117, output_9_6, output_8_117;
mixer gate_output_8_117(.a(output_9_117), .b(output_9_6), .y(output_8_117));
wire output_10_117, output_10_6, output_9_117;
mixer gate_output_9_117(.a(output_10_117), .b(output_10_6), .y(output_9_117));
wire output_11_117, output_11_6, output_10_117;
mixer gate_output_10_117(.a(output_11_117), .b(output_11_6), .y(output_10_117));
wire output_12_117, output_12_6, output_11_117;
mixer gate_output_11_117(.a(output_12_117), .b(output_12_6), .y(output_11_117));
wire output_13_117, output_13_6, output_12_117;
mixer gate_output_12_117(.a(output_13_117), .b(output_13_6), .y(output_12_117));
wire output_14_117, output_14_6, output_13_117;
mixer gate_output_13_117(.a(output_14_117), .b(output_14_6), .y(output_13_117));
wire output_15_117, output_15_6, output_14_117;
mixer gate_output_14_117(.a(output_15_117), .b(output_15_6), .y(output_14_117));
wire output_16_117, output_16_6, output_15_117;
mixer gate_output_15_117(.a(output_16_117), .b(output_16_6), .y(output_15_117));
wire output_1_118, output_1_7, output_0_118;
mixer gate_output_0_118(.a(output_1_118), .b(output_1_7), .y(output_0_118));
wire output_2_118, output_2_7, output_1_118;
mixer gate_output_1_118(.a(output_2_118), .b(output_2_7), .y(output_1_118));
wire output_3_118, output_3_7, output_2_118;
mixer gate_output_2_118(.a(output_3_118), .b(output_3_7), .y(output_2_118));
wire output_4_118, output_4_7, output_3_118;
mixer gate_output_3_118(.a(output_4_118), .b(output_4_7), .y(output_3_118));
wire output_5_118, output_5_7, output_4_118;
mixer gate_output_4_118(.a(output_5_118), .b(output_5_7), .y(output_4_118));
wire output_6_118, output_6_7, output_5_118;
mixer gate_output_5_118(.a(output_6_118), .b(output_6_7), .y(output_5_118));
wire output_7_118, output_7_7, output_6_118;
mixer gate_output_6_118(.a(output_7_118), .b(output_7_7), .y(output_6_118));
wire output_8_118, output_8_7, output_7_118;
mixer gate_output_7_118(.a(output_8_118), .b(output_8_7), .y(output_7_118));
wire output_9_118, output_9_7, output_8_118;
mixer gate_output_8_118(.a(output_9_118), .b(output_9_7), .y(output_8_118));
wire output_10_118, output_10_7, output_9_118;
mixer gate_output_9_118(.a(output_10_118), .b(output_10_7), .y(output_9_118));
wire output_11_118, output_11_7, output_10_118;
mixer gate_output_10_118(.a(output_11_118), .b(output_11_7), .y(output_10_118));
wire output_12_118, output_12_7, output_11_118;
mixer gate_output_11_118(.a(output_12_118), .b(output_12_7), .y(output_11_118));
wire output_13_118, output_13_7, output_12_118;
mixer gate_output_12_118(.a(output_13_118), .b(output_13_7), .y(output_12_118));
wire output_14_118, output_14_7, output_13_118;
mixer gate_output_13_118(.a(output_14_118), .b(output_14_7), .y(output_13_118));
wire output_15_118, output_15_7, output_14_118;
mixer gate_output_14_118(.a(output_15_118), .b(output_15_7), .y(output_14_118));
wire output_16_118, output_16_7, output_15_118;
mixer gate_output_15_118(.a(output_16_118), .b(output_16_7), .y(output_15_118));
wire output_1_119, output_1_8, output_0_119;
mixer gate_output_0_119(.a(output_1_119), .b(output_1_8), .y(output_0_119));
wire output_2_119, output_2_8, output_1_119;
mixer gate_output_1_119(.a(output_2_119), .b(output_2_8), .y(output_1_119));
wire output_3_119, output_3_8, output_2_119;
mixer gate_output_2_119(.a(output_3_119), .b(output_3_8), .y(output_2_119));
wire output_4_119, output_4_8, output_3_119;
mixer gate_output_3_119(.a(output_4_119), .b(output_4_8), .y(output_3_119));
wire output_5_119, output_5_8, output_4_119;
mixer gate_output_4_119(.a(output_5_119), .b(output_5_8), .y(output_4_119));
wire output_6_119, output_6_8, output_5_119;
mixer gate_output_5_119(.a(output_6_119), .b(output_6_8), .y(output_5_119));
wire output_7_119, output_7_8, output_6_119;
mixer gate_output_6_119(.a(output_7_119), .b(output_7_8), .y(output_6_119));
wire output_8_119, output_8_8, output_7_119;
mixer gate_output_7_119(.a(output_8_119), .b(output_8_8), .y(output_7_119));
wire output_9_119, output_9_8, output_8_119;
mixer gate_output_8_119(.a(output_9_119), .b(output_9_8), .y(output_8_119));
wire output_10_119, output_10_8, output_9_119;
mixer gate_output_9_119(.a(output_10_119), .b(output_10_8), .y(output_9_119));
wire output_11_119, output_11_8, output_10_119;
mixer gate_output_10_119(.a(output_11_119), .b(output_11_8), .y(output_10_119));
wire output_12_119, output_12_8, output_11_119;
mixer gate_output_11_119(.a(output_12_119), .b(output_12_8), .y(output_11_119));
wire output_13_119, output_13_8, output_12_119;
mixer gate_output_12_119(.a(output_13_119), .b(output_13_8), .y(output_12_119));
wire output_14_119, output_14_8, output_13_119;
mixer gate_output_13_119(.a(output_14_119), .b(output_14_8), .y(output_13_119));
wire output_15_119, output_15_8, output_14_119;
mixer gate_output_14_119(.a(output_15_119), .b(output_15_8), .y(output_14_119));
wire output_16_119, output_16_8, output_15_119;
mixer gate_output_15_119(.a(output_16_119), .b(output_16_8), .y(output_15_119));
wire output_1_120, output_1_9, output_0_120;
mixer gate_output_0_120(.a(output_1_120), .b(output_1_9), .y(output_0_120));
wire output_2_120, output_2_9, output_1_120;
mixer gate_output_1_120(.a(output_2_120), .b(output_2_9), .y(output_1_120));
wire output_3_120, output_3_9, output_2_120;
mixer gate_output_2_120(.a(output_3_120), .b(output_3_9), .y(output_2_120));
wire output_4_120, output_4_9, output_3_120;
mixer gate_output_3_120(.a(output_4_120), .b(output_4_9), .y(output_3_120));
wire output_5_120, output_5_9, output_4_120;
mixer gate_output_4_120(.a(output_5_120), .b(output_5_9), .y(output_4_120));
wire output_6_120, output_6_9, output_5_120;
mixer gate_output_5_120(.a(output_6_120), .b(output_6_9), .y(output_5_120));
wire output_7_120, output_7_9, output_6_120;
mixer gate_output_6_120(.a(output_7_120), .b(output_7_9), .y(output_6_120));
wire output_8_120, output_8_9, output_7_120;
mixer gate_output_7_120(.a(output_8_120), .b(output_8_9), .y(output_7_120));
wire output_9_120, output_9_9, output_8_120;
mixer gate_output_8_120(.a(output_9_120), .b(output_9_9), .y(output_8_120));
wire output_10_120, output_10_9, output_9_120;
mixer gate_output_9_120(.a(output_10_120), .b(output_10_9), .y(output_9_120));
wire output_11_120, output_11_9, output_10_120;
mixer gate_output_10_120(.a(output_11_120), .b(output_11_9), .y(output_10_120));
wire output_12_120, output_12_9, output_11_120;
mixer gate_output_11_120(.a(output_12_120), .b(output_12_9), .y(output_11_120));
wire output_13_120, output_13_9, output_12_120;
mixer gate_output_12_120(.a(output_13_120), .b(output_13_9), .y(output_12_120));
wire output_14_120, output_14_9, output_13_120;
mixer gate_output_13_120(.a(output_14_120), .b(output_14_9), .y(output_13_120));
wire output_15_120, output_15_9, output_14_120;
mixer gate_output_14_120(.a(output_15_120), .b(output_15_9), .y(output_14_120));
wire output_16_120, output_16_9, output_15_120;
mixer gate_output_15_120(.a(output_16_120), .b(output_16_9), .y(output_15_120));
wire output_1_121, output_1_10, output_0_121;
mixer gate_output_0_121(.a(output_1_121), .b(output_1_10), .y(output_0_121));
wire output_2_121, output_2_10, output_1_121;
mixer gate_output_1_121(.a(output_2_121), .b(output_2_10), .y(output_1_121));
wire output_3_121, output_3_10, output_2_121;
mixer gate_output_2_121(.a(output_3_121), .b(output_3_10), .y(output_2_121));
wire output_4_121, output_4_10, output_3_121;
mixer gate_output_3_121(.a(output_4_121), .b(output_4_10), .y(output_3_121));
wire output_5_121, output_5_10, output_4_121;
mixer gate_output_4_121(.a(output_5_121), .b(output_5_10), .y(output_4_121));
wire output_6_121, output_6_10, output_5_121;
mixer gate_output_5_121(.a(output_6_121), .b(output_6_10), .y(output_5_121));
wire output_7_121, output_7_10, output_6_121;
mixer gate_output_6_121(.a(output_7_121), .b(output_7_10), .y(output_6_121));
wire output_8_121, output_8_10, output_7_121;
mixer gate_output_7_121(.a(output_8_121), .b(output_8_10), .y(output_7_121));
wire output_9_121, output_9_10, output_8_121;
mixer gate_output_8_121(.a(output_9_121), .b(output_9_10), .y(output_8_121));
wire output_10_121, output_10_10, output_9_121;
mixer gate_output_9_121(.a(output_10_121), .b(output_10_10), .y(output_9_121));
wire output_11_121, output_11_10, output_10_121;
mixer gate_output_10_121(.a(output_11_121), .b(output_11_10), .y(output_10_121));
wire output_12_121, output_12_10, output_11_121;
mixer gate_output_11_121(.a(output_12_121), .b(output_12_10), .y(output_11_121));
wire output_13_121, output_13_10, output_12_121;
mixer gate_output_12_121(.a(output_13_121), .b(output_13_10), .y(output_12_121));
wire output_14_121, output_14_10, output_13_121;
mixer gate_output_13_121(.a(output_14_121), .b(output_14_10), .y(output_13_121));
wire output_15_121, output_15_10, output_14_121;
mixer gate_output_14_121(.a(output_15_121), .b(output_15_10), .y(output_14_121));
wire output_16_121, output_16_10, output_15_121;
mixer gate_output_15_121(.a(output_16_121), .b(output_16_10), .y(output_15_121));
wire output_1_122, output_1_11, output_0_122;
mixer gate_output_0_122(.a(output_1_122), .b(output_1_11), .y(output_0_122));
wire output_2_122, output_2_11, output_1_122;
mixer gate_output_1_122(.a(output_2_122), .b(output_2_11), .y(output_1_122));
wire output_3_122, output_3_11, output_2_122;
mixer gate_output_2_122(.a(output_3_122), .b(output_3_11), .y(output_2_122));
wire output_4_122, output_4_11, output_3_122;
mixer gate_output_3_122(.a(output_4_122), .b(output_4_11), .y(output_3_122));
wire output_5_122, output_5_11, output_4_122;
mixer gate_output_4_122(.a(output_5_122), .b(output_5_11), .y(output_4_122));
wire output_6_122, output_6_11, output_5_122;
mixer gate_output_5_122(.a(output_6_122), .b(output_6_11), .y(output_5_122));
wire output_7_122, output_7_11, output_6_122;
mixer gate_output_6_122(.a(output_7_122), .b(output_7_11), .y(output_6_122));
wire output_8_122, output_8_11, output_7_122;
mixer gate_output_7_122(.a(output_8_122), .b(output_8_11), .y(output_7_122));
wire output_9_122, output_9_11, output_8_122;
mixer gate_output_8_122(.a(output_9_122), .b(output_9_11), .y(output_8_122));
wire output_10_122, output_10_11, output_9_122;
mixer gate_output_9_122(.a(output_10_122), .b(output_10_11), .y(output_9_122));
wire output_11_122, output_11_11, output_10_122;
mixer gate_output_10_122(.a(output_11_122), .b(output_11_11), .y(output_10_122));
wire output_12_122, output_12_11, output_11_122;
mixer gate_output_11_122(.a(output_12_122), .b(output_12_11), .y(output_11_122));
wire output_13_122, output_13_11, output_12_122;
mixer gate_output_12_122(.a(output_13_122), .b(output_13_11), .y(output_12_122));
wire output_14_122, output_14_11, output_13_122;
mixer gate_output_13_122(.a(output_14_122), .b(output_14_11), .y(output_13_122));
wire output_15_122, output_15_11, output_14_122;
mixer gate_output_14_122(.a(output_15_122), .b(output_15_11), .y(output_14_122));
wire output_16_122, output_16_11, output_15_122;
mixer gate_output_15_122(.a(output_16_122), .b(output_16_11), .y(output_15_122));
wire output_1_123, output_1_12, output_0_123;
mixer gate_output_0_123(.a(output_1_123), .b(output_1_12), .y(output_0_123));
wire output_2_123, output_2_12, output_1_123;
mixer gate_output_1_123(.a(output_2_123), .b(output_2_12), .y(output_1_123));
wire output_3_123, output_3_12, output_2_123;
mixer gate_output_2_123(.a(output_3_123), .b(output_3_12), .y(output_2_123));
wire output_4_123, output_4_12, output_3_123;
mixer gate_output_3_123(.a(output_4_123), .b(output_4_12), .y(output_3_123));
wire output_5_123, output_5_12, output_4_123;
mixer gate_output_4_123(.a(output_5_123), .b(output_5_12), .y(output_4_123));
wire output_6_123, output_6_12, output_5_123;
mixer gate_output_5_123(.a(output_6_123), .b(output_6_12), .y(output_5_123));
wire output_7_123, output_7_12, output_6_123;
mixer gate_output_6_123(.a(output_7_123), .b(output_7_12), .y(output_6_123));
wire output_8_123, output_8_12, output_7_123;
mixer gate_output_7_123(.a(output_8_123), .b(output_8_12), .y(output_7_123));
wire output_9_123, output_9_12, output_8_123;
mixer gate_output_8_123(.a(output_9_123), .b(output_9_12), .y(output_8_123));
wire output_10_123, output_10_12, output_9_123;
mixer gate_output_9_123(.a(output_10_123), .b(output_10_12), .y(output_9_123));
wire output_11_123, output_11_12, output_10_123;
mixer gate_output_10_123(.a(output_11_123), .b(output_11_12), .y(output_10_123));
wire output_12_123, output_12_12, output_11_123;
mixer gate_output_11_123(.a(output_12_123), .b(output_12_12), .y(output_11_123));
wire output_13_123, output_13_12, output_12_123;
mixer gate_output_12_123(.a(output_13_123), .b(output_13_12), .y(output_12_123));
wire output_14_123, output_14_12, output_13_123;
mixer gate_output_13_123(.a(output_14_123), .b(output_14_12), .y(output_13_123));
wire output_15_123, output_15_12, output_14_123;
mixer gate_output_14_123(.a(output_15_123), .b(output_15_12), .y(output_14_123));
wire output_16_123, output_16_12, output_15_123;
mixer gate_output_15_123(.a(output_16_123), .b(output_16_12), .y(output_15_123));
wire output_1_124, output_1_13, output_0_124;
mixer gate_output_0_124(.a(output_1_124), .b(output_1_13), .y(output_0_124));
wire output_2_124, output_2_13, output_1_124;
mixer gate_output_1_124(.a(output_2_124), .b(output_2_13), .y(output_1_124));
wire output_3_124, output_3_13, output_2_124;
mixer gate_output_2_124(.a(output_3_124), .b(output_3_13), .y(output_2_124));
wire output_4_124, output_4_13, output_3_124;
mixer gate_output_3_124(.a(output_4_124), .b(output_4_13), .y(output_3_124));
wire output_5_124, output_5_13, output_4_124;
mixer gate_output_4_124(.a(output_5_124), .b(output_5_13), .y(output_4_124));
wire output_6_124, output_6_13, output_5_124;
mixer gate_output_5_124(.a(output_6_124), .b(output_6_13), .y(output_5_124));
wire output_7_124, output_7_13, output_6_124;
mixer gate_output_6_124(.a(output_7_124), .b(output_7_13), .y(output_6_124));
wire output_8_124, output_8_13, output_7_124;
mixer gate_output_7_124(.a(output_8_124), .b(output_8_13), .y(output_7_124));
wire output_9_124, output_9_13, output_8_124;
mixer gate_output_8_124(.a(output_9_124), .b(output_9_13), .y(output_8_124));
wire output_10_124, output_10_13, output_9_124;
mixer gate_output_9_124(.a(output_10_124), .b(output_10_13), .y(output_9_124));
wire output_11_124, output_11_13, output_10_124;
mixer gate_output_10_124(.a(output_11_124), .b(output_11_13), .y(output_10_124));
wire output_12_124, output_12_13, output_11_124;
mixer gate_output_11_124(.a(output_12_124), .b(output_12_13), .y(output_11_124));
wire output_13_124, output_13_13, output_12_124;
mixer gate_output_12_124(.a(output_13_124), .b(output_13_13), .y(output_12_124));
wire output_14_124, output_14_13, output_13_124;
mixer gate_output_13_124(.a(output_14_124), .b(output_14_13), .y(output_13_124));
wire output_15_124, output_15_13, output_14_124;
mixer gate_output_14_124(.a(output_15_124), .b(output_15_13), .y(output_14_124));
wire output_16_124, output_16_13, output_15_124;
mixer gate_output_15_124(.a(output_16_124), .b(output_16_13), .y(output_15_124));
wire output_1_125, output_1_14, output_0_125;
mixer gate_output_0_125(.a(output_1_125), .b(output_1_14), .y(output_0_125));
wire output_2_125, output_2_14, output_1_125;
mixer gate_output_1_125(.a(output_2_125), .b(output_2_14), .y(output_1_125));
wire output_3_125, output_3_14, output_2_125;
mixer gate_output_2_125(.a(output_3_125), .b(output_3_14), .y(output_2_125));
wire output_4_125, output_4_14, output_3_125;
mixer gate_output_3_125(.a(output_4_125), .b(output_4_14), .y(output_3_125));
wire output_5_125, output_5_14, output_4_125;
mixer gate_output_4_125(.a(output_5_125), .b(output_5_14), .y(output_4_125));
wire output_6_125, output_6_14, output_5_125;
mixer gate_output_5_125(.a(output_6_125), .b(output_6_14), .y(output_5_125));
wire output_7_125, output_7_14, output_6_125;
mixer gate_output_6_125(.a(output_7_125), .b(output_7_14), .y(output_6_125));
wire output_8_125, output_8_14, output_7_125;
mixer gate_output_7_125(.a(output_8_125), .b(output_8_14), .y(output_7_125));
wire output_9_125, output_9_14, output_8_125;
mixer gate_output_8_125(.a(output_9_125), .b(output_9_14), .y(output_8_125));
wire output_10_125, output_10_14, output_9_125;
mixer gate_output_9_125(.a(output_10_125), .b(output_10_14), .y(output_9_125));
wire output_11_125, output_11_14, output_10_125;
mixer gate_output_10_125(.a(output_11_125), .b(output_11_14), .y(output_10_125));
wire output_12_125, output_12_14, output_11_125;
mixer gate_output_11_125(.a(output_12_125), .b(output_12_14), .y(output_11_125));
wire output_13_125, output_13_14, output_12_125;
mixer gate_output_12_125(.a(output_13_125), .b(output_13_14), .y(output_12_125));
wire output_14_125, output_14_14, output_13_125;
mixer gate_output_13_125(.a(output_14_125), .b(output_14_14), .y(output_13_125));
wire output_15_125, output_15_14, output_14_125;
mixer gate_output_14_125(.a(output_15_125), .b(output_15_14), .y(output_14_125));
wire output_16_125, output_16_14, output_15_125;
mixer gate_output_15_125(.a(output_16_125), .b(output_16_14), .y(output_15_125));
wire output_1_126, output_1_15, output_0_126;
mixer gate_output_0_126(.a(output_1_126), .b(output_1_15), .y(output_0_126));
wire output_2_126, output_2_15, output_1_126;
mixer gate_output_1_126(.a(output_2_126), .b(output_2_15), .y(output_1_126));
wire output_3_126, output_3_15, output_2_126;
mixer gate_output_2_126(.a(output_3_126), .b(output_3_15), .y(output_2_126));
wire output_4_126, output_4_15, output_3_126;
mixer gate_output_3_126(.a(output_4_126), .b(output_4_15), .y(output_3_126));
wire output_5_126, output_5_15, output_4_126;
mixer gate_output_4_126(.a(output_5_126), .b(output_5_15), .y(output_4_126));
wire output_6_126, output_6_15, output_5_126;
mixer gate_output_5_126(.a(output_6_126), .b(output_6_15), .y(output_5_126));
wire output_7_126, output_7_15, output_6_126;
mixer gate_output_6_126(.a(output_7_126), .b(output_7_15), .y(output_6_126));
wire output_8_126, output_8_15, output_7_126;
mixer gate_output_7_126(.a(output_8_126), .b(output_8_15), .y(output_7_126));
wire output_9_126, output_9_15, output_8_126;
mixer gate_output_8_126(.a(output_9_126), .b(output_9_15), .y(output_8_126));
wire output_10_126, output_10_15, output_9_126;
mixer gate_output_9_126(.a(output_10_126), .b(output_10_15), .y(output_9_126));
wire output_11_126, output_11_15, output_10_126;
mixer gate_output_10_126(.a(output_11_126), .b(output_11_15), .y(output_10_126));
wire output_12_126, output_12_15, output_11_126;
mixer gate_output_11_126(.a(output_12_126), .b(output_12_15), .y(output_11_126));
wire output_13_126, output_13_15, output_12_126;
mixer gate_output_12_126(.a(output_13_126), .b(output_13_15), .y(output_12_126));
wire output_14_126, output_14_15, output_13_126;
mixer gate_output_13_126(.a(output_14_126), .b(output_14_15), .y(output_13_126));
wire output_15_126, output_15_15, output_14_126;
mixer gate_output_14_126(.a(output_15_126), .b(output_15_15), .y(output_14_126));
wire output_16_126, output_16_15, output_15_126;
mixer gate_output_15_126(.a(output_16_126), .b(output_16_15), .y(output_15_126));
wire output_1_127, output_1_0, output_0_127;
mixer gate_output_0_127(.a(output_1_127), .b(output_1_0), .y(output_0_127));
wire output_2_127, output_2_0, output_1_127;
mixer gate_output_1_127(.a(output_2_127), .b(output_2_0), .y(output_1_127));
wire output_3_127, output_3_0, output_2_127;
mixer gate_output_2_127(.a(output_3_127), .b(output_3_0), .y(output_2_127));
wire output_4_127, output_4_0, output_3_127;
mixer gate_output_3_127(.a(output_4_127), .b(output_4_0), .y(output_3_127));
wire output_5_127, output_5_0, output_4_127;
mixer gate_output_4_127(.a(output_5_127), .b(output_5_0), .y(output_4_127));
wire output_6_127, output_6_0, output_5_127;
mixer gate_output_5_127(.a(output_6_127), .b(output_6_0), .y(output_5_127));
wire output_7_127, output_7_0, output_6_127;
mixer gate_output_6_127(.a(output_7_127), .b(output_7_0), .y(output_6_127));
wire output_8_127, output_8_0, output_7_127;
mixer gate_output_7_127(.a(output_8_127), .b(output_8_0), .y(output_7_127));
wire output_9_127, output_9_0, output_8_127;
mixer gate_output_8_127(.a(output_9_127), .b(output_9_0), .y(output_8_127));
wire output_10_127, output_10_0, output_9_127;
mixer gate_output_9_127(.a(output_10_127), .b(output_10_0), .y(output_9_127));
wire output_11_127, output_11_0, output_10_127;
mixer gate_output_10_127(.a(output_11_127), .b(output_11_0), .y(output_10_127));
wire output_12_127, output_12_0, output_11_127;
mixer gate_output_11_127(.a(output_12_127), .b(output_12_0), .y(output_11_127));
wire output_13_127, output_13_0, output_12_127;
mixer gate_output_12_127(.a(output_13_127), .b(output_13_0), .y(output_12_127));
wire output_14_127, output_14_0, output_13_127;
mixer gate_output_13_127(.a(output_14_127), .b(output_14_0), .y(output_13_127));
wire output_15_127, output_15_0, output_14_127;
mixer gate_output_14_127(.a(output_15_127), .b(output_15_0), .y(output_14_127));
wire output_16_127, output_16_0, output_15_127;
mixer gate_output_15_127(.a(output_16_127), .b(output_16_0), .y(output_15_127));
wire output_1_128, output_1_1, output_0_128;
mixer gate_output_0_128(.a(output_1_128), .b(output_1_1), .y(output_0_128));
wire output_2_128, output_2_1, output_1_128;
mixer gate_output_1_128(.a(output_2_128), .b(output_2_1), .y(output_1_128));
wire output_3_128, output_3_1, output_2_128;
mixer gate_output_2_128(.a(output_3_128), .b(output_3_1), .y(output_2_128));
wire output_4_128, output_4_1, output_3_128;
mixer gate_output_3_128(.a(output_4_128), .b(output_4_1), .y(output_3_128));
wire output_5_128, output_5_1, output_4_128;
mixer gate_output_4_128(.a(output_5_128), .b(output_5_1), .y(output_4_128));
wire output_6_128, output_6_1, output_5_128;
mixer gate_output_5_128(.a(output_6_128), .b(output_6_1), .y(output_5_128));
wire output_7_128, output_7_1, output_6_128;
mixer gate_output_6_128(.a(output_7_128), .b(output_7_1), .y(output_6_128));
wire output_8_128, output_8_1, output_7_128;
mixer gate_output_7_128(.a(output_8_128), .b(output_8_1), .y(output_7_128));
wire output_9_128, output_9_1, output_8_128;
mixer gate_output_8_128(.a(output_9_128), .b(output_9_1), .y(output_8_128));
wire output_10_128, output_10_1, output_9_128;
mixer gate_output_9_128(.a(output_10_128), .b(output_10_1), .y(output_9_128));
wire output_11_128, output_11_1, output_10_128;
mixer gate_output_10_128(.a(output_11_128), .b(output_11_1), .y(output_10_128));
wire output_12_128, output_12_1, output_11_128;
mixer gate_output_11_128(.a(output_12_128), .b(output_12_1), .y(output_11_128));
wire output_13_128, output_13_1, output_12_128;
mixer gate_output_12_128(.a(output_13_128), .b(output_13_1), .y(output_12_128));
wire output_14_128, output_14_1, output_13_128;
mixer gate_output_13_128(.a(output_14_128), .b(output_14_1), .y(output_13_128));
wire output_15_128, output_15_1, output_14_128;
mixer gate_output_14_128(.a(output_15_128), .b(output_15_1), .y(output_14_128));
wire output_16_128, output_16_1, output_15_128;
mixer gate_output_15_128(.a(output_16_128), .b(output_16_1), .y(output_15_128));
wire output_1_129, output_1_2, output_0_129;
mixer gate_output_0_129(.a(output_1_129), .b(output_1_2), .y(output_0_129));
wire output_2_129, output_2_2, output_1_129;
mixer gate_output_1_129(.a(output_2_129), .b(output_2_2), .y(output_1_129));
wire output_3_129, output_3_2, output_2_129;
mixer gate_output_2_129(.a(output_3_129), .b(output_3_2), .y(output_2_129));
wire output_4_129, output_4_2, output_3_129;
mixer gate_output_3_129(.a(output_4_129), .b(output_4_2), .y(output_3_129));
wire output_5_129, output_5_2, output_4_129;
mixer gate_output_4_129(.a(output_5_129), .b(output_5_2), .y(output_4_129));
wire output_6_129, output_6_2, output_5_129;
mixer gate_output_5_129(.a(output_6_129), .b(output_6_2), .y(output_5_129));
wire output_7_129, output_7_2, output_6_129;
mixer gate_output_6_129(.a(output_7_129), .b(output_7_2), .y(output_6_129));
wire output_8_129, output_8_2, output_7_129;
mixer gate_output_7_129(.a(output_8_129), .b(output_8_2), .y(output_7_129));
wire output_9_129, output_9_2, output_8_129;
mixer gate_output_8_129(.a(output_9_129), .b(output_9_2), .y(output_8_129));
wire output_10_129, output_10_2, output_9_129;
mixer gate_output_9_129(.a(output_10_129), .b(output_10_2), .y(output_9_129));
wire output_11_129, output_11_2, output_10_129;
mixer gate_output_10_129(.a(output_11_129), .b(output_11_2), .y(output_10_129));
wire output_12_129, output_12_2, output_11_129;
mixer gate_output_11_129(.a(output_12_129), .b(output_12_2), .y(output_11_129));
wire output_13_129, output_13_2, output_12_129;
mixer gate_output_12_129(.a(output_13_129), .b(output_13_2), .y(output_12_129));
wire output_14_129, output_14_2, output_13_129;
mixer gate_output_13_129(.a(output_14_129), .b(output_14_2), .y(output_13_129));
wire output_15_129, output_15_2, output_14_129;
mixer gate_output_14_129(.a(output_15_129), .b(output_15_2), .y(output_14_129));
wire output_16_129, output_16_2, output_15_129;
mixer gate_output_15_129(.a(output_16_129), .b(output_16_2), .y(output_15_129));
wire output_1_130, output_1_3, output_0_130;
mixer gate_output_0_130(.a(output_1_130), .b(output_1_3), .y(output_0_130));
wire output_2_130, output_2_3, output_1_130;
mixer gate_output_1_130(.a(output_2_130), .b(output_2_3), .y(output_1_130));
wire output_3_130, output_3_3, output_2_130;
mixer gate_output_2_130(.a(output_3_130), .b(output_3_3), .y(output_2_130));
wire output_4_130, output_4_3, output_3_130;
mixer gate_output_3_130(.a(output_4_130), .b(output_4_3), .y(output_3_130));
wire output_5_130, output_5_3, output_4_130;
mixer gate_output_4_130(.a(output_5_130), .b(output_5_3), .y(output_4_130));
wire output_6_130, output_6_3, output_5_130;
mixer gate_output_5_130(.a(output_6_130), .b(output_6_3), .y(output_5_130));
wire output_7_130, output_7_3, output_6_130;
mixer gate_output_6_130(.a(output_7_130), .b(output_7_3), .y(output_6_130));
wire output_8_130, output_8_3, output_7_130;
mixer gate_output_7_130(.a(output_8_130), .b(output_8_3), .y(output_7_130));
wire output_9_130, output_9_3, output_8_130;
mixer gate_output_8_130(.a(output_9_130), .b(output_9_3), .y(output_8_130));
wire output_10_130, output_10_3, output_9_130;
mixer gate_output_9_130(.a(output_10_130), .b(output_10_3), .y(output_9_130));
wire output_11_130, output_11_3, output_10_130;
mixer gate_output_10_130(.a(output_11_130), .b(output_11_3), .y(output_10_130));
wire output_12_130, output_12_3, output_11_130;
mixer gate_output_11_130(.a(output_12_130), .b(output_12_3), .y(output_11_130));
wire output_13_130, output_13_3, output_12_130;
mixer gate_output_12_130(.a(output_13_130), .b(output_13_3), .y(output_12_130));
wire output_14_130, output_14_3, output_13_130;
mixer gate_output_13_130(.a(output_14_130), .b(output_14_3), .y(output_13_130));
wire output_15_130, output_15_3, output_14_130;
mixer gate_output_14_130(.a(output_15_130), .b(output_15_3), .y(output_14_130));
wire output_16_130, output_16_3, output_15_130;
mixer gate_output_15_130(.a(output_16_130), .b(output_16_3), .y(output_15_130));
wire output_1_131, output_1_4, output_0_131;
mixer gate_output_0_131(.a(output_1_131), .b(output_1_4), .y(output_0_131));
wire output_2_131, output_2_4, output_1_131;
mixer gate_output_1_131(.a(output_2_131), .b(output_2_4), .y(output_1_131));
wire output_3_131, output_3_4, output_2_131;
mixer gate_output_2_131(.a(output_3_131), .b(output_3_4), .y(output_2_131));
wire output_4_131, output_4_4, output_3_131;
mixer gate_output_3_131(.a(output_4_131), .b(output_4_4), .y(output_3_131));
wire output_5_131, output_5_4, output_4_131;
mixer gate_output_4_131(.a(output_5_131), .b(output_5_4), .y(output_4_131));
wire output_6_131, output_6_4, output_5_131;
mixer gate_output_5_131(.a(output_6_131), .b(output_6_4), .y(output_5_131));
wire output_7_131, output_7_4, output_6_131;
mixer gate_output_6_131(.a(output_7_131), .b(output_7_4), .y(output_6_131));
wire output_8_131, output_8_4, output_7_131;
mixer gate_output_7_131(.a(output_8_131), .b(output_8_4), .y(output_7_131));
wire output_9_131, output_9_4, output_8_131;
mixer gate_output_8_131(.a(output_9_131), .b(output_9_4), .y(output_8_131));
wire output_10_131, output_10_4, output_9_131;
mixer gate_output_9_131(.a(output_10_131), .b(output_10_4), .y(output_9_131));
wire output_11_131, output_11_4, output_10_131;
mixer gate_output_10_131(.a(output_11_131), .b(output_11_4), .y(output_10_131));
wire output_12_131, output_12_4, output_11_131;
mixer gate_output_11_131(.a(output_12_131), .b(output_12_4), .y(output_11_131));
wire output_13_131, output_13_4, output_12_131;
mixer gate_output_12_131(.a(output_13_131), .b(output_13_4), .y(output_12_131));
wire output_14_131, output_14_4, output_13_131;
mixer gate_output_13_131(.a(output_14_131), .b(output_14_4), .y(output_13_131));
wire output_15_131, output_15_4, output_14_131;
mixer gate_output_14_131(.a(output_15_131), .b(output_15_4), .y(output_14_131));
wire output_16_131, output_16_4, output_15_131;
mixer gate_output_15_131(.a(output_16_131), .b(output_16_4), .y(output_15_131));
wire output_1_132, output_1_5, output_0_132;
mixer gate_output_0_132(.a(output_1_132), .b(output_1_5), .y(output_0_132));
wire output_2_132, output_2_5, output_1_132;
mixer gate_output_1_132(.a(output_2_132), .b(output_2_5), .y(output_1_132));
wire output_3_132, output_3_5, output_2_132;
mixer gate_output_2_132(.a(output_3_132), .b(output_3_5), .y(output_2_132));
wire output_4_132, output_4_5, output_3_132;
mixer gate_output_3_132(.a(output_4_132), .b(output_4_5), .y(output_3_132));
wire output_5_132, output_5_5, output_4_132;
mixer gate_output_4_132(.a(output_5_132), .b(output_5_5), .y(output_4_132));
wire output_6_132, output_6_5, output_5_132;
mixer gate_output_5_132(.a(output_6_132), .b(output_6_5), .y(output_5_132));
wire output_7_132, output_7_5, output_6_132;
mixer gate_output_6_132(.a(output_7_132), .b(output_7_5), .y(output_6_132));
wire output_8_132, output_8_5, output_7_132;
mixer gate_output_7_132(.a(output_8_132), .b(output_8_5), .y(output_7_132));
wire output_9_132, output_9_5, output_8_132;
mixer gate_output_8_132(.a(output_9_132), .b(output_9_5), .y(output_8_132));
wire output_10_132, output_10_5, output_9_132;
mixer gate_output_9_132(.a(output_10_132), .b(output_10_5), .y(output_9_132));
wire output_11_132, output_11_5, output_10_132;
mixer gate_output_10_132(.a(output_11_132), .b(output_11_5), .y(output_10_132));
wire output_12_132, output_12_5, output_11_132;
mixer gate_output_11_132(.a(output_12_132), .b(output_12_5), .y(output_11_132));
wire output_13_132, output_13_5, output_12_132;
mixer gate_output_12_132(.a(output_13_132), .b(output_13_5), .y(output_12_132));
wire output_14_132, output_14_5, output_13_132;
mixer gate_output_13_132(.a(output_14_132), .b(output_14_5), .y(output_13_132));
wire output_15_132, output_15_5, output_14_132;
mixer gate_output_14_132(.a(output_15_132), .b(output_15_5), .y(output_14_132));
wire output_16_132, output_16_5, output_15_132;
mixer gate_output_15_132(.a(output_16_132), .b(output_16_5), .y(output_15_132));
wire output_1_133, output_1_6, output_0_133;
mixer gate_output_0_133(.a(output_1_133), .b(output_1_6), .y(output_0_133));
wire output_2_133, output_2_6, output_1_133;
mixer gate_output_1_133(.a(output_2_133), .b(output_2_6), .y(output_1_133));
wire output_3_133, output_3_6, output_2_133;
mixer gate_output_2_133(.a(output_3_133), .b(output_3_6), .y(output_2_133));
wire output_4_133, output_4_6, output_3_133;
mixer gate_output_3_133(.a(output_4_133), .b(output_4_6), .y(output_3_133));
wire output_5_133, output_5_6, output_4_133;
mixer gate_output_4_133(.a(output_5_133), .b(output_5_6), .y(output_4_133));
wire output_6_133, output_6_6, output_5_133;
mixer gate_output_5_133(.a(output_6_133), .b(output_6_6), .y(output_5_133));
wire output_7_133, output_7_6, output_6_133;
mixer gate_output_6_133(.a(output_7_133), .b(output_7_6), .y(output_6_133));
wire output_8_133, output_8_6, output_7_133;
mixer gate_output_7_133(.a(output_8_133), .b(output_8_6), .y(output_7_133));
wire output_9_133, output_9_6, output_8_133;
mixer gate_output_8_133(.a(output_9_133), .b(output_9_6), .y(output_8_133));
wire output_10_133, output_10_6, output_9_133;
mixer gate_output_9_133(.a(output_10_133), .b(output_10_6), .y(output_9_133));
wire output_11_133, output_11_6, output_10_133;
mixer gate_output_10_133(.a(output_11_133), .b(output_11_6), .y(output_10_133));
wire output_12_133, output_12_6, output_11_133;
mixer gate_output_11_133(.a(output_12_133), .b(output_12_6), .y(output_11_133));
wire output_13_133, output_13_6, output_12_133;
mixer gate_output_12_133(.a(output_13_133), .b(output_13_6), .y(output_12_133));
wire output_14_133, output_14_6, output_13_133;
mixer gate_output_13_133(.a(output_14_133), .b(output_14_6), .y(output_13_133));
wire output_15_133, output_15_6, output_14_133;
mixer gate_output_14_133(.a(output_15_133), .b(output_15_6), .y(output_14_133));
wire output_16_133, output_16_6, output_15_133;
mixer gate_output_15_133(.a(output_16_133), .b(output_16_6), .y(output_15_133));
wire output_1_134, output_1_7, output_0_134;
mixer gate_output_0_134(.a(output_1_134), .b(output_1_7), .y(output_0_134));
wire output_2_134, output_2_7, output_1_134;
mixer gate_output_1_134(.a(output_2_134), .b(output_2_7), .y(output_1_134));
wire output_3_134, output_3_7, output_2_134;
mixer gate_output_2_134(.a(output_3_134), .b(output_3_7), .y(output_2_134));
wire output_4_134, output_4_7, output_3_134;
mixer gate_output_3_134(.a(output_4_134), .b(output_4_7), .y(output_3_134));
wire output_5_134, output_5_7, output_4_134;
mixer gate_output_4_134(.a(output_5_134), .b(output_5_7), .y(output_4_134));
wire output_6_134, output_6_7, output_5_134;
mixer gate_output_5_134(.a(output_6_134), .b(output_6_7), .y(output_5_134));
wire output_7_134, output_7_7, output_6_134;
mixer gate_output_6_134(.a(output_7_134), .b(output_7_7), .y(output_6_134));
wire output_8_134, output_8_7, output_7_134;
mixer gate_output_7_134(.a(output_8_134), .b(output_8_7), .y(output_7_134));
wire output_9_134, output_9_7, output_8_134;
mixer gate_output_8_134(.a(output_9_134), .b(output_9_7), .y(output_8_134));
wire output_10_134, output_10_7, output_9_134;
mixer gate_output_9_134(.a(output_10_134), .b(output_10_7), .y(output_9_134));
wire output_11_134, output_11_7, output_10_134;
mixer gate_output_10_134(.a(output_11_134), .b(output_11_7), .y(output_10_134));
wire output_12_134, output_12_7, output_11_134;
mixer gate_output_11_134(.a(output_12_134), .b(output_12_7), .y(output_11_134));
wire output_13_134, output_13_7, output_12_134;
mixer gate_output_12_134(.a(output_13_134), .b(output_13_7), .y(output_12_134));
wire output_14_134, output_14_7, output_13_134;
mixer gate_output_13_134(.a(output_14_134), .b(output_14_7), .y(output_13_134));
wire output_15_134, output_15_7, output_14_134;
mixer gate_output_14_134(.a(output_15_134), .b(output_15_7), .y(output_14_134));
wire output_16_134, output_16_7, output_15_134;
mixer gate_output_15_134(.a(output_16_134), .b(output_16_7), .y(output_15_134));
wire output_1_135, output_1_8, output_0_135;
mixer gate_output_0_135(.a(output_1_135), .b(output_1_8), .y(output_0_135));
wire output_2_135, output_2_8, output_1_135;
mixer gate_output_1_135(.a(output_2_135), .b(output_2_8), .y(output_1_135));
wire output_3_135, output_3_8, output_2_135;
mixer gate_output_2_135(.a(output_3_135), .b(output_3_8), .y(output_2_135));
wire output_4_135, output_4_8, output_3_135;
mixer gate_output_3_135(.a(output_4_135), .b(output_4_8), .y(output_3_135));
wire output_5_135, output_5_8, output_4_135;
mixer gate_output_4_135(.a(output_5_135), .b(output_5_8), .y(output_4_135));
wire output_6_135, output_6_8, output_5_135;
mixer gate_output_5_135(.a(output_6_135), .b(output_6_8), .y(output_5_135));
wire output_7_135, output_7_8, output_6_135;
mixer gate_output_6_135(.a(output_7_135), .b(output_7_8), .y(output_6_135));
wire output_8_135, output_8_8, output_7_135;
mixer gate_output_7_135(.a(output_8_135), .b(output_8_8), .y(output_7_135));
wire output_9_135, output_9_8, output_8_135;
mixer gate_output_8_135(.a(output_9_135), .b(output_9_8), .y(output_8_135));
wire output_10_135, output_10_8, output_9_135;
mixer gate_output_9_135(.a(output_10_135), .b(output_10_8), .y(output_9_135));
wire output_11_135, output_11_8, output_10_135;
mixer gate_output_10_135(.a(output_11_135), .b(output_11_8), .y(output_10_135));
wire output_12_135, output_12_8, output_11_135;
mixer gate_output_11_135(.a(output_12_135), .b(output_12_8), .y(output_11_135));
wire output_13_135, output_13_8, output_12_135;
mixer gate_output_12_135(.a(output_13_135), .b(output_13_8), .y(output_12_135));
wire output_14_135, output_14_8, output_13_135;
mixer gate_output_13_135(.a(output_14_135), .b(output_14_8), .y(output_13_135));
wire output_15_135, output_15_8, output_14_135;
mixer gate_output_14_135(.a(output_15_135), .b(output_15_8), .y(output_14_135));
wire output_16_135, output_16_8, output_15_135;
mixer gate_output_15_135(.a(output_16_135), .b(output_16_8), .y(output_15_135));
wire output_1_136, output_1_9, output_0_136;
mixer gate_output_0_136(.a(output_1_136), .b(output_1_9), .y(output_0_136));
wire output_2_136, output_2_9, output_1_136;
mixer gate_output_1_136(.a(output_2_136), .b(output_2_9), .y(output_1_136));
wire output_3_136, output_3_9, output_2_136;
mixer gate_output_2_136(.a(output_3_136), .b(output_3_9), .y(output_2_136));
wire output_4_136, output_4_9, output_3_136;
mixer gate_output_3_136(.a(output_4_136), .b(output_4_9), .y(output_3_136));
wire output_5_136, output_5_9, output_4_136;
mixer gate_output_4_136(.a(output_5_136), .b(output_5_9), .y(output_4_136));
wire output_6_136, output_6_9, output_5_136;
mixer gate_output_5_136(.a(output_6_136), .b(output_6_9), .y(output_5_136));
wire output_7_136, output_7_9, output_6_136;
mixer gate_output_6_136(.a(output_7_136), .b(output_7_9), .y(output_6_136));
wire output_8_136, output_8_9, output_7_136;
mixer gate_output_7_136(.a(output_8_136), .b(output_8_9), .y(output_7_136));
wire output_9_136, output_9_9, output_8_136;
mixer gate_output_8_136(.a(output_9_136), .b(output_9_9), .y(output_8_136));
wire output_10_136, output_10_9, output_9_136;
mixer gate_output_9_136(.a(output_10_136), .b(output_10_9), .y(output_9_136));
wire output_11_136, output_11_9, output_10_136;
mixer gate_output_10_136(.a(output_11_136), .b(output_11_9), .y(output_10_136));
wire output_12_136, output_12_9, output_11_136;
mixer gate_output_11_136(.a(output_12_136), .b(output_12_9), .y(output_11_136));
wire output_13_136, output_13_9, output_12_136;
mixer gate_output_12_136(.a(output_13_136), .b(output_13_9), .y(output_12_136));
wire output_14_136, output_14_9, output_13_136;
mixer gate_output_13_136(.a(output_14_136), .b(output_14_9), .y(output_13_136));
wire output_15_136, output_15_9, output_14_136;
mixer gate_output_14_136(.a(output_15_136), .b(output_15_9), .y(output_14_136));
wire output_16_136, output_16_9, output_15_136;
mixer gate_output_15_136(.a(output_16_136), .b(output_16_9), .y(output_15_136));
wire output_1_137, output_1_10, output_0_137;
mixer gate_output_0_137(.a(output_1_137), .b(output_1_10), .y(output_0_137));
wire output_2_137, output_2_10, output_1_137;
mixer gate_output_1_137(.a(output_2_137), .b(output_2_10), .y(output_1_137));
wire output_3_137, output_3_10, output_2_137;
mixer gate_output_2_137(.a(output_3_137), .b(output_3_10), .y(output_2_137));
wire output_4_137, output_4_10, output_3_137;
mixer gate_output_3_137(.a(output_4_137), .b(output_4_10), .y(output_3_137));
wire output_5_137, output_5_10, output_4_137;
mixer gate_output_4_137(.a(output_5_137), .b(output_5_10), .y(output_4_137));
wire output_6_137, output_6_10, output_5_137;
mixer gate_output_5_137(.a(output_6_137), .b(output_6_10), .y(output_5_137));
wire output_7_137, output_7_10, output_6_137;
mixer gate_output_6_137(.a(output_7_137), .b(output_7_10), .y(output_6_137));
wire output_8_137, output_8_10, output_7_137;
mixer gate_output_7_137(.a(output_8_137), .b(output_8_10), .y(output_7_137));
wire output_9_137, output_9_10, output_8_137;
mixer gate_output_8_137(.a(output_9_137), .b(output_9_10), .y(output_8_137));
wire output_10_137, output_10_10, output_9_137;
mixer gate_output_9_137(.a(output_10_137), .b(output_10_10), .y(output_9_137));
wire output_11_137, output_11_10, output_10_137;
mixer gate_output_10_137(.a(output_11_137), .b(output_11_10), .y(output_10_137));
wire output_12_137, output_12_10, output_11_137;
mixer gate_output_11_137(.a(output_12_137), .b(output_12_10), .y(output_11_137));
wire output_13_137, output_13_10, output_12_137;
mixer gate_output_12_137(.a(output_13_137), .b(output_13_10), .y(output_12_137));
wire output_14_137, output_14_10, output_13_137;
mixer gate_output_13_137(.a(output_14_137), .b(output_14_10), .y(output_13_137));
wire output_15_137, output_15_10, output_14_137;
mixer gate_output_14_137(.a(output_15_137), .b(output_15_10), .y(output_14_137));
wire output_16_137, output_16_10, output_15_137;
mixer gate_output_15_137(.a(output_16_137), .b(output_16_10), .y(output_15_137));
wire output_1_138, output_1_11, output_0_138;
mixer gate_output_0_138(.a(output_1_138), .b(output_1_11), .y(output_0_138));
wire output_2_138, output_2_11, output_1_138;
mixer gate_output_1_138(.a(output_2_138), .b(output_2_11), .y(output_1_138));
wire output_3_138, output_3_11, output_2_138;
mixer gate_output_2_138(.a(output_3_138), .b(output_3_11), .y(output_2_138));
wire output_4_138, output_4_11, output_3_138;
mixer gate_output_3_138(.a(output_4_138), .b(output_4_11), .y(output_3_138));
wire output_5_138, output_5_11, output_4_138;
mixer gate_output_4_138(.a(output_5_138), .b(output_5_11), .y(output_4_138));
wire output_6_138, output_6_11, output_5_138;
mixer gate_output_5_138(.a(output_6_138), .b(output_6_11), .y(output_5_138));
wire output_7_138, output_7_11, output_6_138;
mixer gate_output_6_138(.a(output_7_138), .b(output_7_11), .y(output_6_138));
wire output_8_138, output_8_11, output_7_138;
mixer gate_output_7_138(.a(output_8_138), .b(output_8_11), .y(output_7_138));
wire output_9_138, output_9_11, output_8_138;
mixer gate_output_8_138(.a(output_9_138), .b(output_9_11), .y(output_8_138));
wire output_10_138, output_10_11, output_9_138;
mixer gate_output_9_138(.a(output_10_138), .b(output_10_11), .y(output_9_138));
wire output_11_138, output_11_11, output_10_138;
mixer gate_output_10_138(.a(output_11_138), .b(output_11_11), .y(output_10_138));
wire output_12_138, output_12_11, output_11_138;
mixer gate_output_11_138(.a(output_12_138), .b(output_12_11), .y(output_11_138));
wire output_13_138, output_13_11, output_12_138;
mixer gate_output_12_138(.a(output_13_138), .b(output_13_11), .y(output_12_138));
wire output_14_138, output_14_11, output_13_138;
mixer gate_output_13_138(.a(output_14_138), .b(output_14_11), .y(output_13_138));
wire output_15_138, output_15_11, output_14_138;
mixer gate_output_14_138(.a(output_15_138), .b(output_15_11), .y(output_14_138));
wire output_16_138, output_16_11, output_15_138;
mixer gate_output_15_138(.a(output_16_138), .b(output_16_11), .y(output_15_138));
wire output_1_139, output_1_12, output_0_139;
mixer gate_output_0_139(.a(output_1_139), .b(output_1_12), .y(output_0_139));
wire output_2_139, output_2_12, output_1_139;
mixer gate_output_1_139(.a(output_2_139), .b(output_2_12), .y(output_1_139));
wire output_3_139, output_3_12, output_2_139;
mixer gate_output_2_139(.a(output_3_139), .b(output_3_12), .y(output_2_139));
wire output_4_139, output_4_12, output_3_139;
mixer gate_output_3_139(.a(output_4_139), .b(output_4_12), .y(output_3_139));
wire output_5_139, output_5_12, output_4_139;
mixer gate_output_4_139(.a(output_5_139), .b(output_5_12), .y(output_4_139));
wire output_6_139, output_6_12, output_5_139;
mixer gate_output_5_139(.a(output_6_139), .b(output_6_12), .y(output_5_139));
wire output_7_139, output_7_12, output_6_139;
mixer gate_output_6_139(.a(output_7_139), .b(output_7_12), .y(output_6_139));
wire output_8_139, output_8_12, output_7_139;
mixer gate_output_7_139(.a(output_8_139), .b(output_8_12), .y(output_7_139));
wire output_9_139, output_9_12, output_8_139;
mixer gate_output_8_139(.a(output_9_139), .b(output_9_12), .y(output_8_139));
wire output_10_139, output_10_12, output_9_139;
mixer gate_output_9_139(.a(output_10_139), .b(output_10_12), .y(output_9_139));
wire output_11_139, output_11_12, output_10_139;
mixer gate_output_10_139(.a(output_11_139), .b(output_11_12), .y(output_10_139));
wire output_12_139, output_12_12, output_11_139;
mixer gate_output_11_139(.a(output_12_139), .b(output_12_12), .y(output_11_139));
wire output_13_139, output_13_12, output_12_139;
mixer gate_output_12_139(.a(output_13_139), .b(output_13_12), .y(output_12_139));
wire output_14_139, output_14_12, output_13_139;
mixer gate_output_13_139(.a(output_14_139), .b(output_14_12), .y(output_13_139));
wire output_15_139, output_15_12, output_14_139;
mixer gate_output_14_139(.a(output_15_139), .b(output_15_12), .y(output_14_139));
wire output_16_139, output_16_12, output_15_139;
mixer gate_output_15_139(.a(output_16_139), .b(output_16_12), .y(output_15_139));
wire output_1_140, output_1_13, output_0_140;
mixer gate_output_0_140(.a(output_1_140), .b(output_1_13), .y(output_0_140));
wire output_2_140, output_2_13, output_1_140;
mixer gate_output_1_140(.a(output_2_140), .b(output_2_13), .y(output_1_140));
wire output_3_140, output_3_13, output_2_140;
mixer gate_output_2_140(.a(output_3_140), .b(output_3_13), .y(output_2_140));
wire output_4_140, output_4_13, output_3_140;
mixer gate_output_3_140(.a(output_4_140), .b(output_4_13), .y(output_3_140));
wire output_5_140, output_5_13, output_4_140;
mixer gate_output_4_140(.a(output_5_140), .b(output_5_13), .y(output_4_140));
wire output_6_140, output_6_13, output_5_140;
mixer gate_output_5_140(.a(output_6_140), .b(output_6_13), .y(output_5_140));
wire output_7_140, output_7_13, output_6_140;
mixer gate_output_6_140(.a(output_7_140), .b(output_7_13), .y(output_6_140));
wire output_8_140, output_8_13, output_7_140;
mixer gate_output_7_140(.a(output_8_140), .b(output_8_13), .y(output_7_140));
wire output_9_140, output_9_13, output_8_140;
mixer gate_output_8_140(.a(output_9_140), .b(output_9_13), .y(output_8_140));
wire output_10_140, output_10_13, output_9_140;
mixer gate_output_9_140(.a(output_10_140), .b(output_10_13), .y(output_9_140));
wire output_11_140, output_11_13, output_10_140;
mixer gate_output_10_140(.a(output_11_140), .b(output_11_13), .y(output_10_140));
wire output_12_140, output_12_13, output_11_140;
mixer gate_output_11_140(.a(output_12_140), .b(output_12_13), .y(output_11_140));
wire output_13_140, output_13_13, output_12_140;
mixer gate_output_12_140(.a(output_13_140), .b(output_13_13), .y(output_12_140));
wire output_14_140, output_14_13, output_13_140;
mixer gate_output_13_140(.a(output_14_140), .b(output_14_13), .y(output_13_140));
wire output_15_140, output_15_13, output_14_140;
mixer gate_output_14_140(.a(output_15_140), .b(output_15_13), .y(output_14_140));
wire output_16_140, output_16_13, output_15_140;
mixer gate_output_15_140(.a(output_16_140), .b(output_16_13), .y(output_15_140));
wire output_1_141, output_1_14, output_0_141;
mixer gate_output_0_141(.a(output_1_141), .b(output_1_14), .y(output_0_141));
wire output_2_141, output_2_14, output_1_141;
mixer gate_output_1_141(.a(output_2_141), .b(output_2_14), .y(output_1_141));
wire output_3_141, output_3_14, output_2_141;
mixer gate_output_2_141(.a(output_3_141), .b(output_3_14), .y(output_2_141));
wire output_4_141, output_4_14, output_3_141;
mixer gate_output_3_141(.a(output_4_141), .b(output_4_14), .y(output_3_141));
wire output_5_141, output_5_14, output_4_141;
mixer gate_output_4_141(.a(output_5_141), .b(output_5_14), .y(output_4_141));
wire output_6_141, output_6_14, output_5_141;
mixer gate_output_5_141(.a(output_6_141), .b(output_6_14), .y(output_5_141));
wire output_7_141, output_7_14, output_6_141;
mixer gate_output_6_141(.a(output_7_141), .b(output_7_14), .y(output_6_141));
wire output_8_141, output_8_14, output_7_141;
mixer gate_output_7_141(.a(output_8_141), .b(output_8_14), .y(output_7_141));
wire output_9_141, output_9_14, output_8_141;
mixer gate_output_8_141(.a(output_9_141), .b(output_9_14), .y(output_8_141));
wire output_10_141, output_10_14, output_9_141;
mixer gate_output_9_141(.a(output_10_141), .b(output_10_14), .y(output_9_141));
wire output_11_141, output_11_14, output_10_141;
mixer gate_output_10_141(.a(output_11_141), .b(output_11_14), .y(output_10_141));
wire output_12_141, output_12_14, output_11_141;
mixer gate_output_11_141(.a(output_12_141), .b(output_12_14), .y(output_11_141));
wire output_13_141, output_13_14, output_12_141;
mixer gate_output_12_141(.a(output_13_141), .b(output_13_14), .y(output_12_141));
wire output_14_141, output_14_14, output_13_141;
mixer gate_output_13_141(.a(output_14_141), .b(output_14_14), .y(output_13_141));
wire output_15_141, output_15_14, output_14_141;
mixer gate_output_14_141(.a(output_15_141), .b(output_15_14), .y(output_14_141));
wire output_16_141, output_16_14, output_15_141;
mixer gate_output_15_141(.a(output_16_141), .b(output_16_14), .y(output_15_141));
wire output_1_142, output_1_15, output_0_142;
mixer gate_output_0_142(.a(output_1_142), .b(output_1_15), .y(output_0_142));
wire output_2_142, output_2_15, output_1_142;
mixer gate_output_1_142(.a(output_2_142), .b(output_2_15), .y(output_1_142));
wire output_3_142, output_3_15, output_2_142;
mixer gate_output_2_142(.a(output_3_142), .b(output_3_15), .y(output_2_142));
wire output_4_142, output_4_15, output_3_142;
mixer gate_output_3_142(.a(output_4_142), .b(output_4_15), .y(output_3_142));
wire output_5_142, output_5_15, output_4_142;
mixer gate_output_4_142(.a(output_5_142), .b(output_5_15), .y(output_4_142));
wire output_6_142, output_6_15, output_5_142;
mixer gate_output_5_142(.a(output_6_142), .b(output_6_15), .y(output_5_142));
wire output_7_142, output_7_15, output_6_142;
mixer gate_output_6_142(.a(output_7_142), .b(output_7_15), .y(output_6_142));
wire output_8_142, output_8_15, output_7_142;
mixer gate_output_7_142(.a(output_8_142), .b(output_8_15), .y(output_7_142));
wire output_9_142, output_9_15, output_8_142;
mixer gate_output_8_142(.a(output_9_142), .b(output_9_15), .y(output_8_142));
wire output_10_142, output_10_15, output_9_142;
mixer gate_output_9_142(.a(output_10_142), .b(output_10_15), .y(output_9_142));
wire output_11_142, output_11_15, output_10_142;
mixer gate_output_10_142(.a(output_11_142), .b(output_11_15), .y(output_10_142));
wire output_12_142, output_12_15, output_11_142;
mixer gate_output_11_142(.a(output_12_142), .b(output_12_15), .y(output_11_142));
wire output_13_142, output_13_15, output_12_142;
mixer gate_output_12_142(.a(output_13_142), .b(output_13_15), .y(output_12_142));
wire output_14_142, output_14_15, output_13_142;
mixer gate_output_13_142(.a(output_14_142), .b(output_14_15), .y(output_13_142));
wire output_15_142, output_15_15, output_14_142;
mixer gate_output_14_142(.a(output_15_142), .b(output_15_15), .y(output_14_142));
wire output_16_142, output_16_15, output_15_142;
mixer gate_output_15_142(.a(output_16_142), .b(output_16_15), .y(output_15_142));
wire output_1_143, output_1_0, output_0_143;
mixer gate_output_0_143(.a(output_1_143), .b(output_1_0), .y(output_0_143));
wire output_2_143, output_2_0, output_1_143;
mixer gate_output_1_143(.a(output_2_143), .b(output_2_0), .y(output_1_143));
wire output_3_143, output_3_0, output_2_143;
mixer gate_output_2_143(.a(output_3_143), .b(output_3_0), .y(output_2_143));
wire output_4_143, output_4_0, output_3_143;
mixer gate_output_3_143(.a(output_4_143), .b(output_4_0), .y(output_3_143));
wire output_5_143, output_5_0, output_4_143;
mixer gate_output_4_143(.a(output_5_143), .b(output_5_0), .y(output_4_143));
wire output_6_143, output_6_0, output_5_143;
mixer gate_output_5_143(.a(output_6_143), .b(output_6_0), .y(output_5_143));
wire output_7_143, output_7_0, output_6_143;
mixer gate_output_6_143(.a(output_7_143), .b(output_7_0), .y(output_6_143));
wire output_8_143, output_8_0, output_7_143;
mixer gate_output_7_143(.a(output_8_143), .b(output_8_0), .y(output_7_143));
wire output_9_143, output_9_0, output_8_143;
mixer gate_output_8_143(.a(output_9_143), .b(output_9_0), .y(output_8_143));
wire output_10_143, output_10_0, output_9_143;
mixer gate_output_9_143(.a(output_10_143), .b(output_10_0), .y(output_9_143));
wire output_11_143, output_11_0, output_10_143;
mixer gate_output_10_143(.a(output_11_143), .b(output_11_0), .y(output_10_143));
wire output_12_143, output_12_0, output_11_143;
mixer gate_output_11_143(.a(output_12_143), .b(output_12_0), .y(output_11_143));
wire output_13_143, output_13_0, output_12_143;
mixer gate_output_12_143(.a(output_13_143), .b(output_13_0), .y(output_12_143));
wire output_14_143, output_14_0, output_13_143;
mixer gate_output_13_143(.a(output_14_143), .b(output_14_0), .y(output_13_143));
wire output_15_143, output_15_0, output_14_143;
mixer gate_output_14_143(.a(output_15_143), .b(output_15_0), .y(output_14_143));
wire output_16_143, output_16_0, output_15_143;
mixer gate_output_15_143(.a(output_16_143), .b(output_16_0), .y(output_15_143));
wire output_1_144, output_1_1, output_0_144;
mixer gate_output_0_144(.a(output_1_144), .b(output_1_1), .y(output_0_144));
wire output_2_144, output_2_1, output_1_144;
mixer gate_output_1_144(.a(output_2_144), .b(output_2_1), .y(output_1_144));
wire output_3_144, output_3_1, output_2_144;
mixer gate_output_2_144(.a(output_3_144), .b(output_3_1), .y(output_2_144));
wire output_4_144, output_4_1, output_3_144;
mixer gate_output_3_144(.a(output_4_144), .b(output_4_1), .y(output_3_144));
wire output_5_144, output_5_1, output_4_144;
mixer gate_output_4_144(.a(output_5_144), .b(output_5_1), .y(output_4_144));
wire output_6_144, output_6_1, output_5_144;
mixer gate_output_5_144(.a(output_6_144), .b(output_6_1), .y(output_5_144));
wire output_7_144, output_7_1, output_6_144;
mixer gate_output_6_144(.a(output_7_144), .b(output_7_1), .y(output_6_144));
wire output_8_144, output_8_1, output_7_144;
mixer gate_output_7_144(.a(output_8_144), .b(output_8_1), .y(output_7_144));
wire output_9_144, output_9_1, output_8_144;
mixer gate_output_8_144(.a(output_9_144), .b(output_9_1), .y(output_8_144));
wire output_10_144, output_10_1, output_9_144;
mixer gate_output_9_144(.a(output_10_144), .b(output_10_1), .y(output_9_144));
wire output_11_144, output_11_1, output_10_144;
mixer gate_output_10_144(.a(output_11_144), .b(output_11_1), .y(output_10_144));
wire output_12_144, output_12_1, output_11_144;
mixer gate_output_11_144(.a(output_12_144), .b(output_12_1), .y(output_11_144));
wire output_13_144, output_13_1, output_12_144;
mixer gate_output_12_144(.a(output_13_144), .b(output_13_1), .y(output_12_144));
wire output_14_144, output_14_1, output_13_144;
mixer gate_output_13_144(.a(output_14_144), .b(output_14_1), .y(output_13_144));
wire output_15_144, output_15_1, output_14_144;
mixer gate_output_14_144(.a(output_15_144), .b(output_15_1), .y(output_14_144));
wire output_16_144, output_16_1, output_15_144;
mixer gate_output_15_144(.a(output_16_144), .b(output_16_1), .y(output_15_144));
wire output_1_145, output_1_2, output_0_145;
mixer gate_output_0_145(.a(output_1_145), .b(output_1_2), .y(output_0_145));
wire output_2_145, output_2_2, output_1_145;
mixer gate_output_1_145(.a(output_2_145), .b(output_2_2), .y(output_1_145));
wire output_3_145, output_3_2, output_2_145;
mixer gate_output_2_145(.a(output_3_145), .b(output_3_2), .y(output_2_145));
wire output_4_145, output_4_2, output_3_145;
mixer gate_output_3_145(.a(output_4_145), .b(output_4_2), .y(output_3_145));
wire output_5_145, output_5_2, output_4_145;
mixer gate_output_4_145(.a(output_5_145), .b(output_5_2), .y(output_4_145));
wire output_6_145, output_6_2, output_5_145;
mixer gate_output_5_145(.a(output_6_145), .b(output_6_2), .y(output_5_145));
wire output_7_145, output_7_2, output_6_145;
mixer gate_output_6_145(.a(output_7_145), .b(output_7_2), .y(output_6_145));
wire output_8_145, output_8_2, output_7_145;
mixer gate_output_7_145(.a(output_8_145), .b(output_8_2), .y(output_7_145));
wire output_9_145, output_9_2, output_8_145;
mixer gate_output_8_145(.a(output_9_145), .b(output_9_2), .y(output_8_145));
wire output_10_145, output_10_2, output_9_145;
mixer gate_output_9_145(.a(output_10_145), .b(output_10_2), .y(output_9_145));
wire output_11_145, output_11_2, output_10_145;
mixer gate_output_10_145(.a(output_11_145), .b(output_11_2), .y(output_10_145));
wire output_12_145, output_12_2, output_11_145;
mixer gate_output_11_145(.a(output_12_145), .b(output_12_2), .y(output_11_145));
wire output_13_145, output_13_2, output_12_145;
mixer gate_output_12_145(.a(output_13_145), .b(output_13_2), .y(output_12_145));
wire output_14_145, output_14_2, output_13_145;
mixer gate_output_13_145(.a(output_14_145), .b(output_14_2), .y(output_13_145));
wire output_15_145, output_15_2, output_14_145;
mixer gate_output_14_145(.a(output_15_145), .b(output_15_2), .y(output_14_145));
wire output_16_145, output_16_2, output_15_145;
mixer gate_output_15_145(.a(output_16_145), .b(output_16_2), .y(output_15_145));
wire output_1_146, output_1_3, output_0_146;
mixer gate_output_0_146(.a(output_1_146), .b(output_1_3), .y(output_0_146));
wire output_2_146, output_2_3, output_1_146;
mixer gate_output_1_146(.a(output_2_146), .b(output_2_3), .y(output_1_146));
wire output_3_146, output_3_3, output_2_146;
mixer gate_output_2_146(.a(output_3_146), .b(output_3_3), .y(output_2_146));
wire output_4_146, output_4_3, output_3_146;
mixer gate_output_3_146(.a(output_4_146), .b(output_4_3), .y(output_3_146));
wire output_5_146, output_5_3, output_4_146;
mixer gate_output_4_146(.a(output_5_146), .b(output_5_3), .y(output_4_146));
wire output_6_146, output_6_3, output_5_146;
mixer gate_output_5_146(.a(output_6_146), .b(output_6_3), .y(output_5_146));
wire output_7_146, output_7_3, output_6_146;
mixer gate_output_6_146(.a(output_7_146), .b(output_7_3), .y(output_6_146));
wire output_8_146, output_8_3, output_7_146;
mixer gate_output_7_146(.a(output_8_146), .b(output_8_3), .y(output_7_146));
wire output_9_146, output_9_3, output_8_146;
mixer gate_output_8_146(.a(output_9_146), .b(output_9_3), .y(output_8_146));
wire output_10_146, output_10_3, output_9_146;
mixer gate_output_9_146(.a(output_10_146), .b(output_10_3), .y(output_9_146));
wire output_11_146, output_11_3, output_10_146;
mixer gate_output_10_146(.a(output_11_146), .b(output_11_3), .y(output_10_146));
wire output_12_146, output_12_3, output_11_146;
mixer gate_output_11_146(.a(output_12_146), .b(output_12_3), .y(output_11_146));
wire output_13_146, output_13_3, output_12_146;
mixer gate_output_12_146(.a(output_13_146), .b(output_13_3), .y(output_12_146));
wire output_14_146, output_14_3, output_13_146;
mixer gate_output_13_146(.a(output_14_146), .b(output_14_3), .y(output_13_146));
wire output_15_146, output_15_3, output_14_146;
mixer gate_output_14_146(.a(output_15_146), .b(output_15_3), .y(output_14_146));
wire output_16_146, output_16_3, output_15_146;
mixer gate_output_15_146(.a(output_16_146), .b(output_16_3), .y(output_15_146));
wire output_1_147, output_1_4, output_0_147;
mixer gate_output_0_147(.a(output_1_147), .b(output_1_4), .y(output_0_147));
wire output_2_147, output_2_4, output_1_147;
mixer gate_output_1_147(.a(output_2_147), .b(output_2_4), .y(output_1_147));
wire output_3_147, output_3_4, output_2_147;
mixer gate_output_2_147(.a(output_3_147), .b(output_3_4), .y(output_2_147));
wire output_4_147, output_4_4, output_3_147;
mixer gate_output_3_147(.a(output_4_147), .b(output_4_4), .y(output_3_147));
wire output_5_147, output_5_4, output_4_147;
mixer gate_output_4_147(.a(output_5_147), .b(output_5_4), .y(output_4_147));
wire output_6_147, output_6_4, output_5_147;
mixer gate_output_5_147(.a(output_6_147), .b(output_6_4), .y(output_5_147));
wire output_7_147, output_7_4, output_6_147;
mixer gate_output_6_147(.a(output_7_147), .b(output_7_4), .y(output_6_147));
wire output_8_147, output_8_4, output_7_147;
mixer gate_output_7_147(.a(output_8_147), .b(output_8_4), .y(output_7_147));
wire output_9_147, output_9_4, output_8_147;
mixer gate_output_8_147(.a(output_9_147), .b(output_9_4), .y(output_8_147));
wire output_10_147, output_10_4, output_9_147;
mixer gate_output_9_147(.a(output_10_147), .b(output_10_4), .y(output_9_147));
wire output_11_147, output_11_4, output_10_147;
mixer gate_output_10_147(.a(output_11_147), .b(output_11_4), .y(output_10_147));
wire output_12_147, output_12_4, output_11_147;
mixer gate_output_11_147(.a(output_12_147), .b(output_12_4), .y(output_11_147));
wire output_13_147, output_13_4, output_12_147;
mixer gate_output_12_147(.a(output_13_147), .b(output_13_4), .y(output_12_147));
wire output_14_147, output_14_4, output_13_147;
mixer gate_output_13_147(.a(output_14_147), .b(output_14_4), .y(output_13_147));
wire output_15_147, output_15_4, output_14_147;
mixer gate_output_14_147(.a(output_15_147), .b(output_15_4), .y(output_14_147));
wire output_16_147, output_16_4, output_15_147;
mixer gate_output_15_147(.a(output_16_147), .b(output_16_4), .y(output_15_147));
wire output_1_148, output_1_5, output_0_148;
mixer gate_output_0_148(.a(output_1_148), .b(output_1_5), .y(output_0_148));
wire output_2_148, output_2_5, output_1_148;
mixer gate_output_1_148(.a(output_2_148), .b(output_2_5), .y(output_1_148));
wire output_3_148, output_3_5, output_2_148;
mixer gate_output_2_148(.a(output_3_148), .b(output_3_5), .y(output_2_148));
wire output_4_148, output_4_5, output_3_148;
mixer gate_output_3_148(.a(output_4_148), .b(output_4_5), .y(output_3_148));
wire output_5_148, output_5_5, output_4_148;
mixer gate_output_4_148(.a(output_5_148), .b(output_5_5), .y(output_4_148));
wire output_6_148, output_6_5, output_5_148;
mixer gate_output_5_148(.a(output_6_148), .b(output_6_5), .y(output_5_148));
wire output_7_148, output_7_5, output_6_148;
mixer gate_output_6_148(.a(output_7_148), .b(output_7_5), .y(output_6_148));
wire output_8_148, output_8_5, output_7_148;
mixer gate_output_7_148(.a(output_8_148), .b(output_8_5), .y(output_7_148));
wire output_9_148, output_9_5, output_8_148;
mixer gate_output_8_148(.a(output_9_148), .b(output_9_5), .y(output_8_148));
wire output_10_148, output_10_5, output_9_148;
mixer gate_output_9_148(.a(output_10_148), .b(output_10_5), .y(output_9_148));
wire output_11_148, output_11_5, output_10_148;
mixer gate_output_10_148(.a(output_11_148), .b(output_11_5), .y(output_10_148));
wire output_12_148, output_12_5, output_11_148;
mixer gate_output_11_148(.a(output_12_148), .b(output_12_5), .y(output_11_148));
wire output_13_148, output_13_5, output_12_148;
mixer gate_output_12_148(.a(output_13_148), .b(output_13_5), .y(output_12_148));
wire output_14_148, output_14_5, output_13_148;
mixer gate_output_13_148(.a(output_14_148), .b(output_14_5), .y(output_13_148));
wire output_15_148, output_15_5, output_14_148;
mixer gate_output_14_148(.a(output_15_148), .b(output_15_5), .y(output_14_148));
wire output_16_148, output_16_5, output_15_148;
mixer gate_output_15_148(.a(output_16_148), .b(output_16_5), .y(output_15_148));
wire output_1_149, output_1_6, output_0_149;
mixer gate_output_0_149(.a(output_1_149), .b(output_1_6), .y(output_0_149));
wire output_2_149, output_2_6, output_1_149;
mixer gate_output_1_149(.a(output_2_149), .b(output_2_6), .y(output_1_149));
wire output_3_149, output_3_6, output_2_149;
mixer gate_output_2_149(.a(output_3_149), .b(output_3_6), .y(output_2_149));
wire output_4_149, output_4_6, output_3_149;
mixer gate_output_3_149(.a(output_4_149), .b(output_4_6), .y(output_3_149));
wire output_5_149, output_5_6, output_4_149;
mixer gate_output_4_149(.a(output_5_149), .b(output_5_6), .y(output_4_149));
wire output_6_149, output_6_6, output_5_149;
mixer gate_output_5_149(.a(output_6_149), .b(output_6_6), .y(output_5_149));
wire output_7_149, output_7_6, output_6_149;
mixer gate_output_6_149(.a(output_7_149), .b(output_7_6), .y(output_6_149));
wire output_8_149, output_8_6, output_7_149;
mixer gate_output_7_149(.a(output_8_149), .b(output_8_6), .y(output_7_149));
wire output_9_149, output_9_6, output_8_149;
mixer gate_output_8_149(.a(output_9_149), .b(output_9_6), .y(output_8_149));
wire output_10_149, output_10_6, output_9_149;
mixer gate_output_9_149(.a(output_10_149), .b(output_10_6), .y(output_9_149));
wire output_11_149, output_11_6, output_10_149;
mixer gate_output_10_149(.a(output_11_149), .b(output_11_6), .y(output_10_149));
wire output_12_149, output_12_6, output_11_149;
mixer gate_output_11_149(.a(output_12_149), .b(output_12_6), .y(output_11_149));
wire output_13_149, output_13_6, output_12_149;
mixer gate_output_12_149(.a(output_13_149), .b(output_13_6), .y(output_12_149));
wire output_14_149, output_14_6, output_13_149;
mixer gate_output_13_149(.a(output_14_149), .b(output_14_6), .y(output_13_149));
wire output_15_149, output_15_6, output_14_149;
mixer gate_output_14_149(.a(output_15_149), .b(output_15_6), .y(output_14_149));
wire output_16_149, output_16_6, output_15_149;
mixer gate_output_15_149(.a(output_16_149), .b(output_16_6), .y(output_15_149));
wire output_1_150, output_1_7, output_0_150;
mixer gate_output_0_150(.a(output_1_150), .b(output_1_7), .y(output_0_150));
wire output_2_150, output_2_7, output_1_150;
mixer gate_output_1_150(.a(output_2_150), .b(output_2_7), .y(output_1_150));
wire output_3_150, output_3_7, output_2_150;
mixer gate_output_2_150(.a(output_3_150), .b(output_3_7), .y(output_2_150));
wire output_4_150, output_4_7, output_3_150;
mixer gate_output_3_150(.a(output_4_150), .b(output_4_7), .y(output_3_150));
wire output_5_150, output_5_7, output_4_150;
mixer gate_output_4_150(.a(output_5_150), .b(output_5_7), .y(output_4_150));
wire output_6_150, output_6_7, output_5_150;
mixer gate_output_5_150(.a(output_6_150), .b(output_6_7), .y(output_5_150));
wire output_7_150, output_7_7, output_6_150;
mixer gate_output_6_150(.a(output_7_150), .b(output_7_7), .y(output_6_150));
wire output_8_150, output_8_7, output_7_150;
mixer gate_output_7_150(.a(output_8_150), .b(output_8_7), .y(output_7_150));
wire output_9_150, output_9_7, output_8_150;
mixer gate_output_8_150(.a(output_9_150), .b(output_9_7), .y(output_8_150));
wire output_10_150, output_10_7, output_9_150;
mixer gate_output_9_150(.a(output_10_150), .b(output_10_7), .y(output_9_150));
wire output_11_150, output_11_7, output_10_150;
mixer gate_output_10_150(.a(output_11_150), .b(output_11_7), .y(output_10_150));
wire output_12_150, output_12_7, output_11_150;
mixer gate_output_11_150(.a(output_12_150), .b(output_12_7), .y(output_11_150));
wire output_13_150, output_13_7, output_12_150;
mixer gate_output_12_150(.a(output_13_150), .b(output_13_7), .y(output_12_150));
wire output_14_150, output_14_7, output_13_150;
mixer gate_output_13_150(.a(output_14_150), .b(output_14_7), .y(output_13_150));
wire output_15_150, output_15_7, output_14_150;
mixer gate_output_14_150(.a(output_15_150), .b(output_15_7), .y(output_14_150));
wire output_16_150, output_16_7, output_15_150;
mixer gate_output_15_150(.a(output_16_150), .b(output_16_7), .y(output_15_150));
wire output_1_151, output_1_8, output_0_151;
mixer gate_output_0_151(.a(output_1_151), .b(output_1_8), .y(output_0_151));
wire output_2_151, output_2_8, output_1_151;
mixer gate_output_1_151(.a(output_2_151), .b(output_2_8), .y(output_1_151));
wire output_3_151, output_3_8, output_2_151;
mixer gate_output_2_151(.a(output_3_151), .b(output_3_8), .y(output_2_151));
wire output_4_151, output_4_8, output_3_151;
mixer gate_output_3_151(.a(output_4_151), .b(output_4_8), .y(output_3_151));
wire output_5_151, output_5_8, output_4_151;
mixer gate_output_4_151(.a(output_5_151), .b(output_5_8), .y(output_4_151));
wire output_6_151, output_6_8, output_5_151;
mixer gate_output_5_151(.a(output_6_151), .b(output_6_8), .y(output_5_151));
wire output_7_151, output_7_8, output_6_151;
mixer gate_output_6_151(.a(output_7_151), .b(output_7_8), .y(output_6_151));
wire output_8_151, output_8_8, output_7_151;
mixer gate_output_7_151(.a(output_8_151), .b(output_8_8), .y(output_7_151));
wire output_9_151, output_9_8, output_8_151;
mixer gate_output_8_151(.a(output_9_151), .b(output_9_8), .y(output_8_151));
wire output_10_151, output_10_8, output_9_151;
mixer gate_output_9_151(.a(output_10_151), .b(output_10_8), .y(output_9_151));
wire output_11_151, output_11_8, output_10_151;
mixer gate_output_10_151(.a(output_11_151), .b(output_11_8), .y(output_10_151));
wire output_12_151, output_12_8, output_11_151;
mixer gate_output_11_151(.a(output_12_151), .b(output_12_8), .y(output_11_151));
wire output_13_151, output_13_8, output_12_151;
mixer gate_output_12_151(.a(output_13_151), .b(output_13_8), .y(output_12_151));
wire output_14_151, output_14_8, output_13_151;
mixer gate_output_13_151(.a(output_14_151), .b(output_14_8), .y(output_13_151));
wire output_15_151, output_15_8, output_14_151;
mixer gate_output_14_151(.a(output_15_151), .b(output_15_8), .y(output_14_151));
wire output_16_151, output_16_8, output_15_151;
mixer gate_output_15_151(.a(output_16_151), .b(output_16_8), .y(output_15_151));
wire output_1_152, output_1_9, output_0_152;
mixer gate_output_0_152(.a(output_1_152), .b(output_1_9), .y(output_0_152));
wire output_2_152, output_2_9, output_1_152;
mixer gate_output_1_152(.a(output_2_152), .b(output_2_9), .y(output_1_152));
wire output_3_152, output_3_9, output_2_152;
mixer gate_output_2_152(.a(output_3_152), .b(output_3_9), .y(output_2_152));
wire output_4_152, output_4_9, output_3_152;
mixer gate_output_3_152(.a(output_4_152), .b(output_4_9), .y(output_3_152));
wire output_5_152, output_5_9, output_4_152;
mixer gate_output_4_152(.a(output_5_152), .b(output_5_9), .y(output_4_152));
wire output_6_152, output_6_9, output_5_152;
mixer gate_output_5_152(.a(output_6_152), .b(output_6_9), .y(output_5_152));
wire output_7_152, output_7_9, output_6_152;
mixer gate_output_6_152(.a(output_7_152), .b(output_7_9), .y(output_6_152));
wire output_8_152, output_8_9, output_7_152;
mixer gate_output_7_152(.a(output_8_152), .b(output_8_9), .y(output_7_152));
wire output_9_152, output_9_9, output_8_152;
mixer gate_output_8_152(.a(output_9_152), .b(output_9_9), .y(output_8_152));
wire output_10_152, output_10_9, output_9_152;
mixer gate_output_9_152(.a(output_10_152), .b(output_10_9), .y(output_9_152));
wire output_11_152, output_11_9, output_10_152;
mixer gate_output_10_152(.a(output_11_152), .b(output_11_9), .y(output_10_152));
wire output_12_152, output_12_9, output_11_152;
mixer gate_output_11_152(.a(output_12_152), .b(output_12_9), .y(output_11_152));
wire output_13_152, output_13_9, output_12_152;
mixer gate_output_12_152(.a(output_13_152), .b(output_13_9), .y(output_12_152));
wire output_14_152, output_14_9, output_13_152;
mixer gate_output_13_152(.a(output_14_152), .b(output_14_9), .y(output_13_152));
wire output_15_152, output_15_9, output_14_152;
mixer gate_output_14_152(.a(output_15_152), .b(output_15_9), .y(output_14_152));
wire output_16_152, output_16_9, output_15_152;
mixer gate_output_15_152(.a(output_16_152), .b(output_16_9), .y(output_15_152));
wire output_1_153, output_1_10, output_0_153;
mixer gate_output_0_153(.a(output_1_153), .b(output_1_10), .y(output_0_153));
wire output_2_153, output_2_10, output_1_153;
mixer gate_output_1_153(.a(output_2_153), .b(output_2_10), .y(output_1_153));
wire output_3_153, output_3_10, output_2_153;
mixer gate_output_2_153(.a(output_3_153), .b(output_3_10), .y(output_2_153));
wire output_4_153, output_4_10, output_3_153;
mixer gate_output_3_153(.a(output_4_153), .b(output_4_10), .y(output_3_153));
wire output_5_153, output_5_10, output_4_153;
mixer gate_output_4_153(.a(output_5_153), .b(output_5_10), .y(output_4_153));
wire output_6_153, output_6_10, output_5_153;
mixer gate_output_5_153(.a(output_6_153), .b(output_6_10), .y(output_5_153));
wire output_7_153, output_7_10, output_6_153;
mixer gate_output_6_153(.a(output_7_153), .b(output_7_10), .y(output_6_153));
wire output_8_153, output_8_10, output_7_153;
mixer gate_output_7_153(.a(output_8_153), .b(output_8_10), .y(output_7_153));
wire output_9_153, output_9_10, output_8_153;
mixer gate_output_8_153(.a(output_9_153), .b(output_9_10), .y(output_8_153));
wire output_10_153, output_10_10, output_9_153;
mixer gate_output_9_153(.a(output_10_153), .b(output_10_10), .y(output_9_153));
wire output_11_153, output_11_10, output_10_153;
mixer gate_output_10_153(.a(output_11_153), .b(output_11_10), .y(output_10_153));
wire output_12_153, output_12_10, output_11_153;
mixer gate_output_11_153(.a(output_12_153), .b(output_12_10), .y(output_11_153));
wire output_13_153, output_13_10, output_12_153;
mixer gate_output_12_153(.a(output_13_153), .b(output_13_10), .y(output_12_153));
wire output_14_153, output_14_10, output_13_153;
mixer gate_output_13_153(.a(output_14_153), .b(output_14_10), .y(output_13_153));
wire output_15_153, output_15_10, output_14_153;
mixer gate_output_14_153(.a(output_15_153), .b(output_15_10), .y(output_14_153));
wire output_16_153, output_16_10, output_15_153;
mixer gate_output_15_153(.a(output_16_153), .b(output_16_10), .y(output_15_153));
wire output_1_154, output_1_11, output_0_154;
mixer gate_output_0_154(.a(output_1_154), .b(output_1_11), .y(output_0_154));
wire output_2_154, output_2_11, output_1_154;
mixer gate_output_1_154(.a(output_2_154), .b(output_2_11), .y(output_1_154));
wire output_3_154, output_3_11, output_2_154;
mixer gate_output_2_154(.a(output_3_154), .b(output_3_11), .y(output_2_154));
wire output_4_154, output_4_11, output_3_154;
mixer gate_output_3_154(.a(output_4_154), .b(output_4_11), .y(output_3_154));
wire output_5_154, output_5_11, output_4_154;
mixer gate_output_4_154(.a(output_5_154), .b(output_5_11), .y(output_4_154));
wire output_6_154, output_6_11, output_5_154;
mixer gate_output_5_154(.a(output_6_154), .b(output_6_11), .y(output_5_154));
wire output_7_154, output_7_11, output_6_154;
mixer gate_output_6_154(.a(output_7_154), .b(output_7_11), .y(output_6_154));
wire output_8_154, output_8_11, output_7_154;
mixer gate_output_7_154(.a(output_8_154), .b(output_8_11), .y(output_7_154));
wire output_9_154, output_9_11, output_8_154;
mixer gate_output_8_154(.a(output_9_154), .b(output_9_11), .y(output_8_154));
wire output_10_154, output_10_11, output_9_154;
mixer gate_output_9_154(.a(output_10_154), .b(output_10_11), .y(output_9_154));
wire output_11_154, output_11_11, output_10_154;
mixer gate_output_10_154(.a(output_11_154), .b(output_11_11), .y(output_10_154));
wire output_12_154, output_12_11, output_11_154;
mixer gate_output_11_154(.a(output_12_154), .b(output_12_11), .y(output_11_154));
wire output_13_154, output_13_11, output_12_154;
mixer gate_output_12_154(.a(output_13_154), .b(output_13_11), .y(output_12_154));
wire output_14_154, output_14_11, output_13_154;
mixer gate_output_13_154(.a(output_14_154), .b(output_14_11), .y(output_13_154));
wire output_15_154, output_15_11, output_14_154;
mixer gate_output_14_154(.a(output_15_154), .b(output_15_11), .y(output_14_154));
wire output_16_154, output_16_11, output_15_154;
mixer gate_output_15_154(.a(output_16_154), .b(output_16_11), .y(output_15_154));
wire output_1_155, output_1_12, output_0_155;
mixer gate_output_0_155(.a(output_1_155), .b(output_1_12), .y(output_0_155));
wire output_2_155, output_2_12, output_1_155;
mixer gate_output_1_155(.a(output_2_155), .b(output_2_12), .y(output_1_155));
wire output_3_155, output_3_12, output_2_155;
mixer gate_output_2_155(.a(output_3_155), .b(output_3_12), .y(output_2_155));
wire output_4_155, output_4_12, output_3_155;
mixer gate_output_3_155(.a(output_4_155), .b(output_4_12), .y(output_3_155));
wire output_5_155, output_5_12, output_4_155;
mixer gate_output_4_155(.a(output_5_155), .b(output_5_12), .y(output_4_155));
wire output_6_155, output_6_12, output_5_155;
mixer gate_output_5_155(.a(output_6_155), .b(output_6_12), .y(output_5_155));
wire output_7_155, output_7_12, output_6_155;
mixer gate_output_6_155(.a(output_7_155), .b(output_7_12), .y(output_6_155));
wire output_8_155, output_8_12, output_7_155;
mixer gate_output_7_155(.a(output_8_155), .b(output_8_12), .y(output_7_155));
wire output_9_155, output_9_12, output_8_155;
mixer gate_output_8_155(.a(output_9_155), .b(output_9_12), .y(output_8_155));
wire output_10_155, output_10_12, output_9_155;
mixer gate_output_9_155(.a(output_10_155), .b(output_10_12), .y(output_9_155));
wire output_11_155, output_11_12, output_10_155;
mixer gate_output_10_155(.a(output_11_155), .b(output_11_12), .y(output_10_155));
wire output_12_155, output_12_12, output_11_155;
mixer gate_output_11_155(.a(output_12_155), .b(output_12_12), .y(output_11_155));
wire output_13_155, output_13_12, output_12_155;
mixer gate_output_12_155(.a(output_13_155), .b(output_13_12), .y(output_12_155));
wire output_14_155, output_14_12, output_13_155;
mixer gate_output_13_155(.a(output_14_155), .b(output_14_12), .y(output_13_155));
wire output_15_155, output_15_12, output_14_155;
mixer gate_output_14_155(.a(output_15_155), .b(output_15_12), .y(output_14_155));
wire output_16_155, output_16_12, output_15_155;
mixer gate_output_15_155(.a(output_16_155), .b(output_16_12), .y(output_15_155));
wire output_1_156, output_1_13, output_0_156;
mixer gate_output_0_156(.a(output_1_156), .b(output_1_13), .y(output_0_156));
wire output_2_156, output_2_13, output_1_156;
mixer gate_output_1_156(.a(output_2_156), .b(output_2_13), .y(output_1_156));
wire output_3_156, output_3_13, output_2_156;
mixer gate_output_2_156(.a(output_3_156), .b(output_3_13), .y(output_2_156));
wire output_4_156, output_4_13, output_3_156;
mixer gate_output_3_156(.a(output_4_156), .b(output_4_13), .y(output_3_156));
wire output_5_156, output_5_13, output_4_156;
mixer gate_output_4_156(.a(output_5_156), .b(output_5_13), .y(output_4_156));
wire output_6_156, output_6_13, output_5_156;
mixer gate_output_5_156(.a(output_6_156), .b(output_6_13), .y(output_5_156));
wire output_7_156, output_7_13, output_6_156;
mixer gate_output_6_156(.a(output_7_156), .b(output_7_13), .y(output_6_156));
wire output_8_156, output_8_13, output_7_156;
mixer gate_output_7_156(.a(output_8_156), .b(output_8_13), .y(output_7_156));
wire output_9_156, output_9_13, output_8_156;
mixer gate_output_8_156(.a(output_9_156), .b(output_9_13), .y(output_8_156));
wire output_10_156, output_10_13, output_9_156;
mixer gate_output_9_156(.a(output_10_156), .b(output_10_13), .y(output_9_156));
wire output_11_156, output_11_13, output_10_156;
mixer gate_output_10_156(.a(output_11_156), .b(output_11_13), .y(output_10_156));
wire output_12_156, output_12_13, output_11_156;
mixer gate_output_11_156(.a(output_12_156), .b(output_12_13), .y(output_11_156));
wire output_13_156, output_13_13, output_12_156;
mixer gate_output_12_156(.a(output_13_156), .b(output_13_13), .y(output_12_156));
wire output_14_156, output_14_13, output_13_156;
mixer gate_output_13_156(.a(output_14_156), .b(output_14_13), .y(output_13_156));
wire output_15_156, output_15_13, output_14_156;
mixer gate_output_14_156(.a(output_15_156), .b(output_15_13), .y(output_14_156));
wire output_16_156, output_16_13, output_15_156;
mixer gate_output_15_156(.a(output_16_156), .b(output_16_13), .y(output_15_156));
wire output_1_157, output_1_14, output_0_157;
mixer gate_output_0_157(.a(output_1_157), .b(output_1_14), .y(output_0_157));
wire output_2_157, output_2_14, output_1_157;
mixer gate_output_1_157(.a(output_2_157), .b(output_2_14), .y(output_1_157));
wire output_3_157, output_3_14, output_2_157;
mixer gate_output_2_157(.a(output_3_157), .b(output_3_14), .y(output_2_157));
wire output_4_157, output_4_14, output_3_157;
mixer gate_output_3_157(.a(output_4_157), .b(output_4_14), .y(output_3_157));
wire output_5_157, output_5_14, output_4_157;
mixer gate_output_4_157(.a(output_5_157), .b(output_5_14), .y(output_4_157));
wire output_6_157, output_6_14, output_5_157;
mixer gate_output_5_157(.a(output_6_157), .b(output_6_14), .y(output_5_157));
wire output_7_157, output_7_14, output_6_157;
mixer gate_output_6_157(.a(output_7_157), .b(output_7_14), .y(output_6_157));
wire output_8_157, output_8_14, output_7_157;
mixer gate_output_7_157(.a(output_8_157), .b(output_8_14), .y(output_7_157));
wire output_9_157, output_9_14, output_8_157;
mixer gate_output_8_157(.a(output_9_157), .b(output_9_14), .y(output_8_157));
wire output_10_157, output_10_14, output_9_157;
mixer gate_output_9_157(.a(output_10_157), .b(output_10_14), .y(output_9_157));
wire output_11_157, output_11_14, output_10_157;
mixer gate_output_10_157(.a(output_11_157), .b(output_11_14), .y(output_10_157));
wire output_12_157, output_12_14, output_11_157;
mixer gate_output_11_157(.a(output_12_157), .b(output_12_14), .y(output_11_157));
wire output_13_157, output_13_14, output_12_157;
mixer gate_output_12_157(.a(output_13_157), .b(output_13_14), .y(output_12_157));
wire output_14_157, output_14_14, output_13_157;
mixer gate_output_13_157(.a(output_14_157), .b(output_14_14), .y(output_13_157));
wire output_15_157, output_15_14, output_14_157;
mixer gate_output_14_157(.a(output_15_157), .b(output_15_14), .y(output_14_157));
wire output_16_157, output_16_14, output_15_157;
mixer gate_output_15_157(.a(output_16_157), .b(output_16_14), .y(output_15_157));
wire output_1_158, output_1_15, output_0_158;
mixer gate_output_0_158(.a(output_1_158), .b(output_1_15), .y(output_0_158));
wire output_2_158, output_2_15, output_1_158;
mixer gate_output_1_158(.a(output_2_158), .b(output_2_15), .y(output_1_158));
wire output_3_158, output_3_15, output_2_158;
mixer gate_output_2_158(.a(output_3_158), .b(output_3_15), .y(output_2_158));
wire output_4_158, output_4_15, output_3_158;
mixer gate_output_3_158(.a(output_4_158), .b(output_4_15), .y(output_3_158));
wire output_5_158, output_5_15, output_4_158;
mixer gate_output_4_158(.a(output_5_158), .b(output_5_15), .y(output_4_158));
wire output_6_158, output_6_15, output_5_158;
mixer gate_output_5_158(.a(output_6_158), .b(output_6_15), .y(output_5_158));
wire output_7_158, output_7_15, output_6_158;
mixer gate_output_6_158(.a(output_7_158), .b(output_7_15), .y(output_6_158));
wire output_8_158, output_8_15, output_7_158;
mixer gate_output_7_158(.a(output_8_158), .b(output_8_15), .y(output_7_158));
wire output_9_158, output_9_15, output_8_158;
mixer gate_output_8_158(.a(output_9_158), .b(output_9_15), .y(output_8_158));
wire output_10_158, output_10_15, output_9_158;
mixer gate_output_9_158(.a(output_10_158), .b(output_10_15), .y(output_9_158));
wire output_11_158, output_11_15, output_10_158;
mixer gate_output_10_158(.a(output_11_158), .b(output_11_15), .y(output_10_158));
wire output_12_158, output_12_15, output_11_158;
mixer gate_output_11_158(.a(output_12_158), .b(output_12_15), .y(output_11_158));
wire output_13_158, output_13_15, output_12_158;
mixer gate_output_12_158(.a(output_13_158), .b(output_13_15), .y(output_12_158));
wire output_14_158, output_14_15, output_13_158;
mixer gate_output_13_158(.a(output_14_158), .b(output_14_15), .y(output_13_158));
wire output_15_158, output_15_15, output_14_158;
mixer gate_output_14_158(.a(output_15_158), .b(output_15_15), .y(output_14_158));
wire output_16_158, output_16_15, output_15_158;
mixer gate_output_15_158(.a(output_16_158), .b(output_16_15), .y(output_15_158));
wire output_1_159, output_1_0, output_0_159;
mixer gate_output_0_159(.a(output_1_159), .b(output_1_0), .y(output_0_159));
wire output_2_159, output_2_0, output_1_159;
mixer gate_output_1_159(.a(output_2_159), .b(output_2_0), .y(output_1_159));
wire output_3_159, output_3_0, output_2_159;
mixer gate_output_2_159(.a(output_3_159), .b(output_3_0), .y(output_2_159));
wire output_4_159, output_4_0, output_3_159;
mixer gate_output_3_159(.a(output_4_159), .b(output_4_0), .y(output_3_159));
wire output_5_159, output_5_0, output_4_159;
mixer gate_output_4_159(.a(output_5_159), .b(output_5_0), .y(output_4_159));
wire output_6_159, output_6_0, output_5_159;
mixer gate_output_5_159(.a(output_6_159), .b(output_6_0), .y(output_5_159));
wire output_7_159, output_7_0, output_6_159;
mixer gate_output_6_159(.a(output_7_159), .b(output_7_0), .y(output_6_159));
wire output_8_159, output_8_0, output_7_159;
mixer gate_output_7_159(.a(output_8_159), .b(output_8_0), .y(output_7_159));
wire output_9_159, output_9_0, output_8_159;
mixer gate_output_8_159(.a(output_9_159), .b(output_9_0), .y(output_8_159));
wire output_10_159, output_10_0, output_9_159;
mixer gate_output_9_159(.a(output_10_159), .b(output_10_0), .y(output_9_159));
wire output_11_159, output_11_0, output_10_159;
mixer gate_output_10_159(.a(output_11_159), .b(output_11_0), .y(output_10_159));
wire output_12_159, output_12_0, output_11_159;
mixer gate_output_11_159(.a(output_12_159), .b(output_12_0), .y(output_11_159));
wire output_13_159, output_13_0, output_12_159;
mixer gate_output_12_159(.a(output_13_159), .b(output_13_0), .y(output_12_159));
wire output_14_159, output_14_0, output_13_159;
mixer gate_output_13_159(.a(output_14_159), .b(output_14_0), .y(output_13_159));
wire output_15_159, output_15_0, output_14_159;
mixer gate_output_14_159(.a(output_15_159), .b(output_15_0), .y(output_14_159));
wire output_16_159, output_16_0, output_15_159;
mixer gate_output_15_159(.a(output_16_159), .b(output_16_0), .y(output_15_159));
wire output_1_160, output_1_1, output_0_160;
mixer gate_output_0_160(.a(output_1_160), .b(output_1_1), .y(output_0_160));
wire output_2_160, output_2_1, output_1_160;
mixer gate_output_1_160(.a(output_2_160), .b(output_2_1), .y(output_1_160));
wire output_3_160, output_3_1, output_2_160;
mixer gate_output_2_160(.a(output_3_160), .b(output_3_1), .y(output_2_160));
wire output_4_160, output_4_1, output_3_160;
mixer gate_output_3_160(.a(output_4_160), .b(output_4_1), .y(output_3_160));
wire output_5_160, output_5_1, output_4_160;
mixer gate_output_4_160(.a(output_5_160), .b(output_5_1), .y(output_4_160));
wire output_6_160, output_6_1, output_5_160;
mixer gate_output_5_160(.a(output_6_160), .b(output_6_1), .y(output_5_160));
wire output_7_160, output_7_1, output_6_160;
mixer gate_output_6_160(.a(output_7_160), .b(output_7_1), .y(output_6_160));
wire output_8_160, output_8_1, output_7_160;
mixer gate_output_7_160(.a(output_8_160), .b(output_8_1), .y(output_7_160));
wire output_9_160, output_9_1, output_8_160;
mixer gate_output_8_160(.a(output_9_160), .b(output_9_1), .y(output_8_160));
wire output_10_160, output_10_1, output_9_160;
mixer gate_output_9_160(.a(output_10_160), .b(output_10_1), .y(output_9_160));
wire output_11_160, output_11_1, output_10_160;
mixer gate_output_10_160(.a(output_11_160), .b(output_11_1), .y(output_10_160));
wire output_12_160, output_12_1, output_11_160;
mixer gate_output_11_160(.a(output_12_160), .b(output_12_1), .y(output_11_160));
wire output_13_160, output_13_1, output_12_160;
mixer gate_output_12_160(.a(output_13_160), .b(output_13_1), .y(output_12_160));
wire output_14_160, output_14_1, output_13_160;
mixer gate_output_13_160(.a(output_14_160), .b(output_14_1), .y(output_13_160));
wire output_15_160, output_15_1, output_14_160;
mixer gate_output_14_160(.a(output_15_160), .b(output_15_1), .y(output_14_160));
wire output_16_160, output_16_1, output_15_160;
mixer gate_output_15_160(.a(output_16_160), .b(output_16_1), .y(output_15_160));
wire output_1_161, output_1_2, output_0_161;
mixer gate_output_0_161(.a(output_1_161), .b(output_1_2), .y(output_0_161));
wire output_2_161, output_2_2, output_1_161;
mixer gate_output_1_161(.a(output_2_161), .b(output_2_2), .y(output_1_161));
wire output_3_161, output_3_2, output_2_161;
mixer gate_output_2_161(.a(output_3_161), .b(output_3_2), .y(output_2_161));
wire output_4_161, output_4_2, output_3_161;
mixer gate_output_3_161(.a(output_4_161), .b(output_4_2), .y(output_3_161));
wire output_5_161, output_5_2, output_4_161;
mixer gate_output_4_161(.a(output_5_161), .b(output_5_2), .y(output_4_161));
wire output_6_161, output_6_2, output_5_161;
mixer gate_output_5_161(.a(output_6_161), .b(output_6_2), .y(output_5_161));
wire output_7_161, output_7_2, output_6_161;
mixer gate_output_6_161(.a(output_7_161), .b(output_7_2), .y(output_6_161));
wire output_8_161, output_8_2, output_7_161;
mixer gate_output_7_161(.a(output_8_161), .b(output_8_2), .y(output_7_161));
wire output_9_161, output_9_2, output_8_161;
mixer gate_output_8_161(.a(output_9_161), .b(output_9_2), .y(output_8_161));
wire output_10_161, output_10_2, output_9_161;
mixer gate_output_9_161(.a(output_10_161), .b(output_10_2), .y(output_9_161));
wire output_11_161, output_11_2, output_10_161;
mixer gate_output_10_161(.a(output_11_161), .b(output_11_2), .y(output_10_161));
wire output_12_161, output_12_2, output_11_161;
mixer gate_output_11_161(.a(output_12_161), .b(output_12_2), .y(output_11_161));
wire output_13_161, output_13_2, output_12_161;
mixer gate_output_12_161(.a(output_13_161), .b(output_13_2), .y(output_12_161));
wire output_14_161, output_14_2, output_13_161;
mixer gate_output_13_161(.a(output_14_161), .b(output_14_2), .y(output_13_161));
wire output_15_161, output_15_2, output_14_161;
mixer gate_output_14_161(.a(output_15_161), .b(output_15_2), .y(output_14_161));
wire output_16_161, output_16_2, output_15_161;
mixer gate_output_15_161(.a(output_16_161), .b(output_16_2), .y(output_15_161));
wire output_1_162, output_1_3, output_0_162;
mixer gate_output_0_162(.a(output_1_162), .b(output_1_3), .y(output_0_162));
wire output_2_162, output_2_3, output_1_162;
mixer gate_output_1_162(.a(output_2_162), .b(output_2_3), .y(output_1_162));
wire output_3_162, output_3_3, output_2_162;
mixer gate_output_2_162(.a(output_3_162), .b(output_3_3), .y(output_2_162));
wire output_4_162, output_4_3, output_3_162;
mixer gate_output_3_162(.a(output_4_162), .b(output_4_3), .y(output_3_162));
wire output_5_162, output_5_3, output_4_162;
mixer gate_output_4_162(.a(output_5_162), .b(output_5_3), .y(output_4_162));
wire output_6_162, output_6_3, output_5_162;
mixer gate_output_5_162(.a(output_6_162), .b(output_6_3), .y(output_5_162));
wire output_7_162, output_7_3, output_6_162;
mixer gate_output_6_162(.a(output_7_162), .b(output_7_3), .y(output_6_162));
wire output_8_162, output_8_3, output_7_162;
mixer gate_output_7_162(.a(output_8_162), .b(output_8_3), .y(output_7_162));
wire output_9_162, output_9_3, output_8_162;
mixer gate_output_8_162(.a(output_9_162), .b(output_9_3), .y(output_8_162));
wire output_10_162, output_10_3, output_9_162;
mixer gate_output_9_162(.a(output_10_162), .b(output_10_3), .y(output_9_162));
wire output_11_162, output_11_3, output_10_162;
mixer gate_output_10_162(.a(output_11_162), .b(output_11_3), .y(output_10_162));
wire output_12_162, output_12_3, output_11_162;
mixer gate_output_11_162(.a(output_12_162), .b(output_12_3), .y(output_11_162));
wire output_13_162, output_13_3, output_12_162;
mixer gate_output_12_162(.a(output_13_162), .b(output_13_3), .y(output_12_162));
wire output_14_162, output_14_3, output_13_162;
mixer gate_output_13_162(.a(output_14_162), .b(output_14_3), .y(output_13_162));
wire output_15_162, output_15_3, output_14_162;
mixer gate_output_14_162(.a(output_15_162), .b(output_15_3), .y(output_14_162));
wire output_16_162, output_16_3, output_15_162;
mixer gate_output_15_162(.a(output_16_162), .b(output_16_3), .y(output_15_162));
wire output_1_163, output_1_4, output_0_163;
mixer gate_output_0_163(.a(output_1_163), .b(output_1_4), .y(output_0_163));
wire output_2_163, output_2_4, output_1_163;
mixer gate_output_1_163(.a(output_2_163), .b(output_2_4), .y(output_1_163));
wire output_3_163, output_3_4, output_2_163;
mixer gate_output_2_163(.a(output_3_163), .b(output_3_4), .y(output_2_163));
wire output_4_163, output_4_4, output_3_163;
mixer gate_output_3_163(.a(output_4_163), .b(output_4_4), .y(output_3_163));
wire output_5_163, output_5_4, output_4_163;
mixer gate_output_4_163(.a(output_5_163), .b(output_5_4), .y(output_4_163));
wire output_6_163, output_6_4, output_5_163;
mixer gate_output_5_163(.a(output_6_163), .b(output_6_4), .y(output_5_163));
wire output_7_163, output_7_4, output_6_163;
mixer gate_output_6_163(.a(output_7_163), .b(output_7_4), .y(output_6_163));
wire output_8_163, output_8_4, output_7_163;
mixer gate_output_7_163(.a(output_8_163), .b(output_8_4), .y(output_7_163));
wire output_9_163, output_9_4, output_8_163;
mixer gate_output_8_163(.a(output_9_163), .b(output_9_4), .y(output_8_163));
wire output_10_163, output_10_4, output_9_163;
mixer gate_output_9_163(.a(output_10_163), .b(output_10_4), .y(output_9_163));
wire output_11_163, output_11_4, output_10_163;
mixer gate_output_10_163(.a(output_11_163), .b(output_11_4), .y(output_10_163));
wire output_12_163, output_12_4, output_11_163;
mixer gate_output_11_163(.a(output_12_163), .b(output_12_4), .y(output_11_163));
wire output_13_163, output_13_4, output_12_163;
mixer gate_output_12_163(.a(output_13_163), .b(output_13_4), .y(output_12_163));
wire output_14_163, output_14_4, output_13_163;
mixer gate_output_13_163(.a(output_14_163), .b(output_14_4), .y(output_13_163));
wire output_15_163, output_15_4, output_14_163;
mixer gate_output_14_163(.a(output_15_163), .b(output_15_4), .y(output_14_163));
wire output_16_163, output_16_4, output_15_163;
mixer gate_output_15_163(.a(output_16_163), .b(output_16_4), .y(output_15_163));
wire output_1_164, output_1_5, output_0_164;
mixer gate_output_0_164(.a(output_1_164), .b(output_1_5), .y(output_0_164));
wire output_2_164, output_2_5, output_1_164;
mixer gate_output_1_164(.a(output_2_164), .b(output_2_5), .y(output_1_164));
wire output_3_164, output_3_5, output_2_164;
mixer gate_output_2_164(.a(output_3_164), .b(output_3_5), .y(output_2_164));
wire output_4_164, output_4_5, output_3_164;
mixer gate_output_3_164(.a(output_4_164), .b(output_4_5), .y(output_3_164));
wire output_5_164, output_5_5, output_4_164;
mixer gate_output_4_164(.a(output_5_164), .b(output_5_5), .y(output_4_164));
wire output_6_164, output_6_5, output_5_164;
mixer gate_output_5_164(.a(output_6_164), .b(output_6_5), .y(output_5_164));
wire output_7_164, output_7_5, output_6_164;
mixer gate_output_6_164(.a(output_7_164), .b(output_7_5), .y(output_6_164));
wire output_8_164, output_8_5, output_7_164;
mixer gate_output_7_164(.a(output_8_164), .b(output_8_5), .y(output_7_164));
wire output_9_164, output_9_5, output_8_164;
mixer gate_output_8_164(.a(output_9_164), .b(output_9_5), .y(output_8_164));
wire output_10_164, output_10_5, output_9_164;
mixer gate_output_9_164(.a(output_10_164), .b(output_10_5), .y(output_9_164));
wire output_11_164, output_11_5, output_10_164;
mixer gate_output_10_164(.a(output_11_164), .b(output_11_5), .y(output_10_164));
wire output_12_164, output_12_5, output_11_164;
mixer gate_output_11_164(.a(output_12_164), .b(output_12_5), .y(output_11_164));
wire output_13_164, output_13_5, output_12_164;
mixer gate_output_12_164(.a(output_13_164), .b(output_13_5), .y(output_12_164));
wire output_14_164, output_14_5, output_13_164;
mixer gate_output_13_164(.a(output_14_164), .b(output_14_5), .y(output_13_164));
wire output_15_164, output_15_5, output_14_164;
mixer gate_output_14_164(.a(output_15_164), .b(output_15_5), .y(output_14_164));
wire output_16_164, output_16_5, output_15_164;
mixer gate_output_15_164(.a(output_16_164), .b(output_16_5), .y(output_15_164));
wire output_1_165, output_1_6, output_0_165;
mixer gate_output_0_165(.a(output_1_165), .b(output_1_6), .y(output_0_165));
wire output_2_165, output_2_6, output_1_165;
mixer gate_output_1_165(.a(output_2_165), .b(output_2_6), .y(output_1_165));
wire output_3_165, output_3_6, output_2_165;
mixer gate_output_2_165(.a(output_3_165), .b(output_3_6), .y(output_2_165));
wire output_4_165, output_4_6, output_3_165;
mixer gate_output_3_165(.a(output_4_165), .b(output_4_6), .y(output_3_165));
wire output_5_165, output_5_6, output_4_165;
mixer gate_output_4_165(.a(output_5_165), .b(output_5_6), .y(output_4_165));
wire output_6_165, output_6_6, output_5_165;
mixer gate_output_5_165(.a(output_6_165), .b(output_6_6), .y(output_5_165));
wire output_7_165, output_7_6, output_6_165;
mixer gate_output_6_165(.a(output_7_165), .b(output_7_6), .y(output_6_165));
wire output_8_165, output_8_6, output_7_165;
mixer gate_output_7_165(.a(output_8_165), .b(output_8_6), .y(output_7_165));
wire output_9_165, output_9_6, output_8_165;
mixer gate_output_8_165(.a(output_9_165), .b(output_9_6), .y(output_8_165));
wire output_10_165, output_10_6, output_9_165;
mixer gate_output_9_165(.a(output_10_165), .b(output_10_6), .y(output_9_165));
wire output_11_165, output_11_6, output_10_165;
mixer gate_output_10_165(.a(output_11_165), .b(output_11_6), .y(output_10_165));
wire output_12_165, output_12_6, output_11_165;
mixer gate_output_11_165(.a(output_12_165), .b(output_12_6), .y(output_11_165));
wire output_13_165, output_13_6, output_12_165;
mixer gate_output_12_165(.a(output_13_165), .b(output_13_6), .y(output_12_165));
wire output_14_165, output_14_6, output_13_165;
mixer gate_output_13_165(.a(output_14_165), .b(output_14_6), .y(output_13_165));
wire output_15_165, output_15_6, output_14_165;
mixer gate_output_14_165(.a(output_15_165), .b(output_15_6), .y(output_14_165));
wire output_16_165, output_16_6, output_15_165;
mixer gate_output_15_165(.a(output_16_165), .b(output_16_6), .y(output_15_165));
wire output_1_166, output_1_7, output_0_166;
mixer gate_output_0_166(.a(output_1_166), .b(output_1_7), .y(output_0_166));
wire output_2_166, output_2_7, output_1_166;
mixer gate_output_1_166(.a(output_2_166), .b(output_2_7), .y(output_1_166));
wire output_3_166, output_3_7, output_2_166;
mixer gate_output_2_166(.a(output_3_166), .b(output_3_7), .y(output_2_166));
wire output_4_166, output_4_7, output_3_166;
mixer gate_output_3_166(.a(output_4_166), .b(output_4_7), .y(output_3_166));
wire output_5_166, output_5_7, output_4_166;
mixer gate_output_4_166(.a(output_5_166), .b(output_5_7), .y(output_4_166));
wire output_6_166, output_6_7, output_5_166;
mixer gate_output_5_166(.a(output_6_166), .b(output_6_7), .y(output_5_166));
wire output_7_166, output_7_7, output_6_166;
mixer gate_output_6_166(.a(output_7_166), .b(output_7_7), .y(output_6_166));
wire output_8_166, output_8_7, output_7_166;
mixer gate_output_7_166(.a(output_8_166), .b(output_8_7), .y(output_7_166));
wire output_9_166, output_9_7, output_8_166;
mixer gate_output_8_166(.a(output_9_166), .b(output_9_7), .y(output_8_166));
wire output_10_166, output_10_7, output_9_166;
mixer gate_output_9_166(.a(output_10_166), .b(output_10_7), .y(output_9_166));
wire output_11_166, output_11_7, output_10_166;
mixer gate_output_10_166(.a(output_11_166), .b(output_11_7), .y(output_10_166));
wire output_12_166, output_12_7, output_11_166;
mixer gate_output_11_166(.a(output_12_166), .b(output_12_7), .y(output_11_166));
wire output_13_166, output_13_7, output_12_166;
mixer gate_output_12_166(.a(output_13_166), .b(output_13_7), .y(output_12_166));
wire output_14_166, output_14_7, output_13_166;
mixer gate_output_13_166(.a(output_14_166), .b(output_14_7), .y(output_13_166));
wire output_15_166, output_15_7, output_14_166;
mixer gate_output_14_166(.a(output_15_166), .b(output_15_7), .y(output_14_166));
wire output_16_166, output_16_7, output_15_166;
mixer gate_output_15_166(.a(output_16_166), .b(output_16_7), .y(output_15_166));
wire output_1_167, output_1_8, output_0_167;
mixer gate_output_0_167(.a(output_1_167), .b(output_1_8), .y(output_0_167));
wire output_2_167, output_2_8, output_1_167;
mixer gate_output_1_167(.a(output_2_167), .b(output_2_8), .y(output_1_167));
wire output_3_167, output_3_8, output_2_167;
mixer gate_output_2_167(.a(output_3_167), .b(output_3_8), .y(output_2_167));
wire output_4_167, output_4_8, output_3_167;
mixer gate_output_3_167(.a(output_4_167), .b(output_4_8), .y(output_3_167));
wire output_5_167, output_5_8, output_4_167;
mixer gate_output_4_167(.a(output_5_167), .b(output_5_8), .y(output_4_167));
wire output_6_167, output_6_8, output_5_167;
mixer gate_output_5_167(.a(output_6_167), .b(output_6_8), .y(output_5_167));
wire output_7_167, output_7_8, output_6_167;
mixer gate_output_6_167(.a(output_7_167), .b(output_7_8), .y(output_6_167));
wire output_8_167, output_8_8, output_7_167;
mixer gate_output_7_167(.a(output_8_167), .b(output_8_8), .y(output_7_167));
wire output_9_167, output_9_8, output_8_167;
mixer gate_output_8_167(.a(output_9_167), .b(output_9_8), .y(output_8_167));
wire output_10_167, output_10_8, output_9_167;
mixer gate_output_9_167(.a(output_10_167), .b(output_10_8), .y(output_9_167));
wire output_11_167, output_11_8, output_10_167;
mixer gate_output_10_167(.a(output_11_167), .b(output_11_8), .y(output_10_167));
wire output_12_167, output_12_8, output_11_167;
mixer gate_output_11_167(.a(output_12_167), .b(output_12_8), .y(output_11_167));
wire output_13_167, output_13_8, output_12_167;
mixer gate_output_12_167(.a(output_13_167), .b(output_13_8), .y(output_12_167));
wire output_14_167, output_14_8, output_13_167;
mixer gate_output_13_167(.a(output_14_167), .b(output_14_8), .y(output_13_167));
wire output_15_167, output_15_8, output_14_167;
mixer gate_output_14_167(.a(output_15_167), .b(output_15_8), .y(output_14_167));
wire output_16_167, output_16_8, output_15_167;
mixer gate_output_15_167(.a(output_16_167), .b(output_16_8), .y(output_15_167));
wire output_1_168, output_1_9, output_0_168;
mixer gate_output_0_168(.a(output_1_168), .b(output_1_9), .y(output_0_168));
wire output_2_168, output_2_9, output_1_168;
mixer gate_output_1_168(.a(output_2_168), .b(output_2_9), .y(output_1_168));
wire output_3_168, output_3_9, output_2_168;
mixer gate_output_2_168(.a(output_3_168), .b(output_3_9), .y(output_2_168));
wire output_4_168, output_4_9, output_3_168;
mixer gate_output_3_168(.a(output_4_168), .b(output_4_9), .y(output_3_168));
wire output_5_168, output_5_9, output_4_168;
mixer gate_output_4_168(.a(output_5_168), .b(output_5_9), .y(output_4_168));
wire output_6_168, output_6_9, output_5_168;
mixer gate_output_5_168(.a(output_6_168), .b(output_6_9), .y(output_5_168));
wire output_7_168, output_7_9, output_6_168;
mixer gate_output_6_168(.a(output_7_168), .b(output_7_9), .y(output_6_168));
wire output_8_168, output_8_9, output_7_168;
mixer gate_output_7_168(.a(output_8_168), .b(output_8_9), .y(output_7_168));
wire output_9_168, output_9_9, output_8_168;
mixer gate_output_8_168(.a(output_9_168), .b(output_9_9), .y(output_8_168));
wire output_10_168, output_10_9, output_9_168;
mixer gate_output_9_168(.a(output_10_168), .b(output_10_9), .y(output_9_168));
wire output_11_168, output_11_9, output_10_168;
mixer gate_output_10_168(.a(output_11_168), .b(output_11_9), .y(output_10_168));
wire output_12_168, output_12_9, output_11_168;
mixer gate_output_11_168(.a(output_12_168), .b(output_12_9), .y(output_11_168));
wire output_13_168, output_13_9, output_12_168;
mixer gate_output_12_168(.a(output_13_168), .b(output_13_9), .y(output_12_168));
wire output_14_168, output_14_9, output_13_168;
mixer gate_output_13_168(.a(output_14_168), .b(output_14_9), .y(output_13_168));
wire output_15_168, output_15_9, output_14_168;
mixer gate_output_14_168(.a(output_15_168), .b(output_15_9), .y(output_14_168));
wire output_16_168, output_16_9, output_15_168;
mixer gate_output_15_168(.a(output_16_168), .b(output_16_9), .y(output_15_168));
wire output_1_169, output_1_10, output_0_169;
mixer gate_output_0_169(.a(output_1_169), .b(output_1_10), .y(output_0_169));
wire output_2_169, output_2_10, output_1_169;
mixer gate_output_1_169(.a(output_2_169), .b(output_2_10), .y(output_1_169));
wire output_3_169, output_3_10, output_2_169;
mixer gate_output_2_169(.a(output_3_169), .b(output_3_10), .y(output_2_169));
wire output_4_169, output_4_10, output_3_169;
mixer gate_output_3_169(.a(output_4_169), .b(output_4_10), .y(output_3_169));
wire output_5_169, output_5_10, output_4_169;
mixer gate_output_4_169(.a(output_5_169), .b(output_5_10), .y(output_4_169));
wire output_6_169, output_6_10, output_5_169;
mixer gate_output_5_169(.a(output_6_169), .b(output_6_10), .y(output_5_169));
wire output_7_169, output_7_10, output_6_169;
mixer gate_output_6_169(.a(output_7_169), .b(output_7_10), .y(output_6_169));
wire output_8_169, output_8_10, output_7_169;
mixer gate_output_7_169(.a(output_8_169), .b(output_8_10), .y(output_7_169));
wire output_9_169, output_9_10, output_8_169;
mixer gate_output_8_169(.a(output_9_169), .b(output_9_10), .y(output_8_169));
wire output_10_169, output_10_10, output_9_169;
mixer gate_output_9_169(.a(output_10_169), .b(output_10_10), .y(output_9_169));
wire output_11_169, output_11_10, output_10_169;
mixer gate_output_10_169(.a(output_11_169), .b(output_11_10), .y(output_10_169));
wire output_12_169, output_12_10, output_11_169;
mixer gate_output_11_169(.a(output_12_169), .b(output_12_10), .y(output_11_169));
wire output_13_169, output_13_10, output_12_169;
mixer gate_output_12_169(.a(output_13_169), .b(output_13_10), .y(output_12_169));
wire output_14_169, output_14_10, output_13_169;
mixer gate_output_13_169(.a(output_14_169), .b(output_14_10), .y(output_13_169));
wire output_15_169, output_15_10, output_14_169;
mixer gate_output_14_169(.a(output_15_169), .b(output_15_10), .y(output_14_169));
wire output_16_169, output_16_10, output_15_169;
mixer gate_output_15_169(.a(output_16_169), .b(output_16_10), .y(output_15_169));
wire output_1_170, output_1_11, output_0_170;
mixer gate_output_0_170(.a(output_1_170), .b(output_1_11), .y(output_0_170));
wire output_2_170, output_2_11, output_1_170;
mixer gate_output_1_170(.a(output_2_170), .b(output_2_11), .y(output_1_170));
wire output_3_170, output_3_11, output_2_170;
mixer gate_output_2_170(.a(output_3_170), .b(output_3_11), .y(output_2_170));
wire output_4_170, output_4_11, output_3_170;
mixer gate_output_3_170(.a(output_4_170), .b(output_4_11), .y(output_3_170));
wire output_5_170, output_5_11, output_4_170;
mixer gate_output_4_170(.a(output_5_170), .b(output_5_11), .y(output_4_170));
wire output_6_170, output_6_11, output_5_170;
mixer gate_output_5_170(.a(output_6_170), .b(output_6_11), .y(output_5_170));
wire output_7_170, output_7_11, output_6_170;
mixer gate_output_6_170(.a(output_7_170), .b(output_7_11), .y(output_6_170));
wire output_8_170, output_8_11, output_7_170;
mixer gate_output_7_170(.a(output_8_170), .b(output_8_11), .y(output_7_170));
wire output_9_170, output_9_11, output_8_170;
mixer gate_output_8_170(.a(output_9_170), .b(output_9_11), .y(output_8_170));
wire output_10_170, output_10_11, output_9_170;
mixer gate_output_9_170(.a(output_10_170), .b(output_10_11), .y(output_9_170));
wire output_11_170, output_11_11, output_10_170;
mixer gate_output_10_170(.a(output_11_170), .b(output_11_11), .y(output_10_170));
wire output_12_170, output_12_11, output_11_170;
mixer gate_output_11_170(.a(output_12_170), .b(output_12_11), .y(output_11_170));
wire output_13_170, output_13_11, output_12_170;
mixer gate_output_12_170(.a(output_13_170), .b(output_13_11), .y(output_12_170));
wire output_14_170, output_14_11, output_13_170;
mixer gate_output_13_170(.a(output_14_170), .b(output_14_11), .y(output_13_170));
wire output_15_170, output_15_11, output_14_170;
mixer gate_output_14_170(.a(output_15_170), .b(output_15_11), .y(output_14_170));
wire output_16_170, output_16_11, output_15_170;
mixer gate_output_15_170(.a(output_16_170), .b(output_16_11), .y(output_15_170));
wire output_1_171, output_1_12, output_0_171;
mixer gate_output_0_171(.a(output_1_171), .b(output_1_12), .y(output_0_171));
wire output_2_171, output_2_12, output_1_171;
mixer gate_output_1_171(.a(output_2_171), .b(output_2_12), .y(output_1_171));
wire output_3_171, output_3_12, output_2_171;
mixer gate_output_2_171(.a(output_3_171), .b(output_3_12), .y(output_2_171));
wire output_4_171, output_4_12, output_3_171;
mixer gate_output_3_171(.a(output_4_171), .b(output_4_12), .y(output_3_171));
wire output_5_171, output_5_12, output_4_171;
mixer gate_output_4_171(.a(output_5_171), .b(output_5_12), .y(output_4_171));
wire output_6_171, output_6_12, output_5_171;
mixer gate_output_5_171(.a(output_6_171), .b(output_6_12), .y(output_5_171));
wire output_7_171, output_7_12, output_6_171;
mixer gate_output_6_171(.a(output_7_171), .b(output_7_12), .y(output_6_171));
wire output_8_171, output_8_12, output_7_171;
mixer gate_output_7_171(.a(output_8_171), .b(output_8_12), .y(output_7_171));
wire output_9_171, output_9_12, output_8_171;
mixer gate_output_8_171(.a(output_9_171), .b(output_9_12), .y(output_8_171));
wire output_10_171, output_10_12, output_9_171;
mixer gate_output_9_171(.a(output_10_171), .b(output_10_12), .y(output_9_171));
wire output_11_171, output_11_12, output_10_171;
mixer gate_output_10_171(.a(output_11_171), .b(output_11_12), .y(output_10_171));
wire output_12_171, output_12_12, output_11_171;
mixer gate_output_11_171(.a(output_12_171), .b(output_12_12), .y(output_11_171));
wire output_13_171, output_13_12, output_12_171;
mixer gate_output_12_171(.a(output_13_171), .b(output_13_12), .y(output_12_171));
wire output_14_171, output_14_12, output_13_171;
mixer gate_output_13_171(.a(output_14_171), .b(output_14_12), .y(output_13_171));
wire output_15_171, output_15_12, output_14_171;
mixer gate_output_14_171(.a(output_15_171), .b(output_15_12), .y(output_14_171));
wire output_16_171, output_16_12, output_15_171;
mixer gate_output_15_171(.a(output_16_171), .b(output_16_12), .y(output_15_171));
wire output_1_172, output_1_13, output_0_172;
mixer gate_output_0_172(.a(output_1_172), .b(output_1_13), .y(output_0_172));
wire output_2_172, output_2_13, output_1_172;
mixer gate_output_1_172(.a(output_2_172), .b(output_2_13), .y(output_1_172));
wire output_3_172, output_3_13, output_2_172;
mixer gate_output_2_172(.a(output_3_172), .b(output_3_13), .y(output_2_172));
wire output_4_172, output_4_13, output_3_172;
mixer gate_output_3_172(.a(output_4_172), .b(output_4_13), .y(output_3_172));
wire output_5_172, output_5_13, output_4_172;
mixer gate_output_4_172(.a(output_5_172), .b(output_5_13), .y(output_4_172));
wire output_6_172, output_6_13, output_5_172;
mixer gate_output_5_172(.a(output_6_172), .b(output_6_13), .y(output_5_172));
wire output_7_172, output_7_13, output_6_172;
mixer gate_output_6_172(.a(output_7_172), .b(output_7_13), .y(output_6_172));
wire output_8_172, output_8_13, output_7_172;
mixer gate_output_7_172(.a(output_8_172), .b(output_8_13), .y(output_7_172));
wire output_9_172, output_9_13, output_8_172;
mixer gate_output_8_172(.a(output_9_172), .b(output_9_13), .y(output_8_172));
wire output_10_172, output_10_13, output_9_172;
mixer gate_output_9_172(.a(output_10_172), .b(output_10_13), .y(output_9_172));
wire output_11_172, output_11_13, output_10_172;
mixer gate_output_10_172(.a(output_11_172), .b(output_11_13), .y(output_10_172));
wire output_12_172, output_12_13, output_11_172;
mixer gate_output_11_172(.a(output_12_172), .b(output_12_13), .y(output_11_172));
wire output_13_172, output_13_13, output_12_172;
mixer gate_output_12_172(.a(output_13_172), .b(output_13_13), .y(output_12_172));
wire output_14_172, output_14_13, output_13_172;
mixer gate_output_13_172(.a(output_14_172), .b(output_14_13), .y(output_13_172));
wire output_15_172, output_15_13, output_14_172;
mixer gate_output_14_172(.a(output_15_172), .b(output_15_13), .y(output_14_172));
wire output_16_172, output_16_13, output_15_172;
mixer gate_output_15_172(.a(output_16_172), .b(output_16_13), .y(output_15_172));
wire output_1_173, output_1_14, output_0_173;
mixer gate_output_0_173(.a(output_1_173), .b(output_1_14), .y(output_0_173));
wire output_2_173, output_2_14, output_1_173;
mixer gate_output_1_173(.a(output_2_173), .b(output_2_14), .y(output_1_173));
wire output_3_173, output_3_14, output_2_173;
mixer gate_output_2_173(.a(output_3_173), .b(output_3_14), .y(output_2_173));
wire output_4_173, output_4_14, output_3_173;
mixer gate_output_3_173(.a(output_4_173), .b(output_4_14), .y(output_3_173));
wire output_5_173, output_5_14, output_4_173;
mixer gate_output_4_173(.a(output_5_173), .b(output_5_14), .y(output_4_173));
wire output_6_173, output_6_14, output_5_173;
mixer gate_output_5_173(.a(output_6_173), .b(output_6_14), .y(output_5_173));
wire output_7_173, output_7_14, output_6_173;
mixer gate_output_6_173(.a(output_7_173), .b(output_7_14), .y(output_6_173));
wire output_8_173, output_8_14, output_7_173;
mixer gate_output_7_173(.a(output_8_173), .b(output_8_14), .y(output_7_173));
wire output_9_173, output_9_14, output_8_173;
mixer gate_output_8_173(.a(output_9_173), .b(output_9_14), .y(output_8_173));
wire output_10_173, output_10_14, output_9_173;
mixer gate_output_9_173(.a(output_10_173), .b(output_10_14), .y(output_9_173));
wire output_11_173, output_11_14, output_10_173;
mixer gate_output_10_173(.a(output_11_173), .b(output_11_14), .y(output_10_173));
wire output_12_173, output_12_14, output_11_173;
mixer gate_output_11_173(.a(output_12_173), .b(output_12_14), .y(output_11_173));
wire output_13_173, output_13_14, output_12_173;
mixer gate_output_12_173(.a(output_13_173), .b(output_13_14), .y(output_12_173));
wire output_14_173, output_14_14, output_13_173;
mixer gate_output_13_173(.a(output_14_173), .b(output_14_14), .y(output_13_173));
wire output_15_173, output_15_14, output_14_173;
mixer gate_output_14_173(.a(output_15_173), .b(output_15_14), .y(output_14_173));
wire output_16_173, output_16_14, output_15_173;
mixer gate_output_15_173(.a(output_16_173), .b(output_16_14), .y(output_15_173));
wire output_1_174, output_1_15, output_0_174;
mixer gate_output_0_174(.a(output_1_174), .b(output_1_15), .y(output_0_174));
wire output_2_174, output_2_15, output_1_174;
mixer gate_output_1_174(.a(output_2_174), .b(output_2_15), .y(output_1_174));
wire output_3_174, output_3_15, output_2_174;
mixer gate_output_2_174(.a(output_3_174), .b(output_3_15), .y(output_2_174));
wire output_4_174, output_4_15, output_3_174;
mixer gate_output_3_174(.a(output_4_174), .b(output_4_15), .y(output_3_174));
wire output_5_174, output_5_15, output_4_174;
mixer gate_output_4_174(.a(output_5_174), .b(output_5_15), .y(output_4_174));
wire output_6_174, output_6_15, output_5_174;
mixer gate_output_5_174(.a(output_6_174), .b(output_6_15), .y(output_5_174));
wire output_7_174, output_7_15, output_6_174;
mixer gate_output_6_174(.a(output_7_174), .b(output_7_15), .y(output_6_174));
wire output_8_174, output_8_15, output_7_174;
mixer gate_output_7_174(.a(output_8_174), .b(output_8_15), .y(output_7_174));
wire output_9_174, output_9_15, output_8_174;
mixer gate_output_8_174(.a(output_9_174), .b(output_9_15), .y(output_8_174));
wire output_10_174, output_10_15, output_9_174;
mixer gate_output_9_174(.a(output_10_174), .b(output_10_15), .y(output_9_174));
wire output_11_174, output_11_15, output_10_174;
mixer gate_output_10_174(.a(output_11_174), .b(output_11_15), .y(output_10_174));
wire output_12_174, output_12_15, output_11_174;
mixer gate_output_11_174(.a(output_12_174), .b(output_12_15), .y(output_11_174));
wire output_13_174, output_13_15, output_12_174;
mixer gate_output_12_174(.a(output_13_174), .b(output_13_15), .y(output_12_174));
wire output_14_174, output_14_15, output_13_174;
mixer gate_output_13_174(.a(output_14_174), .b(output_14_15), .y(output_13_174));
wire output_15_174, output_15_15, output_14_174;
mixer gate_output_14_174(.a(output_15_174), .b(output_15_15), .y(output_14_174));
wire output_16_174, output_16_15, output_15_174;
mixer gate_output_15_174(.a(output_16_174), .b(output_16_15), .y(output_15_174));
wire output_1_175, output_1_0, output_0_175;
mixer gate_output_0_175(.a(output_1_175), .b(output_1_0), .y(output_0_175));
wire output_2_175, output_2_0, output_1_175;
mixer gate_output_1_175(.a(output_2_175), .b(output_2_0), .y(output_1_175));
wire output_3_175, output_3_0, output_2_175;
mixer gate_output_2_175(.a(output_3_175), .b(output_3_0), .y(output_2_175));
wire output_4_175, output_4_0, output_3_175;
mixer gate_output_3_175(.a(output_4_175), .b(output_4_0), .y(output_3_175));
wire output_5_175, output_5_0, output_4_175;
mixer gate_output_4_175(.a(output_5_175), .b(output_5_0), .y(output_4_175));
wire output_6_175, output_6_0, output_5_175;
mixer gate_output_5_175(.a(output_6_175), .b(output_6_0), .y(output_5_175));
wire output_7_175, output_7_0, output_6_175;
mixer gate_output_6_175(.a(output_7_175), .b(output_7_0), .y(output_6_175));
wire output_8_175, output_8_0, output_7_175;
mixer gate_output_7_175(.a(output_8_175), .b(output_8_0), .y(output_7_175));
wire output_9_175, output_9_0, output_8_175;
mixer gate_output_8_175(.a(output_9_175), .b(output_9_0), .y(output_8_175));
wire output_10_175, output_10_0, output_9_175;
mixer gate_output_9_175(.a(output_10_175), .b(output_10_0), .y(output_9_175));
wire output_11_175, output_11_0, output_10_175;
mixer gate_output_10_175(.a(output_11_175), .b(output_11_0), .y(output_10_175));
wire output_12_175, output_12_0, output_11_175;
mixer gate_output_11_175(.a(output_12_175), .b(output_12_0), .y(output_11_175));
wire output_13_175, output_13_0, output_12_175;
mixer gate_output_12_175(.a(output_13_175), .b(output_13_0), .y(output_12_175));
wire output_14_175, output_14_0, output_13_175;
mixer gate_output_13_175(.a(output_14_175), .b(output_14_0), .y(output_13_175));
wire output_15_175, output_15_0, output_14_175;
mixer gate_output_14_175(.a(output_15_175), .b(output_15_0), .y(output_14_175));
wire output_16_175, output_16_0, output_15_175;
mixer gate_output_15_175(.a(output_16_175), .b(output_16_0), .y(output_15_175));
wire output_1_176, output_1_1, output_0_176;
mixer gate_output_0_176(.a(output_1_176), .b(output_1_1), .y(output_0_176));
wire output_2_176, output_2_1, output_1_176;
mixer gate_output_1_176(.a(output_2_176), .b(output_2_1), .y(output_1_176));
wire output_3_176, output_3_1, output_2_176;
mixer gate_output_2_176(.a(output_3_176), .b(output_3_1), .y(output_2_176));
wire output_4_176, output_4_1, output_3_176;
mixer gate_output_3_176(.a(output_4_176), .b(output_4_1), .y(output_3_176));
wire output_5_176, output_5_1, output_4_176;
mixer gate_output_4_176(.a(output_5_176), .b(output_5_1), .y(output_4_176));
wire output_6_176, output_6_1, output_5_176;
mixer gate_output_5_176(.a(output_6_176), .b(output_6_1), .y(output_5_176));
wire output_7_176, output_7_1, output_6_176;
mixer gate_output_6_176(.a(output_7_176), .b(output_7_1), .y(output_6_176));
wire output_8_176, output_8_1, output_7_176;
mixer gate_output_7_176(.a(output_8_176), .b(output_8_1), .y(output_7_176));
wire output_9_176, output_9_1, output_8_176;
mixer gate_output_8_176(.a(output_9_176), .b(output_9_1), .y(output_8_176));
wire output_10_176, output_10_1, output_9_176;
mixer gate_output_9_176(.a(output_10_176), .b(output_10_1), .y(output_9_176));
wire output_11_176, output_11_1, output_10_176;
mixer gate_output_10_176(.a(output_11_176), .b(output_11_1), .y(output_10_176));
wire output_12_176, output_12_1, output_11_176;
mixer gate_output_11_176(.a(output_12_176), .b(output_12_1), .y(output_11_176));
wire output_13_176, output_13_1, output_12_176;
mixer gate_output_12_176(.a(output_13_176), .b(output_13_1), .y(output_12_176));
wire output_14_176, output_14_1, output_13_176;
mixer gate_output_13_176(.a(output_14_176), .b(output_14_1), .y(output_13_176));
wire output_15_176, output_15_1, output_14_176;
mixer gate_output_14_176(.a(output_15_176), .b(output_15_1), .y(output_14_176));
wire output_16_176, output_16_1, output_15_176;
mixer gate_output_15_176(.a(output_16_176), .b(output_16_1), .y(output_15_176));
wire output_1_177, output_1_2, output_0_177;
mixer gate_output_0_177(.a(output_1_177), .b(output_1_2), .y(output_0_177));
wire output_2_177, output_2_2, output_1_177;
mixer gate_output_1_177(.a(output_2_177), .b(output_2_2), .y(output_1_177));
wire output_3_177, output_3_2, output_2_177;
mixer gate_output_2_177(.a(output_3_177), .b(output_3_2), .y(output_2_177));
wire output_4_177, output_4_2, output_3_177;
mixer gate_output_3_177(.a(output_4_177), .b(output_4_2), .y(output_3_177));
wire output_5_177, output_5_2, output_4_177;
mixer gate_output_4_177(.a(output_5_177), .b(output_5_2), .y(output_4_177));
wire output_6_177, output_6_2, output_5_177;
mixer gate_output_5_177(.a(output_6_177), .b(output_6_2), .y(output_5_177));
wire output_7_177, output_7_2, output_6_177;
mixer gate_output_6_177(.a(output_7_177), .b(output_7_2), .y(output_6_177));
wire output_8_177, output_8_2, output_7_177;
mixer gate_output_7_177(.a(output_8_177), .b(output_8_2), .y(output_7_177));
wire output_9_177, output_9_2, output_8_177;
mixer gate_output_8_177(.a(output_9_177), .b(output_9_2), .y(output_8_177));
wire output_10_177, output_10_2, output_9_177;
mixer gate_output_9_177(.a(output_10_177), .b(output_10_2), .y(output_9_177));
wire output_11_177, output_11_2, output_10_177;
mixer gate_output_10_177(.a(output_11_177), .b(output_11_2), .y(output_10_177));
wire output_12_177, output_12_2, output_11_177;
mixer gate_output_11_177(.a(output_12_177), .b(output_12_2), .y(output_11_177));
wire output_13_177, output_13_2, output_12_177;
mixer gate_output_12_177(.a(output_13_177), .b(output_13_2), .y(output_12_177));
wire output_14_177, output_14_2, output_13_177;
mixer gate_output_13_177(.a(output_14_177), .b(output_14_2), .y(output_13_177));
wire output_15_177, output_15_2, output_14_177;
mixer gate_output_14_177(.a(output_15_177), .b(output_15_2), .y(output_14_177));
wire output_16_177, output_16_2, output_15_177;
mixer gate_output_15_177(.a(output_16_177), .b(output_16_2), .y(output_15_177));
wire output_1_178, output_1_3, output_0_178;
mixer gate_output_0_178(.a(output_1_178), .b(output_1_3), .y(output_0_178));
wire output_2_178, output_2_3, output_1_178;
mixer gate_output_1_178(.a(output_2_178), .b(output_2_3), .y(output_1_178));
wire output_3_178, output_3_3, output_2_178;
mixer gate_output_2_178(.a(output_3_178), .b(output_3_3), .y(output_2_178));
wire output_4_178, output_4_3, output_3_178;
mixer gate_output_3_178(.a(output_4_178), .b(output_4_3), .y(output_3_178));
wire output_5_178, output_5_3, output_4_178;
mixer gate_output_4_178(.a(output_5_178), .b(output_5_3), .y(output_4_178));
wire output_6_178, output_6_3, output_5_178;
mixer gate_output_5_178(.a(output_6_178), .b(output_6_3), .y(output_5_178));
wire output_7_178, output_7_3, output_6_178;
mixer gate_output_6_178(.a(output_7_178), .b(output_7_3), .y(output_6_178));
wire output_8_178, output_8_3, output_7_178;
mixer gate_output_7_178(.a(output_8_178), .b(output_8_3), .y(output_7_178));
wire output_9_178, output_9_3, output_8_178;
mixer gate_output_8_178(.a(output_9_178), .b(output_9_3), .y(output_8_178));
wire output_10_178, output_10_3, output_9_178;
mixer gate_output_9_178(.a(output_10_178), .b(output_10_3), .y(output_9_178));
wire output_11_178, output_11_3, output_10_178;
mixer gate_output_10_178(.a(output_11_178), .b(output_11_3), .y(output_10_178));
wire output_12_178, output_12_3, output_11_178;
mixer gate_output_11_178(.a(output_12_178), .b(output_12_3), .y(output_11_178));
wire output_13_178, output_13_3, output_12_178;
mixer gate_output_12_178(.a(output_13_178), .b(output_13_3), .y(output_12_178));
wire output_14_178, output_14_3, output_13_178;
mixer gate_output_13_178(.a(output_14_178), .b(output_14_3), .y(output_13_178));
wire output_15_178, output_15_3, output_14_178;
mixer gate_output_14_178(.a(output_15_178), .b(output_15_3), .y(output_14_178));
wire output_16_178, output_16_3, output_15_178;
mixer gate_output_15_178(.a(output_16_178), .b(output_16_3), .y(output_15_178));
wire output_1_179, output_1_4, output_0_179;
mixer gate_output_0_179(.a(output_1_179), .b(output_1_4), .y(output_0_179));
wire output_2_179, output_2_4, output_1_179;
mixer gate_output_1_179(.a(output_2_179), .b(output_2_4), .y(output_1_179));
wire output_3_179, output_3_4, output_2_179;
mixer gate_output_2_179(.a(output_3_179), .b(output_3_4), .y(output_2_179));
wire output_4_179, output_4_4, output_3_179;
mixer gate_output_3_179(.a(output_4_179), .b(output_4_4), .y(output_3_179));
wire output_5_179, output_5_4, output_4_179;
mixer gate_output_4_179(.a(output_5_179), .b(output_5_4), .y(output_4_179));
wire output_6_179, output_6_4, output_5_179;
mixer gate_output_5_179(.a(output_6_179), .b(output_6_4), .y(output_5_179));
wire output_7_179, output_7_4, output_6_179;
mixer gate_output_6_179(.a(output_7_179), .b(output_7_4), .y(output_6_179));
wire output_8_179, output_8_4, output_7_179;
mixer gate_output_7_179(.a(output_8_179), .b(output_8_4), .y(output_7_179));
wire output_9_179, output_9_4, output_8_179;
mixer gate_output_8_179(.a(output_9_179), .b(output_9_4), .y(output_8_179));
wire output_10_179, output_10_4, output_9_179;
mixer gate_output_9_179(.a(output_10_179), .b(output_10_4), .y(output_9_179));
wire output_11_179, output_11_4, output_10_179;
mixer gate_output_10_179(.a(output_11_179), .b(output_11_4), .y(output_10_179));
wire output_12_179, output_12_4, output_11_179;
mixer gate_output_11_179(.a(output_12_179), .b(output_12_4), .y(output_11_179));
wire output_13_179, output_13_4, output_12_179;
mixer gate_output_12_179(.a(output_13_179), .b(output_13_4), .y(output_12_179));
wire output_14_179, output_14_4, output_13_179;
mixer gate_output_13_179(.a(output_14_179), .b(output_14_4), .y(output_13_179));
wire output_15_179, output_15_4, output_14_179;
mixer gate_output_14_179(.a(output_15_179), .b(output_15_4), .y(output_14_179));
wire output_16_179, output_16_4, output_15_179;
mixer gate_output_15_179(.a(output_16_179), .b(output_16_4), .y(output_15_179));
wire output_1_180, output_1_5, output_0_180;
mixer gate_output_0_180(.a(output_1_180), .b(output_1_5), .y(output_0_180));
wire output_2_180, output_2_5, output_1_180;
mixer gate_output_1_180(.a(output_2_180), .b(output_2_5), .y(output_1_180));
wire output_3_180, output_3_5, output_2_180;
mixer gate_output_2_180(.a(output_3_180), .b(output_3_5), .y(output_2_180));
wire output_4_180, output_4_5, output_3_180;
mixer gate_output_3_180(.a(output_4_180), .b(output_4_5), .y(output_3_180));
wire output_5_180, output_5_5, output_4_180;
mixer gate_output_4_180(.a(output_5_180), .b(output_5_5), .y(output_4_180));
wire output_6_180, output_6_5, output_5_180;
mixer gate_output_5_180(.a(output_6_180), .b(output_6_5), .y(output_5_180));
wire output_7_180, output_7_5, output_6_180;
mixer gate_output_6_180(.a(output_7_180), .b(output_7_5), .y(output_6_180));
wire output_8_180, output_8_5, output_7_180;
mixer gate_output_7_180(.a(output_8_180), .b(output_8_5), .y(output_7_180));
wire output_9_180, output_9_5, output_8_180;
mixer gate_output_8_180(.a(output_9_180), .b(output_9_5), .y(output_8_180));
wire output_10_180, output_10_5, output_9_180;
mixer gate_output_9_180(.a(output_10_180), .b(output_10_5), .y(output_9_180));
wire output_11_180, output_11_5, output_10_180;
mixer gate_output_10_180(.a(output_11_180), .b(output_11_5), .y(output_10_180));
wire output_12_180, output_12_5, output_11_180;
mixer gate_output_11_180(.a(output_12_180), .b(output_12_5), .y(output_11_180));
wire output_13_180, output_13_5, output_12_180;
mixer gate_output_12_180(.a(output_13_180), .b(output_13_5), .y(output_12_180));
wire output_14_180, output_14_5, output_13_180;
mixer gate_output_13_180(.a(output_14_180), .b(output_14_5), .y(output_13_180));
wire output_15_180, output_15_5, output_14_180;
mixer gate_output_14_180(.a(output_15_180), .b(output_15_5), .y(output_14_180));
wire output_16_180, output_16_5, output_15_180;
mixer gate_output_15_180(.a(output_16_180), .b(output_16_5), .y(output_15_180));
wire output_1_181, output_1_6, output_0_181;
mixer gate_output_0_181(.a(output_1_181), .b(output_1_6), .y(output_0_181));
wire output_2_181, output_2_6, output_1_181;
mixer gate_output_1_181(.a(output_2_181), .b(output_2_6), .y(output_1_181));
wire output_3_181, output_3_6, output_2_181;
mixer gate_output_2_181(.a(output_3_181), .b(output_3_6), .y(output_2_181));
wire output_4_181, output_4_6, output_3_181;
mixer gate_output_3_181(.a(output_4_181), .b(output_4_6), .y(output_3_181));
wire output_5_181, output_5_6, output_4_181;
mixer gate_output_4_181(.a(output_5_181), .b(output_5_6), .y(output_4_181));
wire output_6_181, output_6_6, output_5_181;
mixer gate_output_5_181(.a(output_6_181), .b(output_6_6), .y(output_5_181));
wire output_7_181, output_7_6, output_6_181;
mixer gate_output_6_181(.a(output_7_181), .b(output_7_6), .y(output_6_181));
wire output_8_181, output_8_6, output_7_181;
mixer gate_output_7_181(.a(output_8_181), .b(output_8_6), .y(output_7_181));
wire output_9_181, output_9_6, output_8_181;
mixer gate_output_8_181(.a(output_9_181), .b(output_9_6), .y(output_8_181));
wire output_10_181, output_10_6, output_9_181;
mixer gate_output_9_181(.a(output_10_181), .b(output_10_6), .y(output_9_181));
wire output_11_181, output_11_6, output_10_181;
mixer gate_output_10_181(.a(output_11_181), .b(output_11_6), .y(output_10_181));
wire output_12_181, output_12_6, output_11_181;
mixer gate_output_11_181(.a(output_12_181), .b(output_12_6), .y(output_11_181));
wire output_13_181, output_13_6, output_12_181;
mixer gate_output_12_181(.a(output_13_181), .b(output_13_6), .y(output_12_181));
wire output_14_181, output_14_6, output_13_181;
mixer gate_output_13_181(.a(output_14_181), .b(output_14_6), .y(output_13_181));
wire output_15_181, output_15_6, output_14_181;
mixer gate_output_14_181(.a(output_15_181), .b(output_15_6), .y(output_14_181));
wire output_16_181, output_16_6, output_15_181;
mixer gate_output_15_181(.a(output_16_181), .b(output_16_6), .y(output_15_181));
wire output_1_182, output_1_7, output_0_182;
mixer gate_output_0_182(.a(output_1_182), .b(output_1_7), .y(output_0_182));
wire output_2_182, output_2_7, output_1_182;
mixer gate_output_1_182(.a(output_2_182), .b(output_2_7), .y(output_1_182));
wire output_3_182, output_3_7, output_2_182;
mixer gate_output_2_182(.a(output_3_182), .b(output_3_7), .y(output_2_182));
wire output_4_182, output_4_7, output_3_182;
mixer gate_output_3_182(.a(output_4_182), .b(output_4_7), .y(output_3_182));
wire output_5_182, output_5_7, output_4_182;
mixer gate_output_4_182(.a(output_5_182), .b(output_5_7), .y(output_4_182));
wire output_6_182, output_6_7, output_5_182;
mixer gate_output_5_182(.a(output_6_182), .b(output_6_7), .y(output_5_182));
wire output_7_182, output_7_7, output_6_182;
mixer gate_output_6_182(.a(output_7_182), .b(output_7_7), .y(output_6_182));
wire output_8_182, output_8_7, output_7_182;
mixer gate_output_7_182(.a(output_8_182), .b(output_8_7), .y(output_7_182));
wire output_9_182, output_9_7, output_8_182;
mixer gate_output_8_182(.a(output_9_182), .b(output_9_7), .y(output_8_182));
wire output_10_182, output_10_7, output_9_182;
mixer gate_output_9_182(.a(output_10_182), .b(output_10_7), .y(output_9_182));
wire output_11_182, output_11_7, output_10_182;
mixer gate_output_10_182(.a(output_11_182), .b(output_11_7), .y(output_10_182));
wire output_12_182, output_12_7, output_11_182;
mixer gate_output_11_182(.a(output_12_182), .b(output_12_7), .y(output_11_182));
wire output_13_182, output_13_7, output_12_182;
mixer gate_output_12_182(.a(output_13_182), .b(output_13_7), .y(output_12_182));
wire output_14_182, output_14_7, output_13_182;
mixer gate_output_13_182(.a(output_14_182), .b(output_14_7), .y(output_13_182));
wire output_15_182, output_15_7, output_14_182;
mixer gate_output_14_182(.a(output_15_182), .b(output_15_7), .y(output_14_182));
wire output_16_182, output_16_7, output_15_182;
mixer gate_output_15_182(.a(output_16_182), .b(output_16_7), .y(output_15_182));
wire output_1_183, output_1_8, output_0_183;
mixer gate_output_0_183(.a(output_1_183), .b(output_1_8), .y(output_0_183));
wire output_2_183, output_2_8, output_1_183;
mixer gate_output_1_183(.a(output_2_183), .b(output_2_8), .y(output_1_183));
wire output_3_183, output_3_8, output_2_183;
mixer gate_output_2_183(.a(output_3_183), .b(output_3_8), .y(output_2_183));
wire output_4_183, output_4_8, output_3_183;
mixer gate_output_3_183(.a(output_4_183), .b(output_4_8), .y(output_3_183));
wire output_5_183, output_5_8, output_4_183;
mixer gate_output_4_183(.a(output_5_183), .b(output_5_8), .y(output_4_183));
wire output_6_183, output_6_8, output_5_183;
mixer gate_output_5_183(.a(output_6_183), .b(output_6_8), .y(output_5_183));
wire output_7_183, output_7_8, output_6_183;
mixer gate_output_6_183(.a(output_7_183), .b(output_7_8), .y(output_6_183));
wire output_8_183, output_8_8, output_7_183;
mixer gate_output_7_183(.a(output_8_183), .b(output_8_8), .y(output_7_183));
wire output_9_183, output_9_8, output_8_183;
mixer gate_output_8_183(.a(output_9_183), .b(output_9_8), .y(output_8_183));
wire output_10_183, output_10_8, output_9_183;
mixer gate_output_9_183(.a(output_10_183), .b(output_10_8), .y(output_9_183));
wire output_11_183, output_11_8, output_10_183;
mixer gate_output_10_183(.a(output_11_183), .b(output_11_8), .y(output_10_183));
wire output_12_183, output_12_8, output_11_183;
mixer gate_output_11_183(.a(output_12_183), .b(output_12_8), .y(output_11_183));
wire output_13_183, output_13_8, output_12_183;
mixer gate_output_12_183(.a(output_13_183), .b(output_13_8), .y(output_12_183));
wire output_14_183, output_14_8, output_13_183;
mixer gate_output_13_183(.a(output_14_183), .b(output_14_8), .y(output_13_183));
wire output_15_183, output_15_8, output_14_183;
mixer gate_output_14_183(.a(output_15_183), .b(output_15_8), .y(output_14_183));
wire output_16_183, output_16_8, output_15_183;
mixer gate_output_15_183(.a(output_16_183), .b(output_16_8), .y(output_15_183));
wire output_1_184, output_1_9, output_0_184;
mixer gate_output_0_184(.a(output_1_184), .b(output_1_9), .y(output_0_184));
wire output_2_184, output_2_9, output_1_184;
mixer gate_output_1_184(.a(output_2_184), .b(output_2_9), .y(output_1_184));
wire output_3_184, output_3_9, output_2_184;
mixer gate_output_2_184(.a(output_3_184), .b(output_3_9), .y(output_2_184));
wire output_4_184, output_4_9, output_3_184;
mixer gate_output_3_184(.a(output_4_184), .b(output_4_9), .y(output_3_184));
wire output_5_184, output_5_9, output_4_184;
mixer gate_output_4_184(.a(output_5_184), .b(output_5_9), .y(output_4_184));
wire output_6_184, output_6_9, output_5_184;
mixer gate_output_5_184(.a(output_6_184), .b(output_6_9), .y(output_5_184));
wire output_7_184, output_7_9, output_6_184;
mixer gate_output_6_184(.a(output_7_184), .b(output_7_9), .y(output_6_184));
wire output_8_184, output_8_9, output_7_184;
mixer gate_output_7_184(.a(output_8_184), .b(output_8_9), .y(output_7_184));
wire output_9_184, output_9_9, output_8_184;
mixer gate_output_8_184(.a(output_9_184), .b(output_9_9), .y(output_8_184));
wire output_10_184, output_10_9, output_9_184;
mixer gate_output_9_184(.a(output_10_184), .b(output_10_9), .y(output_9_184));
wire output_11_184, output_11_9, output_10_184;
mixer gate_output_10_184(.a(output_11_184), .b(output_11_9), .y(output_10_184));
wire output_12_184, output_12_9, output_11_184;
mixer gate_output_11_184(.a(output_12_184), .b(output_12_9), .y(output_11_184));
wire output_13_184, output_13_9, output_12_184;
mixer gate_output_12_184(.a(output_13_184), .b(output_13_9), .y(output_12_184));
wire output_14_184, output_14_9, output_13_184;
mixer gate_output_13_184(.a(output_14_184), .b(output_14_9), .y(output_13_184));
wire output_15_184, output_15_9, output_14_184;
mixer gate_output_14_184(.a(output_15_184), .b(output_15_9), .y(output_14_184));
wire output_16_184, output_16_9, output_15_184;
mixer gate_output_15_184(.a(output_16_184), .b(output_16_9), .y(output_15_184));
wire output_1_185, output_1_10, output_0_185;
mixer gate_output_0_185(.a(output_1_185), .b(output_1_10), .y(output_0_185));
wire output_2_185, output_2_10, output_1_185;
mixer gate_output_1_185(.a(output_2_185), .b(output_2_10), .y(output_1_185));
wire output_3_185, output_3_10, output_2_185;
mixer gate_output_2_185(.a(output_3_185), .b(output_3_10), .y(output_2_185));
wire output_4_185, output_4_10, output_3_185;
mixer gate_output_3_185(.a(output_4_185), .b(output_4_10), .y(output_3_185));
wire output_5_185, output_5_10, output_4_185;
mixer gate_output_4_185(.a(output_5_185), .b(output_5_10), .y(output_4_185));
wire output_6_185, output_6_10, output_5_185;
mixer gate_output_5_185(.a(output_6_185), .b(output_6_10), .y(output_5_185));
wire output_7_185, output_7_10, output_6_185;
mixer gate_output_6_185(.a(output_7_185), .b(output_7_10), .y(output_6_185));
wire output_8_185, output_8_10, output_7_185;
mixer gate_output_7_185(.a(output_8_185), .b(output_8_10), .y(output_7_185));
wire output_9_185, output_9_10, output_8_185;
mixer gate_output_8_185(.a(output_9_185), .b(output_9_10), .y(output_8_185));
wire output_10_185, output_10_10, output_9_185;
mixer gate_output_9_185(.a(output_10_185), .b(output_10_10), .y(output_9_185));
wire output_11_185, output_11_10, output_10_185;
mixer gate_output_10_185(.a(output_11_185), .b(output_11_10), .y(output_10_185));
wire output_12_185, output_12_10, output_11_185;
mixer gate_output_11_185(.a(output_12_185), .b(output_12_10), .y(output_11_185));
wire output_13_185, output_13_10, output_12_185;
mixer gate_output_12_185(.a(output_13_185), .b(output_13_10), .y(output_12_185));
wire output_14_185, output_14_10, output_13_185;
mixer gate_output_13_185(.a(output_14_185), .b(output_14_10), .y(output_13_185));
wire output_15_185, output_15_10, output_14_185;
mixer gate_output_14_185(.a(output_15_185), .b(output_15_10), .y(output_14_185));
wire output_16_185, output_16_10, output_15_185;
mixer gate_output_15_185(.a(output_16_185), .b(output_16_10), .y(output_15_185));
wire output_1_186, output_1_11, output_0_186;
mixer gate_output_0_186(.a(output_1_186), .b(output_1_11), .y(output_0_186));
wire output_2_186, output_2_11, output_1_186;
mixer gate_output_1_186(.a(output_2_186), .b(output_2_11), .y(output_1_186));
wire output_3_186, output_3_11, output_2_186;
mixer gate_output_2_186(.a(output_3_186), .b(output_3_11), .y(output_2_186));
wire output_4_186, output_4_11, output_3_186;
mixer gate_output_3_186(.a(output_4_186), .b(output_4_11), .y(output_3_186));
wire output_5_186, output_5_11, output_4_186;
mixer gate_output_4_186(.a(output_5_186), .b(output_5_11), .y(output_4_186));
wire output_6_186, output_6_11, output_5_186;
mixer gate_output_5_186(.a(output_6_186), .b(output_6_11), .y(output_5_186));
wire output_7_186, output_7_11, output_6_186;
mixer gate_output_6_186(.a(output_7_186), .b(output_7_11), .y(output_6_186));
wire output_8_186, output_8_11, output_7_186;
mixer gate_output_7_186(.a(output_8_186), .b(output_8_11), .y(output_7_186));
wire output_9_186, output_9_11, output_8_186;
mixer gate_output_8_186(.a(output_9_186), .b(output_9_11), .y(output_8_186));
wire output_10_186, output_10_11, output_9_186;
mixer gate_output_9_186(.a(output_10_186), .b(output_10_11), .y(output_9_186));
wire output_11_186, output_11_11, output_10_186;
mixer gate_output_10_186(.a(output_11_186), .b(output_11_11), .y(output_10_186));
wire output_12_186, output_12_11, output_11_186;
mixer gate_output_11_186(.a(output_12_186), .b(output_12_11), .y(output_11_186));
wire output_13_186, output_13_11, output_12_186;
mixer gate_output_12_186(.a(output_13_186), .b(output_13_11), .y(output_12_186));
wire output_14_186, output_14_11, output_13_186;
mixer gate_output_13_186(.a(output_14_186), .b(output_14_11), .y(output_13_186));
wire output_15_186, output_15_11, output_14_186;
mixer gate_output_14_186(.a(output_15_186), .b(output_15_11), .y(output_14_186));
wire output_16_186, output_16_11, output_15_186;
mixer gate_output_15_186(.a(output_16_186), .b(output_16_11), .y(output_15_186));
wire output_1_187, output_1_12, output_0_187;
mixer gate_output_0_187(.a(output_1_187), .b(output_1_12), .y(output_0_187));
wire output_2_187, output_2_12, output_1_187;
mixer gate_output_1_187(.a(output_2_187), .b(output_2_12), .y(output_1_187));
wire output_3_187, output_3_12, output_2_187;
mixer gate_output_2_187(.a(output_3_187), .b(output_3_12), .y(output_2_187));
wire output_4_187, output_4_12, output_3_187;
mixer gate_output_3_187(.a(output_4_187), .b(output_4_12), .y(output_3_187));
wire output_5_187, output_5_12, output_4_187;
mixer gate_output_4_187(.a(output_5_187), .b(output_5_12), .y(output_4_187));
wire output_6_187, output_6_12, output_5_187;
mixer gate_output_5_187(.a(output_6_187), .b(output_6_12), .y(output_5_187));
wire output_7_187, output_7_12, output_6_187;
mixer gate_output_6_187(.a(output_7_187), .b(output_7_12), .y(output_6_187));
wire output_8_187, output_8_12, output_7_187;
mixer gate_output_7_187(.a(output_8_187), .b(output_8_12), .y(output_7_187));
wire output_9_187, output_9_12, output_8_187;
mixer gate_output_8_187(.a(output_9_187), .b(output_9_12), .y(output_8_187));
wire output_10_187, output_10_12, output_9_187;
mixer gate_output_9_187(.a(output_10_187), .b(output_10_12), .y(output_9_187));
wire output_11_187, output_11_12, output_10_187;
mixer gate_output_10_187(.a(output_11_187), .b(output_11_12), .y(output_10_187));
wire output_12_187, output_12_12, output_11_187;
mixer gate_output_11_187(.a(output_12_187), .b(output_12_12), .y(output_11_187));
wire output_13_187, output_13_12, output_12_187;
mixer gate_output_12_187(.a(output_13_187), .b(output_13_12), .y(output_12_187));
wire output_14_187, output_14_12, output_13_187;
mixer gate_output_13_187(.a(output_14_187), .b(output_14_12), .y(output_13_187));
wire output_15_187, output_15_12, output_14_187;
mixer gate_output_14_187(.a(output_15_187), .b(output_15_12), .y(output_14_187));
wire output_16_187, output_16_12, output_15_187;
mixer gate_output_15_187(.a(output_16_187), .b(output_16_12), .y(output_15_187));
wire output_1_188, output_1_13, output_0_188;
mixer gate_output_0_188(.a(output_1_188), .b(output_1_13), .y(output_0_188));
wire output_2_188, output_2_13, output_1_188;
mixer gate_output_1_188(.a(output_2_188), .b(output_2_13), .y(output_1_188));
wire output_3_188, output_3_13, output_2_188;
mixer gate_output_2_188(.a(output_3_188), .b(output_3_13), .y(output_2_188));
wire output_4_188, output_4_13, output_3_188;
mixer gate_output_3_188(.a(output_4_188), .b(output_4_13), .y(output_3_188));
wire output_5_188, output_5_13, output_4_188;
mixer gate_output_4_188(.a(output_5_188), .b(output_5_13), .y(output_4_188));
wire output_6_188, output_6_13, output_5_188;
mixer gate_output_5_188(.a(output_6_188), .b(output_6_13), .y(output_5_188));
wire output_7_188, output_7_13, output_6_188;
mixer gate_output_6_188(.a(output_7_188), .b(output_7_13), .y(output_6_188));
wire output_8_188, output_8_13, output_7_188;
mixer gate_output_7_188(.a(output_8_188), .b(output_8_13), .y(output_7_188));
wire output_9_188, output_9_13, output_8_188;
mixer gate_output_8_188(.a(output_9_188), .b(output_9_13), .y(output_8_188));
wire output_10_188, output_10_13, output_9_188;
mixer gate_output_9_188(.a(output_10_188), .b(output_10_13), .y(output_9_188));
wire output_11_188, output_11_13, output_10_188;
mixer gate_output_10_188(.a(output_11_188), .b(output_11_13), .y(output_10_188));
wire output_12_188, output_12_13, output_11_188;
mixer gate_output_11_188(.a(output_12_188), .b(output_12_13), .y(output_11_188));
wire output_13_188, output_13_13, output_12_188;
mixer gate_output_12_188(.a(output_13_188), .b(output_13_13), .y(output_12_188));
wire output_14_188, output_14_13, output_13_188;
mixer gate_output_13_188(.a(output_14_188), .b(output_14_13), .y(output_13_188));
wire output_15_188, output_15_13, output_14_188;
mixer gate_output_14_188(.a(output_15_188), .b(output_15_13), .y(output_14_188));
wire output_16_188, output_16_13, output_15_188;
mixer gate_output_15_188(.a(output_16_188), .b(output_16_13), .y(output_15_188));
wire output_1_189, output_1_14, output_0_189;
mixer gate_output_0_189(.a(output_1_189), .b(output_1_14), .y(output_0_189));
wire output_2_189, output_2_14, output_1_189;
mixer gate_output_1_189(.a(output_2_189), .b(output_2_14), .y(output_1_189));
wire output_3_189, output_3_14, output_2_189;
mixer gate_output_2_189(.a(output_3_189), .b(output_3_14), .y(output_2_189));
wire output_4_189, output_4_14, output_3_189;
mixer gate_output_3_189(.a(output_4_189), .b(output_4_14), .y(output_3_189));
wire output_5_189, output_5_14, output_4_189;
mixer gate_output_4_189(.a(output_5_189), .b(output_5_14), .y(output_4_189));
wire output_6_189, output_6_14, output_5_189;
mixer gate_output_5_189(.a(output_6_189), .b(output_6_14), .y(output_5_189));
wire output_7_189, output_7_14, output_6_189;
mixer gate_output_6_189(.a(output_7_189), .b(output_7_14), .y(output_6_189));
wire output_8_189, output_8_14, output_7_189;
mixer gate_output_7_189(.a(output_8_189), .b(output_8_14), .y(output_7_189));
wire output_9_189, output_9_14, output_8_189;
mixer gate_output_8_189(.a(output_9_189), .b(output_9_14), .y(output_8_189));
wire output_10_189, output_10_14, output_9_189;
mixer gate_output_9_189(.a(output_10_189), .b(output_10_14), .y(output_9_189));
wire output_11_189, output_11_14, output_10_189;
mixer gate_output_10_189(.a(output_11_189), .b(output_11_14), .y(output_10_189));
wire output_12_189, output_12_14, output_11_189;
mixer gate_output_11_189(.a(output_12_189), .b(output_12_14), .y(output_11_189));
wire output_13_189, output_13_14, output_12_189;
mixer gate_output_12_189(.a(output_13_189), .b(output_13_14), .y(output_12_189));
wire output_14_189, output_14_14, output_13_189;
mixer gate_output_13_189(.a(output_14_189), .b(output_14_14), .y(output_13_189));
wire output_15_189, output_15_14, output_14_189;
mixer gate_output_14_189(.a(output_15_189), .b(output_15_14), .y(output_14_189));
wire output_16_189, output_16_14, output_15_189;
mixer gate_output_15_189(.a(output_16_189), .b(output_16_14), .y(output_15_189));
wire output_1_190, output_1_15, output_0_190;
mixer gate_output_0_190(.a(output_1_190), .b(output_1_15), .y(output_0_190));
wire output_2_190, output_2_15, output_1_190;
mixer gate_output_1_190(.a(output_2_190), .b(output_2_15), .y(output_1_190));
wire output_3_190, output_3_15, output_2_190;
mixer gate_output_2_190(.a(output_3_190), .b(output_3_15), .y(output_2_190));
wire output_4_190, output_4_15, output_3_190;
mixer gate_output_3_190(.a(output_4_190), .b(output_4_15), .y(output_3_190));
wire output_5_190, output_5_15, output_4_190;
mixer gate_output_4_190(.a(output_5_190), .b(output_5_15), .y(output_4_190));
wire output_6_190, output_6_15, output_5_190;
mixer gate_output_5_190(.a(output_6_190), .b(output_6_15), .y(output_5_190));
wire output_7_190, output_7_15, output_6_190;
mixer gate_output_6_190(.a(output_7_190), .b(output_7_15), .y(output_6_190));
wire output_8_190, output_8_15, output_7_190;
mixer gate_output_7_190(.a(output_8_190), .b(output_8_15), .y(output_7_190));
wire output_9_190, output_9_15, output_8_190;
mixer gate_output_8_190(.a(output_9_190), .b(output_9_15), .y(output_8_190));
wire output_10_190, output_10_15, output_9_190;
mixer gate_output_9_190(.a(output_10_190), .b(output_10_15), .y(output_9_190));
wire output_11_190, output_11_15, output_10_190;
mixer gate_output_10_190(.a(output_11_190), .b(output_11_15), .y(output_10_190));
wire output_12_190, output_12_15, output_11_190;
mixer gate_output_11_190(.a(output_12_190), .b(output_12_15), .y(output_11_190));
wire output_13_190, output_13_15, output_12_190;
mixer gate_output_12_190(.a(output_13_190), .b(output_13_15), .y(output_12_190));
wire output_14_190, output_14_15, output_13_190;
mixer gate_output_13_190(.a(output_14_190), .b(output_14_15), .y(output_13_190));
wire output_15_190, output_15_15, output_14_190;
mixer gate_output_14_190(.a(output_15_190), .b(output_15_15), .y(output_14_190));
wire output_16_190, output_16_15, output_15_190;
mixer gate_output_15_190(.a(output_16_190), .b(output_16_15), .y(output_15_190));
wire output_1_191, output_1_0, output_0_191;
mixer gate_output_0_191(.a(output_1_191), .b(output_1_0), .y(output_0_191));
wire output_2_191, output_2_0, output_1_191;
mixer gate_output_1_191(.a(output_2_191), .b(output_2_0), .y(output_1_191));
wire output_3_191, output_3_0, output_2_191;
mixer gate_output_2_191(.a(output_3_191), .b(output_3_0), .y(output_2_191));
wire output_4_191, output_4_0, output_3_191;
mixer gate_output_3_191(.a(output_4_191), .b(output_4_0), .y(output_3_191));
wire output_5_191, output_5_0, output_4_191;
mixer gate_output_4_191(.a(output_5_191), .b(output_5_0), .y(output_4_191));
wire output_6_191, output_6_0, output_5_191;
mixer gate_output_5_191(.a(output_6_191), .b(output_6_0), .y(output_5_191));
wire output_7_191, output_7_0, output_6_191;
mixer gate_output_6_191(.a(output_7_191), .b(output_7_0), .y(output_6_191));
wire output_8_191, output_8_0, output_7_191;
mixer gate_output_7_191(.a(output_8_191), .b(output_8_0), .y(output_7_191));
wire output_9_191, output_9_0, output_8_191;
mixer gate_output_8_191(.a(output_9_191), .b(output_9_0), .y(output_8_191));
wire output_10_191, output_10_0, output_9_191;
mixer gate_output_9_191(.a(output_10_191), .b(output_10_0), .y(output_9_191));
wire output_11_191, output_11_0, output_10_191;
mixer gate_output_10_191(.a(output_11_191), .b(output_11_0), .y(output_10_191));
wire output_12_191, output_12_0, output_11_191;
mixer gate_output_11_191(.a(output_12_191), .b(output_12_0), .y(output_11_191));
wire output_13_191, output_13_0, output_12_191;
mixer gate_output_12_191(.a(output_13_191), .b(output_13_0), .y(output_12_191));
wire output_14_191, output_14_0, output_13_191;
mixer gate_output_13_191(.a(output_14_191), .b(output_14_0), .y(output_13_191));
wire output_15_191, output_15_0, output_14_191;
mixer gate_output_14_191(.a(output_15_191), .b(output_15_0), .y(output_14_191));
wire output_16_191, output_16_0, output_15_191;
mixer gate_output_15_191(.a(output_16_191), .b(output_16_0), .y(output_15_191));
wire output_1_192, output_1_1, output_0_192;
mixer gate_output_0_192(.a(output_1_192), .b(output_1_1), .y(output_0_192));
wire output_2_192, output_2_1, output_1_192;
mixer gate_output_1_192(.a(output_2_192), .b(output_2_1), .y(output_1_192));
wire output_3_192, output_3_1, output_2_192;
mixer gate_output_2_192(.a(output_3_192), .b(output_3_1), .y(output_2_192));
wire output_4_192, output_4_1, output_3_192;
mixer gate_output_3_192(.a(output_4_192), .b(output_4_1), .y(output_3_192));
wire output_5_192, output_5_1, output_4_192;
mixer gate_output_4_192(.a(output_5_192), .b(output_5_1), .y(output_4_192));
wire output_6_192, output_6_1, output_5_192;
mixer gate_output_5_192(.a(output_6_192), .b(output_6_1), .y(output_5_192));
wire output_7_192, output_7_1, output_6_192;
mixer gate_output_6_192(.a(output_7_192), .b(output_7_1), .y(output_6_192));
wire output_8_192, output_8_1, output_7_192;
mixer gate_output_7_192(.a(output_8_192), .b(output_8_1), .y(output_7_192));
wire output_9_192, output_9_1, output_8_192;
mixer gate_output_8_192(.a(output_9_192), .b(output_9_1), .y(output_8_192));
wire output_10_192, output_10_1, output_9_192;
mixer gate_output_9_192(.a(output_10_192), .b(output_10_1), .y(output_9_192));
wire output_11_192, output_11_1, output_10_192;
mixer gate_output_10_192(.a(output_11_192), .b(output_11_1), .y(output_10_192));
wire output_12_192, output_12_1, output_11_192;
mixer gate_output_11_192(.a(output_12_192), .b(output_12_1), .y(output_11_192));
wire output_13_192, output_13_1, output_12_192;
mixer gate_output_12_192(.a(output_13_192), .b(output_13_1), .y(output_12_192));
wire output_14_192, output_14_1, output_13_192;
mixer gate_output_13_192(.a(output_14_192), .b(output_14_1), .y(output_13_192));
wire output_15_192, output_15_1, output_14_192;
mixer gate_output_14_192(.a(output_15_192), .b(output_15_1), .y(output_14_192));
wire output_16_192, output_16_1, output_15_192;
mixer gate_output_15_192(.a(output_16_192), .b(output_16_1), .y(output_15_192));
wire output_1_193, output_1_2, output_0_193;
mixer gate_output_0_193(.a(output_1_193), .b(output_1_2), .y(output_0_193));
wire output_2_193, output_2_2, output_1_193;
mixer gate_output_1_193(.a(output_2_193), .b(output_2_2), .y(output_1_193));
wire output_3_193, output_3_2, output_2_193;
mixer gate_output_2_193(.a(output_3_193), .b(output_3_2), .y(output_2_193));
wire output_4_193, output_4_2, output_3_193;
mixer gate_output_3_193(.a(output_4_193), .b(output_4_2), .y(output_3_193));
wire output_5_193, output_5_2, output_4_193;
mixer gate_output_4_193(.a(output_5_193), .b(output_5_2), .y(output_4_193));
wire output_6_193, output_6_2, output_5_193;
mixer gate_output_5_193(.a(output_6_193), .b(output_6_2), .y(output_5_193));
wire output_7_193, output_7_2, output_6_193;
mixer gate_output_6_193(.a(output_7_193), .b(output_7_2), .y(output_6_193));
wire output_8_193, output_8_2, output_7_193;
mixer gate_output_7_193(.a(output_8_193), .b(output_8_2), .y(output_7_193));
wire output_9_193, output_9_2, output_8_193;
mixer gate_output_8_193(.a(output_9_193), .b(output_9_2), .y(output_8_193));
wire output_10_193, output_10_2, output_9_193;
mixer gate_output_9_193(.a(output_10_193), .b(output_10_2), .y(output_9_193));
wire output_11_193, output_11_2, output_10_193;
mixer gate_output_10_193(.a(output_11_193), .b(output_11_2), .y(output_10_193));
wire output_12_193, output_12_2, output_11_193;
mixer gate_output_11_193(.a(output_12_193), .b(output_12_2), .y(output_11_193));
wire output_13_193, output_13_2, output_12_193;
mixer gate_output_12_193(.a(output_13_193), .b(output_13_2), .y(output_12_193));
wire output_14_193, output_14_2, output_13_193;
mixer gate_output_13_193(.a(output_14_193), .b(output_14_2), .y(output_13_193));
wire output_15_193, output_15_2, output_14_193;
mixer gate_output_14_193(.a(output_15_193), .b(output_15_2), .y(output_14_193));
wire output_16_193, output_16_2, output_15_193;
mixer gate_output_15_193(.a(output_16_193), .b(output_16_2), .y(output_15_193));
wire output_1_194, output_1_3, output_0_194;
mixer gate_output_0_194(.a(output_1_194), .b(output_1_3), .y(output_0_194));
wire output_2_194, output_2_3, output_1_194;
mixer gate_output_1_194(.a(output_2_194), .b(output_2_3), .y(output_1_194));
wire output_3_194, output_3_3, output_2_194;
mixer gate_output_2_194(.a(output_3_194), .b(output_3_3), .y(output_2_194));
wire output_4_194, output_4_3, output_3_194;
mixer gate_output_3_194(.a(output_4_194), .b(output_4_3), .y(output_3_194));
wire output_5_194, output_5_3, output_4_194;
mixer gate_output_4_194(.a(output_5_194), .b(output_5_3), .y(output_4_194));
wire output_6_194, output_6_3, output_5_194;
mixer gate_output_5_194(.a(output_6_194), .b(output_6_3), .y(output_5_194));
wire output_7_194, output_7_3, output_6_194;
mixer gate_output_6_194(.a(output_7_194), .b(output_7_3), .y(output_6_194));
wire output_8_194, output_8_3, output_7_194;
mixer gate_output_7_194(.a(output_8_194), .b(output_8_3), .y(output_7_194));
wire output_9_194, output_9_3, output_8_194;
mixer gate_output_8_194(.a(output_9_194), .b(output_9_3), .y(output_8_194));
wire output_10_194, output_10_3, output_9_194;
mixer gate_output_9_194(.a(output_10_194), .b(output_10_3), .y(output_9_194));
wire output_11_194, output_11_3, output_10_194;
mixer gate_output_10_194(.a(output_11_194), .b(output_11_3), .y(output_10_194));
wire output_12_194, output_12_3, output_11_194;
mixer gate_output_11_194(.a(output_12_194), .b(output_12_3), .y(output_11_194));
wire output_13_194, output_13_3, output_12_194;
mixer gate_output_12_194(.a(output_13_194), .b(output_13_3), .y(output_12_194));
wire output_14_194, output_14_3, output_13_194;
mixer gate_output_13_194(.a(output_14_194), .b(output_14_3), .y(output_13_194));
wire output_15_194, output_15_3, output_14_194;
mixer gate_output_14_194(.a(output_15_194), .b(output_15_3), .y(output_14_194));
wire output_16_194, output_16_3, output_15_194;
mixer gate_output_15_194(.a(output_16_194), .b(output_16_3), .y(output_15_194));
wire output_1_195, output_1_4, output_0_195;
mixer gate_output_0_195(.a(output_1_195), .b(output_1_4), .y(output_0_195));
wire output_2_195, output_2_4, output_1_195;
mixer gate_output_1_195(.a(output_2_195), .b(output_2_4), .y(output_1_195));
wire output_3_195, output_3_4, output_2_195;
mixer gate_output_2_195(.a(output_3_195), .b(output_3_4), .y(output_2_195));
wire output_4_195, output_4_4, output_3_195;
mixer gate_output_3_195(.a(output_4_195), .b(output_4_4), .y(output_3_195));
wire output_5_195, output_5_4, output_4_195;
mixer gate_output_4_195(.a(output_5_195), .b(output_5_4), .y(output_4_195));
wire output_6_195, output_6_4, output_5_195;
mixer gate_output_5_195(.a(output_6_195), .b(output_6_4), .y(output_5_195));
wire output_7_195, output_7_4, output_6_195;
mixer gate_output_6_195(.a(output_7_195), .b(output_7_4), .y(output_6_195));
wire output_8_195, output_8_4, output_7_195;
mixer gate_output_7_195(.a(output_8_195), .b(output_8_4), .y(output_7_195));
wire output_9_195, output_9_4, output_8_195;
mixer gate_output_8_195(.a(output_9_195), .b(output_9_4), .y(output_8_195));
wire output_10_195, output_10_4, output_9_195;
mixer gate_output_9_195(.a(output_10_195), .b(output_10_4), .y(output_9_195));
wire output_11_195, output_11_4, output_10_195;
mixer gate_output_10_195(.a(output_11_195), .b(output_11_4), .y(output_10_195));
wire output_12_195, output_12_4, output_11_195;
mixer gate_output_11_195(.a(output_12_195), .b(output_12_4), .y(output_11_195));
wire output_13_195, output_13_4, output_12_195;
mixer gate_output_12_195(.a(output_13_195), .b(output_13_4), .y(output_12_195));
wire output_14_195, output_14_4, output_13_195;
mixer gate_output_13_195(.a(output_14_195), .b(output_14_4), .y(output_13_195));
wire output_15_195, output_15_4, output_14_195;
mixer gate_output_14_195(.a(output_15_195), .b(output_15_4), .y(output_14_195));
wire output_16_195, output_16_4, output_15_195;
mixer gate_output_15_195(.a(output_16_195), .b(output_16_4), .y(output_15_195));
wire output_1_196, output_1_5, output_0_196;
mixer gate_output_0_196(.a(output_1_196), .b(output_1_5), .y(output_0_196));
wire output_2_196, output_2_5, output_1_196;
mixer gate_output_1_196(.a(output_2_196), .b(output_2_5), .y(output_1_196));
wire output_3_196, output_3_5, output_2_196;
mixer gate_output_2_196(.a(output_3_196), .b(output_3_5), .y(output_2_196));
wire output_4_196, output_4_5, output_3_196;
mixer gate_output_3_196(.a(output_4_196), .b(output_4_5), .y(output_3_196));
wire output_5_196, output_5_5, output_4_196;
mixer gate_output_4_196(.a(output_5_196), .b(output_5_5), .y(output_4_196));
wire output_6_196, output_6_5, output_5_196;
mixer gate_output_5_196(.a(output_6_196), .b(output_6_5), .y(output_5_196));
wire output_7_196, output_7_5, output_6_196;
mixer gate_output_6_196(.a(output_7_196), .b(output_7_5), .y(output_6_196));
wire output_8_196, output_8_5, output_7_196;
mixer gate_output_7_196(.a(output_8_196), .b(output_8_5), .y(output_7_196));
wire output_9_196, output_9_5, output_8_196;
mixer gate_output_8_196(.a(output_9_196), .b(output_9_5), .y(output_8_196));
wire output_10_196, output_10_5, output_9_196;
mixer gate_output_9_196(.a(output_10_196), .b(output_10_5), .y(output_9_196));
wire output_11_196, output_11_5, output_10_196;
mixer gate_output_10_196(.a(output_11_196), .b(output_11_5), .y(output_10_196));
wire output_12_196, output_12_5, output_11_196;
mixer gate_output_11_196(.a(output_12_196), .b(output_12_5), .y(output_11_196));
wire output_13_196, output_13_5, output_12_196;
mixer gate_output_12_196(.a(output_13_196), .b(output_13_5), .y(output_12_196));
wire output_14_196, output_14_5, output_13_196;
mixer gate_output_13_196(.a(output_14_196), .b(output_14_5), .y(output_13_196));
wire output_15_196, output_15_5, output_14_196;
mixer gate_output_14_196(.a(output_15_196), .b(output_15_5), .y(output_14_196));
wire output_16_196, output_16_5, output_15_196;
mixer gate_output_15_196(.a(output_16_196), .b(output_16_5), .y(output_15_196));
wire output_1_197, output_1_6, output_0_197;
mixer gate_output_0_197(.a(output_1_197), .b(output_1_6), .y(output_0_197));
wire output_2_197, output_2_6, output_1_197;
mixer gate_output_1_197(.a(output_2_197), .b(output_2_6), .y(output_1_197));
wire output_3_197, output_3_6, output_2_197;
mixer gate_output_2_197(.a(output_3_197), .b(output_3_6), .y(output_2_197));
wire output_4_197, output_4_6, output_3_197;
mixer gate_output_3_197(.a(output_4_197), .b(output_4_6), .y(output_3_197));
wire output_5_197, output_5_6, output_4_197;
mixer gate_output_4_197(.a(output_5_197), .b(output_5_6), .y(output_4_197));
wire output_6_197, output_6_6, output_5_197;
mixer gate_output_5_197(.a(output_6_197), .b(output_6_6), .y(output_5_197));
wire output_7_197, output_7_6, output_6_197;
mixer gate_output_6_197(.a(output_7_197), .b(output_7_6), .y(output_6_197));
wire output_8_197, output_8_6, output_7_197;
mixer gate_output_7_197(.a(output_8_197), .b(output_8_6), .y(output_7_197));
wire output_9_197, output_9_6, output_8_197;
mixer gate_output_8_197(.a(output_9_197), .b(output_9_6), .y(output_8_197));
wire output_10_197, output_10_6, output_9_197;
mixer gate_output_9_197(.a(output_10_197), .b(output_10_6), .y(output_9_197));
wire output_11_197, output_11_6, output_10_197;
mixer gate_output_10_197(.a(output_11_197), .b(output_11_6), .y(output_10_197));
wire output_12_197, output_12_6, output_11_197;
mixer gate_output_11_197(.a(output_12_197), .b(output_12_6), .y(output_11_197));
wire output_13_197, output_13_6, output_12_197;
mixer gate_output_12_197(.a(output_13_197), .b(output_13_6), .y(output_12_197));
wire output_14_197, output_14_6, output_13_197;
mixer gate_output_13_197(.a(output_14_197), .b(output_14_6), .y(output_13_197));
wire output_15_197, output_15_6, output_14_197;
mixer gate_output_14_197(.a(output_15_197), .b(output_15_6), .y(output_14_197));
wire output_16_197, output_16_6, output_15_197;
mixer gate_output_15_197(.a(output_16_197), .b(output_16_6), .y(output_15_197));
wire output_1_198, output_1_7, output_0_198;
mixer gate_output_0_198(.a(output_1_198), .b(output_1_7), .y(output_0_198));
wire output_2_198, output_2_7, output_1_198;
mixer gate_output_1_198(.a(output_2_198), .b(output_2_7), .y(output_1_198));
wire output_3_198, output_3_7, output_2_198;
mixer gate_output_2_198(.a(output_3_198), .b(output_3_7), .y(output_2_198));
wire output_4_198, output_4_7, output_3_198;
mixer gate_output_3_198(.a(output_4_198), .b(output_4_7), .y(output_3_198));
wire output_5_198, output_5_7, output_4_198;
mixer gate_output_4_198(.a(output_5_198), .b(output_5_7), .y(output_4_198));
wire output_6_198, output_6_7, output_5_198;
mixer gate_output_5_198(.a(output_6_198), .b(output_6_7), .y(output_5_198));
wire output_7_198, output_7_7, output_6_198;
mixer gate_output_6_198(.a(output_7_198), .b(output_7_7), .y(output_6_198));
wire output_8_198, output_8_7, output_7_198;
mixer gate_output_7_198(.a(output_8_198), .b(output_8_7), .y(output_7_198));
wire output_9_198, output_9_7, output_8_198;
mixer gate_output_8_198(.a(output_9_198), .b(output_9_7), .y(output_8_198));
wire output_10_198, output_10_7, output_9_198;
mixer gate_output_9_198(.a(output_10_198), .b(output_10_7), .y(output_9_198));
wire output_11_198, output_11_7, output_10_198;
mixer gate_output_10_198(.a(output_11_198), .b(output_11_7), .y(output_10_198));
wire output_12_198, output_12_7, output_11_198;
mixer gate_output_11_198(.a(output_12_198), .b(output_12_7), .y(output_11_198));
wire output_13_198, output_13_7, output_12_198;
mixer gate_output_12_198(.a(output_13_198), .b(output_13_7), .y(output_12_198));
wire output_14_198, output_14_7, output_13_198;
mixer gate_output_13_198(.a(output_14_198), .b(output_14_7), .y(output_13_198));
wire output_15_198, output_15_7, output_14_198;
mixer gate_output_14_198(.a(output_15_198), .b(output_15_7), .y(output_14_198));
wire output_16_198, output_16_7, output_15_198;
mixer gate_output_15_198(.a(output_16_198), .b(output_16_7), .y(output_15_198));
wire output_1_199, output_1_8, output_0_199;
mixer gate_output_0_199(.a(output_1_199), .b(output_1_8), .y(output_0_199));
wire output_2_199, output_2_8, output_1_199;
mixer gate_output_1_199(.a(output_2_199), .b(output_2_8), .y(output_1_199));
wire output_3_199, output_3_8, output_2_199;
mixer gate_output_2_199(.a(output_3_199), .b(output_3_8), .y(output_2_199));
wire output_4_199, output_4_8, output_3_199;
mixer gate_output_3_199(.a(output_4_199), .b(output_4_8), .y(output_3_199));
wire output_5_199, output_5_8, output_4_199;
mixer gate_output_4_199(.a(output_5_199), .b(output_5_8), .y(output_4_199));
wire output_6_199, output_6_8, output_5_199;
mixer gate_output_5_199(.a(output_6_199), .b(output_6_8), .y(output_5_199));
wire output_7_199, output_7_8, output_6_199;
mixer gate_output_6_199(.a(output_7_199), .b(output_7_8), .y(output_6_199));
wire output_8_199, output_8_8, output_7_199;
mixer gate_output_7_199(.a(output_8_199), .b(output_8_8), .y(output_7_199));
wire output_9_199, output_9_8, output_8_199;
mixer gate_output_8_199(.a(output_9_199), .b(output_9_8), .y(output_8_199));
wire output_10_199, output_10_8, output_9_199;
mixer gate_output_9_199(.a(output_10_199), .b(output_10_8), .y(output_9_199));
wire output_11_199, output_11_8, output_10_199;
mixer gate_output_10_199(.a(output_11_199), .b(output_11_8), .y(output_10_199));
wire output_12_199, output_12_8, output_11_199;
mixer gate_output_11_199(.a(output_12_199), .b(output_12_8), .y(output_11_199));
wire output_13_199, output_13_8, output_12_199;
mixer gate_output_12_199(.a(output_13_199), .b(output_13_8), .y(output_12_199));
wire output_14_199, output_14_8, output_13_199;
mixer gate_output_13_199(.a(output_14_199), .b(output_14_8), .y(output_13_199));
wire output_15_199, output_15_8, output_14_199;
mixer gate_output_14_199(.a(output_15_199), .b(output_15_8), .y(output_14_199));
wire output_16_199, output_16_8, output_15_199;
mixer gate_output_15_199(.a(output_16_199), .b(output_16_8), .y(output_15_199));
wire output_1_200, output_1_9, output_0_200;
mixer gate_output_0_200(.a(output_1_200), .b(output_1_9), .y(output_0_200));
wire output_2_200, output_2_9, output_1_200;
mixer gate_output_1_200(.a(output_2_200), .b(output_2_9), .y(output_1_200));
wire output_3_200, output_3_9, output_2_200;
mixer gate_output_2_200(.a(output_3_200), .b(output_3_9), .y(output_2_200));
wire output_4_200, output_4_9, output_3_200;
mixer gate_output_3_200(.a(output_4_200), .b(output_4_9), .y(output_3_200));
wire output_5_200, output_5_9, output_4_200;
mixer gate_output_4_200(.a(output_5_200), .b(output_5_9), .y(output_4_200));
wire output_6_200, output_6_9, output_5_200;
mixer gate_output_5_200(.a(output_6_200), .b(output_6_9), .y(output_5_200));
wire output_7_200, output_7_9, output_6_200;
mixer gate_output_6_200(.a(output_7_200), .b(output_7_9), .y(output_6_200));
wire output_8_200, output_8_9, output_7_200;
mixer gate_output_7_200(.a(output_8_200), .b(output_8_9), .y(output_7_200));
wire output_9_200, output_9_9, output_8_200;
mixer gate_output_8_200(.a(output_9_200), .b(output_9_9), .y(output_8_200));
wire output_10_200, output_10_9, output_9_200;
mixer gate_output_9_200(.a(output_10_200), .b(output_10_9), .y(output_9_200));
wire output_11_200, output_11_9, output_10_200;
mixer gate_output_10_200(.a(output_11_200), .b(output_11_9), .y(output_10_200));
wire output_12_200, output_12_9, output_11_200;
mixer gate_output_11_200(.a(output_12_200), .b(output_12_9), .y(output_11_200));
wire output_13_200, output_13_9, output_12_200;
mixer gate_output_12_200(.a(output_13_200), .b(output_13_9), .y(output_12_200));
wire output_14_200, output_14_9, output_13_200;
mixer gate_output_13_200(.a(output_14_200), .b(output_14_9), .y(output_13_200));
wire output_15_200, output_15_9, output_14_200;
mixer gate_output_14_200(.a(output_15_200), .b(output_15_9), .y(output_14_200));
wire output_16_200, output_16_9, output_15_200;
mixer gate_output_15_200(.a(output_16_200), .b(output_16_9), .y(output_15_200));
wire output_1_201, output_1_10, output_0_201;
mixer gate_output_0_201(.a(output_1_201), .b(output_1_10), .y(output_0_201));
wire output_2_201, output_2_10, output_1_201;
mixer gate_output_1_201(.a(output_2_201), .b(output_2_10), .y(output_1_201));
wire output_3_201, output_3_10, output_2_201;
mixer gate_output_2_201(.a(output_3_201), .b(output_3_10), .y(output_2_201));
wire output_4_201, output_4_10, output_3_201;
mixer gate_output_3_201(.a(output_4_201), .b(output_4_10), .y(output_3_201));
wire output_5_201, output_5_10, output_4_201;
mixer gate_output_4_201(.a(output_5_201), .b(output_5_10), .y(output_4_201));
wire output_6_201, output_6_10, output_5_201;
mixer gate_output_5_201(.a(output_6_201), .b(output_6_10), .y(output_5_201));
wire output_7_201, output_7_10, output_6_201;
mixer gate_output_6_201(.a(output_7_201), .b(output_7_10), .y(output_6_201));
wire output_8_201, output_8_10, output_7_201;
mixer gate_output_7_201(.a(output_8_201), .b(output_8_10), .y(output_7_201));
wire output_9_201, output_9_10, output_8_201;
mixer gate_output_8_201(.a(output_9_201), .b(output_9_10), .y(output_8_201));
wire output_10_201, output_10_10, output_9_201;
mixer gate_output_9_201(.a(output_10_201), .b(output_10_10), .y(output_9_201));
wire output_11_201, output_11_10, output_10_201;
mixer gate_output_10_201(.a(output_11_201), .b(output_11_10), .y(output_10_201));
wire output_12_201, output_12_10, output_11_201;
mixer gate_output_11_201(.a(output_12_201), .b(output_12_10), .y(output_11_201));
wire output_13_201, output_13_10, output_12_201;
mixer gate_output_12_201(.a(output_13_201), .b(output_13_10), .y(output_12_201));
wire output_14_201, output_14_10, output_13_201;
mixer gate_output_13_201(.a(output_14_201), .b(output_14_10), .y(output_13_201));
wire output_15_201, output_15_10, output_14_201;
mixer gate_output_14_201(.a(output_15_201), .b(output_15_10), .y(output_14_201));
wire output_16_201, output_16_10, output_15_201;
mixer gate_output_15_201(.a(output_16_201), .b(output_16_10), .y(output_15_201));
wire output_1_202, output_1_11, output_0_202;
mixer gate_output_0_202(.a(output_1_202), .b(output_1_11), .y(output_0_202));
wire output_2_202, output_2_11, output_1_202;
mixer gate_output_1_202(.a(output_2_202), .b(output_2_11), .y(output_1_202));
wire output_3_202, output_3_11, output_2_202;
mixer gate_output_2_202(.a(output_3_202), .b(output_3_11), .y(output_2_202));
wire output_4_202, output_4_11, output_3_202;
mixer gate_output_3_202(.a(output_4_202), .b(output_4_11), .y(output_3_202));
wire output_5_202, output_5_11, output_4_202;
mixer gate_output_4_202(.a(output_5_202), .b(output_5_11), .y(output_4_202));
wire output_6_202, output_6_11, output_5_202;
mixer gate_output_5_202(.a(output_6_202), .b(output_6_11), .y(output_5_202));
wire output_7_202, output_7_11, output_6_202;
mixer gate_output_6_202(.a(output_7_202), .b(output_7_11), .y(output_6_202));
wire output_8_202, output_8_11, output_7_202;
mixer gate_output_7_202(.a(output_8_202), .b(output_8_11), .y(output_7_202));
wire output_9_202, output_9_11, output_8_202;
mixer gate_output_8_202(.a(output_9_202), .b(output_9_11), .y(output_8_202));
wire output_10_202, output_10_11, output_9_202;
mixer gate_output_9_202(.a(output_10_202), .b(output_10_11), .y(output_9_202));
wire output_11_202, output_11_11, output_10_202;
mixer gate_output_10_202(.a(output_11_202), .b(output_11_11), .y(output_10_202));
wire output_12_202, output_12_11, output_11_202;
mixer gate_output_11_202(.a(output_12_202), .b(output_12_11), .y(output_11_202));
wire output_13_202, output_13_11, output_12_202;
mixer gate_output_12_202(.a(output_13_202), .b(output_13_11), .y(output_12_202));
wire output_14_202, output_14_11, output_13_202;
mixer gate_output_13_202(.a(output_14_202), .b(output_14_11), .y(output_13_202));
wire output_15_202, output_15_11, output_14_202;
mixer gate_output_14_202(.a(output_15_202), .b(output_15_11), .y(output_14_202));
wire output_16_202, output_16_11, output_15_202;
mixer gate_output_15_202(.a(output_16_202), .b(output_16_11), .y(output_15_202));
wire output_1_203, output_1_12, output_0_203;
mixer gate_output_0_203(.a(output_1_203), .b(output_1_12), .y(output_0_203));
wire output_2_203, output_2_12, output_1_203;
mixer gate_output_1_203(.a(output_2_203), .b(output_2_12), .y(output_1_203));
wire output_3_203, output_3_12, output_2_203;
mixer gate_output_2_203(.a(output_3_203), .b(output_3_12), .y(output_2_203));
wire output_4_203, output_4_12, output_3_203;
mixer gate_output_3_203(.a(output_4_203), .b(output_4_12), .y(output_3_203));
wire output_5_203, output_5_12, output_4_203;
mixer gate_output_4_203(.a(output_5_203), .b(output_5_12), .y(output_4_203));
wire output_6_203, output_6_12, output_5_203;
mixer gate_output_5_203(.a(output_6_203), .b(output_6_12), .y(output_5_203));
wire output_7_203, output_7_12, output_6_203;
mixer gate_output_6_203(.a(output_7_203), .b(output_7_12), .y(output_6_203));
wire output_8_203, output_8_12, output_7_203;
mixer gate_output_7_203(.a(output_8_203), .b(output_8_12), .y(output_7_203));
wire output_9_203, output_9_12, output_8_203;
mixer gate_output_8_203(.a(output_9_203), .b(output_9_12), .y(output_8_203));
wire output_10_203, output_10_12, output_9_203;
mixer gate_output_9_203(.a(output_10_203), .b(output_10_12), .y(output_9_203));
wire output_11_203, output_11_12, output_10_203;
mixer gate_output_10_203(.a(output_11_203), .b(output_11_12), .y(output_10_203));
wire output_12_203, output_12_12, output_11_203;
mixer gate_output_11_203(.a(output_12_203), .b(output_12_12), .y(output_11_203));
wire output_13_203, output_13_12, output_12_203;
mixer gate_output_12_203(.a(output_13_203), .b(output_13_12), .y(output_12_203));
wire output_14_203, output_14_12, output_13_203;
mixer gate_output_13_203(.a(output_14_203), .b(output_14_12), .y(output_13_203));
wire output_15_203, output_15_12, output_14_203;
mixer gate_output_14_203(.a(output_15_203), .b(output_15_12), .y(output_14_203));
wire output_16_203, output_16_12, output_15_203;
mixer gate_output_15_203(.a(output_16_203), .b(output_16_12), .y(output_15_203));
wire output_1_204, output_1_13, output_0_204;
mixer gate_output_0_204(.a(output_1_204), .b(output_1_13), .y(output_0_204));
wire output_2_204, output_2_13, output_1_204;
mixer gate_output_1_204(.a(output_2_204), .b(output_2_13), .y(output_1_204));
wire output_3_204, output_3_13, output_2_204;
mixer gate_output_2_204(.a(output_3_204), .b(output_3_13), .y(output_2_204));
wire output_4_204, output_4_13, output_3_204;
mixer gate_output_3_204(.a(output_4_204), .b(output_4_13), .y(output_3_204));
wire output_5_204, output_5_13, output_4_204;
mixer gate_output_4_204(.a(output_5_204), .b(output_5_13), .y(output_4_204));
wire output_6_204, output_6_13, output_5_204;
mixer gate_output_5_204(.a(output_6_204), .b(output_6_13), .y(output_5_204));
wire output_7_204, output_7_13, output_6_204;
mixer gate_output_6_204(.a(output_7_204), .b(output_7_13), .y(output_6_204));
wire output_8_204, output_8_13, output_7_204;
mixer gate_output_7_204(.a(output_8_204), .b(output_8_13), .y(output_7_204));
wire output_9_204, output_9_13, output_8_204;
mixer gate_output_8_204(.a(output_9_204), .b(output_9_13), .y(output_8_204));
wire output_10_204, output_10_13, output_9_204;
mixer gate_output_9_204(.a(output_10_204), .b(output_10_13), .y(output_9_204));
wire output_11_204, output_11_13, output_10_204;
mixer gate_output_10_204(.a(output_11_204), .b(output_11_13), .y(output_10_204));
wire output_12_204, output_12_13, output_11_204;
mixer gate_output_11_204(.a(output_12_204), .b(output_12_13), .y(output_11_204));
wire output_13_204, output_13_13, output_12_204;
mixer gate_output_12_204(.a(output_13_204), .b(output_13_13), .y(output_12_204));
wire output_14_204, output_14_13, output_13_204;
mixer gate_output_13_204(.a(output_14_204), .b(output_14_13), .y(output_13_204));
wire output_15_204, output_15_13, output_14_204;
mixer gate_output_14_204(.a(output_15_204), .b(output_15_13), .y(output_14_204));
wire output_16_204, output_16_13, output_15_204;
mixer gate_output_15_204(.a(output_16_204), .b(output_16_13), .y(output_15_204));
wire output_1_205, output_1_14, output_0_205;
mixer gate_output_0_205(.a(output_1_205), .b(output_1_14), .y(output_0_205));
wire output_2_205, output_2_14, output_1_205;
mixer gate_output_1_205(.a(output_2_205), .b(output_2_14), .y(output_1_205));
wire output_3_205, output_3_14, output_2_205;
mixer gate_output_2_205(.a(output_3_205), .b(output_3_14), .y(output_2_205));
wire output_4_205, output_4_14, output_3_205;
mixer gate_output_3_205(.a(output_4_205), .b(output_4_14), .y(output_3_205));
wire output_5_205, output_5_14, output_4_205;
mixer gate_output_4_205(.a(output_5_205), .b(output_5_14), .y(output_4_205));
wire output_6_205, output_6_14, output_5_205;
mixer gate_output_5_205(.a(output_6_205), .b(output_6_14), .y(output_5_205));
wire output_7_205, output_7_14, output_6_205;
mixer gate_output_6_205(.a(output_7_205), .b(output_7_14), .y(output_6_205));
wire output_8_205, output_8_14, output_7_205;
mixer gate_output_7_205(.a(output_8_205), .b(output_8_14), .y(output_7_205));
wire output_9_205, output_9_14, output_8_205;
mixer gate_output_8_205(.a(output_9_205), .b(output_9_14), .y(output_8_205));
wire output_10_205, output_10_14, output_9_205;
mixer gate_output_9_205(.a(output_10_205), .b(output_10_14), .y(output_9_205));
wire output_11_205, output_11_14, output_10_205;
mixer gate_output_10_205(.a(output_11_205), .b(output_11_14), .y(output_10_205));
wire output_12_205, output_12_14, output_11_205;
mixer gate_output_11_205(.a(output_12_205), .b(output_12_14), .y(output_11_205));
wire output_13_205, output_13_14, output_12_205;
mixer gate_output_12_205(.a(output_13_205), .b(output_13_14), .y(output_12_205));
wire output_14_205, output_14_14, output_13_205;
mixer gate_output_13_205(.a(output_14_205), .b(output_14_14), .y(output_13_205));
wire output_15_205, output_15_14, output_14_205;
mixer gate_output_14_205(.a(output_15_205), .b(output_15_14), .y(output_14_205));
wire output_16_205, output_16_14, output_15_205;
mixer gate_output_15_205(.a(output_16_205), .b(output_16_14), .y(output_15_205));
wire output_1_206, output_1_15, output_0_206;
mixer gate_output_0_206(.a(output_1_206), .b(output_1_15), .y(output_0_206));
wire output_2_206, output_2_15, output_1_206;
mixer gate_output_1_206(.a(output_2_206), .b(output_2_15), .y(output_1_206));
wire output_3_206, output_3_15, output_2_206;
mixer gate_output_2_206(.a(output_3_206), .b(output_3_15), .y(output_2_206));
wire output_4_206, output_4_15, output_3_206;
mixer gate_output_3_206(.a(output_4_206), .b(output_4_15), .y(output_3_206));
wire output_5_206, output_5_15, output_4_206;
mixer gate_output_4_206(.a(output_5_206), .b(output_5_15), .y(output_4_206));
wire output_6_206, output_6_15, output_5_206;
mixer gate_output_5_206(.a(output_6_206), .b(output_6_15), .y(output_5_206));
wire output_7_206, output_7_15, output_6_206;
mixer gate_output_6_206(.a(output_7_206), .b(output_7_15), .y(output_6_206));
wire output_8_206, output_8_15, output_7_206;
mixer gate_output_7_206(.a(output_8_206), .b(output_8_15), .y(output_7_206));
wire output_9_206, output_9_15, output_8_206;
mixer gate_output_8_206(.a(output_9_206), .b(output_9_15), .y(output_8_206));
wire output_10_206, output_10_15, output_9_206;
mixer gate_output_9_206(.a(output_10_206), .b(output_10_15), .y(output_9_206));
wire output_11_206, output_11_15, output_10_206;
mixer gate_output_10_206(.a(output_11_206), .b(output_11_15), .y(output_10_206));
wire output_12_206, output_12_15, output_11_206;
mixer gate_output_11_206(.a(output_12_206), .b(output_12_15), .y(output_11_206));
wire output_13_206, output_13_15, output_12_206;
mixer gate_output_12_206(.a(output_13_206), .b(output_13_15), .y(output_12_206));
wire output_14_206, output_14_15, output_13_206;
mixer gate_output_13_206(.a(output_14_206), .b(output_14_15), .y(output_13_206));
wire output_15_206, output_15_15, output_14_206;
mixer gate_output_14_206(.a(output_15_206), .b(output_15_15), .y(output_14_206));
wire output_16_206, output_16_15, output_15_206;
mixer gate_output_15_206(.a(output_16_206), .b(output_16_15), .y(output_15_206));
wire output_1_207, output_1_0, output_0_207;
mixer gate_output_0_207(.a(output_1_207), .b(output_1_0), .y(output_0_207));
wire output_2_207, output_2_0, output_1_207;
mixer gate_output_1_207(.a(output_2_207), .b(output_2_0), .y(output_1_207));
wire output_3_207, output_3_0, output_2_207;
mixer gate_output_2_207(.a(output_3_207), .b(output_3_0), .y(output_2_207));
wire output_4_207, output_4_0, output_3_207;
mixer gate_output_3_207(.a(output_4_207), .b(output_4_0), .y(output_3_207));
wire output_5_207, output_5_0, output_4_207;
mixer gate_output_4_207(.a(output_5_207), .b(output_5_0), .y(output_4_207));
wire output_6_207, output_6_0, output_5_207;
mixer gate_output_5_207(.a(output_6_207), .b(output_6_0), .y(output_5_207));
wire output_7_207, output_7_0, output_6_207;
mixer gate_output_6_207(.a(output_7_207), .b(output_7_0), .y(output_6_207));
wire output_8_207, output_8_0, output_7_207;
mixer gate_output_7_207(.a(output_8_207), .b(output_8_0), .y(output_7_207));
wire output_9_207, output_9_0, output_8_207;
mixer gate_output_8_207(.a(output_9_207), .b(output_9_0), .y(output_8_207));
wire output_10_207, output_10_0, output_9_207;
mixer gate_output_9_207(.a(output_10_207), .b(output_10_0), .y(output_9_207));
wire output_11_207, output_11_0, output_10_207;
mixer gate_output_10_207(.a(output_11_207), .b(output_11_0), .y(output_10_207));
wire output_12_207, output_12_0, output_11_207;
mixer gate_output_11_207(.a(output_12_207), .b(output_12_0), .y(output_11_207));
wire output_13_207, output_13_0, output_12_207;
mixer gate_output_12_207(.a(output_13_207), .b(output_13_0), .y(output_12_207));
wire output_14_207, output_14_0, output_13_207;
mixer gate_output_13_207(.a(output_14_207), .b(output_14_0), .y(output_13_207));
wire output_15_207, output_15_0, output_14_207;
mixer gate_output_14_207(.a(output_15_207), .b(output_15_0), .y(output_14_207));
wire output_16_207, output_16_0, output_15_207;
mixer gate_output_15_207(.a(output_16_207), .b(output_16_0), .y(output_15_207));
wire output_1_208, output_1_1, output_0_208;
mixer gate_output_0_208(.a(output_1_208), .b(output_1_1), .y(output_0_208));
wire output_2_208, output_2_1, output_1_208;
mixer gate_output_1_208(.a(output_2_208), .b(output_2_1), .y(output_1_208));
wire output_3_208, output_3_1, output_2_208;
mixer gate_output_2_208(.a(output_3_208), .b(output_3_1), .y(output_2_208));
wire output_4_208, output_4_1, output_3_208;
mixer gate_output_3_208(.a(output_4_208), .b(output_4_1), .y(output_3_208));
wire output_5_208, output_5_1, output_4_208;
mixer gate_output_4_208(.a(output_5_208), .b(output_5_1), .y(output_4_208));
wire output_6_208, output_6_1, output_5_208;
mixer gate_output_5_208(.a(output_6_208), .b(output_6_1), .y(output_5_208));
wire output_7_208, output_7_1, output_6_208;
mixer gate_output_6_208(.a(output_7_208), .b(output_7_1), .y(output_6_208));
wire output_8_208, output_8_1, output_7_208;
mixer gate_output_7_208(.a(output_8_208), .b(output_8_1), .y(output_7_208));
wire output_9_208, output_9_1, output_8_208;
mixer gate_output_8_208(.a(output_9_208), .b(output_9_1), .y(output_8_208));
wire output_10_208, output_10_1, output_9_208;
mixer gate_output_9_208(.a(output_10_208), .b(output_10_1), .y(output_9_208));
wire output_11_208, output_11_1, output_10_208;
mixer gate_output_10_208(.a(output_11_208), .b(output_11_1), .y(output_10_208));
wire output_12_208, output_12_1, output_11_208;
mixer gate_output_11_208(.a(output_12_208), .b(output_12_1), .y(output_11_208));
wire output_13_208, output_13_1, output_12_208;
mixer gate_output_12_208(.a(output_13_208), .b(output_13_1), .y(output_12_208));
wire output_14_208, output_14_1, output_13_208;
mixer gate_output_13_208(.a(output_14_208), .b(output_14_1), .y(output_13_208));
wire output_15_208, output_15_1, output_14_208;
mixer gate_output_14_208(.a(output_15_208), .b(output_15_1), .y(output_14_208));
wire output_16_208, output_16_1, output_15_208;
mixer gate_output_15_208(.a(output_16_208), .b(output_16_1), .y(output_15_208));
wire output_1_209, output_1_2, output_0_209;
mixer gate_output_0_209(.a(output_1_209), .b(output_1_2), .y(output_0_209));
wire output_2_209, output_2_2, output_1_209;
mixer gate_output_1_209(.a(output_2_209), .b(output_2_2), .y(output_1_209));
wire output_3_209, output_3_2, output_2_209;
mixer gate_output_2_209(.a(output_3_209), .b(output_3_2), .y(output_2_209));
wire output_4_209, output_4_2, output_3_209;
mixer gate_output_3_209(.a(output_4_209), .b(output_4_2), .y(output_3_209));
wire output_5_209, output_5_2, output_4_209;
mixer gate_output_4_209(.a(output_5_209), .b(output_5_2), .y(output_4_209));
wire output_6_209, output_6_2, output_5_209;
mixer gate_output_5_209(.a(output_6_209), .b(output_6_2), .y(output_5_209));
wire output_7_209, output_7_2, output_6_209;
mixer gate_output_6_209(.a(output_7_209), .b(output_7_2), .y(output_6_209));
wire output_8_209, output_8_2, output_7_209;
mixer gate_output_7_209(.a(output_8_209), .b(output_8_2), .y(output_7_209));
wire output_9_209, output_9_2, output_8_209;
mixer gate_output_8_209(.a(output_9_209), .b(output_9_2), .y(output_8_209));
wire output_10_209, output_10_2, output_9_209;
mixer gate_output_9_209(.a(output_10_209), .b(output_10_2), .y(output_9_209));
wire output_11_209, output_11_2, output_10_209;
mixer gate_output_10_209(.a(output_11_209), .b(output_11_2), .y(output_10_209));
wire output_12_209, output_12_2, output_11_209;
mixer gate_output_11_209(.a(output_12_209), .b(output_12_2), .y(output_11_209));
wire output_13_209, output_13_2, output_12_209;
mixer gate_output_12_209(.a(output_13_209), .b(output_13_2), .y(output_12_209));
wire output_14_209, output_14_2, output_13_209;
mixer gate_output_13_209(.a(output_14_209), .b(output_14_2), .y(output_13_209));
wire output_15_209, output_15_2, output_14_209;
mixer gate_output_14_209(.a(output_15_209), .b(output_15_2), .y(output_14_209));
wire output_16_209, output_16_2, output_15_209;
mixer gate_output_15_209(.a(output_16_209), .b(output_16_2), .y(output_15_209));
wire output_1_210, output_1_3, output_0_210;
mixer gate_output_0_210(.a(output_1_210), .b(output_1_3), .y(output_0_210));
wire output_2_210, output_2_3, output_1_210;
mixer gate_output_1_210(.a(output_2_210), .b(output_2_3), .y(output_1_210));
wire output_3_210, output_3_3, output_2_210;
mixer gate_output_2_210(.a(output_3_210), .b(output_3_3), .y(output_2_210));
wire output_4_210, output_4_3, output_3_210;
mixer gate_output_3_210(.a(output_4_210), .b(output_4_3), .y(output_3_210));
wire output_5_210, output_5_3, output_4_210;
mixer gate_output_4_210(.a(output_5_210), .b(output_5_3), .y(output_4_210));
wire output_6_210, output_6_3, output_5_210;
mixer gate_output_5_210(.a(output_6_210), .b(output_6_3), .y(output_5_210));
wire output_7_210, output_7_3, output_6_210;
mixer gate_output_6_210(.a(output_7_210), .b(output_7_3), .y(output_6_210));
wire output_8_210, output_8_3, output_7_210;
mixer gate_output_7_210(.a(output_8_210), .b(output_8_3), .y(output_7_210));
wire output_9_210, output_9_3, output_8_210;
mixer gate_output_8_210(.a(output_9_210), .b(output_9_3), .y(output_8_210));
wire output_10_210, output_10_3, output_9_210;
mixer gate_output_9_210(.a(output_10_210), .b(output_10_3), .y(output_9_210));
wire output_11_210, output_11_3, output_10_210;
mixer gate_output_10_210(.a(output_11_210), .b(output_11_3), .y(output_10_210));
wire output_12_210, output_12_3, output_11_210;
mixer gate_output_11_210(.a(output_12_210), .b(output_12_3), .y(output_11_210));
wire output_13_210, output_13_3, output_12_210;
mixer gate_output_12_210(.a(output_13_210), .b(output_13_3), .y(output_12_210));
wire output_14_210, output_14_3, output_13_210;
mixer gate_output_13_210(.a(output_14_210), .b(output_14_3), .y(output_13_210));
wire output_15_210, output_15_3, output_14_210;
mixer gate_output_14_210(.a(output_15_210), .b(output_15_3), .y(output_14_210));
wire output_16_210, output_16_3, output_15_210;
mixer gate_output_15_210(.a(output_16_210), .b(output_16_3), .y(output_15_210));
wire output_1_211, output_1_4, output_0_211;
mixer gate_output_0_211(.a(output_1_211), .b(output_1_4), .y(output_0_211));
wire output_2_211, output_2_4, output_1_211;
mixer gate_output_1_211(.a(output_2_211), .b(output_2_4), .y(output_1_211));
wire output_3_211, output_3_4, output_2_211;
mixer gate_output_2_211(.a(output_3_211), .b(output_3_4), .y(output_2_211));
wire output_4_211, output_4_4, output_3_211;
mixer gate_output_3_211(.a(output_4_211), .b(output_4_4), .y(output_3_211));
wire output_5_211, output_5_4, output_4_211;
mixer gate_output_4_211(.a(output_5_211), .b(output_5_4), .y(output_4_211));
wire output_6_211, output_6_4, output_5_211;
mixer gate_output_5_211(.a(output_6_211), .b(output_6_4), .y(output_5_211));
wire output_7_211, output_7_4, output_6_211;
mixer gate_output_6_211(.a(output_7_211), .b(output_7_4), .y(output_6_211));
wire output_8_211, output_8_4, output_7_211;
mixer gate_output_7_211(.a(output_8_211), .b(output_8_4), .y(output_7_211));
wire output_9_211, output_9_4, output_8_211;
mixer gate_output_8_211(.a(output_9_211), .b(output_9_4), .y(output_8_211));
wire output_10_211, output_10_4, output_9_211;
mixer gate_output_9_211(.a(output_10_211), .b(output_10_4), .y(output_9_211));
wire output_11_211, output_11_4, output_10_211;
mixer gate_output_10_211(.a(output_11_211), .b(output_11_4), .y(output_10_211));
wire output_12_211, output_12_4, output_11_211;
mixer gate_output_11_211(.a(output_12_211), .b(output_12_4), .y(output_11_211));
wire output_13_211, output_13_4, output_12_211;
mixer gate_output_12_211(.a(output_13_211), .b(output_13_4), .y(output_12_211));
wire output_14_211, output_14_4, output_13_211;
mixer gate_output_13_211(.a(output_14_211), .b(output_14_4), .y(output_13_211));
wire output_15_211, output_15_4, output_14_211;
mixer gate_output_14_211(.a(output_15_211), .b(output_15_4), .y(output_14_211));
wire output_16_211, output_16_4, output_15_211;
mixer gate_output_15_211(.a(output_16_211), .b(output_16_4), .y(output_15_211));
wire output_1_212, output_1_5, output_0_212;
mixer gate_output_0_212(.a(output_1_212), .b(output_1_5), .y(output_0_212));
wire output_2_212, output_2_5, output_1_212;
mixer gate_output_1_212(.a(output_2_212), .b(output_2_5), .y(output_1_212));
wire output_3_212, output_3_5, output_2_212;
mixer gate_output_2_212(.a(output_3_212), .b(output_3_5), .y(output_2_212));
wire output_4_212, output_4_5, output_3_212;
mixer gate_output_3_212(.a(output_4_212), .b(output_4_5), .y(output_3_212));
wire output_5_212, output_5_5, output_4_212;
mixer gate_output_4_212(.a(output_5_212), .b(output_5_5), .y(output_4_212));
wire output_6_212, output_6_5, output_5_212;
mixer gate_output_5_212(.a(output_6_212), .b(output_6_5), .y(output_5_212));
wire output_7_212, output_7_5, output_6_212;
mixer gate_output_6_212(.a(output_7_212), .b(output_7_5), .y(output_6_212));
wire output_8_212, output_8_5, output_7_212;
mixer gate_output_7_212(.a(output_8_212), .b(output_8_5), .y(output_7_212));
wire output_9_212, output_9_5, output_8_212;
mixer gate_output_8_212(.a(output_9_212), .b(output_9_5), .y(output_8_212));
wire output_10_212, output_10_5, output_9_212;
mixer gate_output_9_212(.a(output_10_212), .b(output_10_5), .y(output_9_212));
wire output_11_212, output_11_5, output_10_212;
mixer gate_output_10_212(.a(output_11_212), .b(output_11_5), .y(output_10_212));
wire output_12_212, output_12_5, output_11_212;
mixer gate_output_11_212(.a(output_12_212), .b(output_12_5), .y(output_11_212));
wire output_13_212, output_13_5, output_12_212;
mixer gate_output_12_212(.a(output_13_212), .b(output_13_5), .y(output_12_212));
wire output_14_212, output_14_5, output_13_212;
mixer gate_output_13_212(.a(output_14_212), .b(output_14_5), .y(output_13_212));
wire output_15_212, output_15_5, output_14_212;
mixer gate_output_14_212(.a(output_15_212), .b(output_15_5), .y(output_14_212));
wire output_16_212, output_16_5, output_15_212;
mixer gate_output_15_212(.a(output_16_212), .b(output_16_5), .y(output_15_212));
wire output_1_213, output_1_6, output_0_213;
mixer gate_output_0_213(.a(output_1_213), .b(output_1_6), .y(output_0_213));
wire output_2_213, output_2_6, output_1_213;
mixer gate_output_1_213(.a(output_2_213), .b(output_2_6), .y(output_1_213));
wire output_3_213, output_3_6, output_2_213;
mixer gate_output_2_213(.a(output_3_213), .b(output_3_6), .y(output_2_213));
wire output_4_213, output_4_6, output_3_213;
mixer gate_output_3_213(.a(output_4_213), .b(output_4_6), .y(output_3_213));
wire output_5_213, output_5_6, output_4_213;
mixer gate_output_4_213(.a(output_5_213), .b(output_5_6), .y(output_4_213));
wire output_6_213, output_6_6, output_5_213;
mixer gate_output_5_213(.a(output_6_213), .b(output_6_6), .y(output_5_213));
wire output_7_213, output_7_6, output_6_213;
mixer gate_output_6_213(.a(output_7_213), .b(output_7_6), .y(output_6_213));
wire output_8_213, output_8_6, output_7_213;
mixer gate_output_7_213(.a(output_8_213), .b(output_8_6), .y(output_7_213));
wire output_9_213, output_9_6, output_8_213;
mixer gate_output_8_213(.a(output_9_213), .b(output_9_6), .y(output_8_213));
wire output_10_213, output_10_6, output_9_213;
mixer gate_output_9_213(.a(output_10_213), .b(output_10_6), .y(output_9_213));
wire output_11_213, output_11_6, output_10_213;
mixer gate_output_10_213(.a(output_11_213), .b(output_11_6), .y(output_10_213));
wire output_12_213, output_12_6, output_11_213;
mixer gate_output_11_213(.a(output_12_213), .b(output_12_6), .y(output_11_213));
wire output_13_213, output_13_6, output_12_213;
mixer gate_output_12_213(.a(output_13_213), .b(output_13_6), .y(output_12_213));
wire output_14_213, output_14_6, output_13_213;
mixer gate_output_13_213(.a(output_14_213), .b(output_14_6), .y(output_13_213));
wire output_15_213, output_15_6, output_14_213;
mixer gate_output_14_213(.a(output_15_213), .b(output_15_6), .y(output_14_213));
wire output_16_213, output_16_6, output_15_213;
mixer gate_output_15_213(.a(output_16_213), .b(output_16_6), .y(output_15_213));
wire output_1_214, output_1_7, output_0_214;
mixer gate_output_0_214(.a(output_1_214), .b(output_1_7), .y(output_0_214));
wire output_2_214, output_2_7, output_1_214;
mixer gate_output_1_214(.a(output_2_214), .b(output_2_7), .y(output_1_214));
wire output_3_214, output_3_7, output_2_214;
mixer gate_output_2_214(.a(output_3_214), .b(output_3_7), .y(output_2_214));
wire output_4_214, output_4_7, output_3_214;
mixer gate_output_3_214(.a(output_4_214), .b(output_4_7), .y(output_3_214));
wire output_5_214, output_5_7, output_4_214;
mixer gate_output_4_214(.a(output_5_214), .b(output_5_7), .y(output_4_214));
wire output_6_214, output_6_7, output_5_214;
mixer gate_output_5_214(.a(output_6_214), .b(output_6_7), .y(output_5_214));
wire output_7_214, output_7_7, output_6_214;
mixer gate_output_6_214(.a(output_7_214), .b(output_7_7), .y(output_6_214));
wire output_8_214, output_8_7, output_7_214;
mixer gate_output_7_214(.a(output_8_214), .b(output_8_7), .y(output_7_214));
wire output_9_214, output_9_7, output_8_214;
mixer gate_output_8_214(.a(output_9_214), .b(output_9_7), .y(output_8_214));
wire output_10_214, output_10_7, output_9_214;
mixer gate_output_9_214(.a(output_10_214), .b(output_10_7), .y(output_9_214));
wire output_11_214, output_11_7, output_10_214;
mixer gate_output_10_214(.a(output_11_214), .b(output_11_7), .y(output_10_214));
wire output_12_214, output_12_7, output_11_214;
mixer gate_output_11_214(.a(output_12_214), .b(output_12_7), .y(output_11_214));
wire output_13_214, output_13_7, output_12_214;
mixer gate_output_12_214(.a(output_13_214), .b(output_13_7), .y(output_12_214));
wire output_14_214, output_14_7, output_13_214;
mixer gate_output_13_214(.a(output_14_214), .b(output_14_7), .y(output_13_214));
wire output_15_214, output_15_7, output_14_214;
mixer gate_output_14_214(.a(output_15_214), .b(output_15_7), .y(output_14_214));
wire output_16_214, output_16_7, output_15_214;
mixer gate_output_15_214(.a(output_16_214), .b(output_16_7), .y(output_15_214));
wire output_1_215, output_1_8, output_0_215;
mixer gate_output_0_215(.a(output_1_215), .b(output_1_8), .y(output_0_215));
wire output_2_215, output_2_8, output_1_215;
mixer gate_output_1_215(.a(output_2_215), .b(output_2_8), .y(output_1_215));
wire output_3_215, output_3_8, output_2_215;
mixer gate_output_2_215(.a(output_3_215), .b(output_3_8), .y(output_2_215));
wire output_4_215, output_4_8, output_3_215;
mixer gate_output_3_215(.a(output_4_215), .b(output_4_8), .y(output_3_215));
wire output_5_215, output_5_8, output_4_215;
mixer gate_output_4_215(.a(output_5_215), .b(output_5_8), .y(output_4_215));
wire output_6_215, output_6_8, output_5_215;
mixer gate_output_5_215(.a(output_6_215), .b(output_6_8), .y(output_5_215));
wire output_7_215, output_7_8, output_6_215;
mixer gate_output_6_215(.a(output_7_215), .b(output_7_8), .y(output_6_215));
wire output_8_215, output_8_8, output_7_215;
mixer gate_output_7_215(.a(output_8_215), .b(output_8_8), .y(output_7_215));
wire output_9_215, output_9_8, output_8_215;
mixer gate_output_8_215(.a(output_9_215), .b(output_9_8), .y(output_8_215));
wire output_10_215, output_10_8, output_9_215;
mixer gate_output_9_215(.a(output_10_215), .b(output_10_8), .y(output_9_215));
wire output_11_215, output_11_8, output_10_215;
mixer gate_output_10_215(.a(output_11_215), .b(output_11_8), .y(output_10_215));
wire output_12_215, output_12_8, output_11_215;
mixer gate_output_11_215(.a(output_12_215), .b(output_12_8), .y(output_11_215));
wire output_13_215, output_13_8, output_12_215;
mixer gate_output_12_215(.a(output_13_215), .b(output_13_8), .y(output_12_215));
wire output_14_215, output_14_8, output_13_215;
mixer gate_output_13_215(.a(output_14_215), .b(output_14_8), .y(output_13_215));
wire output_15_215, output_15_8, output_14_215;
mixer gate_output_14_215(.a(output_15_215), .b(output_15_8), .y(output_14_215));
wire output_16_215, output_16_8, output_15_215;
mixer gate_output_15_215(.a(output_16_215), .b(output_16_8), .y(output_15_215));
wire output_1_216, output_1_9, output_0_216;
mixer gate_output_0_216(.a(output_1_216), .b(output_1_9), .y(output_0_216));
wire output_2_216, output_2_9, output_1_216;
mixer gate_output_1_216(.a(output_2_216), .b(output_2_9), .y(output_1_216));
wire output_3_216, output_3_9, output_2_216;
mixer gate_output_2_216(.a(output_3_216), .b(output_3_9), .y(output_2_216));
wire output_4_216, output_4_9, output_3_216;
mixer gate_output_3_216(.a(output_4_216), .b(output_4_9), .y(output_3_216));
wire output_5_216, output_5_9, output_4_216;
mixer gate_output_4_216(.a(output_5_216), .b(output_5_9), .y(output_4_216));
wire output_6_216, output_6_9, output_5_216;
mixer gate_output_5_216(.a(output_6_216), .b(output_6_9), .y(output_5_216));
wire output_7_216, output_7_9, output_6_216;
mixer gate_output_6_216(.a(output_7_216), .b(output_7_9), .y(output_6_216));
wire output_8_216, output_8_9, output_7_216;
mixer gate_output_7_216(.a(output_8_216), .b(output_8_9), .y(output_7_216));
wire output_9_216, output_9_9, output_8_216;
mixer gate_output_8_216(.a(output_9_216), .b(output_9_9), .y(output_8_216));
wire output_10_216, output_10_9, output_9_216;
mixer gate_output_9_216(.a(output_10_216), .b(output_10_9), .y(output_9_216));
wire output_11_216, output_11_9, output_10_216;
mixer gate_output_10_216(.a(output_11_216), .b(output_11_9), .y(output_10_216));
wire output_12_216, output_12_9, output_11_216;
mixer gate_output_11_216(.a(output_12_216), .b(output_12_9), .y(output_11_216));
wire output_13_216, output_13_9, output_12_216;
mixer gate_output_12_216(.a(output_13_216), .b(output_13_9), .y(output_12_216));
wire output_14_216, output_14_9, output_13_216;
mixer gate_output_13_216(.a(output_14_216), .b(output_14_9), .y(output_13_216));
wire output_15_216, output_15_9, output_14_216;
mixer gate_output_14_216(.a(output_15_216), .b(output_15_9), .y(output_14_216));
wire output_16_216, output_16_9, output_15_216;
mixer gate_output_15_216(.a(output_16_216), .b(output_16_9), .y(output_15_216));
wire output_1_217, output_1_10, output_0_217;
mixer gate_output_0_217(.a(output_1_217), .b(output_1_10), .y(output_0_217));
wire output_2_217, output_2_10, output_1_217;
mixer gate_output_1_217(.a(output_2_217), .b(output_2_10), .y(output_1_217));
wire output_3_217, output_3_10, output_2_217;
mixer gate_output_2_217(.a(output_3_217), .b(output_3_10), .y(output_2_217));
wire output_4_217, output_4_10, output_3_217;
mixer gate_output_3_217(.a(output_4_217), .b(output_4_10), .y(output_3_217));
wire output_5_217, output_5_10, output_4_217;
mixer gate_output_4_217(.a(output_5_217), .b(output_5_10), .y(output_4_217));
wire output_6_217, output_6_10, output_5_217;
mixer gate_output_5_217(.a(output_6_217), .b(output_6_10), .y(output_5_217));
wire output_7_217, output_7_10, output_6_217;
mixer gate_output_6_217(.a(output_7_217), .b(output_7_10), .y(output_6_217));
wire output_8_217, output_8_10, output_7_217;
mixer gate_output_7_217(.a(output_8_217), .b(output_8_10), .y(output_7_217));
wire output_9_217, output_9_10, output_8_217;
mixer gate_output_8_217(.a(output_9_217), .b(output_9_10), .y(output_8_217));
wire output_10_217, output_10_10, output_9_217;
mixer gate_output_9_217(.a(output_10_217), .b(output_10_10), .y(output_9_217));
wire output_11_217, output_11_10, output_10_217;
mixer gate_output_10_217(.a(output_11_217), .b(output_11_10), .y(output_10_217));
wire output_12_217, output_12_10, output_11_217;
mixer gate_output_11_217(.a(output_12_217), .b(output_12_10), .y(output_11_217));
wire output_13_217, output_13_10, output_12_217;
mixer gate_output_12_217(.a(output_13_217), .b(output_13_10), .y(output_12_217));
wire output_14_217, output_14_10, output_13_217;
mixer gate_output_13_217(.a(output_14_217), .b(output_14_10), .y(output_13_217));
wire output_15_217, output_15_10, output_14_217;
mixer gate_output_14_217(.a(output_15_217), .b(output_15_10), .y(output_14_217));
wire output_16_217, output_16_10, output_15_217;
mixer gate_output_15_217(.a(output_16_217), .b(output_16_10), .y(output_15_217));
wire output_1_218, output_1_11, output_0_218;
mixer gate_output_0_218(.a(output_1_218), .b(output_1_11), .y(output_0_218));
wire output_2_218, output_2_11, output_1_218;
mixer gate_output_1_218(.a(output_2_218), .b(output_2_11), .y(output_1_218));
wire output_3_218, output_3_11, output_2_218;
mixer gate_output_2_218(.a(output_3_218), .b(output_3_11), .y(output_2_218));
wire output_4_218, output_4_11, output_3_218;
mixer gate_output_3_218(.a(output_4_218), .b(output_4_11), .y(output_3_218));
wire output_5_218, output_5_11, output_4_218;
mixer gate_output_4_218(.a(output_5_218), .b(output_5_11), .y(output_4_218));
wire output_6_218, output_6_11, output_5_218;
mixer gate_output_5_218(.a(output_6_218), .b(output_6_11), .y(output_5_218));
wire output_7_218, output_7_11, output_6_218;
mixer gate_output_6_218(.a(output_7_218), .b(output_7_11), .y(output_6_218));
wire output_8_218, output_8_11, output_7_218;
mixer gate_output_7_218(.a(output_8_218), .b(output_8_11), .y(output_7_218));
wire output_9_218, output_9_11, output_8_218;
mixer gate_output_8_218(.a(output_9_218), .b(output_9_11), .y(output_8_218));
wire output_10_218, output_10_11, output_9_218;
mixer gate_output_9_218(.a(output_10_218), .b(output_10_11), .y(output_9_218));
wire output_11_218, output_11_11, output_10_218;
mixer gate_output_10_218(.a(output_11_218), .b(output_11_11), .y(output_10_218));
wire output_12_218, output_12_11, output_11_218;
mixer gate_output_11_218(.a(output_12_218), .b(output_12_11), .y(output_11_218));
wire output_13_218, output_13_11, output_12_218;
mixer gate_output_12_218(.a(output_13_218), .b(output_13_11), .y(output_12_218));
wire output_14_218, output_14_11, output_13_218;
mixer gate_output_13_218(.a(output_14_218), .b(output_14_11), .y(output_13_218));
wire output_15_218, output_15_11, output_14_218;
mixer gate_output_14_218(.a(output_15_218), .b(output_15_11), .y(output_14_218));
wire output_16_218, output_16_11, output_15_218;
mixer gate_output_15_218(.a(output_16_218), .b(output_16_11), .y(output_15_218));
wire output_1_219, output_1_12, output_0_219;
mixer gate_output_0_219(.a(output_1_219), .b(output_1_12), .y(output_0_219));
wire output_2_219, output_2_12, output_1_219;
mixer gate_output_1_219(.a(output_2_219), .b(output_2_12), .y(output_1_219));
wire output_3_219, output_3_12, output_2_219;
mixer gate_output_2_219(.a(output_3_219), .b(output_3_12), .y(output_2_219));
wire output_4_219, output_4_12, output_3_219;
mixer gate_output_3_219(.a(output_4_219), .b(output_4_12), .y(output_3_219));
wire output_5_219, output_5_12, output_4_219;
mixer gate_output_4_219(.a(output_5_219), .b(output_5_12), .y(output_4_219));
wire output_6_219, output_6_12, output_5_219;
mixer gate_output_5_219(.a(output_6_219), .b(output_6_12), .y(output_5_219));
wire output_7_219, output_7_12, output_6_219;
mixer gate_output_6_219(.a(output_7_219), .b(output_7_12), .y(output_6_219));
wire output_8_219, output_8_12, output_7_219;
mixer gate_output_7_219(.a(output_8_219), .b(output_8_12), .y(output_7_219));
wire output_9_219, output_9_12, output_8_219;
mixer gate_output_8_219(.a(output_9_219), .b(output_9_12), .y(output_8_219));
wire output_10_219, output_10_12, output_9_219;
mixer gate_output_9_219(.a(output_10_219), .b(output_10_12), .y(output_9_219));
wire output_11_219, output_11_12, output_10_219;
mixer gate_output_10_219(.a(output_11_219), .b(output_11_12), .y(output_10_219));
wire output_12_219, output_12_12, output_11_219;
mixer gate_output_11_219(.a(output_12_219), .b(output_12_12), .y(output_11_219));
wire output_13_219, output_13_12, output_12_219;
mixer gate_output_12_219(.a(output_13_219), .b(output_13_12), .y(output_12_219));
wire output_14_219, output_14_12, output_13_219;
mixer gate_output_13_219(.a(output_14_219), .b(output_14_12), .y(output_13_219));
wire output_15_219, output_15_12, output_14_219;
mixer gate_output_14_219(.a(output_15_219), .b(output_15_12), .y(output_14_219));
wire output_16_219, output_16_12, output_15_219;
mixer gate_output_15_219(.a(output_16_219), .b(output_16_12), .y(output_15_219));
wire output_1_220, output_1_13, output_0_220;
mixer gate_output_0_220(.a(output_1_220), .b(output_1_13), .y(output_0_220));
wire output_2_220, output_2_13, output_1_220;
mixer gate_output_1_220(.a(output_2_220), .b(output_2_13), .y(output_1_220));
wire output_3_220, output_3_13, output_2_220;
mixer gate_output_2_220(.a(output_3_220), .b(output_3_13), .y(output_2_220));
wire output_4_220, output_4_13, output_3_220;
mixer gate_output_3_220(.a(output_4_220), .b(output_4_13), .y(output_3_220));
wire output_5_220, output_5_13, output_4_220;
mixer gate_output_4_220(.a(output_5_220), .b(output_5_13), .y(output_4_220));
wire output_6_220, output_6_13, output_5_220;
mixer gate_output_5_220(.a(output_6_220), .b(output_6_13), .y(output_5_220));
wire output_7_220, output_7_13, output_6_220;
mixer gate_output_6_220(.a(output_7_220), .b(output_7_13), .y(output_6_220));
wire output_8_220, output_8_13, output_7_220;
mixer gate_output_7_220(.a(output_8_220), .b(output_8_13), .y(output_7_220));
wire output_9_220, output_9_13, output_8_220;
mixer gate_output_8_220(.a(output_9_220), .b(output_9_13), .y(output_8_220));
wire output_10_220, output_10_13, output_9_220;
mixer gate_output_9_220(.a(output_10_220), .b(output_10_13), .y(output_9_220));
wire output_11_220, output_11_13, output_10_220;
mixer gate_output_10_220(.a(output_11_220), .b(output_11_13), .y(output_10_220));
wire output_12_220, output_12_13, output_11_220;
mixer gate_output_11_220(.a(output_12_220), .b(output_12_13), .y(output_11_220));
wire output_13_220, output_13_13, output_12_220;
mixer gate_output_12_220(.a(output_13_220), .b(output_13_13), .y(output_12_220));
wire output_14_220, output_14_13, output_13_220;
mixer gate_output_13_220(.a(output_14_220), .b(output_14_13), .y(output_13_220));
wire output_15_220, output_15_13, output_14_220;
mixer gate_output_14_220(.a(output_15_220), .b(output_15_13), .y(output_14_220));
wire output_16_220, output_16_13, output_15_220;
mixer gate_output_15_220(.a(output_16_220), .b(output_16_13), .y(output_15_220));
wire output_1_221, output_1_14, output_0_221;
mixer gate_output_0_221(.a(output_1_221), .b(output_1_14), .y(output_0_221));
wire output_2_221, output_2_14, output_1_221;
mixer gate_output_1_221(.a(output_2_221), .b(output_2_14), .y(output_1_221));
wire output_3_221, output_3_14, output_2_221;
mixer gate_output_2_221(.a(output_3_221), .b(output_3_14), .y(output_2_221));
wire output_4_221, output_4_14, output_3_221;
mixer gate_output_3_221(.a(output_4_221), .b(output_4_14), .y(output_3_221));
wire output_5_221, output_5_14, output_4_221;
mixer gate_output_4_221(.a(output_5_221), .b(output_5_14), .y(output_4_221));
wire output_6_221, output_6_14, output_5_221;
mixer gate_output_5_221(.a(output_6_221), .b(output_6_14), .y(output_5_221));
wire output_7_221, output_7_14, output_6_221;
mixer gate_output_6_221(.a(output_7_221), .b(output_7_14), .y(output_6_221));
wire output_8_221, output_8_14, output_7_221;
mixer gate_output_7_221(.a(output_8_221), .b(output_8_14), .y(output_7_221));
wire output_9_221, output_9_14, output_8_221;
mixer gate_output_8_221(.a(output_9_221), .b(output_9_14), .y(output_8_221));
wire output_10_221, output_10_14, output_9_221;
mixer gate_output_9_221(.a(output_10_221), .b(output_10_14), .y(output_9_221));
wire output_11_221, output_11_14, output_10_221;
mixer gate_output_10_221(.a(output_11_221), .b(output_11_14), .y(output_10_221));
wire output_12_221, output_12_14, output_11_221;
mixer gate_output_11_221(.a(output_12_221), .b(output_12_14), .y(output_11_221));
wire output_13_221, output_13_14, output_12_221;
mixer gate_output_12_221(.a(output_13_221), .b(output_13_14), .y(output_12_221));
wire output_14_221, output_14_14, output_13_221;
mixer gate_output_13_221(.a(output_14_221), .b(output_14_14), .y(output_13_221));
wire output_15_221, output_15_14, output_14_221;
mixer gate_output_14_221(.a(output_15_221), .b(output_15_14), .y(output_14_221));
wire output_16_221, output_16_14, output_15_221;
mixer gate_output_15_221(.a(output_16_221), .b(output_16_14), .y(output_15_221));
wire output_1_222, output_1_15, output_0_222;
mixer gate_output_0_222(.a(output_1_222), .b(output_1_15), .y(output_0_222));
wire output_2_222, output_2_15, output_1_222;
mixer gate_output_1_222(.a(output_2_222), .b(output_2_15), .y(output_1_222));
wire output_3_222, output_3_15, output_2_222;
mixer gate_output_2_222(.a(output_3_222), .b(output_3_15), .y(output_2_222));
wire output_4_222, output_4_15, output_3_222;
mixer gate_output_3_222(.a(output_4_222), .b(output_4_15), .y(output_3_222));
wire output_5_222, output_5_15, output_4_222;
mixer gate_output_4_222(.a(output_5_222), .b(output_5_15), .y(output_4_222));
wire output_6_222, output_6_15, output_5_222;
mixer gate_output_5_222(.a(output_6_222), .b(output_6_15), .y(output_5_222));
wire output_7_222, output_7_15, output_6_222;
mixer gate_output_6_222(.a(output_7_222), .b(output_7_15), .y(output_6_222));
wire output_8_222, output_8_15, output_7_222;
mixer gate_output_7_222(.a(output_8_222), .b(output_8_15), .y(output_7_222));
wire output_9_222, output_9_15, output_8_222;
mixer gate_output_8_222(.a(output_9_222), .b(output_9_15), .y(output_8_222));
wire output_10_222, output_10_15, output_9_222;
mixer gate_output_9_222(.a(output_10_222), .b(output_10_15), .y(output_9_222));
wire output_11_222, output_11_15, output_10_222;
mixer gate_output_10_222(.a(output_11_222), .b(output_11_15), .y(output_10_222));
wire output_12_222, output_12_15, output_11_222;
mixer gate_output_11_222(.a(output_12_222), .b(output_12_15), .y(output_11_222));
wire output_13_222, output_13_15, output_12_222;
mixer gate_output_12_222(.a(output_13_222), .b(output_13_15), .y(output_12_222));
wire output_14_222, output_14_15, output_13_222;
mixer gate_output_13_222(.a(output_14_222), .b(output_14_15), .y(output_13_222));
wire output_15_222, output_15_15, output_14_222;
mixer gate_output_14_222(.a(output_15_222), .b(output_15_15), .y(output_14_222));
wire output_16_222, output_16_15, output_15_222;
mixer gate_output_15_222(.a(output_16_222), .b(output_16_15), .y(output_15_222));
wire output_1_223, output_1_0, output_0_223;
mixer gate_output_0_223(.a(output_1_223), .b(output_1_0), .y(output_0_223));
wire output_2_223, output_2_0, output_1_223;
mixer gate_output_1_223(.a(output_2_223), .b(output_2_0), .y(output_1_223));
wire output_3_223, output_3_0, output_2_223;
mixer gate_output_2_223(.a(output_3_223), .b(output_3_0), .y(output_2_223));
wire output_4_223, output_4_0, output_3_223;
mixer gate_output_3_223(.a(output_4_223), .b(output_4_0), .y(output_3_223));
wire output_5_223, output_5_0, output_4_223;
mixer gate_output_4_223(.a(output_5_223), .b(output_5_0), .y(output_4_223));
wire output_6_223, output_6_0, output_5_223;
mixer gate_output_5_223(.a(output_6_223), .b(output_6_0), .y(output_5_223));
wire output_7_223, output_7_0, output_6_223;
mixer gate_output_6_223(.a(output_7_223), .b(output_7_0), .y(output_6_223));
wire output_8_223, output_8_0, output_7_223;
mixer gate_output_7_223(.a(output_8_223), .b(output_8_0), .y(output_7_223));
wire output_9_223, output_9_0, output_8_223;
mixer gate_output_8_223(.a(output_9_223), .b(output_9_0), .y(output_8_223));
wire output_10_223, output_10_0, output_9_223;
mixer gate_output_9_223(.a(output_10_223), .b(output_10_0), .y(output_9_223));
wire output_11_223, output_11_0, output_10_223;
mixer gate_output_10_223(.a(output_11_223), .b(output_11_0), .y(output_10_223));
wire output_12_223, output_12_0, output_11_223;
mixer gate_output_11_223(.a(output_12_223), .b(output_12_0), .y(output_11_223));
wire output_13_223, output_13_0, output_12_223;
mixer gate_output_12_223(.a(output_13_223), .b(output_13_0), .y(output_12_223));
wire output_14_223, output_14_0, output_13_223;
mixer gate_output_13_223(.a(output_14_223), .b(output_14_0), .y(output_13_223));
wire output_15_223, output_15_0, output_14_223;
mixer gate_output_14_223(.a(output_15_223), .b(output_15_0), .y(output_14_223));
wire output_16_223, output_16_0, output_15_223;
mixer gate_output_15_223(.a(output_16_223), .b(output_16_0), .y(output_15_223));
wire output_1_224, output_1_1, output_0_224;
mixer gate_output_0_224(.a(output_1_224), .b(output_1_1), .y(output_0_224));
wire output_2_224, output_2_1, output_1_224;
mixer gate_output_1_224(.a(output_2_224), .b(output_2_1), .y(output_1_224));
wire output_3_224, output_3_1, output_2_224;
mixer gate_output_2_224(.a(output_3_224), .b(output_3_1), .y(output_2_224));
wire output_4_224, output_4_1, output_3_224;
mixer gate_output_3_224(.a(output_4_224), .b(output_4_1), .y(output_3_224));
wire output_5_224, output_5_1, output_4_224;
mixer gate_output_4_224(.a(output_5_224), .b(output_5_1), .y(output_4_224));
wire output_6_224, output_6_1, output_5_224;
mixer gate_output_5_224(.a(output_6_224), .b(output_6_1), .y(output_5_224));
wire output_7_224, output_7_1, output_6_224;
mixer gate_output_6_224(.a(output_7_224), .b(output_7_1), .y(output_6_224));
wire output_8_224, output_8_1, output_7_224;
mixer gate_output_7_224(.a(output_8_224), .b(output_8_1), .y(output_7_224));
wire output_9_224, output_9_1, output_8_224;
mixer gate_output_8_224(.a(output_9_224), .b(output_9_1), .y(output_8_224));
wire output_10_224, output_10_1, output_9_224;
mixer gate_output_9_224(.a(output_10_224), .b(output_10_1), .y(output_9_224));
wire output_11_224, output_11_1, output_10_224;
mixer gate_output_10_224(.a(output_11_224), .b(output_11_1), .y(output_10_224));
wire output_12_224, output_12_1, output_11_224;
mixer gate_output_11_224(.a(output_12_224), .b(output_12_1), .y(output_11_224));
wire output_13_224, output_13_1, output_12_224;
mixer gate_output_12_224(.a(output_13_224), .b(output_13_1), .y(output_12_224));
wire output_14_224, output_14_1, output_13_224;
mixer gate_output_13_224(.a(output_14_224), .b(output_14_1), .y(output_13_224));
wire output_15_224, output_15_1, output_14_224;
mixer gate_output_14_224(.a(output_15_224), .b(output_15_1), .y(output_14_224));
wire output_16_224, output_16_1, output_15_224;
mixer gate_output_15_224(.a(output_16_224), .b(output_16_1), .y(output_15_224));
wire output_1_225, output_1_2, output_0_225;
mixer gate_output_0_225(.a(output_1_225), .b(output_1_2), .y(output_0_225));
wire output_2_225, output_2_2, output_1_225;
mixer gate_output_1_225(.a(output_2_225), .b(output_2_2), .y(output_1_225));
wire output_3_225, output_3_2, output_2_225;
mixer gate_output_2_225(.a(output_3_225), .b(output_3_2), .y(output_2_225));
wire output_4_225, output_4_2, output_3_225;
mixer gate_output_3_225(.a(output_4_225), .b(output_4_2), .y(output_3_225));
wire output_5_225, output_5_2, output_4_225;
mixer gate_output_4_225(.a(output_5_225), .b(output_5_2), .y(output_4_225));
wire output_6_225, output_6_2, output_5_225;
mixer gate_output_5_225(.a(output_6_225), .b(output_6_2), .y(output_5_225));
wire output_7_225, output_7_2, output_6_225;
mixer gate_output_6_225(.a(output_7_225), .b(output_7_2), .y(output_6_225));
wire output_8_225, output_8_2, output_7_225;
mixer gate_output_7_225(.a(output_8_225), .b(output_8_2), .y(output_7_225));
wire output_9_225, output_9_2, output_8_225;
mixer gate_output_8_225(.a(output_9_225), .b(output_9_2), .y(output_8_225));
wire output_10_225, output_10_2, output_9_225;
mixer gate_output_9_225(.a(output_10_225), .b(output_10_2), .y(output_9_225));
wire output_11_225, output_11_2, output_10_225;
mixer gate_output_10_225(.a(output_11_225), .b(output_11_2), .y(output_10_225));
wire output_12_225, output_12_2, output_11_225;
mixer gate_output_11_225(.a(output_12_225), .b(output_12_2), .y(output_11_225));
wire output_13_225, output_13_2, output_12_225;
mixer gate_output_12_225(.a(output_13_225), .b(output_13_2), .y(output_12_225));
wire output_14_225, output_14_2, output_13_225;
mixer gate_output_13_225(.a(output_14_225), .b(output_14_2), .y(output_13_225));
wire output_15_225, output_15_2, output_14_225;
mixer gate_output_14_225(.a(output_15_225), .b(output_15_2), .y(output_14_225));
wire output_16_225, output_16_2, output_15_225;
mixer gate_output_15_225(.a(output_16_225), .b(output_16_2), .y(output_15_225));
wire output_1_226, output_1_3, output_0_226;
mixer gate_output_0_226(.a(output_1_226), .b(output_1_3), .y(output_0_226));
wire output_2_226, output_2_3, output_1_226;
mixer gate_output_1_226(.a(output_2_226), .b(output_2_3), .y(output_1_226));
wire output_3_226, output_3_3, output_2_226;
mixer gate_output_2_226(.a(output_3_226), .b(output_3_3), .y(output_2_226));
wire output_4_226, output_4_3, output_3_226;
mixer gate_output_3_226(.a(output_4_226), .b(output_4_3), .y(output_3_226));
wire output_5_226, output_5_3, output_4_226;
mixer gate_output_4_226(.a(output_5_226), .b(output_5_3), .y(output_4_226));
wire output_6_226, output_6_3, output_5_226;
mixer gate_output_5_226(.a(output_6_226), .b(output_6_3), .y(output_5_226));
wire output_7_226, output_7_3, output_6_226;
mixer gate_output_6_226(.a(output_7_226), .b(output_7_3), .y(output_6_226));
wire output_8_226, output_8_3, output_7_226;
mixer gate_output_7_226(.a(output_8_226), .b(output_8_3), .y(output_7_226));
wire output_9_226, output_9_3, output_8_226;
mixer gate_output_8_226(.a(output_9_226), .b(output_9_3), .y(output_8_226));
wire output_10_226, output_10_3, output_9_226;
mixer gate_output_9_226(.a(output_10_226), .b(output_10_3), .y(output_9_226));
wire output_11_226, output_11_3, output_10_226;
mixer gate_output_10_226(.a(output_11_226), .b(output_11_3), .y(output_10_226));
wire output_12_226, output_12_3, output_11_226;
mixer gate_output_11_226(.a(output_12_226), .b(output_12_3), .y(output_11_226));
wire output_13_226, output_13_3, output_12_226;
mixer gate_output_12_226(.a(output_13_226), .b(output_13_3), .y(output_12_226));
wire output_14_226, output_14_3, output_13_226;
mixer gate_output_13_226(.a(output_14_226), .b(output_14_3), .y(output_13_226));
wire output_15_226, output_15_3, output_14_226;
mixer gate_output_14_226(.a(output_15_226), .b(output_15_3), .y(output_14_226));
wire output_16_226, output_16_3, output_15_226;
mixer gate_output_15_226(.a(output_16_226), .b(output_16_3), .y(output_15_226));
wire output_1_227, output_1_4, output_0_227;
mixer gate_output_0_227(.a(output_1_227), .b(output_1_4), .y(output_0_227));
wire output_2_227, output_2_4, output_1_227;
mixer gate_output_1_227(.a(output_2_227), .b(output_2_4), .y(output_1_227));
wire output_3_227, output_3_4, output_2_227;
mixer gate_output_2_227(.a(output_3_227), .b(output_3_4), .y(output_2_227));
wire output_4_227, output_4_4, output_3_227;
mixer gate_output_3_227(.a(output_4_227), .b(output_4_4), .y(output_3_227));
wire output_5_227, output_5_4, output_4_227;
mixer gate_output_4_227(.a(output_5_227), .b(output_5_4), .y(output_4_227));
wire output_6_227, output_6_4, output_5_227;
mixer gate_output_5_227(.a(output_6_227), .b(output_6_4), .y(output_5_227));
wire output_7_227, output_7_4, output_6_227;
mixer gate_output_6_227(.a(output_7_227), .b(output_7_4), .y(output_6_227));
wire output_8_227, output_8_4, output_7_227;
mixer gate_output_7_227(.a(output_8_227), .b(output_8_4), .y(output_7_227));
wire output_9_227, output_9_4, output_8_227;
mixer gate_output_8_227(.a(output_9_227), .b(output_9_4), .y(output_8_227));
wire output_10_227, output_10_4, output_9_227;
mixer gate_output_9_227(.a(output_10_227), .b(output_10_4), .y(output_9_227));
wire output_11_227, output_11_4, output_10_227;
mixer gate_output_10_227(.a(output_11_227), .b(output_11_4), .y(output_10_227));
wire output_12_227, output_12_4, output_11_227;
mixer gate_output_11_227(.a(output_12_227), .b(output_12_4), .y(output_11_227));
wire output_13_227, output_13_4, output_12_227;
mixer gate_output_12_227(.a(output_13_227), .b(output_13_4), .y(output_12_227));
wire output_14_227, output_14_4, output_13_227;
mixer gate_output_13_227(.a(output_14_227), .b(output_14_4), .y(output_13_227));
wire output_15_227, output_15_4, output_14_227;
mixer gate_output_14_227(.a(output_15_227), .b(output_15_4), .y(output_14_227));
wire output_16_227, output_16_4, output_15_227;
mixer gate_output_15_227(.a(output_16_227), .b(output_16_4), .y(output_15_227));
wire output_1_228, output_1_5, output_0_228;
mixer gate_output_0_228(.a(output_1_228), .b(output_1_5), .y(output_0_228));
wire output_2_228, output_2_5, output_1_228;
mixer gate_output_1_228(.a(output_2_228), .b(output_2_5), .y(output_1_228));
wire output_3_228, output_3_5, output_2_228;
mixer gate_output_2_228(.a(output_3_228), .b(output_3_5), .y(output_2_228));
wire output_4_228, output_4_5, output_3_228;
mixer gate_output_3_228(.a(output_4_228), .b(output_4_5), .y(output_3_228));
wire output_5_228, output_5_5, output_4_228;
mixer gate_output_4_228(.a(output_5_228), .b(output_5_5), .y(output_4_228));
wire output_6_228, output_6_5, output_5_228;
mixer gate_output_5_228(.a(output_6_228), .b(output_6_5), .y(output_5_228));
wire output_7_228, output_7_5, output_6_228;
mixer gate_output_6_228(.a(output_7_228), .b(output_7_5), .y(output_6_228));
wire output_8_228, output_8_5, output_7_228;
mixer gate_output_7_228(.a(output_8_228), .b(output_8_5), .y(output_7_228));
wire output_9_228, output_9_5, output_8_228;
mixer gate_output_8_228(.a(output_9_228), .b(output_9_5), .y(output_8_228));
wire output_10_228, output_10_5, output_9_228;
mixer gate_output_9_228(.a(output_10_228), .b(output_10_5), .y(output_9_228));
wire output_11_228, output_11_5, output_10_228;
mixer gate_output_10_228(.a(output_11_228), .b(output_11_5), .y(output_10_228));
wire output_12_228, output_12_5, output_11_228;
mixer gate_output_11_228(.a(output_12_228), .b(output_12_5), .y(output_11_228));
wire output_13_228, output_13_5, output_12_228;
mixer gate_output_12_228(.a(output_13_228), .b(output_13_5), .y(output_12_228));
wire output_14_228, output_14_5, output_13_228;
mixer gate_output_13_228(.a(output_14_228), .b(output_14_5), .y(output_13_228));
wire output_15_228, output_15_5, output_14_228;
mixer gate_output_14_228(.a(output_15_228), .b(output_15_5), .y(output_14_228));
wire output_16_228, output_16_5, output_15_228;
mixer gate_output_15_228(.a(output_16_228), .b(output_16_5), .y(output_15_228));
wire output_1_229, output_1_6, output_0_229;
mixer gate_output_0_229(.a(output_1_229), .b(output_1_6), .y(output_0_229));
wire output_2_229, output_2_6, output_1_229;
mixer gate_output_1_229(.a(output_2_229), .b(output_2_6), .y(output_1_229));
wire output_3_229, output_3_6, output_2_229;
mixer gate_output_2_229(.a(output_3_229), .b(output_3_6), .y(output_2_229));
wire output_4_229, output_4_6, output_3_229;
mixer gate_output_3_229(.a(output_4_229), .b(output_4_6), .y(output_3_229));
wire output_5_229, output_5_6, output_4_229;
mixer gate_output_4_229(.a(output_5_229), .b(output_5_6), .y(output_4_229));
wire output_6_229, output_6_6, output_5_229;
mixer gate_output_5_229(.a(output_6_229), .b(output_6_6), .y(output_5_229));
wire output_7_229, output_7_6, output_6_229;
mixer gate_output_6_229(.a(output_7_229), .b(output_7_6), .y(output_6_229));
wire output_8_229, output_8_6, output_7_229;
mixer gate_output_7_229(.a(output_8_229), .b(output_8_6), .y(output_7_229));
wire output_9_229, output_9_6, output_8_229;
mixer gate_output_8_229(.a(output_9_229), .b(output_9_6), .y(output_8_229));
wire output_10_229, output_10_6, output_9_229;
mixer gate_output_9_229(.a(output_10_229), .b(output_10_6), .y(output_9_229));
wire output_11_229, output_11_6, output_10_229;
mixer gate_output_10_229(.a(output_11_229), .b(output_11_6), .y(output_10_229));
wire output_12_229, output_12_6, output_11_229;
mixer gate_output_11_229(.a(output_12_229), .b(output_12_6), .y(output_11_229));
wire output_13_229, output_13_6, output_12_229;
mixer gate_output_12_229(.a(output_13_229), .b(output_13_6), .y(output_12_229));
wire output_14_229, output_14_6, output_13_229;
mixer gate_output_13_229(.a(output_14_229), .b(output_14_6), .y(output_13_229));
wire output_15_229, output_15_6, output_14_229;
mixer gate_output_14_229(.a(output_15_229), .b(output_15_6), .y(output_14_229));
wire output_16_229, output_16_6, output_15_229;
mixer gate_output_15_229(.a(output_16_229), .b(output_16_6), .y(output_15_229));
wire output_1_230, output_1_7, output_0_230;
mixer gate_output_0_230(.a(output_1_230), .b(output_1_7), .y(output_0_230));
wire output_2_230, output_2_7, output_1_230;
mixer gate_output_1_230(.a(output_2_230), .b(output_2_7), .y(output_1_230));
wire output_3_230, output_3_7, output_2_230;
mixer gate_output_2_230(.a(output_3_230), .b(output_3_7), .y(output_2_230));
wire output_4_230, output_4_7, output_3_230;
mixer gate_output_3_230(.a(output_4_230), .b(output_4_7), .y(output_3_230));
wire output_5_230, output_5_7, output_4_230;
mixer gate_output_4_230(.a(output_5_230), .b(output_5_7), .y(output_4_230));
wire output_6_230, output_6_7, output_5_230;
mixer gate_output_5_230(.a(output_6_230), .b(output_6_7), .y(output_5_230));
wire output_7_230, output_7_7, output_6_230;
mixer gate_output_6_230(.a(output_7_230), .b(output_7_7), .y(output_6_230));
wire output_8_230, output_8_7, output_7_230;
mixer gate_output_7_230(.a(output_8_230), .b(output_8_7), .y(output_7_230));
wire output_9_230, output_9_7, output_8_230;
mixer gate_output_8_230(.a(output_9_230), .b(output_9_7), .y(output_8_230));
wire output_10_230, output_10_7, output_9_230;
mixer gate_output_9_230(.a(output_10_230), .b(output_10_7), .y(output_9_230));
wire output_11_230, output_11_7, output_10_230;
mixer gate_output_10_230(.a(output_11_230), .b(output_11_7), .y(output_10_230));
wire output_12_230, output_12_7, output_11_230;
mixer gate_output_11_230(.a(output_12_230), .b(output_12_7), .y(output_11_230));
wire output_13_230, output_13_7, output_12_230;
mixer gate_output_12_230(.a(output_13_230), .b(output_13_7), .y(output_12_230));
wire output_14_230, output_14_7, output_13_230;
mixer gate_output_13_230(.a(output_14_230), .b(output_14_7), .y(output_13_230));
wire output_15_230, output_15_7, output_14_230;
mixer gate_output_14_230(.a(output_15_230), .b(output_15_7), .y(output_14_230));
wire output_16_230, output_16_7, output_15_230;
mixer gate_output_15_230(.a(output_16_230), .b(output_16_7), .y(output_15_230));
wire output_1_231, output_1_8, output_0_231;
mixer gate_output_0_231(.a(output_1_231), .b(output_1_8), .y(output_0_231));
wire output_2_231, output_2_8, output_1_231;
mixer gate_output_1_231(.a(output_2_231), .b(output_2_8), .y(output_1_231));
wire output_3_231, output_3_8, output_2_231;
mixer gate_output_2_231(.a(output_3_231), .b(output_3_8), .y(output_2_231));
wire output_4_231, output_4_8, output_3_231;
mixer gate_output_3_231(.a(output_4_231), .b(output_4_8), .y(output_3_231));
wire output_5_231, output_5_8, output_4_231;
mixer gate_output_4_231(.a(output_5_231), .b(output_5_8), .y(output_4_231));
wire output_6_231, output_6_8, output_5_231;
mixer gate_output_5_231(.a(output_6_231), .b(output_6_8), .y(output_5_231));
wire output_7_231, output_7_8, output_6_231;
mixer gate_output_6_231(.a(output_7_231), .b(output_7_8), .y(output_6_231));
wire output_8_231, output_8_8, output_7_231;
mixer gate_output_7_231(.a(output_8_231), .b(output_8_8), .y(output_7_231));
wire output_9_231, output_9_8, output_8_231;
mixer gate_output_8_231(.a(output_9_231), .b(output_9_8), .y(output_8_231));
wire output_10_231, output_10_8, output_9_231;
mixer gate_output_9_231(.a(output_10_231), .b(output_10_8), .y(output_9_231));
wire output_11_231, output_11_8, output_10_231;
mixer gate_output_10_231(.a(output_11_231), .b(output_11_8), .y(output_10_231));
wire output_12_231, output_12_8, output_11_231;
mixer gate_output_11_231(.a(output_12_231), .b(output_12_8), .y(output_11_231));
wire output_13_231, output_13_8, output_12_231;
mixer gate_output_12_231(.a(output_13_231), .b(output_13_8), .y(output_12_231));
wire output_14_231, output_14_8, output_13_231;
mixer gate_output_13_231(.a(output_14_231), .b(output_14_8), .y(output_13_231));
wire output_15_231, output_15_8, output_14_231;
mixer gate_output_14_231(.a(output_15_231), .b(output_15_8), .y(output_14_231));
wire output_16_231, output_16_8, output_15_231;
mixer gate_output_15_231(.a(output_16_231), .b(output_16_8), .y(output_15_231));
wire output_1_232, output_1_9, output_0_232;
mixer gate_output_0_232(.a(output_1_232), .b(output_1_9), .y(output_0_232));
wire output_2_232, output_2_9, output_1_232;
mixer gate_output_1_232(.a(output_2_232), .b(output_2_9), .y(output_1_232));
wire output_3_232, output_3_9, output_2_232;
mixer gate_output_2_232(.a(output_3_232), .b(output_3_9), .y(output_2_232));
wire output_4_232, output_4_9, output_3_232;
mixer gate_output_3_232(.a(output_4_232), .b(output_4_9), .y(output_3_232));
wire output_5_232, output_5_9, output_4_232;
mixer gate_output_4_232(.a(output_5_232), .b(output_5_9), .y(output_4_232));
wire output_6_232, output_6_9, output_5_232;
mixer gate_output_5_232(.a(output_6_232), .b(output_6_9), .y(output_5_232));
wire output_7_232, output_7_9, output_6_232;
mixer gate_output_6_232(.a(output_7_232), .b(output_7_9), .y(output_6_232));
wire output_8_232, output_8_9, output_7_232;
mixer gate_output_7_232(.a(output_8_232), .b(output_8_9), .y(output_7_232));
wire output_9_232, output_9_9, output_8_232;
mixer gate_output_8_232(.a(output_9_232), .b(output_9_9), .y(output_8_232));
wire output_10_232, output_10_9, output_9_232;
mixer gate_output_9_232(.a(output_10_232), .b(output_10_9), .y(output_9_232));
wire output_11_232, output_11_9, output_10_232;
mixer gate_output_10_232(.a(output_11_232), .b(output_11_9), .y(output_10_232));
wire output_12_232, output_12_9, output_11_232;
mixer gate_output_11_232(.a(output_12_232), .b(output_12_9), .y(output_11_232));
wire output_13_232, output_13_9, output_12_232;
mixer gate_output_12_232(.a(output_13_232), .b(output_13_9), .y(output_12_232));
wire output_14_232, output_14_9, output_13_232;
mixer gate_output_13_232(.a(output_14_232), .b(output_14_9), .y(output_13_232));
wire output_15_232, output_15_9, output_14_232;
mixer gate_output_14_232(.a(output_15_232), .b(output_15_9), .y(output_14_232));
wire output_16_232, output_16_9, output_15_232;
mixer gate_output_15_232(.a(output_16_232), .b(output_16_9), .y(output_15_232));
wire output_1_233, output_1_10, output_0_233;
mixer gate_output_0_233(.a(output_1_233), .b(output_1_10), .y(output_0_233));
wire output_2_233, output_2_10, output_1_233;
mixer gate_output_1_233(.a(output_2_233), .b(output_2_10), .y(output_1_233));
wire output_3_233, output_3_10, output_2_233;
mixer gate_output_2_233(.a(output_3_233), .b(output_3_10), .y(output_2_233));
wire output_4_233, output_4_10, output_3_233;
mixer gate_output_3_233(.a(output_4_233), .b(output_4_10), .y(output_3_233));
wire output_5_233, output_5_10, output_4_233;
mixer gate_output_4_233(.a(output_5_233), .b(output_5_10), .y(output_4_233));
wire output_6_233, output_6_10, output_5_233;
mixer gate_output_5_233(.a(output_6_233), .b(output_6_10), .y(output_5_233));
wire output_7_233, output_7_10, output_6_233;
mixer gate_output_6_233(.a(output_7_233), .b(output_7_10), .y(output_6_233));
wire output_8_233, output_8_10, output_7_233;
mixer gate_output_7_233(.a(output_8_233), .b(output_8_10), .y(output_7_233));
wire output_9_233, output_9_10, output_8_233;
mixer gate_output_8_233(.a(output_9_233), .b(output_9_10), .y(output_8_233));
wire output_10_233, output_10_10, output_9_233;
mixer gate_output_9_233(.a(output_10_233), .b(output_10_10), .y(output_9_233));
wire output_11_233, output_11_10, output_10_233;
mixer gate_output_10_233(.a(output_11_233), .b(output_11_10), .y(output_10_233));
wire output_12_233, output_12_10, output_11_233;
mixer gate_output_11_233(.a(output_12_233), .b(output_12_10), .y(output_11_233));
wire output_13_233, output_13_10, output_12_233;
mixer gate_output_12_233(.a(output_13_233), .b(output_13_10), .y(output_12_233));
wire output_14_233, output_14_10, output_13_233;
mixer gate_output_13_233(.a(output_14_233), .b(output_14_10), .y(output_13_233));
wire output_15_233, output_15_10, output_14_233;
mixer gate_output_14_233(.a(output_15_233), .b(output_15_10), .y(output_14_233));
wire output_16_233, output_16_10, output_15_233;
mixer gate_output_15_233(.a(output_16_233), .b(output_16_10), .y(output_15_233));
wire output_1_234, output_1_11, output_0_234;
mixer gate_output_0_234(.a(output_1_234), .b(output_1_11), .y(output_0_234));
wire output_2_234, output_2_11, output_1_234;
mixer gate_output_1_234(.a(output_2_234), .b(output_2_11), .y(output_1_234));
wire output_3_234, output_3_11, output_2_234;
mixer gate_output_2_234(.a(output_3_234), .b(output_3_11), .y(output_2_234));
wire output_4_234, output_4_11, output_3_234;
mixer gate_output_3_234(.a(output_4_234), .b(output_4_11), .y(output_3_234));
wire output_5_234, output_5_11, output_4_234;
mixer gate_output_4_234(.a(output_5_234), .b(output_5_11), .y(output_4_234));
wire output_6_234, output_6_11, output_5_234;
mixer gate_output_5_234(.a(output_6_234), .b(output_6_11), .y(output_5_234));
wire output_7_234, output_7_11, output_6_234;
mixer gate_output_6_234(.a(output_7_234), .b(output_7_11), .y(output_6_234));
wire output_8_234, output_8_11, output_7_234;
mixer gate_output_7_234(.a(output_8_234), .b(output_8_11), .y(output_7_234));
wire output_9_234, output_9_11, output_8_234;
mixer gate_output_8_234(.a(output_9_234), .b(output_9_11), .y(output_8_234));
wire output_10_234, output_10_11, output_9_234;
mixer gate_output_9_234(.a(output_10_234), .b(output_10_11), .y(output_9_234));
wire output_11_234, output_11_11, output_10_234;
mixer gate_output_10_234(.a(output_11_234), .b(output_11_11), .y(output_10_234));
wire output_12_234, output_12_11, output_11_234;
mixer gate_output_11_234(.a(output_12_234), .b(output_12_11), .y(output_11_234));
wire output_13_234, output_13_11, output_12_234;
mixer gate_output_12_234(.a(output_13_234), .b(output_13_11), .y(output_12_234));
wire output_14_234, output_14_11, output_13_234;
mixer gate_output_13_234(.a(output_14_234), .b(output_14_11), .y(output_13_234));
wire output_15_234, output_15_11, output_14_234;
mixer gate_output_14_234(.a(output_15_234), .b(output_15_11), .y(output_14_234));
wire output_16_234, output_16_11, output_15_234;
mixer gate_output_15_234(.a(output_16_234), .b(output_16_11), .y(output_15_234));
wire output_1_235, output_1_12, output_0_235;
mixer gate_output_0_235(.a(output_1_235), .b(output_1_12), .y(output_0_235));
wire output_2_235, output_2_12, output_1_235;
mixer gate_output_1_235(.a(output_2_235), .b(output_2_12), .y(output_1_235));
wire output_3_235, output_3_12, output_2_235;
mixer gate_output_2_235(.a(output_3_235), .b(output_3_12), .y(output_2_235));
wire output_4_235, output_4_12, output_3_235;
mixer gate_output_3_235(.a(output_4_235), .b(output_4_12), .y(output_3_235));
wire output_5_235, output_5_12, output_4_235;
mixer gate_output_4_235(.a(output_5_235), .b(output_5_12), .y(output_4_235));
wire output_6_235, output_6_12, output_5_235;
mixer gate_output_5_235(.a(output_6_235), .b(output_6_12), .y(output_5_235));
wire output_7_235, output_7_12, output_6_235;
mixer gate_output_6_235(.a(output_7_235), .b(output_7_12), .y(output_6_235));
wire output_8_235, output_8_12, output_7_235;
mixer gate_output_7_235(.a(output_8_235), .b(output_8_12), .y(output_7_235));
wire output_9_235, output_9_12, output_8_235;
mixer gate_output_8_235(.a(output_9_235), .b(output_9_12), .y(output_8_235));
wire output_10_235, output_10_12, output_9_235;
mixer gate_output_9_235(.a(output_10_235), .b(output_10_12), .y(output_9_235));
wire output_11_235, output_11_12, output_10_235;
mixer gate_output_10_235(.a(output_11_235), .b(output_11_12), .y(output_10_235));
wire output_12_235, output_12_12, output_11_235;
mixer gate_output_11_235(.a(output_12_235), .b(output_12_12), .y(output_11_235));
wire output_13_235, output_13_12, output_12_235;
mixer gate_output_12_235(.a(output_13_235), .b(output_13_12), .y(output_12_235));
wire output_14_235, output_14_12, output_13_235;
mixer gate_output_13_235(.a(output_14_235), .b(output_14_12), .y(output_13_235));
wire output_15_235, output_15_12, output_14_235;
mixer gate_output_14_235(.a(output_15_235), .b(output_15_12), .y(output_14_235));
wire output_16_235, output_16_12, output_15_235;
mixer gate_output_15_235(.a(output_16_235), .b(output_16_12), .y(output_15_235));
wire output_1_236, output_1_13, output_0_236;
mixer gate_output_0_236(.a(output_1_236), .b(output_1_13), .y(output_0_236));
wire output_2_236, output_2_13, output_1_236;
mixer gate_output_1_236(.a(output_2_236), .b(output_2_13), .y(output_1_236));
wire output_3_236, output_3_13, output_2_236;
mixer gate_output_2_236(.a(output_3_236), .b(output_3_13), .y(output_2_236));
wire output_4_236, output_4_13, output_3_236;
mixer gate_output_3_236(.a(output_4_236), .b(output_4_13), .y(output_3_236));
wire output_5_236, output_5_13, output_4_236;
mixer gate_output_4_236(.a(output_5_236), .b(output_5_13), .y(output_4_236));
wire output_6_236, output_6_13, output_5_236;
mixer gate_output_5_236(.a(output_6_236), .b(output_6_13), .y(output_5_236));
wire output_7_236, output_7_13, output_6_236;
mixer gate_output_6_236(.a(output_7_236), .b(output_7_13), .y(output_6_236));
wire output_8_236, output_8_13, output_7_236;
mixer gate_output_7_236(.a(output_8_236), .b(output_8_13), .y(output_7_236));
wire output_9_236, output_9_13, output_8_236;
mixer gate_output_8_236(.a(output_9_236), .b(output_9_13), .y(output_8_236));
wire output_10_236, output_10_13, output_9_236;
mixer gate_output_9_236(.a(output_10_236), .b(output_10_13), .y(output_9_236));
wire output_11_236, output_11_13, output_10_236;
mixer gate_output_10_236(.a(output_11_236), .b(output_11_13), .y(output_10_236));
wire output_12_236, output_12_13, output_11_236;
mixer gate_output_11_236(.a(output_12_236), .b(output_12_13), .y(output_11_236));
wire output_13_236, output_13_13, output_12_236;
mixer gate_output_12_236(.a(output_13_236), .b(output_13_13), .y(output_12_236));
wire output_14_236, output_14_13, output_13_236;
mixer gate_output_13_236(.a(output_14_236), .b(output_14_13), .y(output_13_236));
wire output_15_236, output_15_13, output_14_236;
mixer gate_output_14_236(.a(output_15_236), .b(output_15_13), .y(output_14_236));
wire output_16_236, output_16_13, output_15_236;
mixer gate_output_15_236(.a(output_16_236), .b(output_16_13), .y(output_15_236));
wire output_1_237, output_1_14, output_0_237;
mixer gate_output_0_237(.a(output_1_237), .b(output_1_14), .y(output_0_237));
wire output_2_237, output_2_14, output_1_237;
mixer gate_output_1_237(.a(output_2_237), .b(output_2_14), .y(output_1_237));
wire output_3_237, output_3_14, output_2_237;
mixer gate_output_2_237(.a(output_3_237), .b(output_3_14), .y(output_2_237));
wire output_4_237, output_4_14, output_3_237;
mixer gate_output_3_237(.a(output_4_237), .b(output_4_14), .y(output_3_237));
wire output_5_237, output_5_14, output_4_237;
mixer gate_output_4_237(.a(output_5_237), .b(output_5_14), .y(output_4_237));
wire output_6_237, output_6_14, output_5_237;
mixer gate_output_5_237(.a(output_6_237), .b(output_6_14), .y(output_5_237));
wire output_7_237, output_7_14, output_6_237;
mixer gate_output_6_237(.a(output_7_237), .b(output_7_14), .y(output_6_237));
wire output_8_237, output_8_14, output_7_237;
mixer gate_output_7_237(.a(output_8_237), .b(output_8_14), .y(output_7_237));
wire output_9_237, output_9_14, output_8_237;
mixer gate_output_8_237(.a(output_9_237), .b(output_9_14), .y(output_8_237));
wire output_10_237, output_10_14, output_9_237;
mixer gate_output_9_237(.a(output_10_237), .b(output_10_14), .y(output_9_237));
wire output_11_237, output_11_14, output_10_237;
mixer gate_output_10_237(.a(output_11_237), .b(output_11_14), .y(output_10_237));
wire output_12_237, output_12_14, output_11_237;
mixer gate_output_11_237(.a(output_12_237), .b(output_12_14), .y(output_11_237));
wire output_13_237, output_13_14, output_12_237;
mixer gate_output_12_237(.a(output_13_237), .b(output_13_14), .y(output_12_237));
wire output_14_237, output_14_14, output_13_237;
mixer gate_output_13_237(.a(output_14_237), .b(output_14_14), .y(output_13_237));
wire output_15_237, output_15_14, output_14_237;
mixer gate_output_14_237(.a(output_15_237), .b(output_15_14), .y(output_14_237));
wire output_16_237, output_16_14, output_15_237;
mixer gate_output_15_237(.a(output_16_237), .b(output_16_14), .y(output_15_237));
wire output_1_238, output_1_15, output_0_238;
mixer gate_output_0_238(.a(output_1_238), .b(output_1_15), .y(output_0_238));
wire output_2_238, output_2_15, output_1_238;
mixer gate_output_1_238(.a(output_2_238), .b(output_2_15), .y(output_1_238));
wire output_3_238, output_3_15, output_2_238;
mixer gate_output_2_238(.a(output_3_238), .b(output_3_15), .y(output_2_238));
wire output_4_238, output_4_15, output_3_238;
mixer gate_output_3_238(.a(output_4_238), .b(output_4_15), .y(output_3_238));
wire output_5_238, output_5_15, output_4_238;
mixer gate_output_4_238(.a(output_5_238), .b(output_5_15), .y(output_4_238));
wire output_6_238, output_6_15, output_5_238;
mixer gate_output_5_238(.a(output_6_238), .b(output_6_15), .y(output_5_238));
wire output_7_238, output_7_15, output_6_238;
mixer gate_output_6_238(.a(output_7_238), .b(output_7_15), .y(output_6_238));
wire output_8_238, output_8_15, output_7_238;
mixer gate_output_7_238(.a(output_8_238), .b(output_8_15), .y(output_7_238));
wire output_9_238, output_9_15, output_8_238;
mixer gate_output_8_238(.a(output_9_238), .b(output_9_15), .y(output_8_238));
wire output_10_238, output_10_15, output_9_238;
mixer gate_output_9_238(.a(output_10_238), .b(output_10_15), .y(output_9_238));
wire output_11_238, output_11_15, output_10_238;
mixer gate_output_10_238(.a(output_11_238), .b(output_11_15), .y(output_10_238));
wire output_12_238, output_12_15, output_11_238;
mixer gate_output_11_238(.a(output_12_238), .b(output_12_15), .y(output_11_238));
wire output_13_238, output_13_15, output_12_238;
mixer gate_output_12_238(.a(output_13_238), .b(output_13_15), .y(output_12_238));
wire output_14_238, output_14_15, output_13_238;
mixer gate_output_13_238(.a(output_14_238), .b(output_14_15), .y(output_13_238));
wire output_15_238, output_15_15, output_14_238;
mixer gate_output_14_238(.a(output_15_238), .b(output_15_15), .y(output_14_238));
wire output_16_238, output_16_15, output_15_238;
mixer gate_output_15_238(.a(output_16_238), .b(output_16_15), .y(output_15_238));
wire output_1_239, output_1_0, output_0_239;
mixer gate_output_0_239(.a(output_1_239), .b(output_1_0), .y(output_0_239));
wire output_2_239, output_2_0, output_1_239;
mixer gate_output_1_239(.a(output_2_239), .b(output_2_0), .y(output_1_239));
wire output_3_239, output_3_0, output_2_239;
mixer gate_output_2_239(.a(output_3_239), .b(output_3_0), .y(output_2_239));
wire output_4_239, output_4_0, output_3_239;
mixer gate_output_3_239(.a(output_4_239), .b(output_4_0), .y(output_3_239));
wire output_5_239, output_5_0, output_4_239;
mixer gate_output_4_239(.a(output_5_239), .b(output_5_0), .y(output_4_239));
wire output_6_239, output_6_0, output_5_239;
mixer gate_output_5_239(.a(output_6_239), .b(output_6_0), .y(output_5_239));
wire output_7_239, output_7_0, output_6_239;
mixer gate_output_6_239(.a(output_7_239), .b(output_7_0), .y(output_6_239));
wire output_8_239, output_8_0, output_7_239;
mixer gate_output_7_239(.a(output_8_239), .b(output_8_0), .y(output_7_239));
wire output_9_239, output_9_0, output_8_239;
mixer gate_output_8_239(.a(output_9_239), .b(output_9_0), .y(output_8_239));
wire output_10_239, output_10_0, output_9_239;
mixer gate_output_9_239(.a(output_10_239), .b(output_10_0), .y(output_9_239));
wire output_11_239, output_11_0, output_10_239;
mixer gate_output_10_239(.a(output_11_239), .b(output_11_0), .y(output_10_239));
wire output_12_239, output_12_0, output_11_239;
mixer gate_output_11_239(.a(output_12_239), .b(output_12_0), .y(output_11_239));
wire output_13_239, output_13_0, output_12_239;
mixer gate_output_12_239(.a(output_13_239), .b(output_13_0), .y(output_12_239));
wire output_14_239, output_14_0, output_13_239;
mixer gate_output_13_239(.a(output_14_239), .b(output_14_0), .y(output_13_239));
wire output_15_239, output_15_0, output_14_239;
mixer gate_output_14_239(.a(output_15_239), .b(output_15_0), .y(output_14_239));
wire output_16_239, output_16_0, output_15_239;
mixer gate_output_15_239(.a(output_16_239), .b(output_16_0), .y(output_15_239));
wire output_1_240, output_1_1, output_0_240;
mixer gate_output_0_240(.a(output_1_240), .b(output_1_1), .y(output_0_240));
wire output_2_240, output_2_1, output_1_240;
mixer gate_output_1_240(.a(output_2_240), .b(output_2_1), .y(output_1_240));
wire output_3_240, output_3_1, output_2_240;
mixer gate_output_2_240(.a(output_3_240), .b(output_3_1), .y(output_2_240));
wire output_4_240, output_4_1, output_3_240;
mixer gate_output_3_240(.a(output_4_240), .b(output_4_1), .y(output_3_240));
wire output_5_240, output_5_1, output_4_240;
mixer gate_output_4_240(.a(output_5_240), .b(output_5_1), .y(output_4_240));
wire output_6_240, output_6_1, output_5_240;
mixer gate_output_5_240(.a(output_6_240), .b(output_6_1), .y(output_5_240));
wire output_7_240, output_7_1, output_6_240;
mixer gate_output_6_240(.a(output_7_240), .b(output_7_1), .y(output_6_240));
wire output_8_240, output_8_1, output_7_240;
mixer gate_output_7_240(.a(output_8_240), .b(output_8_1), .y(output_7_240));
wire output_9_240, output_9_1, output_8_240;
mixer gate_output_8_240(.a(output_9_240), .b(output_9_1), .y(output_8_240));
wire output_10_240, output_10_1, output_9_240;
mixer gate_output_9_240(.a(output_10_240), .b(output_10_1), .y(output_9_240));
wire output_11_240, output_11_1, output_10_240;
mixer gate_output_10_240(.a(output_11_240), .b(output_11_1), .y(output_10_240));
wire output_12_240, output_12_1, output_11_240;
mixer gate_output_11_240(.a(output_12_240), .b(output_12_1), .y(output_11_240));
wire output_13_240, output_13_1, output_12_240;
mixer gate_output_12_240(.a(output_13_240), .b(output_13_1), .y(output_12_240));
wire output_14_240, output_14_1, output_13_240;
mixer gate_output_13_240(.a(output_14_240), .b(output_14_1), .y(output_13_240));
wire output_15_240, output_15_1, output_14_240;
mixer gate_output_14_240(.a(output_15_240), .b(output_15_1), .y(output_14_240));
wire output_16_240, output_16_1, output_15_240;
mixer gate_output_15_240(.a(output_16_240), .b(output_16_1), .y(output_15_240));
wire output_1_241, output_1_2, output_0_241;
mixer gate_output_0_241(.a(output_1_241), .b(output_1_2), .y(output_0_241));
wire output_2_241, output_2_2, output_1_241;
mixer gate_output_1_241(.a(output_2_241), .b(output_2_2), .y(output_1_241));
wire output_3_241, output_3_2, output_2_241;
mixer gate_output_2_241(.a(output_3_241), .b(output_3_2), .y(output_2_241));
wire output_4_241, output_4_2, output_3_241;
mixer gate_output_3_241(.a(output_4_241), .b(output_4_2), .y(output_3_241));
wire output_5_241, output_5_2, output_4_241;
mixer gate_output_4_241(.a(output_5_241), .b(output_5_2), .y(output_4_241));
wire output_6_241, output_6_2, output_5_241;
mixer gate_output_5_241(.a(output_6_241), .b(output_6_2), .y(output_5_241));
wire output_7_241, output_7_2, output_6_241;
mixer gate_output_6_241(.a(output_7_241), .b(output_7_2), .y(output_6_241));
wire output_8_241, output_8_2, output_7_241;
mixer gate_output_7_241(.a(output_8_241), .b(output_8_2), .y(output_7_241));
wire output_9_241, output_9_2, output_8_241;
mixer gate_output_8_241(.a(output_9_241), .b(output_9_2), .y(output_8_241));
wire output_10_241, output_10_2, output_9_241;
mixer gate_output_9_241(.a(output_10_241), .b(output_10_2), .y(output_9_241));
wire output_11_241, output_11_2, output_10_241;
mixer gate_output_10_241(.a(output_11_241), .b(output_11_2), .y(output_10_241));
wire output_12_241, output_12_2, output_11_241;
mixer gate_output_11_241(.a(output_12_241), .b(output_12_2), .y(output_11_241));
wire output_13_241, output_13_2, output_12_241;
mixer gate_output_12_241(.a(output_13_241), .b(output_13_2), .y(output_12_241));
wire output_14_241, output_14_2, output_13_241;
mixer gate_output_13_241(.a(output_14_241), .b(output_14_2), .y(output_13_241));
wire output_15_241, output_15_2, output_14_241;
mixer gate_output_14_241(.a(output_15_241), .b(output_15_2), .y(output_14_241));
wire output_16_241, output_16_2, output_15_241;
mixer gate_output_15_241(.a(output_16_241), .b(output_16_2), .y(output_15_241));
wire output_1_242, output_1_3, output_0_242;
mixer gate_output_0_242(.a(output_1_242), .b(output_1_3), .y(output_0_242));
wire output_2_242, output_2_3, output_1_242;
mixer gate_output_1_242(.a(output_2_242), .b(output_2_3), .y(output_1_242));
wire output_3_242, output_3_3, output_2_242;
mixer gate_output_2_242(.a(output_3_242), .b(output_3_3), .y(output_2_242));
wire output_4_242, output_4_3, output_3_242;
mixer gate_output_3_242(.a(output_4_242), .b(output_4_3), .y(output_3_242));
wire output_5_242, output_5_3, output_4_242;
mixer gate_output_4_242(.a(output_5_242), .b(output_5_3), .y(output_4_242));
wire output_6_242, output_6_3, output_5_242;
mixer gate_output_5_242(.a(output_6_242), .b(output_6_3), .y(output_5_242));
wire output_7_242, output_7_3, output_6_242;
mixer gate_output_6_242(.a(output_7_242), .b(output_7_3), .y(output_6_242));
wire output_8_242, output_8_3, output_7_242;
mixer gate_output_7_242(.a(output_8_242), .b(output_8_3), .y(output_7_242));
wire output_9_242, output_9_3, output_8_242;
mixer gate_output_8_242(.a(output_9_242), .b(output_9_3), .y(output_8_242));
wire output_10_242, output_10_3, output_9_242;
mixer gate_output_9_242(.a(output_10_242), .b(output_10_3), .y(output_9_242));
wire output_11_242, output_11_3, output_10_242;
mixer gate_output_10_242(.a(output_11_242), .b(output_11_3), .y(output_10_242));
wire output_12_242, output_12_3, output_11_242;
mixer gate_output_11_242(.a(output_12_242), .b(output_12_3), .y(output_11_242));
wire output_13_242, output_13_3, output_12_242;
mixer gate_output_12_242(.a(output_13_242), .b(output_13_3), .y(output_12_242));
wire output_14_242, output_14_3, output_13_242;
mixer gate_output_13_242(.a(output_14_242), .b(output_14_3), .y(output_13_242));
wire output_15_242, output_15_3, output_14_242;
mixer gate_output_14_242(.a(output_15_242), .b(output_15_3), .y(output_14_242));
wire output_16_242, output_16_3, output_15_242;
mixer gate_output_15_242(.a(output_16_242), .b(output_16_3), .y(output_15_242));
wire output_1_243, output_1_4, output_0_243;
mixer gate_output_0_243(.a(output_1_243), .b(output_1_4), .y(output_0_243));
wire output_2_243, output_2_4, output_1_243;
mixer gate_output_1_243(.a(output_2_243), .b(output_2_4), .y(output_1_243));
wire output_3_243, output_3_4, output_2_243;
mixer gate_output_2_243(.a(output_3_243), .b(output_3_4), .y(output_2_243));
wire output_4_243, output_4_4, output_3_243;
mixer gate_output_3_243(.a(output_4_243), .b(output_4_4), .y(output_3_243));
wire output_5_243, output_5_4, output_4_243;
mixer gate_output_4_243(.a(output_5_243), .b(output_5_4), .y(output_4_243));
wire output_6_243, output_6_4, output_5_243;
mixer gate_output_5_243(.a(output_6_243), .b(output_6_4), .y(output_5_243));
wire output_7_243, output_7_4, output_6_243;
mixer gate_output_6_243(.a(output_7_243), .b(output_7_4), .y(output_6_243));
wire output_8_243, output_8_4, output_7_243;
mixer gate_output_7_243(.a(output_8_243), .b(output_8_4), .y(output_7_243));
wire output_9_243, output_9_4, output_8_243;
mixer gate_output_8_243(.a(output_9_243), .b(output_9_4), .y(output_8_243));
wire output_10_243, output_10_4, output_9_243;
mixer gate_output_9_243(.a(output_10_243), .b(output_10_4), .y(output_9_243));
wire output_11_243, output_11_4, output_10_243;
mixer gate_output_10_243(.a(output_11_243), .b(output_11_4), .y(output_10_243));
wire output_12_243, output_12_4, output_11_243;
mixer gate_output_11_243(.a(output_12_243), .b(output_12_4), .y(output_11_243));
wire output_13_243, output_13_4, output_12_243;
mixer gate_output_12_243(.a(output_13_243), .b(output_13_4), .y(output_12_243));
wire output_14_243, output_14_4, output_13_243;
mixer gate_output_13_243(.a(output_14_243), .b(output_14_4), .y(output_13_243));
wire output_15_243, output_15_4, output_14_243;
mixer gate_output_14_243(.a(output_15_243), .b(output_15_4), .y(output_14_243));
wire output_16_243, output_16_4, output_15_243;
mixer gate_output_15_243(.a(output_16_243), .b(output_16_4), .y(output_15_243));
wire output_1_244, output_1_5, output_0_244;
mixer gate_output_0_244(.a(output_1_244), .b(output_1_5), .y(output_0_244));
wire output_2_244, output_2_5, output_1_244;
mixer gate_output_1_244(.a(output_2_244), .b(output_2_5), .y(output_1_244));
wire output_3_244, output_3_5, output_2_244;
mixer gate_output_2_244(.a(output_3_244), .b(output_3_5), .y(output_2_244));
wire output_4_244, output_4_5, output_3_244;
mixer gate_output_3_244(.a(output_4_244), .b(output_4_5), .y(output_3_244));
wire output_5_244, output_5_5, output_4_244;
mixer gate_output_4_244(.a(output_5_244), .b(output_5_5), .y(output_4_244));
wire output_6_244, output_6_5, output_5_244;
mixer gate_output_5_244(.a(output_6_244), .b(output_6_5), .y(output_5_244));
wire output_7_244, output_7_5, output_6_244;
mixer gate_output_6_244(.a(output_7_244), .b(output_7_5), .y(output_6_244));
wire output_8_244, output_8_5, output_7_244;
mixer gate_output_7_244(.a(output_8_244), .b(output_8_5), .y(output_7_244));
wire output_9_244, output_9_5, output_8_244;
mixer gate_output_8_244(.a(output_9_244), .b(output_9_5), .y(output_8_244));
wire output_10_244, output_10_5, output_9_244;
mixer gate_output_9_244(.a(output_10_244), .b(output_10_5), .y(output_9_244));
wire output_11_244, output_11_5, output_10_244;
mixer gate_output_10_244(.a(output_11_244), .b(output_11_5), .y(output_10_244));
wire output_12_244, output_12_5, output_11_244;
mixer gate_output_11_244(.a(output_12_244), .b(output_12_5), .y(output_11_244));
wire output_13_244, output_13_5, output_12_244;
mixer gate_output_12_244(.a(output_13_244), .b(output_13_5), .y(output_12_244));
wire output_14_244, output_14_5, output_13_244;
mixer gate_output_13_244(.a(output_14_244), .b(output_14_5), .y(output_13_244));
wire output_15_244, output_15_5, output_14_244;
mixer gate_output_14_244(.a(output_15_244), .b(output_15_5), .y(output_14_244));
wire output_16_244, output_16_5, output_15_244;
mixer gate_output_15_244(.a(output_16_244), .b(output_16_5), .y(output_15_244));
wire output_1_245, output_1_6, output_0_245;
mixer gate_output_0_245(.a(output_1_245), .b(output_1_6), .y(output_0_245));
wire output_2_245, output_2_6, output_1_245;
mixer gate_output_1_245(.a(output_2_245), .b(output_2_6), .y(output_1_245));
wire output_3_245, output_3_6, output_2_245;
mixer gate_output_2_245(.a(output_3_245), .b(output_3_6), .y(output_2_245));
wire output_4_245, output_4_6, output_3_245;
mixer gate_output_3_245(.a(output_4_245), .b(output_4_6), .y(output_3_245));
wire output_5_245, output_5_6, output_4_245;
mixer gate_output_4_245(.a(output_5_245), .b(output_5_6), .y(output_4_245));
wire output_6_245, output_6_6, output_5_245;
mixer gate_output_5_245(.a(output_6_245), .b(output_6_6), .y(output_5_245));
wire output_7_245, output_7_6, output_6_245;
mixer gate_output_6_245(.a(output_7_245), .b(output_7_6), .y(output_6_245));
wire output_8_245, output_8_6, output_7_245;
mixer gate_output_7_245(.a(output_8_245), .b(output_8_6), .y(output_7_245));
wire output_9_245, output_9_6, output_8_245;
mixer gate_output_8_245(.a(output_9_245), .b(output_9_6), .y(output_8_245));
wire output_10_245, output_10_6, output_9_245;
mixer gate_output_9_245(.a(output_10_245), .b(output_10_6), .y(output_9_245));
wire output_11_245, output_11_6, output_10_245;
mixer gate_output_10_245(.a(output_11_245), .b(output_11_6), .y(output_10_245));
wire output_12_245, output_12_6, output_11_245;
mixer gate_output_11_245(.a(output_12_245), .b(output_12_6), .y(output_11_245));
wire output_13_245, output_13_6, output_12_245;
mixer gate_output_12_245(.a(output_13_245), .b(output_13_6), .y(output_12_245));
wire output_14_245, output_14_6, output_13_245;
mixer gate_output_13_245(.a(output_14_245), .b(output_14_6), .y(output_13_245));
wire output_15_245, output_15_6, output_14_245;
mixer gate_output_14_245(.a(output_15_245), .b(output_15_6), .y(output_14_245));
wire output_16_245, output_16_6, output_15_245;
mixer gate_output_15_245(.a(output_16_245), .b(output_16_6), .y(output_15_245));
wire output_1_246, output_1_7, output_0_246;
mixer gate_output_0_246(.a(output_1_246), .b(output_1_7), .y(output_0_246));
wire output_2_246, output_2_7, output_1_246;
mixer gate_output_1_246(.a(output_2_246), .b(output_2_7), .y(output_1_246));
wire output_3_246, output_3_7, output_2_246;
mixer gate_output_2_246(.a(output_3_246), .b(output_3_7), .y(output_2_246));
wire output_4_246, output_4_7, output_3_246;
mixer gate_output_3_246(.a(output_4_246), .b(output_4_7), .y(output_3_246));
wire output_5_246, output_5_7, output_4_246;
mixer gate_output_4_246(.a(output_5_246), .b(output_5_7), .y(output_4_246));
wire output_6_246, output_6_7, output_5_246;
mixer gate_output_5_246(.a(output_6_246), .b(output_6_7), .y(output_5_246));
wire output_7_246, output_7_7, output_6_246;
mixer gate_output_6_246(.a(output_7_246), .b(output_7_7), .y(output_6_246));
wire output_8_246, output_8_7, output_7_246;
mixer gate_output_7_246(.a(output_8_246), .b(output_8_7), .y(output_7_246));
wire output_9_246, output_9_7, output_8_246;
mixer gate_output_8_246(.a(output_9_246), .b(output_9_7), .y(output_8_246));
wire output_10_246, output_10_7, output_9_246;
mixer gate_output_9_246(.a(output_10_246), .b(output_10_7), .y(output_9_246));
wire output_11_246, output_11_7, output_10_246;
mixer gate_output_10_246(.a(output_11_246), .b(output_11_7), .y(output_10_246));
wire output_12_246, output_12_7, output_11_246;
mixer gate_output_11_246(.a(output_12_246), .b(output_12_7), .y(output_11_246));
wire output_13_246, output_13_7, output_12_246;
mixer gate_output_12_246(.a(output_13_246), .b(output_13_7), .y(output_12_246));
wire output_14_246, output_14_7, output_13_246;
mixer gate_output_13_246(.a(output_14_246), .b(output_14_7), .y(output_13_246));
wire output_15_246, output_15_7, output_14_246;
mixer gate_output_14_246(.a(output_15_246), .b(output_15_7), .y(output_14_246));
wire output_16_246, output_16_7, output_15_246;
mixer gate_output_15_246(.a(output_16_246), .b(output_16_7), .y(output_15_246));
wire output_1_247, output_1_8, output_0_247;
mixer gate_output_0_247(.a(output_1_247), .b(output_1_8), .y(output_0_247));
wire output_2_247, output_2_8, output_1_247;
mixer gate_output_1_247(.a(output_2_247), .b(output_2_8), .y(output_1_247));
wire output_3_247, output_3_8, output_2_247;
mixer gate_output_2_247(.a(output_3_247), .b(output_3_8), .y(output_2_247));
wire output_4_247, output_4_8, output_3_247;
mixer gate_output_3_247(.a(output_4_247), .b(output_4_8), .y(output_3_247));
wire output_5_247, output_5_8, output_4_247;
mixer gate_output_4_247(.a(output_5_247), .b(output_5_8), .y(output_4_247));
wire output_6_247, output_6_8, output_5_247;
mixer gate_output_5_247(.a(output_6_247), .b(output_6_8), .y(output_5_247));
wire output_7_247, output_7_8, output_6_247;
mixer gate_output_6_247(.a(output_7_247), .b(output_7_8), .y(output_6_247));
wire output_8_247, output_8_8, output_7_247;
mixer gate_output_7_247(.a(output_8_247), .b(output_8_8), .y(output_7_247));
wire output_9_247, output_9_8, output_8_247;
mixer gate_output_8_247(.a(output_9_247), .b(output_9_8), .y(output_8_247));
wire output_10_247, output_10_8, output_9_247;
mixer gate_output_9_247(.a(output_10_247), .b(output_10_8), .y(output_9_247));
wire output_11_247, output_11_8, output_10_247;
mixer gate_output_10_247(.a(output_11_247), .b(output_11_8), .y(output_10_247));
wire output_12_247, output_12_8, output_11_247;
mixer gate_output_11_247(.a(output_12_247), .b(output_12_8), .y(output_11_247));
wire output_13_247, output_13_8, output_12_247;
mixer gate_output_12_247(.a(output_13_247), .b(output_13_8), .y(output_12_247));
wire output_14_247, output_14_8, output_13_247;
mixer gate_output_13_247(.a(output_14_247), .b(output_14_8), .y(output_13_247));
wire output_15_247, output_15_8, output_14_247;
mixer gate_output_14_247(.a(output_15_247), .b(output_15_8), .y(output_14_247));
wire output_16_247, output_16_8, output_15_247;
mixer gate_output_15_247(.a(output_16_247), .b(output_16_8), .y(output_15_247));
wire output_1_248, output_1_9, output_0_248;
mixer gate_output_0_248(.a(output_1_248), .b(output_1_9), .y(output_0_248));
wire output_2_248, output_2_9, output_1_248;
mixer gate_output_1_248(.a(output_2_248), .b(output_2_9), .y(output_1_248));
wire output_3_248, output_3_9, output_2_248;
mixer gate_output_2_248(.a(output_3_248), .b(output_3_9), .y(output_2_248));
wire output_4_248, output_4_9, output_3_248;
mixer gate_output_3_248(.a(output_4_248), .b(output_4_9), .y(output_3_248));
wire output_5_248, output_5_9, output_4_248;
mixer gate_output_4_248(.a(output_5_248), .b(output_5_9), .y(output_4_248));
wire output_6_248, output_6_9, output_5_248;
mixer gate_output_5_248(.a(output_6_248), .b(output_6_9), .y(output_5_248));
wire output_7_248, output_7_9, output_6_248;
mixer gate_output_6_248(.a(output_7_248), .b(output_7_9), .y(output_6_248));
wire output_8_248, output_8_9, output_7_248;
mixer gate_output_7_248(.a(output_8_248), .b(output_8_9), .y(output_7_248));
wire output_9_248, output_9_9, output_8_248;
mixer gate_output_8_248(.a(output_9_248), .b(output_9_9), .y(output_8_248));
wire output_10_248, output_10_9, output_9_248;
mixer gate_output_9_248(.a(output_10_248), .b(output_10_9), .y(output_9_248));
wire output_11_248, output_11_9, output_10_248;
mixer gate_output_10_248(.a(output_11_248), .b(output_11_9), .y(output_10_248));
wire output_12_248, output_12_9, output_11_248;
mixer gate_output_11_248(.a(output_12_248), .b(output_12_9), .y(output_11_248));
wire output_13_248, output_13_9, output_12_248;
mixer gate_output_12_248(.a(output_13_248), .b(output_13_9), .y(output_12_248));
wire output_14_248, output_14_9, output_13_248;
mixer gate_output_13_248(.a(output_14_248), .b(output_14_9), .y(output_13_248));
wire output_15_248, output_15_9, output_14_248;
mixer gate_output_14_248(.a(output_15_248), .b(output_15_9), .y(output_14_248));
wire output_16_248, output_16_9, output_15_248;
mixer gate_output_15_248(.a(output_16_248), .b(output_16_9), .y(output_15_248));
wire output_1_249, output_1_10, output_0_249;
mixer gate_output_0_249(.a(output_1_249), .b(output_1_10), .y(output_0_249));
wire output_2_249, output_2_10, output_1_249;
mixer gate_output_1_249(.a(output_2_249), .b(output_2_10), .y(output_1_249));
wire output_3_249, output_3_10, output_2_249;
mixer gate_output_2_249(.a(output_3_249), .b(output_3_10), .y(output_2_249));
wire output_4_249, output_4_10, output_3_249;
mixer gate_output_3_249(.a(output_4_249), .b(output_4_10), .y(output_3_249));
wire output_5_249, output_5_10, output_4_249;
mixer gate_output_4_249(.a(output_5_249), .b(output_5_10), .y(output_4_249));
wire output_6_249, output_6_10, output_5_249;
mixer gate_output_5_249(.a(output_6_249), .b(output_6_10), .y(output_5_249));
wire output_7_249, output_7_10, output_6_249;
mixer gate_output_6_249(.a(output_7_249), .b(output_7_10), .y(output_6_249));
wire output_8_249, output_8_10, output_7_249;
mixer gate_output_7_249(.a(output_8_249), .b(output_8_10), .y(output_7_249));
wire output_9_249, output_9_10, output_8_249;
mixer gate_output_8_249(.a(output_9_249), .b(output_9_10), .y(output_8_249));
wire output_10_249, output_10_10, output_9_249;
mixer gate_output_9_249(.a(output_10_249), .b(output_10_10), .y(output_9_249));
wire output_11_249, output_11_10, output_10_249;
mixer gate_output_10_249(.a(output_11_249), .b(output_11_10), .y(output_10_249));
wire output_12_249, output_12_10, output_11_249;
mixer gate_output_11_249(.a(output_12_249), .b(output_12_10), .y(output_11_249));
wire output_13_249, output_13_10, output_12_249;
mixer gate_output_12_249(.a(output_13_249), .b(output_13_10), .y(output_12_249));
wire output_14_249, output_14_10, output_13_249;
mixer gate_output_13_249(.a(output_14_249), .b(output_14_10), .y(output_13_249));
wire output_15_249, output_15_10, output_14_249;
mixer gate_output_14_249(.a(output_15_249), .b(output_15_10), .y(output_14_249));
wire output_16_249, output_16_10, output_15_249;
mixer gate_output_15_249(.a(output_16_249), .b(output_16_10), .y(output_15_249));
wire output_1_250, output_1_11, output_0_250;
mixer gate_output_0_250(.a(output_1_250), .b(output_1_11), .y(output_0_250));
wire output_2_250, output_2_11, output_1_250;
mixer gate_output_1_250(.a(output_2_250), .b(output_2_11), .y(output_1_250));
wire output_3_250, output_3_11, output_2_250;
mixer gate_output_2_250(.a(output_3_250), .b(output_3_11), .y(output_2_250));
wire output_4_250, output_4_11, output_3_250;
mixer gate_output_3_250(.a(output_4_250), .b(output_4_11), .y(output_3_250));
wire output_5_250, output_5_11, output_4_250;
mixer gate_output_4_250(.a(output_5_250), .b(output_5_11), .y(output_4_250));
wire output_6_250, output_6_11, output_5_250;
mixer gate_output_5_250(.a(output_6_250), .b(output_6_11), .y(output_5_250));
wire output_7_250, output_7_11, output_6_250;
mixer gate_output_6_250(.a(output_7_250), .b(output_7_11), .y(output_6_250));
wire output_8_250, output_8_11, output_7_250;
mixer gate_output_7_250(.a(output_8_250), .b(output_8_11), .y(output_7_250));
wire output_9_250, output_9_11, output_8_250;
mixer gate_output_8_250(.a(output_9_250), .b(output_9_11), .y(output_8_250));
wire output_10_250, output_10_11, output_9_250;
mixer gate_output_9_250(.a(output_10_250), .b(output_10_11), .y(output_9_250));
wire output_11_250, output_11_11, output_10_250;
mixer gate_output_10_250(.a(output_11_250), .b(output_11_11), .y(output_10_250));
wire output_12_250, output_12_11, output_11_250;
mixer gate_output_11_250(.a(output_12_250), .b(output_12_11), .y(output_11_250));
wire output_13_250, output_13_11, output_12_250;
mixer gate_output_12_250(.a(output_13_250), .b(output_13_11), .y(output_12_250));
wire output_14_250, output_14_11, output_13_250;
mixer gate_output_13_250(.a(output_14_250), .b(output_14_11), .y(output_13_250));
wire output_15_250, output_15_11, output_14_250;
mixer gate_output_14_250(.a(output_15_250), .b(output_15_11), .y(output_14_250));
wire output_16_250, output_16_11, output_15_250;
mixer gate_output_15_250(.a(output_16_250), .b(output_16_11), .y(output_15_250));
wire output_1_251, output_1_12, output_0_251;
mixer gate_output_0_251(.a(output_1_251), .b(output_1_12), .y(output_0_251));
wire output_2_251, output_2_12, output_1_251;
mixer gate_output_1_251(.a(output_2_251), .b(output_2_12), .y(output_1_251));
wire output_3_251, output_3_12, output_2_251;
mixer gate_output_2_251(.a(output_3_251), .b(output_3_12), .y(output_2_251));
wire output_4_251, output_4_12, output_3_251;
mixer gate_output_3_251(.a(output_4_251), .b(output_4_12), .y(output_3_251));
wire output_5_251, output_5_12, output_4_251;
mixer gate_output_4_251(.a(output_5_251), .b(output_5_12), .y(output_4_251));
wire output_6_251, output_6_12, output_5_251;
mixer gate_output_5_251(.a(output_6_251), .b(output_6_12), .y(output_5_251));
wire output_7_251, output_7_12, output_6_251;
mixer gate_output_6_251(.a(output_7_251), .b(output_7_12), .y(output_6_251));
wire output_8_251, output_8_12, output_7_251;
mixer gate_output_7_251(.a(output_8_251), .b(output_8_12), .y(output_7_251));
wire output_9_251, output_9_12, output_8_251;
mixer gate_output_8_251(.a(output_9_251), .b(output_9_12), .y(output_8_251));
wire output_10_251, output_10_12, output_9_251;
mixer gate_output_9_251(.a(output_10_251), .b(output_10_12), .y(output_9_251));
wire output_11_251, output_11_12, output_10_251;
mixer gate_output_10_251(.a(output_11_251), .b(output_11_12), .y(output_10_251));
wire output_12_251, output_12_12, output_11_251;
mixer gate_output_11_251(.a(output_12_251), .b(output_12_12), .y(output_11_251));
wire output_13_251, output_13_12, output_12_251;
mixer gate_output_12_251(.a(output_13_251), .b(output_13_12), .y(output_12_251));
wire output_14_251, output_14_12, output_13_251;
mixer gate_output_13_251(.a(output_14_251), .b(output_14_12), .y(output_13_251));
wire output_15_251, output_15_12, output_14_251;
mixer gate_output_14_251(.a(output_15_251), .b(output_15_12), .y(output_14_251));
wire output_16_251, output_16_12, output_15_251;
mixer gate_output_15_251(.a(output_16_251), .b(output_16_12), .y(output_15_251));
wire output_1_252, output_1_13, output_0_252;
mixer gate_output_0_252(.a(output_1_252), .b(output_1_13), .y(output_0_252));
wire output_2_252, output_2_13, output_1_252;
mixer gate_output_1_252(.a(output_2_252), .b(output_2_13), .y(output_1_252));
wire output_3_252, output_3_13, output_2_252;
mixer gate_output_2_252(.a(output_3_252), .b(output_3_13), .y(output_2_252));
wire output_4_252, output_4_13, output_3_252;
mixer gate_output_3_252(.a(output_4_252), .b(output_4_13), .y(output_3_252));
wire output_5_252, output_5_13, output_4_252;
mixer gate_output_4_252(.a(output_5_252), .b(output_5_13), .y(output_4_252));
wire output_6_252, output_6_13, output_5_252;
mixer gate_output_5_252(.a(output_6_252), .b(output_6_13), .y(output_5_252));
wire output_7_252, output_7_13, output_6_252;
mixer gate_output_6_252(.a(output_7_252), .b(output_7_13), .y(output_6_252));
wire output_8_252, output_8_13, output_7_252;
mixer gate_output_7_252(.a(output_8_252), .b(output_8_13), .y(output_7_252));
wire output_9_252, output_9_13, output_8_252;
mixer gate_output_8_252(.a(output_9_252), .b(output_9_13), .y(output_8_252));
wire output_10_252, output_10_13, output_9_252;
mixer gate_output_9_252(.a(output_10_252), .b(output_10_13), .y(output_9_252));
wire output_11_252, output_11_13, output_10_252;
mixer gate_output_10_252(.a(output_11_252), .b(output_11_13), .y(output_10_252));
wire output_12_252, output_12_13, output_11_252;
mixer gate_output_11_252(.a(output_12_252), .b(output_12_13), .y(output_11_252));
wire output_13_252, output_13_13, output_12_252;
mixer gate_output_12_252(.a(output_13_252), .b(output_13_13), .y(output_12_252));
wire output_14_252, output_14_13, output_13_252;
mixer gate_output_13_252(.a(output_14_252), .b(output_14_13), .y(output_13_252));
wire output_15_252, output_15_13, output_14_252;
mixer gate_output_14_252(.a(output_15_252), .b(output_15_13), .y(output_14_252));
wire output_16_252, output_16_13, output_15_252;
mixer gate_output_15_252(.a(output_16_252), .b(output_16_13), .y(output_15_252));
wire output_1_253, output_1_14, output_0_253;
mixer gate_output_0_253(.a(output_1_253), .b(output_1_14), .y(output_0_253));
wire output_2_253, output_2_14, output_1_253;
mixer gate_output_1_253(.a(output_2_253), .b(output_2_14), .y(output_1_253));
wire output_3_253, output_3_14, output_2_253;
mixer gate_output_2_253(.a(output_3_253), .b(output_3_14), .y(output_2_253));
wire output_4_253, output_4_14, output_3_253;
mixer gate_output_3_253(.a(output_4_253), .b(output_4_14), .y(output_3_253));
wire output_5_253, output_5_14, output_4_253;
mixer gate_output_4_253(.a(output_5_253), .b(output_5_14), .y(output_4_253));
wire output_6_253, output_6_14, output_5_253;
mixer gate_output_5_253(.a(output_6_253), .b(output_6_14), .y(output_5_253));
wire output_7_253, output_7_14, output_6_253;
mixer gate_output_6_253(.a(output_7_253), .b(output_7_14), .y(output_6_253));
wire output_8_253, output_8_14, output_7_253;
mixer gate_output_7_253(.a(output_8_253), .b(output_8_14), .y(output_7_253));
wire output_9_253, output_9_14, output_8_253;
mixer gate_output_8_253(.a(output_9_253), .b(output_9_14), .y(output_8_253));
wire output_10_253, output_10_14, output_9_253;
mixer gate_output_9_253(.a(output_10_253), .b(output_10_14), .y(output_9_253));
wire output_11_253, output_11_14, output_10_253;
mixer gate_output_10_253(.a(output_11_253), .b(output_11_14), .y(output_10_253));
wire output_12_253, output_12_14, output_11_253;
mixer gate_output_11_253(.a(output_12_253), .b(output_12_14), .y(output_11_253));
wire output_13_253, output_13_14, output_12_253;
mixer gate_output_12_253(.a(output_13_253), .b(output_13_14), .y(output_12_253));
wire output_14_253, output_14_14, output_13_253;
mixer gate_output_13_253(.a(output_14_253), .b(output_14_14), .y(output_13_253));
wire output_15_253, output_15_14, output_14_253;
mixer gate_output_14_253(.a(output_15_253), .b(output_15_14), .y(output_14_253));
wire output_16_253, output_16_14, output_15_253;
mixer gate_output_15_253(.a(output_16_253), .b(output_16_14), .y(output_15_253));
wire output_1_254, output_1_15, output_0_254;
mixer gate_output_0_254(.a(output_1_254), .b(output_1_15), .y(output_0_254));
wire output_2_254, output_2_15, output_1_254;
mixer gate_output_1_254(.a(output_2_254), .b(output_2_15), .y(output_1_254));
wire output_3_254, output_3_15, output_2_254;
mixer gate_output_2_254(.a(output_3_254), .b(output_3_15), .y(output_2_254));
wire output_4_254, output_4_15, output_3_254;
mixer gate_output_3_254(.a(output_4_254), .b(output_4_15), .y(output_3_254));
wire output_5_254, output_5_15, output_4_254;
mixer gate_output_4_254(.a(output_5_254), .b(output_5_15), .y(output_4_254));
wire output_6_254, output_6_15, output_5_254;
mixer gate_output_5_254(.a(output_6_254), .b(output_6_15), .y(output_5_254));
wire output_7_254, output_7_15, output_6_254;
mixer gate_output_6_254(.a(output_7_254), .b(output_7_15), .y(output_6_254));
wire output_8_254, output_8_15, output_7_254;
mixer gate_output_7_254(.a(output_8_254), .b(output_8_15), .y(output_7_254));
wire output_9_254, output_9_15, output_8_254;
mixer gate_output_8_254(.a(output_9_254), .b(output_9_15), .y(output_8_254));
wire output_10_254, output_10_15, output_9_254;
mixer gate_output_9_254(.a(output_10_254), .b(output_10_15), .y(output_9_254));
wire output_11_254, output_11_15, output_10_254;
mixer gate_output_10_254(.a(output_11_254), .b(output_11_15), .y(output_10_254));
wire output_12_254, output_12_15, output_11_254;
mixer gate_output_11_254(.a(output_12_254), .b(output_12_15), .y(output_11_254));
wire output_13_254, output_13_15, output_12_254;
mixer gate_output_12_254(.a(output_13_254), .b(output_13_15), .y(output_12_254));
wire output_14_254, output_14_15, output_13_254;
mixer gate_output_13_254(.a(output_14_254), .b(output_14_15), .y(output_13_254));
wire output_15_254, output_15_15, output_14_254;
mixer gate_output_14_254(.a(output_15_254), .b(output_15_15), .y(output_14_254));
wire output_16_254, output_16_15, output_15_254;
mixer gate_output_15_254(.a(output_16_254), .b(output_16_15), .y(output_15_254));
wire output_1_255, output_1_0, output_0_255;
mixer gate_output_0_255(.a(output_1_255), .b(output_1_0), .y(output_0_255));
wire output_2_255, output_2_0, output_1_255;
mixer gate_output_1_255(.a(output_2_255), .b(output_2_0), .y(output_1_255));
wire output_3_255, output_3_0, output_2_255;
mixer gate_output_2_255(.a(output_3_255), .b(output_3_0), .y(output_2_255));
wire output_4_255, output_4_0, output_3_255;
mixer gate_output_3_255(.a(output_4_255), .b(output_4_0), .y(output_3_255));
wire output_5_255, output_5_0, output_4_255;
mixer gate_output_4_255(.a(output_5_255), .b(output_5_0), .y(output_4_255));
wire output_6_255, output_6_0, output_5_255;
mixer gate_output_5_255(.a(output_6_255), .b(output_6_0), .y(output_5_255));
wire output_7_255, output_7_0, output_6_255;
mixer gate_output_6_255(.a(output_7_255), .b(output_7_0), .y(output_6_255));
wire output_8_255, output_8_0, output_7_255;
mixer gate_output_7_255(.a(output_8_255), .b(output_8_0), .y(output_7_255));
wire output_9_255, output_9_0, output_8_255;
mixer gate_output_8_255(.a(output_9_255), .b(output_9_0), .y(output_8_255));
wire output_10_255, output_10_0, output_9_255;
mixer gate_output_9_255(.a(output_10_255), .b(output_10_0), .y(output_9_255));
wire output_11_255, output_11_0, output_10_255;
mixer gate_output_10_255(.a(output_11_255), .b(output_11_0), .y(output_10_255));
wire output_12_255, output_12_0, output_11_255;
mixer gate_output_11_255(.a(output_12_255), .b(output_12_0), .y(output_11_255));
wire output_13_255, output_13_0, output_12_255;
mixer gate_output_12_255(.a(output_13_255), .b(output_13_0), .y(output_12_255));
wire output_14_255, output_14_0, output_13_255;
mixer gate_output_13_255(.a(output_14_255), .b(output_14_0), .y(output_13_255));
wire output_15_255, output_15_0, output_14_255;
mixer gate_output_14_255(.a(output_15_255), .b(output_15_0), .y(output_14_255));
wire output_16_255, output_16_0, output_15_255;
mixer gate_output_15_255(.a(output_16_255), .b(output_16_0), .y(output_15_255));
assign output_0 = output_0_0;
wire output_0_256;
assign output_0_256 = input_0;
assign output_1 = output_1_0;
wire output_1_256;
assign output_1_256 = input_1;
assign output_2 = output_2_0;
wire output_2_256;
assign output_2_256 = input_2;
assign output_3 = output_3_0;
wire output_3_256;
assign output_3_256 = input_3;
assign output_4 = output_4_0;
wire output_4_256;
assign output_4_256 = input_4;
assign output_5 = output_5_0;
wire output_5_256;
assign output_5_256 = input_5;
assign output_6 = output_6_0;
wire output_6_256;
assign output_6_256 = input_6;
assign output_7 = output_7_0;
wire output_7_256;
assign output_7_256 = input_7;
assign output_8 = output_8_0;
wire output_8_256;
assign output_8_256 = input_8;
assign output_9 = output_9_0;
wire output_9_256;
assign output_9_256 = input_9;
assign output_10 = output_10_0;
wire output_10_256;
assign output_10_256 = input_10;
assign output_11 = output_11_0;
wire output_11_256;
assign output_11_256 = input_11;
assign output_12 = output_12_0;
wire output_12_256;
assign output_12_256 = input_12;
assign output_13 = output_13_0;
wire output_13_256;
assign output_13_256 = input_13;
assign output_14 = output_14_0;
wire output_14_256;
assign output_14_256 = input_14;
assign output_15 = output_15_0;
wire output_15_256;
assign output_15_256 = input_15;
endmodule
