module chain_8 (
inout k0, k8
);
wire {wires};
chamber ch0 (.in(k0), .out(k1)
chamber ch1 (.in(k1), .out(k2)
chamber ch2 (.in(k2), .out(k3)
chamber ch3 (.in(k3), .out(k4)
chamber ch4 (.in(k4), .out(k5)
chamber ch5 (.in(k5), .out(k6)
chamber ch6 (.in(k6), .out(k7)
chamber ch7 (.in(k7), .out(k8)
endmodule
