module binary_tree_1_6 (
output out_0,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_000000 (.a(t0_0000000), .b(t0_0000001), .y(t0_000000));
wire t0_0000000, t0_0000001;
mixer mix_t0_000001 (.a(t0_0000010), .b(t0_0000011), .y(t0_000001));
wire t0_0000010, t0_0000011;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_000010 (.a(t0_0000100), .b(t0_0000101), .y(t0_000010));
wire t0_0000100, t0_0000101;
mixer mix_t0_000011 (.a(t0_0000110), .b(t0_0000111), .y(t0_000011));
wire t0_0000110, t0_0000111;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_000100 (.a(t0_0001000), .b(t0_0001001), .y(t0_000100));
wire t0_0001000, t0_0001001;
mixer mix_t0_000101 (.a(t0_0001010), .b(t0_0001011), .y(t0_000101));
wire t0_0001010, t0_0001011;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_000110 (.a(t0_0001100), .b(t0_0001101), .y(t0_000110));
wire t0_0001100, t0_0001101;
mixer mix_t0_000111 (.a(t0_0001110), .b(t0_0001111), .y(t0_000111));
wire t0_0001110, t0_0001111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_001000 (.a(t0_0010000), .b(t0_0010001), .y(t0_001000));
wire t0_0010000, t0_0010001;
mixer mix_t0_001001 (.a(t0_0010010), .b(t0_0010011), .y(t0_001001));
wire t0_0010010, t0_0010011;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_001010 (.a(t0_0010100), .b(t0_0010101), .y(t0_001010));
wire t0_0010100, t0_0010101;
mixer mix_t0_001011 (.a(t0_0010110), .b(t0_0010111), .y(t0_001011));
wire t0_0010110, t0_0010111;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_001100 (.a(t0_0011000), .b(t0_0011001), .y(t0_001100));
wire t0_0011000, t0_0011001;
mixer mix_t0_001101 (.a(t0_0011010), .b(t0_0011011), .y(t0_001101));
wire t0_0011010, t0_0011011;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_001110 (.a(t0_0011100), .b(t0_0011101), .y(t0_001110));
wire t0_0011100, t0_0011101;
mixer mix_t0_001111 (.a(t0_0011110), .b(t0_0011111), .y(t0_001111));
wire t0_0011110, t0_0011111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_010000 (.a(t0_0100000), .b(t0_0100001), .y(t0_010000));
wire t0_0100000, t0_0100001;
mixer mix_t0_010001 (.a(t0_0100010), .b(t0_0100011), .y(t0_010001));
wire t0_0100010, t0_0100011;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_010010 (.a(t0_0100100), .b(t0_0100101), .y(t0_010010));
wire t0_0100100, t0_0100101;
mixer mix_t0_010011 (.a(t0_0100110), .b(t0_0100111), .y(t0_010011));
wire t0_0100110, t0_0100111;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_010100 (.a(t0_0101000), .b(t0_0101001), .y(t0_010100));
wire t0_0101000, t0_0101001;
mixer mix_t0_010101 (.a(t0_0101010), .b(t0_0101011), .y(t0_010101));
wire t0_0101010, t0_0101011;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_010110 (.a(t0_0101100), .b(t0_0101101), .y(t0_010110));
wire t0_0101100, t0_0101101;
mixer mix_t0_010111 (.a(t0_0101110), .b(t0_0101111), .y(t0_010111));
wire t0_0101110, t0_0101111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_011000 (.a(t0_0110000), .b(t0_0110001), .y(t0_011000));
wire t0_0110000, t0_0110001;
mixer mix_t0_011001 (.a(t0_0110010), .b(t0_0110011), .y(t0_011001));
wire t0_0110010, t0_0110011;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_011010 (.a(t0_0110100), .b(t0_0110101), .y(t0_011010));
wire t0_0110100, t0_0110101;
mixer mix_t0_011011 (.a(t0_0110110), .b(t0_0110111), .y(t0_011011));
wire t0_0110110, t0_0110111;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_011100 (.a(t0_0111000), .b(t0_0111001), .y(t0_011100));
wire t0_0111000, t0_0111001;
mixer mix_t0_011101 (.a(t0_0111010), .b(t0_0111011), .y(t0_011101));
wire t0_0111010, t0_0111011;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
mixer mix_t0_011110 (.a(t0_0111100), .b(t0_0111101), .y(t0_011110));
wire t0_0111100, t0_0111101;
mixer mix_t0_011111 (.a(t0_0111110), .b(t0_0111111), .y(t0_011111));
wire t0_0111110, t0_0111111;
wire t0_0;
assign out_0 = t0_0;
assign input_0 = t0_0000000;
assign input_1 = t0_0000001;
assign input_2 = t0_0000010;
assign input_3 = t0_0000011;
assign input_4 = t0_0000100;
assign input_5 = t0_0000101;
assign input_6 = t0_0000110;
assign input_7 = t0_0000111;
assign input_8 = t0_0001000;
assign input_9 = t0_0001001;
assign input_10 = t0_0001010;
assign input_11 = t0_0001011;
assign input_12 = t0_0001100;
assign input_13 = t0_0001101;
assign input_14 = t0_0001110;
assign input_15 = t0_0001111;
assign input_16 = t0_0010000;
assign input_17 = t0_0010001;
assign input_18 = t0_0010010;
assign input_19 = t0_0010011;
assign input_20 = t0_0010100;
assign input_21 = t0_0010101;
assign input_22 = t0_0010110;
assign input_23 = t0_0010111;
assign input_24 = t0_0011000;
assign input_25 = t0_0011001;
assign input_26 = t0_0011010;
assign input_27 = t0_0011011;
assign input_28 = t0_0011100;
assign input_29 = t0_0011101;
assign input_30 = t0_0011110;
assign input_31 = t0_0011111;
assign input_32 = t0_0100000;
assign input_33 = t0_0100001;
assign input_34 = t0_0100010;
assign input_35 = t0_0100011;
assign input_36 = t0_0100100;
assign input_37 = t0_0100101;
assign input_38 = t0_0100110;
assign input_39 = t0_0100111;
assign input_40 = t0_0101000;
assign input_41 = t0_0101001;
assign input_42 = t0_0101010;
assign input_43 = t0_0101011;
assign input_44 = t0_0101100;
assign input_45 = t0_0101101;
assign input_46 = t0_0101110;
assign input_47 = t0_0101111;
assign input_48 = t0_0110000;
assign input_49 = t0_0110001;
assign input_50 = t0_0110010;
assign input_51 = t0_0110011;
assign input_52 = t0_0110100;
assign input_53 = t0_0110101;
assign input_54 = t0_0110110;
assign input_55 = t0_0110111;
assign input_56 = t0_0111000;
assign input_57 = t0_0111001;
assign input_58 = t0_0111010;
assign input_59 = t0_0111011;
assign input_60 = t0_0111100;
assign input_61 = t0_0111101;
assign input_62 = t0_0111110;
assign input_63 = t0_0111111;
endmodule
