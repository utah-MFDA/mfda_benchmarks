module galaban10();
	mixer m_0(.a(e_0_1), .b(e_0_2), .y(e_0_3));
	mixer m_1(.a(e_0_1), .b(e_1_64), .y(e_1_69));
	mixer m_2(.a(e_0_2), .b(e_2_65), .y(e_2_66));
	mixer m_3(.a(e_0_3), .b(e_3_67), .y(e_3_68));
	mixer m_4(.a(e_4_8), .b(e_4_12), .y(e_4_16));
	mixer m_5(.a(e_5_9), .b(e_5_15), .y(e_5_17));
	mixer m_6(.a(e_6_11), .b(e_6_13), .y(e_6_19));
	mixer m_7(.a(e_7_10), .b(e_7_14), .y(e_7_18));
	mixer m_8(.a(e_4_8), .b(e_8_35), .y(e_8_39));
	mixer m_9(.a(e_5_9), .b(e_9_34), .y(e_9_40));
	mixer m_10(.a(e_7_10), .b(e_10_36), .y(e_10_38));
	mixer m_11(.a(e_6_11), .b(e_11_37), .y(e_11_41));
	mixer m_12(.a(e_4_12), .b(e_12_32), .y(e_12_43));
	mixer m_13(.a(e_6_13), .b(e_13_30), .y(e_13_45));
	mixer m_14(.a(e_7_14), .b(e_14_31), .y(e_14_42));
	mixer m_15(.a(e_5_15), .b(e_15_33), .y(e_15_44));
	mixer m_16(.a(e_4_16), .b(e_16_28), .y(e_16_30));
	mixer m_17(.a(e_5_17), .b(e_17_28), .y(e_17_31));
	mixer m_18(.a(e_7_18), .b(e_18_29), .y(e_18_32));
	mixer m_19(.a(e_6_19), .b(e_19_29), .y(e_19_33));
	mixer m_20(.a(e_20_37), .b(e_20_46), .y(e_20_48));
	mixer m_21(.a(e_21_36), .b(e_21_46), .y(e_21_49));
	mixer m_22(.a(e_22_35), .b(e_22_47), .y(e_22_51));
	mixer m_23(.a(e_23_34), .b(e_23_47), .y(e_23_50));
	mixer m_24(.a(e_24_39), .b(e_24_42), .y(e_24_48));
	mixer m_25(.a(e_25_40), .b(e_25_45), .y(e_25_49));
	mixer m_26(.a(e_26_38), .b(e_26_44), .y(e_26_51));
	mixer m_27(.a(e_27_41), .b(e_27_43), .y(e_27_50));
	mixer m_28(.a(e_16_28), .b(e_17_28), .y(e_28_63));
	mixer m_29(.a(e_18_29), .b(e_19_29), .y(e_29_62));
	mixer m_30(.a(e_13_30), .b(e_16_30), .y(e_30_58));
	mixer m_31(.a(e_14_31), .b(e_17_31), .y(e_31_59));
	mixer m_32(.a(e_12_32), .b(e_18_32), .y(e_32_60));
	mixer m_33(.a(e_15_33), .b(e_19_33), .y(e_33_61));
	mixer m_34(.a(e_9_34), .b(e_23_34), .y(e_34_52));
	mixer m_35(.a(e_8_35), .b(e_22_35), .y(e_35_53));
	mixer m_36(.a(e_10_36), .b(e_21_36), .y(e_36_55));
	mixer m_37(.a(e_11_37), .b(e_20_37), .y(e_37_54));
	mixer m_38(.a(e_10_38), .b(e_26_38), .y(e_38_58));
	mixer m_39(.a(e_8_39), .b(e_24_39), .y(e_39_61));
	mixer m_40(.a(e_9_40), .b(e_25_40), .y(e_40_60));
	mixer m_41(.a(e_11_41), .b(e_27_41), .y(e_41_59));
	mixer m_42(.a(e_14_42), .b(e_24_42), .y(e_42_56));
	mixer m_43(.a(e_12_43), .b(e_27_43), .y(e_43_57));
	mixer m_44(.a(e_15_44), .b(e_26_44), .y(e_44_57));
	mixer m_45(.a(e_13_45), .b(e_25_45), .y(e_45_56));
	mixer m_46(.a(e_20_46), .b(e_21_46), .y(e_46_63));
	mixer m_47(.a(e_22_47), .b(e_23_47), .y(e_47_62));
	mixer m_48(.a(e_20_48), .b(e_24_48), .y(e_48_52));
	mixer m_49(.a(e_21_49), .b(e_25_49), .y(e_49_53));
	mixer m_50(.a(e_23_50), .b(e_27_50), .y(e_50_55));
	mixer m_51(.a(e_22_51), .b(e_26_51), .y(e_51_54));
	mixer m_52(.a(e_34_52), .b(e_48_52), .y(e_52_65));
	mixer m_53(.a(e_35_53), .b(e_49_53), .y(e_53_66));
	mixer m_54(.a(e_37_54), .b(e_51_54), .y(e_54_68));
	mixer m_55(.a(e_36_55), .b(e_50_55), .y(e_55_67));
	mixer m_56(.a(e_42_56), .b(e_45_56), .y(e_56_69));
	mixer m_57(.a(e_43_57), .b(e_44_57), .y(e_57_69));
	mixer m_58(.a(e_30_58), .b(e_38_58), .y(e_58_65));
	mixer m_59(.a(e_31_59), .b(e_41_59), .y(e_59_66));
	mixer m_60(.a(e_32_60), .b(e_40_60), .y(e_60_68));
	mixer m_61(.a(e_33_61), .b(e_39_61), .y(e_61_67));
	mixer m_62(.a(e_29_62), .b(e_47_62), .y(e_62_64));
	mixer m_63(.a(e_28_63), .b(e_46_63), .y(e_63_64));
	mixer m_64(.a(e_1_64), .b(e_62_64), .y(e_63_64));
	mixer m_65(.a(e_2_65), .b(e_52_65), .y(e_58_65));
	mixer m_66(.a(e_2_66), .b(e_53_66), .y(e_59_66));
	mixer m_67(.a(e_3_67), .b(e_55_67), .y(e_61_67));
	mixer m_68(.a(e_3_68), .b(e_54_68), .y(e_60_68));
	mixer m_69(.a(e_1_69), .b(e_56_69), .y(e_57_69));
wire e_0_1,
	e_0_2,
	e_0_3,
	e_1_64,
	e_1_69,
	e_2_65,
	e_2_66,
	e_3_67,
	e_3_68,
	e_4_8,
	e_4_12,
	e_4_16,
	e_5_9,
	e_5_15,
	e_5_17,
	e_6_11,
	e_6_13,
	e_6_19,
	e_7_10,
	e_7_14,
	e_7_18,
	e_8_35,
	e_8_39,
	e_9_34,
	e_9_40,
	e_10_36,
	e_10_38,
	e_11_37,
	e_11_41,
	e_12_32,
	e_12_43,
	e_13_30,
	e_13_45,
	e_14_31,
	e_14_42,
	e_15_33,
	e_15_44,
	e_16_28,
	e_16_30,
	e_17_28,
	e_17_31,
	e_18_29,
	e_18_32,
	e_19_29,
	e_19_33,
	e_20_37,
	e_20_46,
	e_20_48,
	e_21_36,
	e_21_46,
	e_21_49,
	e_22_35,
	e_22_47,
	e_22_51,
	e_23_34,
	e_23_47,
	e_23_50,
	e_24_39,
	e_24_42,
	e_24_48,
	e_25_40,
	e_25_45,
	e_25_49,
	e_26_38,
	e_26_44,
	e_26_51,
	e_27_41,
	e_27_43,
	e_27_50,
	e_28_63,
	e_29_62,
	e_30_58,
	e_31_59,
	e_32_60,
	e_33_61,
	e_34_52,
	e_35_53,
	e_36_55,
	e_37_54,
	e_38_58,
	e_39_61,
	e_40_60,
	e_41_59,
	e_42_56,
	e_43_57,
	e_44_57,
	e_45_56,
	e_46_63,
	e_47_62,
	e_48_52,
	e_49_53,
	e_50_55,
	e_51_54,
	e_52_65,
	e_53_66,
	e_54_68,
	e_55_67,
	e_56_69,
	e_57_69,
	e_58_65,
	e_59_66,
	e_60_68,
	e_61_67,
	e_62_64,
	e_63_64;
endmodule
