module binary_tree_1_7 (
output out_0,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63,input input_64,input input_65,input input_66,input input_67,input input_68,input input_69,input input_70,input input_71,input input_72,input input_73,input input_74,input input_75,input input_76,input input_77,input input_78,input input_79,input input_80,input input_81,input input_82,input input_83,input input_84,input input_85,input input_86,input input_87,input input_88,input input_89,input input_90,input input_91,input input_92,input input_93,input input_94,input input_95,input input_96,input input_97,input input_98,input input_99,input input_100,input input_101,input input_102,input input_103,input input_104,input input_105,input input_106,input input_107,input input_108,input input_109,input input_110,input input_111,input input_112,input input_113,input input_114,input input_115,input input_116,input input_117,input input_118,input input_119,input input_120,input input_121,input input_122,input input_123,input input_124,input input_125,input input_126,input input_127
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_000000 (.a(t0_0000000), .b(t0_0000001), .y(t0_000000));
wire t0_0000000, t0_0000001;
mixer mix_t0_0000000 (.a(t0_00000000), .b(t0_00000001), .y(t0_0000000));
wire t0_00000000, t0_00000001;
mixer mix_t0_0000001 (.a(t0_00000010), .b(t0_00000011), .y(t0_0000001));
wire t0_00000010, t0_00000011;
mixer mix_t0_000001 (.a(t0_0000010), .b(t0_0000011), .y(t0_000001));
wire t0_0000010, t0_0000011;
mixer mix_t0_0000010 (.a(t0_00000100), .b(t0_00000101), .y(t0_0000010));
wire t0_00000100, t0_00000101;
mixer mix_t0_0000011 (.a(t0_00000110), .b(t0_00000111), .y(t0_0000011));
wire t0_00000110, t0_00000111;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_000010 (.a(t0_0000100), .b(t0_0000101), .y(t0_000010));
wire t0_0000100, t0_0000101;
mixer mix_t0_0000100 (.a(t0_00001000), .b(t0_00001001), .y(t0_0000100));
wire t0_00001000, t0_00001001;
mixer mix_t0_0000101 (.a(t0_00001010), .b(t0_00001011), .y(t0_0000101));
wire t0_00001010, t0_00001011;
mixer mix_t0_000011 (.a(t0_0000110), .b(t0_0000111), .y(t0_000011));
wire t0_0000110, t0_0000111;
mixer mix_t0_0000110 (.a(t0_00001100), .b(t0_00001101), .y(t0_0000110));
wire t0_00001100, t0_00001101;
mixer mix_t0_0000111 (.a(t0_00001110), .b(t0_00001111), .y(t0_0000111));
wire t0_00001110, t0_00001111;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_000100 (.a(t0_0001000), .b(t0_0001001), .y(t0_000100));
wire t0_0001000, t0_0001001;
mixer mix_t0_0001000 (.a(t0_00010000), .b(t0_00010001), .y(t0_0001000));
wire t0_00010000, t0_00010001;
mixer mix_t0_0001001 (.a(t0_00010010), .b(t0_00010011), .y(t0_0001001));
wire t0_00010010, t0_00010011;
mixer mix_t0_000101 (.a(t0_0001010), .b(t0_0001011), .y(t0_000101));
wire t0_0001010, t0_0001011;
mixer mix_t0_0001010 (.a(t0_00010100), .b(t0_00010101), .y(t0_0001010));
wire t0_00010100, t0_00010101;
mixer mix_t0_0001011 (.a(t0_00010110), .b(t0_00010111), .y(t0_0001011));
wire t0_00010110, t0_00010111;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_000110 (.a(t0_0001100), .b(t0_0001101), .y(t0_000110));
wire t0_0001100, t0_0001101;
mixer mix_t0_0001100 (.a(t0_00011000), .b(t0_00011001), .y(t0_0001100));
wire t0_00011000, t0_00011001;
mixer mix_t0_0001101 (.a(t0_00011010), .b(t0_00011011), .y(t0_0001101));
wire t0_00011010, t0_00011011;
mixer mix_t0_000111 (.a(t0_0001110), .b(t0_0001111), .y(t0_000111));
wire t0_0001110, t0_0001111;
mixer mix_t0_0001110 (.a(t0_00011100), .b(t0_00011101), .y(t0_0001110));
wire t0_00011100, t0_00011101;
mixer mix_t0_0001111 (.a(t0_00011110), .b(t0_00011111), .y(t0_0001111));
wire t0_00011110, t0_00011111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_001000 (.a(t0_0010000), .b(t0_0010001), .y(t0_001000));
wire t0_0010000, t0_0010001;
mixer mix_t0_0010000 (.a(t0_00100000), .b(t0_00100001), .y(t0_0010000));
wire t0_00100000, t0_00100001;
mixer mix_t0_0010001 (.a(t0_00100010), .b(t0_00100011), .y(t0_0010001));
wire t0_00100010, t0_00100011;
mixer mix_t0_001001 (.a(t0_0010010), .b(t0_0010011), .y(t0_001001));
wire t0_0010010, t0_0010011;
mixer mix_t0_0010010 (.a(t0_00100100), .b(t0_00100101), .y(t0_0010010));
wire t0_00100100, t0_00100101;
mixer mix_t0_0010011 (.a(t0_00100110), .b(t0_00100111), .y(t0_0010011));
wire t0_00100110, t0_00100111;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_001010 (.a(t0_0010100), .b(t0_0010101), .y(t0_001010));
wire t0_0010100, t0_0010101;
mixer mix_t0_0010100 (.a(t0_00101000), .b(t0_00101001), .y(t0_0010100));
wire t0_00101000, t0_00101001;
mixer mix_t0_0010101 (.a(t0_00101010), .b(t0_00101011), .y(t0_0010101));
wire t0_00101010, t0_00101011;
mixer mix_t0_001011 (.a(t0_0010110), .b(t0_0010111), .y(t0_001011));
wire t0_0010110, t0_0010111;
mixer mix_t0_0010110 (.a(t0_00101100), .b(t0_00101101), .y(t0_0010110));
wire t0_00101100, t0_00101101;
mixer mix_t0_0010111 (.a(t0_00101110), .b(t0_00101111), .y(t0_0010111));
wire t0_00101110, t0_00101111;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_001100 (.a(t0_0011000), .b(t0_0011001), .y(t0_001100));
wire t0_0011000, t0_0011001;
mixer mix_t0_0011000 (.a(t0_00110000), .b(t0_00110001), .y(t0_0011000));
wire t0_00110000, t0_00110001;
mixer mix_t0_0011001 (.a(t0_00110010), .b(t0_00110011), .y(t0_0011001));
wire t0_00110010, t0_00110011;
mixer mix_t0_001101 (.a(t0_0011010), .b(t0_0011011), .y(t0_001101));
wire t0_0011010, t0_0011011;
mixer mix_t0_0011010 (.a(t0_00110100), .b(t0_00110101), .y(t0_0011010));
wire t0_00110100, t0_00110101;
mixer mix_t0_0011011 (.a(t0_00110110), .b(t0_00110111), .y(t0_0011011));
wire t0_00110110, t0_00110111;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_001110 (.a(t0_0011100), .b(t0_0011101), .y(t0_001110));
wire t0_0011100, t0_0011101;
mixer mix_t0_0011100 (.a(t0_00111000), .b(t0_00111001), .y(t0_0011100));
wire t0_00111000, t0_00111001;
mixer mix_t0_0011101 (.a(t0_00111010), .b(t0_00111011), .y(t0_0011101));
wire t0_00111010, t0_00111011;
mixer mix_t0_001111 (.a(t0_0011110), .b(t0_0011111), .y(t0_001111));
wire t0_0011110, t0_0011111;
mixer mix_t0_0011110 (.a(t0_00111100), .b(t0_00111101), .y(t0_0011110));
wire t0_00111100, t0_00111101;
mixer mix_t0_0011111 (.a(t0_00111110), .b(t0_00111111), .y(t0_0011111));
wire t0_00111110, t0_00111111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_010000 (.a(t0_0100000), .b(t0_0100001), .y(t0_010000));
wire t0_0100000, t0_0100001;
mixer mix_t0_0100000 (.a(t0_01000000), .b(t0_01000001), .y(t0_0100000));
wire t0_01000000, t0_01000001;
mixer mix_t0_0100001 (.a(t0_01000010), .b(t0_01000011), .y(t0_0100001));
wire t0_01000010, t0_01000011;
mixer mix_t0_010001 (.a(t0_0100010), .b(t0_0100011), .y(t0_010001));
wire t0_0100010, t0_0100011;
mixer mix_t0_0100010 (.a(t0_01000100), .b(t0_01000101), .y(t0_0100010));
wire t0_01000100, t0_01000101;
mixer mix_t0_0100011 (.a(t0_01000110), .b(t0_01000111), .y(t0_0100011));
wire t0_01000110, t0_01000111;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_010010 (.a(t0_0100100), .b(t0_0100101), .y(t0_010010));
wire t0_0100100, t0_0100101;
mixer mix_t0_0100100 (.a(t0_01001000), .b(t0_01001001), .y(t0_0100100));
wire t0_01001000, t0_01001001;
mixer mix_t0_0100101 (.a(t0_01001010), .b(t0_01001011), .y(t0_0100101));
wire t0_01001010, t0_01001011;
mixer mix_t0_010011 (.a(t0_0100110), .b(t0_0100111), .y(t0_010011));
wire t0_0100110, t0_0100111;
mixer mix_t0_0100110 (.a(t0_01001100), .b(t0_01001101), .y(t0_0100110));
wire t0_01001100, t0_01001101;
mixer mix_t0_0100111 (.a(t0_01001110), .b(t0_01001111), .y(t0_0100111));
wire t0_01001110, t0_01001111;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_010100 (.a(t0_0101000), .b(t0_0101001), .y(t0_010100));
wire t0_0101000, t0_0101001;
mixer mix_t0_0101000 (.a(t0_01010000), .b(t0_01010001), .y(t0_0101000));
wire t0_01010000, t0_01010001;
mixer mix_t0_0101001 (.a(t0_01010010), .b(t0_01010011), .y(t0_0101001));
wire t0_01010010, t0_01010011;
mixer mix_t0_010101 (.a(t0_0101010), .b(t0_0101011), .y(t0_010101));
wire t0_0101010, t0_0101011;
mixer mix_t0_0101010 (.a(t0_01010100), .b(t0_01010101), .y(t0_0101010));
wire t0_01010100, t0_01010101;
mixer mix_t0_0101011 (.a(t0_01010110), .b(t0_01010111), .y(t0_0101011));
wire t0_01010110, t0_01010111;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_010110 (.a(t0_0101100), .b(t0_0101101), .y(t0_010110));
wire t0_0101100, t0_0101101;
mixer mix_t0_0101100 (.a(t0_01011000), .b(t0_01011001), .y(t0_0101100));
wire t0_01011000, t0_01011001;
mixer mix_t0_0101101 (.a(t0_01011010), .b(t0_01011011), .y(t0_0101101));
wire t0_01011010, t0_01011011;
mixer mix_t0_010111 (.a(t0_0101110), .b(t0_0101111), .y(t0_010111));
wire t0_0101110, t0_0101111;
mixer mix_t0_0101110 (.a(t0_01011100), .b(t0_01011101), .y(t0_0101110));
wire t0_01011100, t0_01011101;
mixer mix_t0_0101111 (.a(t0_01011110), .b(t0_01011111), .y(t0_0101111));
wire t0_01011110, t0_01011111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_011000 (.a(t0_0110000), .b(t0_0110001), .y(t0_011000));
wire t0_0110000, t0_0110001;
mixer mix_t0_0110000 (.a(t0_01100000), .b(t0_01100001), .y(t0_0110000));
wire t0_01100000, t0_01100001;
mixer mix_t0_0110001 (.a(t0_01100010), .b(t0_01100011), .y(t0_0110001));
wire t0_01100010, t0_01100011;
mixer mix_t0_011001 (.a(t0_0110010), .b(t0_0110011), .y(t0_011001));
wire t0_0110010, t0_0110011;
mixer mix_t0_0110010 (.a(t0_01100100), .b(t0_01100101), .y(t0_0110010));
wire t0_01100100, t0_01100101;
mixer mix_t0_0110011 (.a(t0_01100110), .b(t0_01100111), .y(t0_0110011));
wire t0_01100110, t0_01100111;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_011010 (.a(t0_0110100), .b(t0_0110101), .y(t0_011010));
wire t0_0110100, t0_0110101;
mixer mix_t0_0110100 (.a(t0_01101000), .b(t0_01101001), .y(t0_0110100));
wire t0_01101000, t0_01101001;
mixer mix_t0_0110101 (.a(t0_01101010), .b(t0_01101011), .y(t0_0110101));
wire t0_01101010, t0_01101011;
mixer mix_t0_011011 (.a(t0_0110110), .b(t0_0110111), .y(t0_011011));
wire t0_0110110, t0_0110111;
mixer mix_t0_0110110 (.a(t0_01101100), .b(t0_01101101), .y(t0_0110110));
wire t0_01101100, t0_01101101;
mixer mix_t0_0110111 (.a(t0_01101110), .b(t0_01101111), .y(t0_0110111));
wire t0_01101110, t0_01101111;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_011100 (.a(t0_0111000), .b(t0_0111001), .y(t0_011100));
wire t0_0111000, t0_0111001;
mixer mix_t0_0111000 (.a(t0_01110000), .b(t0_01110001), .y(t0_0111000));
wire t0_01110000, t0_01110001;
mixer mix_t0_0111001 (.a(t0_01110010), .b(t0_01110011), .y(t0_0111001));
wire t0_01110010, t0_01110011;
mixer mix_t0_011101 (.a(t0_0111010), .b(t0_0111011), .y(t0_011101));
wire t0_0111010, t0_0111011;
mixer mix_t0_0111010 (.a(t0_01110100), .b(t0_01110101), .y(t0_0111010));
wire t0_01110100, t0_01110101;
mixer mix_t0_0111011 (.a(t0_01110110), .b(t0_01110111), .y(t0_0111011));
wire t0_01110110, t0_01110111;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
mixer mix_t0_011110 (.a(t0_0111100), .b(t0_0111101), .y(t0_011110));
wire t0_0111100, t0_0111101;
mixer mix_t0_0111100 (.a(t0_01111000), .b(t0_01111001), .y(t0_0111100));
wire t0_01111000, t0_01111001;
mixer mix_t0_0111101 (.a(t0_01111010), .b(t0_01111011), .y(t0_0111101));
wire t0_01111010, t0_01111011;
mixer mix_t0_011111 (.a(t0_0111110), .b(t0_0111111), .y(t0_011111));
wire t0_0111110, t0_0111111;
mixer mix_t0_0111110 (.a(t0_01111100), .b(t0_01111101), .y(t0_0111110));
wire t0_01111100, t0_01111101;
mixer mix_t0_0111111 (.a(t0_01111110), .b(t0_01111111), .y(t0_0111111));
wire t0_01111110, t0_01111111;
wire t0_0;
assign out_0 = t0_0;
assign input_0 = t0_00000000;
assign input_1 = t0_00000001;
assign input_2 = t0_00000010;
assign input_3 = t0_00000011;
assign input_4 = t0_00000100;
assign input_5 = t0_00000101;
assign input_6 = t0_00000110;
assign input_7 = t0_00000111;
assign input_8 = t0_00001000;
assign input_9 = t0_00001001;
assign input_10 = t0_00001010;
assign input_11 = t0_00001011;
assign input_12 = t0_00001100;
assign input_13 = t0_00001101;
assign input_14 = t0_00001110;
assign input_15 = t0_00001111;
assign input_16 = t0_00010000;
assign input_17 = t0_00010001;
assign input_18 = t0_00010010;
assign input_19 = t0_00010011;
assign input_20 = t0_00010100;
assign input_21 = t0_00010101;
assign input_22 = t0_00010110;
assign input_23 = t0_00010111;
assign input_24 = t0_00011000;
assign input_25 = t0_00011001;
assign input_26 = t0_00011010;
assign input_27 = t0_00011011;
assign input_28 = t0_00011100;
assign input_29 = t0_00011101;
assign input_30 = t0_00011110;
assign input_31 = t0_00011111;
assign input_32 = t0_00100000;
assign input_33 = t0_00100001;
assign input_34 = t0_00100010;
assign input_35 = t0_00100011;
assign input_36 = t0_00100100;
assign input_37 = t0_00100101;
assign input_38 = t0_00100110;
assign input_39 = t0_00100111;
assign input_40 = t0_00101000;
assign input_41 = t0_00101001;
assign input_42 = t0_00101010;
assign input_43 = t0_00101011;
assign input_44 = t0_00101100;
assign input_45 = t0_00101101;
assign input_46 = t0_00101110;
assign input_47 = t0_00101111;
assign input_48 = t0_00110000;
assign input_49 = t0_00110001;
assign input_50 = t0_00110010;
assign input_51 = t0_00110011;
assign input_52 = t0_00110100;
assign input_53 = t0_00110101;
assign input_54 = t0_00110110;
assign input_55 = t0_00110111;
assign input_56 = t0_00111000;
assign input_57 = t0_00111001;
assign input_58 = t0_00111010;
assign input_59 = t0_00111011;
assign input_60 = t0_00111100;
assign input_61 = t0_00111101;
assign input_62 = t0_00111110;
assign input_63 = t0_00111111;
assign input_64 = t0_01000000;
assign input_65 = t0_01000001;
assign input_66 = t0_01000010;
assign input_67 = t0_01000011;
assign input_68 = t0_01000100;
assign input_69 = t0_01000101;
assign input_70 = t0_01000110;
assign input_71 = t0_01000111;
assign input_72 = t0_01001000;
assign input_73 = t0_01001001;
assign input_74 = t0_01001010;
assign input_75 = t0_01001011;
assign input_76 = t0_01001100;
assign input_77 = t0_01001101;
assign input_78 = t0_01001110;
assign input_79 = t0_01001111;
assign input_80 = t0_01010000;
assign input_81 = t0_01010001;
assign input_82 = t0_01010010;
assign input_83 = t0_01010011;
assign input_84 = t0_01010100;
assign input_85 = t0_01010101;
assign input_86 = t0_01010110;
assign input_87 = t0_01010111;
assign input_88 = t0_01011000;
assign input_89 = t0_01011001;
assign input_90 = t0_01011010;
assign input_91 = t0_01011011;
assign input_92 = t0_01011100;
assign input_93 = t0_01011101;
assign input_94 = t0_01011110;
assign input_95 = t0_01011111;
assign input_96 = t0_01100000;
assign input_97 = t0_01100001;
assign input_98 = t0_01100010;
assign input_99 = t0_01100011;
assign input_100 = t0_01100100;
assign input_101 = t0_01100101;
assign input_102 = t0_01100110;
assign input_103 = t0_01100111;
assign input_104 = t0_01101000;
assign input_105 = t0_01101001;
assign input_106 = t0_01101010;
assign input_107 = t0_01101011;
assign input_108 = t0_01101100;
assign input_109 = t0_01101101;
assign input_110 = t0_01101110;
assign input_111 = t0_01101111;
assign input_112 = t0_01110000;
assign input_113 = t0_01110001;
assign input_114 = t0_01110010;
assign input_115 = t0_01110011;
assign input_116 = t0_01110100;
assign input_117 = t0_01110101;
assign input_118 = t0_01110110;
assign input_119 = t0_01110111;
assign input_120 = t0_01111000;
assign input_121 = t0_01111001;
assign input_122 = t0_01111010;
assign input_123 = t0_01111011;
assign input_124 = t0_01111100;
assign input_125 = t0_01111101;
assign input_126 = t0_01111110;
assign input_127 = t0_01111111;
endmodule
