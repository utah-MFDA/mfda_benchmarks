module chain_mixer_64 (
output j64,input j0,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64,input k64
);
mixer m0(.a(in), .b(k0), .y(j1));
wire j1;
wire j2;
wire j3;
wire j4;
wire j5;
wire j6;
wire j7;
wire j8;
wire j9;
wire j10;
wire j11;
wire j12;
wire j13;
wire j14;
wire j15;
wire j16;
wire j17;
wire j18;
wire j19;
wire j20;
wire j21;
wire j22;
wire j23;
wire j24;
wire j25;
wire j26;
wire j27;
wire j28;
wire j29;
wire j30;
wire j31;
wire j32;
wire j33;
wire j34;
wire j35;
wire j36;
wire j37;
wire j38;
wire j39;
wire j40;
wire j41;
wire j42;
wire j43;
wire j44;
wire j45;
wire j46;
wire j47;
wire j48;
wire j49;
wire j50;
wire j51;
wire j52;
wire j53;
wire j54;
wire j55;
wire j56;
wire j57;
wire j58;
wire j59;
wire j60;
wire j61;
wire j62;
wire j63;
mixer m0(.a(j0), .b(k0), .y(j1));
mixer m1(.a(j1), .b(k1), .y(j2));
mixer m2(.a(j2), .b(k2), .y(j3));
mixer m3(.a(j3), .b(k3), .y(j4));
mixer m4(.a(j4), .b(k4), .y(j5));
mixer m5(.a(j5), .b(k5), .y(j6));
mixer m6(.a(j6), .b(k6), .y(j7));
mixer m7(.a(j7), .b(k7), .y(j8));
mixer m8(.a(j8), .b(k8), .y(j9));
mixer m9(.a(j9), .b(k9), .y(j10));
mixer m10(.a(j10), .b(k10), .y(j11));
mixer m11(.a(j11), .b(k11), .y(j12));
mixer m12(.a(j12), .b(k12), .y(j13));
mixer m13(.a(j13), .b(k13), .y(j14));
mixer m14(.a(j14), .b(k14), .y(j15));
mixer m15(.a(j15), .b(k15), .y(j16));
mixer m16(.a(j16), .b(k16), .y(j17));
mixer m17(.a(j17), .b(k17), .y(j18));
mixer m18(.a(j18), .b(k18), .y(j19));
mixer m19(.a(j19), .b(k19), .y(j20));
mixer m20(.a(j20), .b(k20), .y(j21));
mixer m21(.a(j21), .b(k21), .y(j22));
mixer m22(.a(j22), .b(k22), .y(j23));
mixer m23(.a(j23), .b(k23), .y(j24));
mixer m24(.a(j24), .b(k24), .y(j25));
mixer m25(.a(j25), .b(k25), .y(j26));
mixer m26(.a(j26), .b(k26), .y(j27));
mixer m27(.a(j27), .b(k27), .y(j28));
mixer m28(.a(j28), .b(k28), .y(j29));
mixer m29(.a(j29), .b(k29), .y(j30));
mixer m30(.a(j30), .b(k30), .y(j31));
mixer m31(.a(j31), .b(k31), .y(j32));
mixer m32(.a(j32), .b(k32), .y(j33));
mixer m33(.a(j33), .b(k33), .y(j34));
mixer m34(.a(j34), .b(k34), .y(j35));
mixer m35(.a(j35), .b(k35), .y(j36));
mixer m36(.a(j36), .b(k36), .y(j37));
mixer m37(.a(j37), .b(k37), .y(j38));
mixer m38(.a(j38), .b(k38), .y(j39));
mixer m39(.a(j39), .b(k39), .y(j40));
mixer m40(.a(j40), .b(k40), .y(j41));
mixer m41(.a(j41), .b(k41), .y(j42));
mixer m42(.a(j42), .b(k42), .y(j43));
mixer m43(.a(j43), .b(k43), .y(j44));
mixer m44(.a(j44), .b(k44), .y(j45));
mixer m45(.a(j45), .b(k45), .y(j46));
mixer m46(.a(j46), .b(k46), .y(j47));
mixer m47(.a(j47), .b(k47), .y(j48));
mixer m48(.a(j48), .b(k48), .y(j49));
mixer m49(.a(j49), .b(k49), .y(j50));
mixer m50(.a(j50), .b(k50), .y(j51));
mixer m51(.a(j51), .b(k51), .y(j52));
mixer m52(.a(j52), .b(k52), .y(j53));
mixer m53(.a(j53), .b(k53), .y(j54));
mixer m54(.a(j54), .b(k54), .y(j55));
mixer m55(.a(j55), .b(k55), .y(j56));
mixer m56(.a(j56), .b(k56), .y(j57));
mixer m57(.a(j57), .b(k57), .y(j58));
mixer m58(.a(j58), .b(k58), .y(j59));
mixer m59(.a(j59), .b(k59), .y(j60));
mixer m60(.a(j60), .b(k60), .y(j61));
mixer m61(.a(j61), .b(k61), .y(j62));
mixer m62(.a(j62), .b(k62), .y(j63));
mixer m63(.a(j63), .b(k63), .y(j64));
endmodule
