module galaban11();
	mixer m_0(.a(e_0_1), .b(e_0_2), .y(e_0_3));
	mixer m_1(.a(e_0_1), .b(e_1_106), .y(e_1_108));
	mixer m_2(.a(e_0_2), .b(e_2_107), .y(e_2_109));
	mixer m_3(.a(e_0_3), .b(e_3_110), .y(e_3_111));
	mixer m_4(.a(e_4_7), .b(e_4_64), .y(e_4_66));
	mixer m_5(.a(e_5_6), .b(e_5_62), .y(e_5_67));
	mixer m_6(.a(e_5_6), .b(e_6_68), .y(e_6_69));
	mixer m_7(.a(e_4_7), .b(e_7_63), .y(e_7_65));
	mixer m_8(.a(e_8_16), .b(e_8_46), .y(e_8_47));
	mixer m_9(.a(e_9_17), .b(e_9_48), .y(e_9_52));
	mixer m_10(.a(e_10_17), .b(e_10_49), .y(e_10_51));
	mixer m_11(.a(e_11_16), .b(e_11_50), .y(e_11_53));
	mixer m_12(.a(e_12_18), .b(e_12_54), .y(e_12_61));
	mixer m_13(.a(e_13_19), .b(e_13_55), .y(e_13_60));
	mixer m_14(.a(e_14_19), .b(e_14_57), .y(e_14_59));
	mixer m_15(.a(e_15_18), .b(e_15_56), .y(e_15_58));
	mixer m_16(.a(e_8_16), .b(e_11_16), .y(e_16_20));
	mixer m_17(.a(e_9_17), .b(e_10_17), .y(e_17_20));
	mixer m_18(.a(e_12_18), .b(e_15_18), .y(e_18_21));
	mixer m_19(.a(e_13_19), .b(e_14_19), .y(e_19_21));
	mixer m_20(.a(e_16_20), .b(e_17_20), .y(e_20_21));
	mixer m_21(.a(e_18_21), .b(e_19_21), .y(e_20_21));
	mixer m_22(.a(e_22_24), .b(e_22_38), .y(e_22_92));
	mixer m_23(.a(e_23_25), .b(e_23_43), .y(e_23_87));
	mixer m_24(.a(e_22_24), .b(e_24_40), .y(e_24_90));
	mixer m_25(.a(e_23_25), .b(e_25_42), .y(e_25_89));
	mixer m_26(.a(e_26_28), .b(e_26_39), .y(e_26_91));
	mixer m_27(.a(e_27_29), .b(e_27_41), .y(e_27_86));
	mixer m_28(.a(e_26_28), .b(e_28_45), .y(e_28_93));
	mixer m_29(.a(e_27_29), .b(e_29_44), .y(e_29_88));
	mixer m_30(.a(e_30_46), .b(e_30_62), .y(e_30_70));
	mixer m_31(.a(e_31_47), .b(e_31_64), .y(e_31_74));
	mixer m_32(.a(e_32_52), .b(e_32_67), .y(e_32_77));
	mixer m_33(.a(e_33_48), .b(e_33_66), .y(e_33_71));
	mixer m_34(.a(e_34_49), .b(e_34_65), .y(e_34_72));
	mixer m_35(.a(e_35_53), .b(e_35_69), .y(e_35_73));
	mixer m_36(.a(e_36_50), .b(e_36_63), .y(e_36_76));
	mixer m_37(.a(e_37_51), .b(e_37_68), .y(e_37_75));
	mixer m_38(.a(e_22_38), .b(e_38_54), .y(e_38_70));
	mixer m_39(.a(e_26_39), .b(e_39_61), .y(e_39_74));
	mixer m_40(.a(e_24_40), .b(e_40_55), .y(e_40_77));
	mixer m_41(.a(e_27_41), .b(e_41_57), .y(e_41_73));
	mixer m_42(.a(e_25_42), .b(e_42_59), .y(e_42_76));
	mixer m_43(.a(e_23_43), .b(e_43_58), .y(e_43_72));
	mixer m_44(.a(e_29_44), .b(e_44_56), .y(e_44_75));
	mixer m_45(.a(e_28_45), .b(e_45_60), .y(e_45_71));
	mixer m_46(.a(e_8_46), .b(e_30_46), .y(e_46_88));
	mixer m_47(.a(e_8_47), .b(e_31_47), .y(e_47_87));
	mixer m_48(.a(e_9_48), .b(e_33_48), .y(e_48_89));
	mixer m_49(.a(e_10_49), .b(e_34_49), .y(e_49_91));
	mixer m_50(.a(e_11_50), .b(e_36_50), .y(e_50_93));
	mixer m_51(.a(e_10_51), .b(e_37_51), .y(e_51_92));
	mixer m_52(.a(e_9_52), .b(e_32_52), .y(e_52_86));
	mixer m_53(.a(e_11_53), .b(e_35_53), .y(e_53_90));
	mixer m_54(.a(e_12_54), .b(e_38_54), .y(e_54_78));
	mixer m_55(.a(e_13_55), .b(e_40_55), .y(e_55_80));
	mixer m_56(.a(e_15_56), .b(e_44_56), .y(e_56_82));
	mixer m_57(.a(e_14_57), .b(e_41_57), .y(e_57_84));
	mixer m_58(.a(e_15_58), .b(e_43_58), .y(e_58_85));
	mixer m_59(.a(e_14_59), .b(e_42_59), .y(e_59_83));
	mixer m_60(.a(e_13_60), .b(e_45_60), .y(e_60_79));
	mixer m_61(.a(e_12_61), .b(e_39_61), .y(e_61_81));
	mixer m_62(.a(e_5_62), .b(e_30_62), .y(e_62_83));
	mixer m_63(.a(e_7_63), .b(e_36_63), .y(e_63_78));
	mixer m_64(.a(e_4_64), .b(e_31_64), .y(e_64_84));
	mixer m_65(.a(e_7_65), .b(e_34_65), .y(e_65_80));
	mixer m_66(.a(e_4_66), .b(e_33_66), .y(e_66_82));
	mixer m_67(.a(e_5_67), .b(e_32_67), .y(e_67_85));
	mixer m_68(.a(e_6_68), .b(e_37_68), .y(e_68_79));
	mixer m_69(.a(e_6_69), .b(e_35_69), .y(e_69_81));
	mixer m_70(.a(e_30_70), .b(e_38_70), .y(e_70_102));
	mixer m_71(.a(e_33_71), .b(e_45_71), .y(e_71_102));
	mixer m_72(.a(e_34_72), .b(e_43_72), .y(e_72_105));
	mixer m_73(.a(e_35_73), .b(e_41_73), .y(e_73_105));
	mixer m_74(.a(e_31_74), .b(e_39_74), .y(e_74_103));
	mixer m_75(.a(e_37_75), .b(e_44_75), .y(e_75_104));
	mixer m_76(.a(e_36_76), .b(e_42_76), .y(e_76_104));
	mixer m_77(.a(e_32_77), .b(e_40_77), .y(e_77_103));
	mixer m_78(.a(e_54_78), .b(e_63_78), .y(e_78_94));
	mixer m_79(.a(e_60_79), .b(e_68_79), .y(e_79_95));
	mixer m_80(.a(e_55_80), .b(e_65_80), .y(e_80_96));
	mixer m_81(.a(e_61_81), .b(e_69_81), .y(e_81_97));
	mixer m_82(.a(e_56_82), .b(e_66_82), .y(e_82_98));
	mixer m_83(.a(e_59_83), .b(e_62_83), .y(e_83_101));
	mixer m_84(.a(e_57_84), .b(e_64_84), .y(e_84_100));
	mixer m_85(.a(e_58_85), .b(e_67_85), .y(e_85_99));
	mixer m_86(.a(e_27_86), .b(e_52_86), .y(e_86_94));
	mixer m_87(.a(e_23_87), .b(e_47_87), .y(e_87_95));
	mixer m_88(.a(e_29_88), .b(e_46_88), .y(e_88_96));
	mixer m_89(.a(e_25_89), .b(e_48_89), .y(e_89_97));
	mixer m_90(.a(e_24_90), .b(e_53_90), .y(e_90_98));
	mixer m_91(.a(e_26_91), .b(e_49_91), .y(e_91_101));
	mixer m_92(.a(e_22_92), .b(e_51_92), .y(e_92_100));
	mixer m_93(.a(e_28_93), .b(e_50_93), .y(e_93_99));
	mixer m_94(.a(e_78_94), .b(e_86_94), .y(e_94_106));
	mixer m_95(.a(e_79_95), .b(e_87_95), .y(e_95_106));
	mixer m_96(.a(e_80_96), .b(e_88_96), .y(e_96_107));
	mixer m_97(.a(e_81_97), .b(e_89_97), .y(e_97_107));
	mixer m_98(.a(e_82_98), .b(e_90_98), .y(e_98_108));
	mixer m_99(.a(e_85_99), .b(e_93_99), .y(e_99_109));
	mixer m_100(.a(e_84_100), .b(e_92_100), .y(e_100_109));
	mixer m_101(.a(e_83_101), .b(e_91_101), .y(e_101_108));
	mixer m_102(.a(e_70_102), .b(e_71_102), .y(e_102_110));
	mixer m_103(.a(e_74_103), .b(e_77_103), .y(e_103_111));
	mixer m_104(.a(e_75_104), .b(e_76_104), .y(e_104_111));
	mixer m_105(.a(e_72_105), .b(e_73_105), .y(e_105_110));
	mixer m_106(.a(e_1_106), .b(e_94_106), .y(e_95_106));
	mixer m_107(.a(e_2_107), .b(e_96_107), .y(e_97_107));
	mixer m_108(.a(e_1_108), .b(e_98_108), .y(e_101_108));
	mixer m_109(.a(e_2_109), .b(e_99_109), .y(e_100_109));
	mixer m_110(.a(e_3_110), .b(e_102_110), .y(e_105_110));
	mixer m_111(.a(e_3_111), .b(e_103_111), .y(e_104_111));
wire e_0_1,
	e_0_2,
	e_0_3,
	e_1_106,
	e_1_108,
	e_2_107,
	e_2_109,
	e_3_110,
	e_3_111,
	e_4_7,
	e_4_64,
	e_4_66,
	e_5_6,
	e_5_62,
	e_5_67,
	e_6_68,
	e_6_69,
	e_7_63,
	e_7_65,
	e_8_16,
	e_8_46,
	e_8_47,
	e_9_17,
	e_9_48,
	e_9_52,
	e_10_17,
	e_10_49,
	e_10_51,
	e_11_16,
	e_11_50,
	e_11_53,
	e_12_18,
	e_12_54,
	e_12_61,
	e_13_19,
	e_13_55,
	e_13_60,
	e_14_19,
	e_14_57,
	e_14_59,
	e_15_18,
	e_15_56,
	e_15_58,
	e_16_20,
	e_17_20,
	e_18_21,
	e_19_21,
	e_20_21,
	e_22_24,
	e_22_38,
	e_22_92,
	e_23_25,
	e_23_43,
	e_23_87,
	e_24_40,
	e_24_90,
	e_25_42,
	e_25_89,
	e_26_28,
	e_26_39,
	e_26_91,
	e_27_29,
	e_27_41,
	e_27_86,
	e_28_45,
	e_28_93,
	e_29_44,
	e_29_88,
	e_30_46,
	e_30_62,
	e_30_70,
	e_31_47,
	e_31_64,
	e_31_74,
	e_32_52,
	e_32_67,
	e_32_77,
	e_33_48,
	e_33_66,
	e_33_71,
	e_34_49,
	e_34_65,
	e_34_72,
	e_35_53,
	e_35_69,
	e_35_73,
	e_36_50,
	e_36_63,
	e_36_76,
	e_37_51,
	e_37_68,
	e_37_75,
	e_38_54,
	e_38_70,
	e_39_61,
	e_39_74,
	e_40_55,
	e_40_77,
	e_41_57,
	e_41_73,
	e_42_59,
	e_42_76,
	e_43_58,
	e_43_72,
	e_44_56,
	e_44_75,
	e_45_60,
	e_45_71,
	e_46_88,
	e_47_87,
	e_48_89,
	e_49_91,
	e_50_93,
	e_51_92,
	e_52_86,
	e_53_90,
	e_54_78,
	e_55_80,
	e_56_82,
	e_57_84,
	e_58_85,
	e_59_83,
	e_60_79,
	e_61_81,
	e_62_83,
	e_63_78,
	e_64_84,
	e_65_80,
	e_66_82,
	e_67_85,
	e_68_79,
	e_69_81,
	e_70_102,
	e_71_102,
	e_72_105,
	e_73_105,
	e_74_103,
	e_75_104,
	e_76_104,
	e_77_103,
	e_78_94,
	e_79_95,
	e_80_96,
	e_81_97,
	e_82_98,
	e_83_101,
	e_84_100,
	e_85_99,
	e_86_94,
	e_87_95,
	e_88_96,
	e_89_97,
	e_90_98,
	e_91_101,
	e_92_100,
	e_93_99,
	e_94_106,
	e_95_106,
	e_96_107,
	e_97_107,
	e_98_108,
	e_99_109,
	e_100_109,
	e_101_108,
	e_102_110,
	e_103_111,
	e_104_111,
	e_105_110;
endmodule
