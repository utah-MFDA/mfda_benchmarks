module complete_64 (
inout io_0,inout io_1,inout io_2,inout io_3,inout io_4,inout io_5,inout io_6,inout io_7,inout io_8,inout io_9,inout io_10,inout io_11,inout io_12,inout io_13,inout io_14,inout io_15,inout io_16,inout io_17,inout io_18,inout io_19,inout io_20,inout io_21,inout io_22,inout io_23,inout io_24,inout io_25,inout io_26,inout io_27,inout io_28,inout io_29,inout io_30,inout io_31,inout io_32,inout io_33,inout io_34,inout io_35,inout io_36,inout io_37,inout io_38,inout io_39,inout io_40,inout io_41,inout io_42,inout io_43,inout io_44,inout io_45,inout io_46,inout io_47,inout io_48,inout io_49,inout io_50,inout io_51,inout io_52,inout io_53,inout io_54,inout io_55,inout io_56,inout io_57,inout io_58,inout io_59,inout io_60,inout io_61,inout io_62,inout io_63
);
assign io_0 = input_0;
assign io_0 = input_1;
assign io_0 = input_2;
assign io_0 = input_3;
assign io_0 = input_4;
assign io_0 = input_5;
assign io_0 = input_6;
assign io_0 = input_7;
assign io_0 = input_8;
assign io_0 = input_9;
assign io_0 = input_10;
assign io_0 = input_11;
assign io_0 = input_12;
assign io_0 = input_13;
assign io_0 = input_14;
assign io_0 = input_15;
assign io_0 = input_16;
assign io_0 = input_17;
assign io_0 = input_18;
assign io_0 = input_19;
assign io_0 = input_20;
assign io_0 = input_21;
assign io_0 = input_22;
assign io_0 = input_23;
assign io_0 = input_24;
assign io_0 = input_25;
assign io_0 = input_26;
assign io_0 = input_27;
assign io_0 = input_28;
assign io_0 = input_29;
assign io_0 = input_30;
assign io_0 = input_31;
assign io_0 = input_32;
assign io_0 = input_33;
assign io_0 = input_34;
assign io_0 = input_35;
assign io_0 = input_36;
assign io_0 = input_37;
assign io_0 = input_38;
assign io_0 = input_39;
assign io_0 = input_40;
assign io_0 = input_41;
assign io_0 = input_42;
assign io_0 = input_43;
assign io_0 = input_44;
assign io_0 = input_45;
assign io_0 = input_46;
assign io_0 = input_47;
assign io_0 = input_48;
assign io_0 = input_49;
assign io_0 = input_50;
assign io_0 = input_51;
assign io_0 = input_52;
assign io_0 = input_53;
assign io_0 = input_54;
assign io_0 = input_55;
assign io_0 = input_56;
assign io_0 = input_57;
assign io_0 = input_58;
assign io_0 = input_59;
assign io_0 = input_60;
assign io_0 = input_61;
assign io_0 = input_62;
assign io_0 = input_63;
assign io_1 = input_1;
assign io_1 = input_2;
assign io_1 = input_3;
assign io_1 = input_4;
assign io_1 = input_5;
assign io_1 = input_6;
assign io_1 = input_7;
assign io_1 = input_8;
assign io_1 = input_9;
assign io_1 = input_10;
assign io_1 = input_11;
assign io_1 = input_12;
assign io_1 = input_13;
assign io_1 = input_14;
assign io_1 = input_15;
assign io_1 = input_16;
assign io_1 = input_17;
assign io_1 = input_18;
assign io_1 = input_19;
assign io_1 = input_20;
assign io_1 = input_21;
assign io_1 = input_22;
assign io_1 = input_23;
assign io_1 = input_24;
assign io_1 = input_25;
assign io_1 = input_26;
assign io_1 = input_27;
assign io_1 = input_28;
assign io_1 = input_29;
assign io_1 = input_30;
assign io_1 = input_31;
assign io_1 = input_32;
assign io_1 = input_33;
assign io_1 = input_34;
assign io_1 = input_35;
assign io_1 = input_36;
assign io_1 = input_37;
assign io_1 = input_38;
assign io_1 = input_39;
assign io_1 = input_40;
assign io_1 = input_41;
assign io_1 = input_42;
assign io_1 = input_43;
assign io_1 = input_44;
assign io_1 = input_45;
assign io_1 = input_46;
assign io_1 = input_47;
assign io_1 = input_48;
assign io_1 = input_49;
assign io_1 = input_50;
assign io_1 = input_51;
assign io_1 = input_52;
assign io_1 = input_53;
assign io_1 = input_54;
assign io_1 = input_55;
assign io_1 = input_56;
assign io_1 = input_57;
assign io_1 = input_58;
assign io_1 = input_59;
assign io_1 = input_60;
assign io_1 = input_61;
assign io_1 = input_62;
assign io_1 = input_63;
assign io_2 = input_2;
assign io_2 = input_3;
assign io_2 = input_4;
assign io_2 = input_5;
assign io_2 = input_6;
assign io_2 = input_7;
assign io_2 = input_8;
assign io_2 = input_9;
assign io_2 = input_10;
assign io_2 = input_11;
assign io_2 = input_12;
assign io_2 = input_13;
assign io_2 = input_14;
assign io_2 = input_15;
assign io_2 = input_16;
assign io_2 = input_17;
assign io_2 = input_18;
assign io_2 = input_19;
assign io_2 = input_20;
assign io_2 = input_21;
assign io_2 = input_22;
assign io_2 = input_23;
assign io_2 = input_24;
assign io_2 = input_25;
assign io_2 = input_26;
assign io_2 = input_27;
assign io_2 = input_28;
assign io_2 = input_29;
assign io_2 = input_30;
assign io_2 = input_31;
assign io_2 = input_32;
assign io_2 = input_33;
assign io_2 = input_34;
assign io_2 = input_35;
assign io_2 = input_36;
assign io_2 = input_37;
assign io_2 = input_38;
assign io_2 = input_39;
assign io_2 = input_40;
assign io_2 = input_41;
assign io_2 = input_42;
assign io_2 = input_43;
assign io_2 = input_44;
assign io_2 = input_45;
assign io_2 = input_46;
assign io_2 = input_47;
assign io_2 = input_48;
assign io_2 = input_49;
assign io_2 = input_50;
assign io_2 = input_51;
assign io_2 = input_52;
assign io_2 = input_53;
assign io_2 = input_54;
assign io_2 = input_55;
assign io_2 = input_56;
assign io_2 = input_57;
assign io_2 = input_58;
assign io_2 = input_59;
assign io_2 = input_60;
assign io_2 = input_61;
assign io_2 = input_62;
assign io_2 = input_63;
assign io_3 = input_3;
assign io_3 = input_4;
assign io_3 = input_5;
assign io_3 = input_6;
assign io_3 = input_7;
assign io_3 = input_8;
assign io_3 = input_9;
assign io_3 = input_10;
assign io_3 = input_11;
assign io_3 = input_12;
assign io_3 = input_13;
assign io_3 = input_14;
assign io_3 = input_15;
assign io_3 = input_16;
assign io_3 = input_17;
assign io_3 = input_18;
assign io_3 = input_19;
assign io_3 = input_20;
assign io_3 = input_21;
assign io_3 = input_22;
assign io_3 = input_23;
assign io_3 = input_24;
assign io_3 = input_25;
assign io_3 = input_26;
assign io_3 = input_27;
assign io_3 = input_28;
assign io_3 = input_29;
assign io_3 = input_30;
assign io_3 = input_31;
assign io_3 = input_32;
assign io_3 = input_33;
assign io_3 = input_34;
assign io_3 = input_35;
assign io_3 = input_36;
assign io_3 = input_37;
assign io_3 = input_38;
assign io_3 = input_39;
assign io_3 = input_40;
assign io_3 = input_41;
assign io_3 = input_42;
assign io_3 = input_43;
assign io_3 = input_44;
assign io_3 = input_45;
assign io_3 = input_46;
assign io_3 = input_47;
assign io_3 = input_48;
assign io_3 = input_49;
assign io_3 = input_50;
assign io_3 = input_51;
assign io_3 = input_52;
assign io_3 = input_53;
assign io_3 = input_54;
assign io_3 = input_55;
assign io_3 = input_56;
assign io_3 = input_57;
assign io_3 = input_58;
assign io_3 = input_59;
assign io_3 = input_60;
assign io_3 = input_61;
assign io_3 = input_62;
assign io_3 = input_63;
assign io_4 = input_4;
assign io_4 = input_5;
assign io_4 = input_6;
assign io_4 = input_7;
assign io_4 = input_8;
assign io_4 = input_9;
assign io_4 = input_10;
assign io_4 = input_11;
assign io_4 = input_12;
assign io_4 = input_13;
assign io_4 = input_14;
assign io_4 = input_15;
assign io_4 = input_16;
assign io_4 = input_17;
assign io_4 = input_18;
assign io_4 = input_19;
assign io_4 = input_20;
assign io_4 = input_21;
assign io_4 = input_22;
assign io_4 = input_23;
assign io_4 = input_24;
assign io_4 = input_25;
assign io_4 = input_26;
assign io_4 = input_27;
assign io_4 = input_28;
assign io_4 = input_29;
assign io_4 = input_30;
assign io_4 = input_31;
assign io_4 = input_32;
assign io_4 = input_33;
assign io_4 = input_34;
assign io_4 = input_35;
assign io_4 = input_36;
assign io_4 = input_37;
assign io_4 = input_38;
assign io_4 = input_39;
assign io_4 = input_40;
assign io_4 = input_41;
assign io_4 = input_42;
assign io_4 = input_43;
assign io_4 = input_44;
assign io_4 = input_45;
assign io_4 = input_46;
assign io_4 = input_47;
assign io_4 = input_48;
assign io_4 = input_49;
assign io_4 = input_50;
assign io_4 = input_51;
assign io_4 = input_52;
assign io_4 = input_53;
assign io_4 = input_54;
assign io_4 = input_55;
assign io_4 = input_56;
assign io_4 = input_57;
assign io_4 = input_58;
assign io_4 = input_59;
assign io_4 = input_60;
assign io_4 = input_61;
assign io_4 = input_62;
assign io_4 = input_63;
assign io_5 = input_5;
assign io_5 = input_6;
assign io_5 = input_7;
assign io_5 = input_8;
assign io_5 = input_9;
assign io_5 = input_10;
assign io_5 = input_11;
assign io_5 = input_12;
assign io_5 = input_13;
assign io_5 = input_14;
assign io_5 = input_15;
assign io_5 = input_16;
assign io_5 = input_17;
assign io_5 = input_18;
assign io_5 = input_19;
assign io_5 = input_20;
assign io_5 = input_21;
assign io_5 = input_22;
assign io_5 = input_23;
assign io_5 = input_24;
assign io_5 = input_25;
assign io_5 = input_26;
assign io_5 = input_27;
assign io_5 = input_28;
assign io_5 = input_29;
assign io_5 = input_30;
assign io_5 = input_31;
assign io_5 = input_32;
assign io_5 = input_33;
assign io_5 = input_34;
assign io_5 = input_35;
assign io_5 = input_36;
assign io_5 = input_37;
assign io_5 = input_38;
assign io_5 = input_39;
assign io_5 = input_40;
assign io_5 = input_41;
assign io_5 = input_42;
assign io_5 = input_43;
assign io_5 = input_44;
assign io_5 = input_45;
assign io_5 = input_46;
assign io_5 = input_47;
assign io_5 = input_48;
assign io_5 = input_49;
assign io_5 = input_50;
assign io_5 = input_51;
assign io_5 = input_52;
assign io_5 = input_53;
assign io_5 = input_54;
assign io_5 = input_55;
assign io_5 = input_56;
assign io_5 = input_57;
assign io_5 = input_58;
assign io_5 = input_59;
assign io_5 = input_60;
assign io_5 = input_61;
assign io_5 = input_62;
assign io_5 = input_63;
assign io_6 = input_6;
assign io_6 = input_7;
assign io_6 = input_8;
assign io_6 = input_9;
assign io_6 = input_10;
assign io_6 = input_11;
assign io_6 = input_12;
assign io_6 = input_13;
assign io_6 = input_14;
assign io_6 = input_15;
assign io_6 = input_16;
assign io_6 = input_17;
assign io_6 = input_18;
assign io_6 = input_19;
assign io_6 = input_20;
assign io_6 = input_21;
assign io_6 = input_22;
assign io_6 = input_23;
assign io_6 = input_24;
assign io_6 = input_25;
assign io_6 = input_26;
assign io_6 = input_27;
assign io_6 = input_28;
assign io_6 = input_29;
assign io_6 = input_30;
assign io_6 = input_31;
assign io_6 = input_32;
assign io_6 = input_33;
assign io_6 = input_34;
assign io_6 = input_35;
assign io_6 = input_36;
assign io_6 = input_37;
assign io_6 = input_38;
assign io_6 = input_39;
assign io_6 = input_40;
assign io_6 = input_41;
assign io_6 = input_42;
assign io_6 = input_43;
assign io_6 = input_44;
assign io_6 = input_45;
assign io_6 = input_46;
assign io_6 = input_47;
assign io_6 = input_48;
assign io_6 = input_49;
assign io_6 = input_50;
assign io_6 = input_51;
assign io_6 = input_52;
assign io_6 = input_53;
assign io_6 = input_54;
assign io_6 = input_55;
assign io_6 = input_56;
assign io_6 = input_57;
assign io_6 = input_58;
assign io_6 = input_59;
assign io_6 = input_60;
assign io_6 = input_61;
assign io_6 = input_62;
assign io_6 = input_63;
assign io_7 = input_7;
assign io_7 = input_8;
assign io_7 = input_9;
assign io_7 = input_10;
assign io_7 = input_11;
assign io_7 = input_12;
assign io_7 = input_13;
assign io_7 = input_14;
assign io_7 = input_15;
assign io_7 = input_16;
assign io_7 = input_17;
assign io_7 = input_18;
assign io_7 = input_19;
assign io_7 = input_20;
assign io_7 = input_21;
assign io_7 = input_22;
assign io_7 = input_23;
assign io_7 = input_24;
assign io_7 = input_25;
assign io_7 = input_26;
assign io_7 = input_27;
assign io_7 = input_28;
assign io_7 = input_29;
assign io_7 = input_30;
assign io_7 = input_31;
assign io_7 = input_32;
assign io_7 = input_33;
assign io_7 = input_34;
assign io_7 = input_35;
assign io_7 = input_36;
assign io_7 = input_37;
assign io_7 = input_38;
assign io_7 = input_39;
assign io_7 = input_40;
assign io_7 = input_41;
assign io_7 = input_42;
assign io_7 = input_43;
assign io_7 = input_44;
assign io_7 = input_45;
assign io_7 = input_46;
assign io_7 = input_47;
assign io_7 = input_48;
assign io_7 = input_49;
assign io_7 = input_50;
assign io_7 = input_51;
assign io_7 = input_52;
assign io_7 = input_53;
assign io_7 = input_54;
assign io_7 = input_55;
assign io_7 = input_56;
assign io_7 = input_57;
assign io_7 = input_58;
assign io_7 = input_59;
assign io_7 = input_60;
assign io_7 = input_61;
assign io_7 = input_62;
assign io_7 = input_63;
assign io_8 = input_8;
assign io_8 = input_9;
assign io_8 = input_10;
assign io_8 = input_11;
assign io_8 = input_12;
assign io_8 = input_13;
assign io_8 = input_14;
assign io_8 = input_15;
assign io_8 = input_16;
assign io_8 = input_17;
assign io_8 = input_18;
assign io_8 = input_19;
assign io_8 = input_20;
assign io_8 = input_21;
assign io_8 = input_22;
assign io_8 = input_23;
assign io_8 = input_24;
assign io_8 = input_25;
assign io_8 = input_26;
assign io_8 = input_27;
assign io_8 = input_28;
assign io_8 = input_29;
assign io_8 = input_30;
assign io_8 = input_31;
assign io_8 = input_32;
assign io_8 = input_33;
assign io_8 = input_34;
assign io_8 = input_35;
assign io_8 = input_36;
assign io_8 = input_37;
assign io_8 = input_38;
assign io_8 = input_39;
assign io_8 = input_40;
assign io_8 = input_41;
assign io_8 = input_42;
assign io_8 = input_43;
assign io_8 = input_44;
assign io_8 = input_45;
assign io_8 = input_46;
assign io_8 = input_47;
assign io_8 = input_48;
assign io_8 = input_49;
assign io_8 = input_50;
assign io_8 = input_51;
assign io_8 = input_52;
assign io_8 = input_53;
assign io_8 = input_54;
assign io_8 = input_55;
assign io_8 = input_56;
assign io_8 = input_57;
assign io_8 = input_58;
assign io_8 = input_59;
assign io_8 = input_60;
assign io_8 = input_61;
assign io_8 = input_62;
assign io_8 = input_63;
assign io_9 = input_9;
assign io_9 = input_10;
assign io_9 = input_11;
assign io_9 = input_12;
assign io_9 = input_13;
assign io_9 = input_14;
assign io_9 = input_15;
assign io_9 = input_16;
assign io_9 = input_17;
assign io_9 = input_18;
assign io_9 = input_19;
assign io_9 = input_20;
assign io_9 = input_21;
assign io_9 = input_22;
assign io_9 = input_23;
assign io_9 = input_24;
assign io_9 = input_25;
assign io_9 = input_26;
assign io_9 = input_27;
assign io_9 = input_28;
assign io_9 = input_29;
assign io_9 = input_30;
assign io_9 = input_31;
assign io_9 = input_32;
assign io_9 = input_33;
assign io_9 = input_34;
assign io_9 = input_35;
assign io_9 = input_36;
assign io_9 = input_37;
assign io_9 = input_38;
assign io_9 = input_39;
assign io_9 = input_40;
assign io_9 = input_41;
assign io_9 = input_42;
assign io_9 = input_43;
assign io_9 = input_44;
assign io_9 = input_45;
assign io_9 = input_46;
assign io_9 = input_47;
assign io_9 = input_48;
assign io_9 = input_49;
assign io_9 = input_50;
assign io_9 = input_51;
assign io_9 = input_52;
assign io_9 = input_53;
assign io_9 = input_54;
assign io_9 = input_55;
assign io_9 = input_56;
assign io_9 = input_57;
assign io_9 = input_58;
assign io_9 = input_59;
assign io_9 = input_60;
assign io_9 = input_61;
assign io_9 = input_62;
assign io_9 = input_63;
assign io_10 = input_10;
assign io_10 = input_11;
assign io_10 = input_12;
assign io_10 = input_13;
assign io_10 = input_14;
assign io_10 = input_15;
assign io_10 = input_16;
assign io_10 = input_17;
assign io_10 = input_18;
assign io_10 = input_19;
assign io_10 = input_20;
assign io_10 = input_21;
assign io_10 = input_22;
assign io_10 = input_23;
assign io_10 = input_24;
assign io_10 = input_25;
assign io_10 = input_26;
assign io_10 = input_27;
assign io_10 = input_28;
assign io_10 = input_29;
assign io_10 = input_30;
assign io_10 = input_31;
assign io_10 = input_32;
assign io_10 = input_33;
assign io_10 = input_34;
assign io_10 = input_35;
assign io_10 = input_36;
assign io_10 = input_37;
assign io_10 = input_38;
assign io_10 = input_39;
assign io_10 = input_40;
assign io_10 = input_41;
assign io_10 = input_42;
assign io_10 = input_43;
assign io_10 = input_44;
assign io_10 = input_45;
assign io_10 = input_46;
assign io_10 = input_47;
assign io_10 = input_48;
assign io_10 = input_49;
assign io_10 = input_50;
assign io_10 = input_51;
assign io_10 = input_52;
assign io_10 = input_53;
assign io_10 = input_54;
assign io_10 = input_55;
assign io_10 = input_56;
assign io_10 = input_57;
assign io_10 = input_58;
assign io_10 = input_59;
assign io_10 = input_60;
assign io_10 = input_61;
assign io_10 = input_62;
assign io_10 = input_63;
assign io_11 = input_11;
assign io_11 = input_12;
assign io_11 = input_13;
assign io_11 = input_14;
assign io_11 = input_15;
assign io_11 = input_16;
assign io_11 = input_17;
assign io_11 = input_18;
assign io_11 = input_19;
assign io_11 = input_20;
assign io_11 = input_21;
assign io_11 = input_22;
assign io_11 = input_23;
assign io_11 = input_24;
assign io_11 = input_25;
assign io_11 = input_26;
assign io_11 = input_27;
assign io_11 = input_28;
assign io_11 = input_29;
assign io_11 = input_30;
assign io_11 = input_31;
assign io_11 = input_32;
assign io_11 = input_33;
assign io_11 = input_34;
assign io_11 = input_35;
assign io_11 = input_36;
assign io_11 = input_37;
assign io_11 = input_38;
assign io_11 = input_39;
assign io_11 = input_40;
assign io_11 = input_41;
assign io_11 = input_42;
assign io_11 = input_43;
assign io_11 = input_44;
assign io_11 = input_45;
assign io_11 = input_46;
assign io_11 = input_47;
assign io_11 = input_48;
assign io_11 = input_49;
assign io_11 = input_50;
assign io_11 = input_51;
assign io_11 = input_52;
assign io_11 = input_53;
assign io_11 = input_54;
assign io_11 = input_55;
assign io_11 = input_56;
assign io_11 = input_57;
assign io_11 = input_58;
assign io_11 = input_59;
assign io_11 = input_60;
assign io_11 = input_61;
assign io_11 = input_62;
assign io_11 = input_63;
assign io_12 = input_12;
assign io_12 = input_13;
assign io_12 = input_14;
assign io_12 = input_15;
assign io_12 = input_16;
assign io_12 = input_17;
assign io_12 = input_18;
assign io_12 = input_19;
assign io_12 = input_20;
assign io_12 = input_21;
assign io_12 = input_22;
assign io_12 = input_23;
assign io_12 = input_24;
assign io_12 = input_25;
assign io_12 = input_26;
assign io_12 = input_27;
assign io_12 = input_28;
assign io_12 = input_29;
assign io_12 = input_30;
assign io_12 = input_31;
assign io_12 = input_32;
assign io_12 = input_33;
assign io_12 = input_34;
assign io_12 = input_35;
assign io_12 = input_36;
assign io_12 = input_37;
assign io_12 = input_38;
assign io_12 = input_39;
assign io_12 = input_40;
assign io_12 = input_41;
assign io_12 = input_42;
assign io_12 = input_43;
assign io_12 = input_44;
assign io_12 = input_45;
assign io_12 = input_46;
assign io_12 = input_47;
assign io_12 = input_48;
assign io_12 = input_49;
assign io_12 = input_50;
assign io_12 = input_51;
assign io_12 = input_52;
assign io_12 = input_53;
assign io_12 = input_54;
assign io_12 = input_55;
assign io_12 = input_56;
assign io_12 = input_57;
assign io_12 = input_58;
assign io_12 = input_59;
assign io_12 = input_60;
assign io_12 = input_61;
assign io_12 = input_62;
assign io_12 = input_63;
assign io_13 = input_13;
assign io_13 = input_14;
assign io_13 = input_15;
assign io_13 = input_16;
assign io_13 = input_17;
assign io_13 = input_18;
assign io_13 = input_19;
assign io_13 = input_20;
assign io_13 = input_21;
assign io_13 = input_22;
assign io_13 = input_23;
assign io_13 = input_24;
assign io_13 = input_25;
assign io_13 = input_26;
assign io_13 = input_27;
assign io_13 = input_28;
assign io_13 = input_29;
assign io_13 = input_30;
assign io_13 = input_31;
assign io_13 = input_32;
assign io_13 = input_33;
assign io_13 = input_34;
assign io_13 = input_35;
assign io_13 = input_36;
assign io_13 = input_37;
assign io_13 = input_38;
assign io_13 = input_39;
assign io_13 = input_40;
assign io_13 = input_41;
assign io_13 = input_42;
assign io_13 = input_43;
assign io_13 = input_44;
assign io_13 = input_45;
assign io_13 = input_46;
assign io_13 = input_47;
assign io_13 = input_48;
assign io_13 = input_49;
assign io_13 = input_50;
assign io_13 = input_51;
assign io_13 = input_52;
assign io_13 = input_53;
assign io_13 = input_54;
assign io_13 = input_55;
assign io_13 = input_56;
assign io_13 = input_57;
assign io_13 = input_58;
assign io_13 = input_59;
assign io_13 = input_60;
assign io_13 = input_61;
assign io_13 = input_62;
assign io_13 = input_63;
assign io_14 = input_14;
assign io_14 = input_15;
assign io_14 = input_16;
assign io_14 = input_17;
assign io_14 = input_18;
assign io_14 = input_19;
assign io_14 = input_20;
assign io_14 = input_21;
assign io_14 = input_22;
assign io_14 = input_23;
assign io_14 = input_24;
assign io_14 = input_25;
assign io_14 = input_26;
assign io_14 = input_27;
assign io_14 = input_28;
assign io_14 = input_29;
assign io_14 = input_30;
assign io_14 = input_31;
assign io_14 = input_32;
assign io_14 = input_33;
assign io_14 = input_34;
assign io_14 = input_35;
assign io_14 = input_36;
assign io_14 = input_37;
assign io_14 = input_38;
assign io_14 = input_39;
assign io_14 = input_40;
assign io_14 = input_41;
assign io_14 = input_42;
assign io_14 = input_43;
assign io_14 = input_44;
assign io_14 = input_45;
assign io_14 = input_46;
assign io_14 = input_47;
assign io_14 = input_48;
assign io_14 = input_49;
assign io_14 = input_50;
assign io_14 = input_51;
assign io_14 = input_52;
assign io_14 = input_53;
assign io_14 = input_54;
assign io_14 = input_55;
assign io_14 = input_56;
assign io_14 = input_57;
assign io_14 = input_58;
assign io_14 = input_59;
assign io_14 = input_60;
assign io_14 = input_61;
assign io_14 = input_62;
assign io_14 = input_63;
assign io_15 = input_15;
assign io_15 = input_16;
assign io_15 = input_17;
assign io_15 = input_18;
assign io_15 = input_19;
assign io_15 = input_20;
assign io_15 = input_21;
assign io_15 = input_22;
assign io_15 = input_23;
assign io_15 = input_24;
assign io_15 = input_25;
assign io_15 = input_26;
assign io_15 = input_27;
assign io_15 = input_28;
assign io_15 = input_29;
assign io_15 = input_30;
assign io_15 = input_31;
assign io_15 = input_32;
assign io_15 = input_33;
assign io_15 = input_34;
assign io_15 = input_35;
assign io_15 = input_36;
assign io_15 = input_37;
assign io_15 = input_38;
assign io_15 = input_39;
assign io_15 = input_40;
assign io_15 = input_41;
assign io_15 = input_42;
assign io_15 = input_43;
assign io_15 = input_44;
assign io_15 = input_45;
assign io_15 = input_46;
assign io_15 = input_47;
assign io_15 = input_48;
assign io_15 = input_49;
assign io_15 = input_50;
assign io_15 = input_51;
assign io_15 = input_52;
assign io_15 = input_53;
assign io_15 = input_54;
assign io_15 = input_55;
assign io_15 = input_56;
assign io_15 = input_57;
assign io_15 = input_58;
assign io_15 = input_59;
assign io_15 = input_60;
assign io_15 = input_61;
assign io_15 = input_62;
assign io_15 = input_63;
assign io_16 = input_16;
assign io_16 = input_17;
assign io_16 = input_18;
assign io_16 = input_19;
assign io_16 = input_20;
assign io_16 = input_21;
assign io_16 = input_22;
assign io_16 = input_23;
assign io_16 = input_24;
assign io_16 = input_25;
assign io_16 = input_26;
assign io_16 = input_27;
assign io_16 = input_28;
assign io_16 = input_29;
assign io_16 = input_30;
assign io_16 = input_31;
assign io_16 = input_32;
assign io_16 = input_33;
assign io_16 = input_34;
assign io_16 = input_35;
assign io_16 = input_36;
assign io_16 = input_37;
assign io_16 = input_38;
assign io_16 = input_39;
assign io_16 = input_40;
assign io_16 = input_41;
assign io_16 = input_42;
assign io_16 = input_43;
assign io_16 = input_44;
assign io_16 = input_45;
assign io_16 = input_46;
assign io_16 = input_47;
assign io_16 = input_48;
assign io_16 = input_49;
assign io_16 = input_50;
assign io_16 = input_51;
assign io_16 = input_52;
assign io_16 = input_53;
assign io_16 = input_54;
assign io_16 = input_55;
assign io_16 = input_56;
assign io_16 = input_57;
assign io_16 = input_58;
assign io_16 = input_59;
assign io_16 = input_60;
assign io_16 = input_61;
assign io_16 = input_62;
assign io_16 = input_63;
assign io_17 = input_17;
assign io_17 = input_18;
assign io_17 = input_19;
assign io_17 = input_20;
assign io_17 = input_21;
assign io_17 = input_22;
assign io_17 = input_23;
assign io_17 = input_24;
assign io_17 = input_25;
assign io_17 = input_26;
assign io_17 = input_27;
assign io_17 = input_28;
assign io_17 = input_29;
assign io_17 = input_30;
assign io_17 = input_31;
assign io_17 = input_32;
assign io_17 = input_33;
assign io_17 = input_34;
assign io_17 = input_35;
assign io_17 = input_36;
assign io_17 = input_37;
assign io_17 = input_38;
assign io_17 = input_39;
assign io_17 = input_40;
assign io_17 = input_41;
assign io_17 = input_42;
assign io_17 = input_43;
assign io_17 = input_44;
assign io_17 = input_45;
assign io_17 = input_46;
assign io_17 = input_47;
assign io_17 = input_48;
assign io_17 = input_49;
assign io_17 = input_50;
assign io_17 = input_51;
assign io_17 = input_52;
assign io_17 = input_53;
assign io_17 = input_54;
assign io_17 = input_55;
assign io_17 = input_56;
assign io_17 = input_57;
assign io_17 = input_58;
assign io_17 = input_59;
assign io_17 = input_60;
assign io_17 = input_61;
assign io_17 = input_62;
assign io_17 = input_63;
assign io_18 = input_18;
assign io_18 = input_19;
assign io_18 = input_20;
assign io_18 = input_21;
assign io_18 = input_22;
assign io_18 = input_23;
assign io_18 = input_24;
assign io_18 = input_25;
assign io_18 = input_26;
assign io_18 = input_27;
assign io_18 = input_28;
assign io_18 = input_29;
assign io_18 = input_30;
assign io_18 = input_31;
assign io_18 = input_32;
assign io_18 = input_33;
assign io_18 = input_34;
assign io_18 = input_35;
assign io_18 = input_36;
assign io_18 = input_37;
assign io_18 = input_38;
assign io_18 = input_39;
assign io_18 = input_40;
assign io_18 = input_41;
assign io_18 = input_42;
assign io_18 = input_43;
assign io_18 = input_44;
assign io_18 = input_45;
assign io_18 = input_46;
assign io_18 = input_47;
assign io_18 = input_48;
assign io_18 = input_49;
assign io_18 = input_50;
assign io_18 = input_51;
assign io_18 = input_52;
assign io_18 = input_53;
assign io_18 = input_54;
assign io_18 = input_55;
assign io_18 = input_56;
assign io_18 = input_57;
assign io_18 = input_58;
assign io_18 = input_59;
assign io_18 = input_60;
assign io_18 = input_61;
assign io_18 = input_62;
assign io_18 = input_63;
assign io_19 = input_19;
assign io_19 = input_20;
assign io_19 = input_21;
assign io_19 = input_22;
assign io_19 = input_23;
assign io_19 = input_24;
assign io_19 = input_25;
assign io_19 = input_26;
assign io_19 = input_27;
assign io_19 = input_28;
assign io_19 = input_29;
assign io_19 = input_30;
assign io_19 = input_31;
assign io_19 = input_32;
assign io_19 = input_33;
assign io_19 = input_34;
assign io_19 = input_35;
assign io_19 = input_36;
assign io_19 = input_37;
assign io_19 = input_38;
assign io_19 = input_39;
assign io_19 = input_40;
assign io_19 = input_41;
assign io_19 = input_42;
assign io_19 = input_43;
assign io_19 = input_44;
assign io_19 = input_45;
assign io_19 = input_46;
assign io_19 = input_47;
assign io_19 = input_48;
assign io_19 = input_49;
assign io_19 = input_50;
assign io_19 = input_51;
assign io_19 = input_52;
assign io_19 = input_53;
assign io_19 = input_54;
assign io_19 = input_55;
assign io_19 = input_56;
assign io_19 = input_57;
assign io_19 = input_58;
assign io_19 = input_59;
assign io_19 = input_60;
assign io_19 = input_61;
assign io_19 = input_62;
assign io_19 = input_63;
assign io_20 = input_20;
assign io_20 = input_21;
assign io_20 = input_22;
assign io_20 = input_23;
assign io_20 = input_24;
assign io_20 = input_25;
assign io_20 = input_26;
assign io_20 = input_27;
assign io_20 = input_28;
assign io_20 = input_29;
assign io_20 = input_30;
assign io_20 = input_31;
assign io_20 = input_32;
assign io_20 = input_33;
assign io_20 = input_34;
assign io_20 = input_35;
assign io_20 = input_36;
assign io_20 = input_37;
assign io_20 = input_38;
assign io_20 = input_39;
assign io_20 = input_40;
assign io_20 = input_41;
assign io_20 = input_42;
assign io_20 = input_43;
assign io_20 = input_44;
assign io_20 = input_45;
assign io_20 = input_46;
assign io_20 = input_47;
assign io_20 = input_48;
assign io_20 = input_49;
assign io_20 = input_50;
assign io_20 = input_51;
assign io_20 = input_52;
assign io_20 = input_53;
assign io_20 = input_54;
assign io_20 = input_55;
assign io_20 = input_56;
assign io_20 = input_57;
assign io_20 = input_58;
assign io_20 = input_59;
assign io_20 = input_60;
assign io_20 = input_61;
assign io_20 = input_62;
assign io_20 = input_63;
assign io_21 = input_21;
assign io_21 = input_22;
assign io_21 = input_23;
assign io_21 = input_24;
assign io_21 = input_25;
assign io_21 = input_26;
assign io_21 = input_27;
assign io_21 = input_28;
assign io_21 = input_29;
assign io_21 = input_30;
assign io_21 = input_31;
assign io_21 = input_32;
assign io_21 = input_33;
assign io_21 = input_34;
assign io_21 = input_35;
assign io_21 = input_36;
assign io_21 = input_37;
assign io_21 = input_38;
assign io_21 = input_39;
assign io_21 = input_40;
assign io_21 = input_41;
assign io_21 = input_42;
assign io_21 = input_43;
assign io_21 = input_44;
assign io_21 = input_45;
assign io_21 = input_46;
assign io_21 = input_47;
assign io_21 = input_48;
assign io_21 = input_49;
assign io_21 = input_50;
assign io_21 = input_51;
assign io_21 = input_52;
assign io_21 = input_53;
assign io_21 = input_54;
assign io_21 = input_55;
assign io_21 = input_56;
assign io_21 = input_57;
assign io_21 = input_58;
assign io_21 = input_59;
assign io_21 = input_60;
assign io_21 = input_61;
assign io_21 = input_62;
assign io_21 = input_63;
assign io_22 = input_22;
assign io_22 = input_23;
assign io_22 = input_24;
assign io_22 = input_25;
assign io_22 = input_26;
assign io_22 = input_27;
assign io_22 = input_28;
assign io_22 = input_29;
assign io_22 = input_30;
assign io_22 = input_31;
assign io_22 = input_32;
assign io_22 = input_33;
assign io_22 = input_34;
assign io_22 = input_35;
assign io_22 = input_36;
assign io_22 = input_37;
assign io_22 = input_38;
assign io_22 = input_39;
assign io_22 = input_40;
assign io_22 = input_41;
assign io_22 = input_42;
assign io_22 = input_43;
assign io_22 = input_44;
assign io_22 = input_45;
assign io_22 = input_46;
assign io_22 = input_47;
assign io_22 = input_48;
assign io_22 = input_49;
assign io_22 = input_50;
assign io_22 = input_51;
assign io_22 = input_52;
assign io_22 = input_53;
assign io_22 = input_54;
assign io_22 = input_55;
assign io_22 = input_56;
assign io_22 = input_57;
assign io_22 = input_58;
assign io_22 = input_59;
assign io_22 = input_60;
assign io_22 = input_61;
assign io_22 = input_62;
assign io_22 = input_63;
assign io_23 = input_23;
assign io_23 = input_24;
assign io_23 = input_25;
assign io_23 = input_26;
assign io_23 = input_27;
assign io_23 = input_28;
assign io_23 = input_29;
assign io_23 = input_30;
assign io_23 = input_31;
assign io_23 = input_32;
assign io_23 = input_33;
assign io_23 = input_34;
assign io_23 = input_35;
assign io_23 = input_36;
assign io_23 = input_37;
assign io_23 = input_38;
assign io_23 = input_39;
assign io_23 = input_40;
assign io_23 = input_41;
assign io_23 = input_42;
assign io_23 = input_43;
assign io_23 = input_44;
assign io_23 = input_45;
assign io_23 = input_46;
assign io_23 = input_47;
assign io_23 = input_48;
assign io_23 = input_49;
assign io_23 = input_50;
assign io_23 = input_51;
assign io_23 = input_52;
assign io_23 = input_53;
assign io_23 = input_54;
assign io_23 = input_55;
assign io_23 = input_56;
assign io_23 = input_57;
assign io_23 = input_58;
assign io_23 = input_59;
assign io_23 = input_60;
assign io_23 = input_61;
assign io_23 = input_62;
assign io_23 = input_63;
assign io_24 = input_24;
assign io_24 = input_25;
assign io_24 = input_26;
assign io_24 = input_27;
assign io_24 = input_28;
assign io_24 = input_29;
assign io_24 = input_30;
assign io_24 = input_31;
assign io_24 = input_32;
assign io_24 = input_33;
assign io_24 = input_34;
assign io_24 = input_35;
assign io_24 = input_36;
assign io_24 = input_37;
assign io_24 = input_38;
assign io_24 = input_39;
assign io_24 = input_40;
assign io_24 = input_41;
assign io_24 = input_42;
assign io_24 = input_43;
assign io_24 = input_44;
assign io_24 = input_45;
assign io_24 = input_46;
assign io_24 = input_47;
assign io_24 = input_48;
assign io_24 = input_49;
assign io_24 = input_50;
assign io_24 = input_51;
assign io_24 = input_52;
assign io_24 = input_53;
assign io_24 = input_54;
assign io_24 = input_55;
assign io_24 = input_56;
assign io_24 = input_57;
assign io_24 = input_58;
assign io_24 = input_59;
assign io_24 = input_60;
assign io_24 = input_61;
assign io_24 = input_62;
assign io_24 = input_63;
assign io_25 = input_25;
assign io_25 = input_26;
assign io_25 = input_27;
assign io_25 = input_28;
assign io_25 = input_29;
assign io_25 = input_30;
assign io_25 = input_31;
assign io_25 = input_32;
assign io_25 = input_33;
assign io_25 = input_34;
assign io_25 = input_35;
assign io_25 = input_36;
assign io_25 = input_37;
assign io_25 = input_38;
assign io_25 = input_39;
assign io_25 = input_40;
assign io_25 = input_41;
assign io_25 = input_42;
assign io_25 = input_43;
assign io_25 = input_44;
assign io_25 = input_45;
assign io_25 = input_46;
assign io_25 = input_47;
assign io_25 = input_48;
assign io_25 = input_49;
assign io_25 = input_50;
assign io_25 = input_51;
assign io_25 = input_52;
assign io_25 = input_53;
assign io_25 = input_54;
assign io_25 = input_55;
assign io_25 = input_56;
assign io_25 = input_57;
assign io_25 = input_58;
assign io_25 = input_59;
assign io_25 = input_60;
assign io_25 = input_61;
assign io_25 = input_62;
assign io_25 = input_63;
assign io_26 = input_26;
assign io_26 = input_27;
assign io_26 = input_28;
assign io_26 = input_29;
assign io_26 = input_30;
assign io_26 = input_31;
assign io_26 = input_32;
assign io_26 = input_33;
assign io_26 = input_34;
assign io_26 = input_35;
assign io_26 = input_36;
assign io_26 = input_37;
assign io_26 = input_38;
assign io_26 = input_39;
assign io_26 = input_40;
assign io_26 = input_41;
assign io_26 = input_42;
assign io_26 = input_43;
assign io_26 = input_44;
assign io_26 = input_45;
assign io_26 = input_46;
assign io_26 = input_47;
assign io_26 = input_48;
assign io_26 = input_49;
assign io_26 = input_50;
assign io_26 = input_51;
assign io_26 = input_52;
assign io_26 = input_53;
assign io_26 = input_54;
assign io_26 = input_55;
assign io_26 = input_56;
assign io_26 = input_57;
assign io_26 = input_58;
assign io_26 = input_59;
assign io_26 = input_60;
assign io_26 = input_61;
assign io_26 = input_62;
assign io_26 = input_63;
assign io_27 = input_27;
assign io_27 = input_28;
assign io_27 = input_29;
assign io_27 = input_30;
assign io_27 = input_31;
assign io_27 = input_32;
assign io_27 = input_33;
assign io_27 = input_34;
assign io_27 = input_35;
assign io_27 = input_36;
assign io_27 = input_37;
assign io_27 = input_38;
assign io_27 = input_39;
assign io_27 = input_40;
assign io_27 = input_41;
assign io_27 = input_42;
assign io_27 = input_43;
assign io_27 = input_44;
assign io_27 = input_45;
assign io_27 = input_46;
assign io_27 = input_47;
assign io_27 = input_48;
assign io_27 = input_49;
assign io_27 = input_50;
assign io_27 = input_51;
assign io_27 = input_52;
assign io_27 = input_53;
assign io_27 = input_54;
assign io_27 = input_55;
assign io_27 = input_56;
assign io_27 = input_57;
assign io_27 = input_58;
assign io_27 = input_59;
assign io_27 = input_60;
assign io_27 = input_61;
assign io_27 = input_62;
assign io_27 = input_63;
assign io_28 = input_28;
assign io_28 = input_29;
assign io_28 = input_30;
assign io_28 = input_31;
assign io_28 = input_32;
assign io_28 = input_33;
assign io_28 = input_34;
assign io_28 = input_35;
assign io_28 = input_36;
assign io_28 = input_37;
assign io_28 = input_38;
assign io_28 = input_39;
assign io_28 = input_40;
assign io_28 = input_41;
assign io_28 = input_42;
assign io_28 = input_43;
assign io_28 = input_44;
assign io_28 = input_45;
assign io_28 = input_46;
assign io_28 = input_47;
assign io_28 = input_48;
assign io_28 = input_49;
assign io_28 = input_50;
assign io_28 = input_51;
assign io_28 = input_52;
assign io_28 = input_53;
assign io_28 = input_54;
assign io_28 = input_55;
assign io_28 = input_56;
assign io_28 = input_57;
assign io_28 = input_58;
assign io_28 = input_59;
assign io_28 = input_60;
assign io_28 = input_61;
assign io_28 = input_62;
assign io_28 = input_63;
assign io_29 = input_29;
assign io_29 = input_30;
assign io_29 = input_31;
assign io_29 = input_32;
assign io_29 = input_33;
assign io_29 = input_34;
assign io_29 = input_35;
assign io_29 = input_36;
assign io_29 = input_37;
assign io_29 = input_38;
assign io_29 = input_39;
assign io_29 = input_40;
assign io_29 = input_41;
assign io_29 = input_42;
assign io_29 = input_43;
assign io_29 = input_44;
assign io_29 = input_45;
assign io_29 = input_46;
assign io_29 = input_47;
assign io_29 = input_48;
assign io_29 = input_49;
assign io_29 = input_50;
assign io_29 = input_51;
assign io_29 = input_52;
assign io_29 = input_53;
assign io_29 = input_54;
assign io_29 = input_55;
assign io_29 = input_56;
assign io_29 = input_57;
assign io_29 = input_58;
assign io_29 = input_59;
assign io_29 = input_60;
assign io_29 = input_61;
assign io_29 = input_62;
assign io_29 = input_63;
assign io_30 = input_30;
assign io_30 = input_31;
assign io_30 = input_32;
assign io_30 = input_33;
assign io_30 = input_34;
assign io_30 = input_35;
assign io_30 = input_36;
assign io_30 = input_37;
assign io_30 = input_38;
assign io_30 = input_39;
assign io_30 = input_40;
assign io_30 = input_41;
assign io_30 = input_42;
assign io_30 = input_43;
assign io_30 = input_44;
assign io_30 = input_45;
assign io_30 = input_46;
assign io_30 = input_47;
assign io_30 = input_48;
assign io_30 = input_49;
assign io_30 = input_50;
assign io_30 = input_51;
assign io_30 = input_52;
assign io_30 = input_53;
assign io_30 = input_54;
assign io_30 = input_55;
assign io_30 = input_56;
assign io_30 = input_57;
assign io_30 = input_58;
assign io_30 = input_59;
assign io_30 = input_60;
assign io_30 = input_61;
assign io_30 = input_62;
assign io_30 = input_63;
assign io_31 = input_31;
assign io_31 = input_32;
assign io_31 = input_33;
assign io_31 = input_34;
assign io_31 = input_35;
assign io_31 = input_36;
assign io_31 = input_37;
assign io_31 = input_38;
assign io_31 = input_39;
assign io_31 = input_40;
assign io_31 = input_41;
assign io_31 = input_42;
assign io_31 = input_43;
assign io_31 = input_44;
assign io_31 = input_45;
assign io_31 = input_46;
assign io_31 = input_47;
assign io_31 = input_48;
assign io_31 = input_49;
assign io_31 = input_50;
assign io_31 = input_51;
assign io_31 = input_52;
assign io_31 = input_53;
assign io_31 = input_54;
assign io_31 = input_55;
assign io_31 = input_56;
assign io_31 = input_57;
assign io_31 = input_58;
assign io_31 = input_59;
assign io_31 = input_60;
assign io_31 = input_61;
assign io_31 = input_62;
assign io_31 = input_63;
assign io_32 = input_32;
assign io_32 = input_33;
assign io_32 = input_34;
assign io_32 = input_35;
assign io_32 = input_36;
assign io_32 = input_37;
assign io_32 = input_38;
assign io_32 = input_39;
assign io_32 = input_40;
assign io_32 = input_41;
assign io_32 = input_42;
assign io_32 = input_43;
assign io_32 = input_44;
assign io_32 = input_45;
assign io_32 = input_46;
assign io_32 = input_47;
assign io_32 = input_48;
assign io_32 = input_49;
assign io_32 = input_50;
assign io_32 = input_51;
assign io_32 = input_52;
assign io_32 = input_53;
assign io_32 = input_54;
assign io_32 = input_55;
assign io_32 = input_56;
assign io_32 = input_57;
assign io_32 = input_58;
assign io_32 = input_59;
assign io_32 = input_60;
assign io_32 = input_61;
assign io_32 = input_62;
assign io_32 = input_63;
assign io_33 = input_33;
assign io_33 = input_34;
assign io_33 = input_35;
assign io_33 = input_36;
assign io_33 = input_37;
assign io_33 = input_38;
assign io_33 = input_39;
assign io_33 = input_40;
assign io_33 = input_41;
assign io_33 = input_42;
assign io_33 = input_43;
assign io_33 = input_44;
assign io_33 = input_45;
assign io_33 = input_46;
assign io_33 = input_47;
assign io_33 = input_48;
assign io_33 = input_49;
assign io_33 = input_50;
assign io_33 = input_51;
assign io_33 = input_52;
assign io_33 = input_53;
assign io_33 = input_54;
assign io_33 = input_55;
assign io_33 = input_56;
assign io_33 = input_57;
assign io_33 = input_58;
assign io_33 = input_59;
assign io_33 = input_60;
assign io_33 = input_61;
assign io_33 = input_62;
assign io_33 = input_63;
assign io_34 = input_34;
assign io_34 = input_35;
assign io_34 = input_36;
assign io_34 = input_37;
assign io_34 = input_38;
assign io_34 = input_39;
assign io_34 = input_40;
assign io_34 = input_41;
assign io_34 = input_42;
assign io_34 = input_43;
assign io_34 = input_44;
assign io_34 = input_45;
assign io_34 = input_46;
assign io_34 = input_47;
assign io_34 = input_48;
assign io_34 = input_49;
assign io_34 = input_50;
assign io_34 = input_51;
assign io_34 = input_52;
assign io_34 = input_53;
assign io_34 = input_54;
assign io_34 = input_55;
assign io_34 = input_56;
assign io_34 = input_57;
assign io_34 = input_58;
assign io_34 = input_59;
assign io_34 = input_60;
assign io_34 = input_61;
assign io_34 = input_62;
assign io_34 = input_63;
assign io_35 = input_35;
assign io_35 = input_36;
assign io_35 = input_37;
assign io_35 = input_38;
assign io_35 = input_39;
assign io_35 = input_40;
assign io_35 = input_41;
assign io_35 = input_42;
assign io_35 = input_43;
assign io_35 = input_44;
assign io_35 = input_45;
assign io_35 = input_46;
assign io_35 = input_47;
assign io_35 = input_48;
assign io_35 = input_49;
assign io_35 = input_50;
assign io_35 = input_51;
assign io_35 = input_52;
assign io_35 = input_53;
assign io_35 = input_54;
assign io_35 = input_55;
assign io_35 = input_56;
assign io_35 = input_57;
assign io_35 = input_58;
assign io_35 = input_59;
assign io_35 = input_60;
assign io_35 = input_61;
assign io_35 = input_62;
assign io_35 = input_63;
assign io_36 = input_36;
assign io_36 = input_37;
assign io_36 = input_38;
assign io_36 = input_39;
assign io_36 = input_40;
assign io_36 = input_41;
assign io_36 = input_42;
assign io_36 = input_43;
assign io_36 = input_44;
assign io_36 = input_45;
assign io_36 = input_46;
assign io_36 = input_47;
assign io_36 = input_48;
assign io_36 = input_49;
assign io_36 = input_50;
assign io_36 = input_51;
assign io_36 = input_52;
assign io_36 = input_53;
assign io_36 = input_54;
assign io_36 = input_55;
assign io_36 = input_56;
assign io_36 = input_57;
assign io_36 = input_58;
assign io_36 = input_59;
assign io_36 = input_60;
assign io_36 = input_61;
assign io_36 = input_62;
assign io_36 = input_63;
assign io_37 = input_37;
assign io_37 = input_38;
assign io_37 = input_39;
assign io_37 = input_40;
assign io_37 = input_41;
assign io_37 = input_42;
assign io_37 = input_43;
assign io_37 = input_44;
assign io_37 = input_45;
assign io_37 = input_46;
assign io_37 = input_47;
assign io_37 = input_48;
assign io_37 = input_49;
assign io_37 = input_50;
assign io_37 = input_51;
assign io_37 = input_52;
assign io_37 = input_53;
assign io_37 = input_54;
assign io_37 = input_55;
assign io_37 = input_56;
assign io_37 = input_57;
assign io_37 = input_58;
assign io_37 = input_59;
assign io_37 = input_60;
assign io_37 = input_61;
assign io_37 = input_62;
assign io_37 = input_63;
assign io_38 = input_38;
assign io_38 = input_39;
assign io_38 = input_40;
assign io_38 = input_41;
assign io_38 = input_42;
assign io_38 = input_43;
assign io_38 = input_44;
assign io_38 = input_45;
assign io_38 = input_46;
assign io_38 = input_47;
assign io_38 = input_48;
assign io_38 = input_49;
assign io_38 = input_50;
assign io_38 = input_51;
assign io_38 = input_52;
assign io_38 = input_53;
assign io_38 = input_54;
assign io_38 = input_55;
assign io_38 = input_56;
assign io_38 = input_57;
assign io_38 = input_58;
assign io_38 = input_59;
assign io_38 = input_60;
assign io_38 = input_61;
assign io_38 = input_62;
assign io_38 = input_63;
assign io_39 = input_39;
assign io_39 = input_40;
assign io_39 = input_41;
assign io_39 = input_42;
assign io_39 = input_43;
assign io_39 = input_44;
assign io_39 = input_45;
assign io_39 = input_46;
assign io_39 = input_47;
assign io_39 = input_48;
assign io_39 = input_49;
assign io_39 = input_50;
assign io_39 = input_51;
assign io_39 = input_52;
assign io_39 = input_53;
assign io_39 = input_54;
assign io_39 = input_55;
assign io_39 = input_56;
assign io_39 = input_57;
assign io_39 = input_58;
assign io_39 = input_59;
assign io_39 = input_60;
assign io_39 = input_61;
assign io_39 = input_62;
assign io_39 = input_63;
assign io_40 = input_40;
assign io_40 = input_41;
assign io_40 = input_42;
assign io_40 = input_43;
assign io_40 = input_44;
assign io_40 = input_45;
assign io_40 = input_46;
assign io_40 = input_47;
assign io_40 = input_48;
assign io_40 = input_49;
assign io_40 = input_50;
assign io_40 = input_51;
assign io_40 = input_52;
assign io_40 = input_53;
assign io_40 = input_54;
assign io_40 = input_55;
assign io_40 = input_56;
assign io_40 = input_57;
assign io_40 = input_58;
assign io_40 = input_59;
assign io_40 = input_60;
assign io_40 = input_61;
assign io_40 = input_62;
assign io_40 = input_63;
assign io_41 = input_41;
assign io_41 = input_42;
assign io_41 = input_43;
assign io_41 = input_44;
assign io_41 = input_45;
assign io_41 = input_46;
assign io_41 = input_47;
assign io_41 = input_48;
assign io_41 = input_49;
assign io_41 = input_50;
assign io_41 = input_51;
assign io_41 = input_52;
assign io_41 = input_53;
assign io_41 = input_54;
assign io_41 = input_55;
assign io_41 = input_56;
assign io_41 = input_57;
assign io_41 = input_58;
assign io_41 = input_59;
assign io_41 = input_60;
assign io_41 = input_61;
assign io_41 = input_62;
assign io_41 = input_63;
assign io_42 = input_42;
assign io_42 = input_43;
assign io_42 = input_44;
assign io_42 = input_45;
assign io_42 = input_46;
assign io_42 = input_47;
assign io_42 = input_48;
assign io_42 = input_49;
assign io_42 = input_50;
assign io_42 = input_51;
assign io_42 = input_52;
assign io_42 = input_53;
assign io_42 = input_54;
assign io_42 = input_55;
assign io_42 = input_56;
assign io_42 = input_57;
assign io_42 = input_58;
assign io_42 = input_59;
assign io_42 = input_60;
assign io_42 = input_61;
assign io_42 = input_62;
assign io_42 = input_63;
assign io_43 = input_43;
assign io_43 = input_44;
assign io_43 = input_45;
assign io_43 = input_46;
assign io_43 = input_47;
assign io_43 = input_48;
assign io_43 = input_49;
assign io_43 = input_50;
assign io_43 = input_51;
assign io_43 = input_52;
assign io_43 = input_53;
assign io_43 = input_54;
assign io_43 = input_55;
assign io_43 = input_56;
assign io_43 = input_57;
assign io_43 = input_58;
assign io_43 = input_59;
assign io_43 = input_60;
assign io_43 = input_61;
assign io_43 = input_62;
assign io_43 = input_63;
assign io_44 = input_44;
assign io_44 = input_45;
assign io_44 = input_46;
assign io_44 = input_47;
assign io_44 = input_48;
assign io_44 = input_49;
assign io_44 = input_50;
assign io_44 = input_51;
assign io_44 = input_52;
assign io_44 = input_53;
assign io_44 = input_54;
assign io_44 = input_55;
assign io_44 = input_56;
assign io_44 = input_57;
assign io_44 = input_58;
assign io_44 = input_59;
assign io_44 = input_60;
assign io_44 = input_61;
assign io_44 = input_62;
assign io_44 = input_63;
assign io_45 = input_45;
assign io_45 = input_46;
assign io_45 = input_47;
assign io_45 = input_48;
assign io_45 = input_49;
assign io_45 = input_50;
assign io_45 = input_51;
assign io_45 = input_52;
assign io_45 = input_53;
assign io_45 = input_54;
assign io_45 = input_55;
assign io_45 = input_56;
assign io_45 = input_57;
assign io_45 = input_58;
assign io_45 = input_59;
assign io_45 = input_60;
assign io_45 = input_61;
assign io_45 = input_62;
assign io_45 = input_63;
assign io_46 = input_46;
assign io_46 = input_47;
assign io_46 = input_48;
assign io_46 = input_49;
assign io_46 = input_50;
assign io_46 = input_51;
assign io_46 = input_52;
assign io_46 = input_53;
assign io_46 = input_54;
assign io_46 = input_55;
assign io_46 = input_56;
assign io_46 = input_57;
assign io_46 = input_58;
assign io_46 = input_59;
assign io_46 = input_60;
assign io_46 = input_61;
assign io_46 = input_62;
assign io_46 = input_63;
assign io_47 = input_47;
assign io_47 = input_48;
assign io_47 = input_49;
assign io_47 = input_50;
assign io_47 = input_51;
assign io_47 = input_52;
assign io_47 = input_53;
assign io_47 = input_54;
assign io_47 = input_55;
assign io_47 = input_56;
assign io_47 = input_57;
assign io_47 = input_58;
assign io_47 = input_59;
assign io_47 = input_60;
assign io_47 = input_61;
assign io_47 = input_62;
assign io_47 = input_63;
assign io_48 = input_48;
assign io_48 = input_49;
assign io_48 = input_50;
assign io_48 = input_51;
assign io_48 = input_52;
assign io_48 = input_53;
assign io_48 = input_54;
assign io_48 = input_55;
assign io_48 = input_56;
assign io_48 = input_57;
assign io_48 = input_58;
assign io_48 = input_59;
assign io_48 = input_60;
assign io_48 = input_61;
assign io_48 = input_62;
assign io_48 = input_63;
assign io_49 = input_49;
assign io_49 = input_50;
assign io_49 = input_51;
assign io_49 = input_52;
assign io_49 = input_53;
assign io_49 = input_54;
assign io_49 = input_55;
assign io_49 = input_56;
assign io_49 = input_57;
assign io_49 = input_58;
assign io_49 = input_59;
assign io_49 = input_60;
assign io_49 = input_61;
assign io_49 = input_62;
assign io_49 = input_63;
assign io_50 = input_50;
assign io_50 = input_51;
assign io_50 = input_52;
assign io_50 = input_53;
assign io_50 = input_54;
assign io_50 = input_55;
assign io_50 = input_56;
assign io_50 = input_57;
assign io_50 = input_58;
assign io_50 = input_59;
assign io_50 = input_60;
assign io_50 = input_61;
assign io_50 = input_62;
assign io_50 = input_63;
assign io_51 = input_51;
assign io_51 = input_52;
assign io_51 = input_53;
assign io_51 = input_54;
assign io_51 = input_55;
assign io_51 = input_56;
assign io_51 = input_57;
assign io_51 = input_58;
assign io_51 = input_59;
assign io_51 = input_60;
assign io_51 = input_61;
assign io_51 = input_62;
assign io_51 = input_63;
assign io_52 = input_52;
assign io_52 = input_53;
assign io_52 = input_54;
assign io_52 = input_55;
assign io_52 = input_56;
assign io_52 = input_57;
assign io_52 = input_58;
assign io_52 = input_59;
assign io_52 = input_60;
assign io_52 = input_61;
assign io_52 = input_62;
assign io_52 = input_63;
assign io_53 = input_53;
assign io_53 = input_54;
assign io_53 = input_55;
assign io_53 = input_56;
assign io_53 = input_57;
assign io_53 = input_58;
assign io_53 = input_59;
assign io_53 = input_60;
assign io_53 = input_61;
assign io_53 = input_62;
assign io_53 = input_63;
assign io_54 = input_54;
assign io_54 = input_55;
assign io_54 = input_56;
assign io_54 = input_57;
assign io_54 = input_58;
assign io_54 = input_59;
assign io_54 = input_60;
assign io_54 = input_61;
assign io_54 = input_62;
assign io_54 = input_63;
assign io_55 = input_55;
assign io_55 = input_56;
assign io_55 = input_57;
assign io_55 = input_58;
assign io_55 = input_59;
assign io_55 = input_60;
assign io_55 = input_61;
assign io_55 = input_62;
assign io_55 = input_63;
assign io_56 = input_56;
assign io_56 = input_57;
assign io_56 = input_58;
assign io_56 = input_59;
assign io_56 = input_60;
assign io_56 = input_61;
assign io_56 = input_62;
assign io_56 = input_63;
assign io_57 = input_57;
assign io_57 = input_58;
assign io_57 = input_59;
assign io_57 = input_60;
assign io_57 = input_61;
assign io_57 = input_62;
assign io_57 = input_63;
assign io_58 = input_58;
assign io_58 = input_59;
assign io_58 = input_60;
assign io_58 = input_61;
assign io_58 = input_62;
assign io_58 = input_63;
assign io_59 = input_59;
assign io_59 = input_60;
assign io_59 = input_61;
assign io_59 = input_62;
assign io_59 = input_63;
assign io_60 = input_60;
assign io_60 = input_61;
assign io_60 = input_62;
assign io_60 = input_63;
assign io_61 = input_61;
assign io_61 = input_62;
assign io_61 = input_63;
assign io_62 = input_62;
assign io_62 = input_63;
assign io_63 = input_63;
endmodule
