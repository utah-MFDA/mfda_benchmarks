module fanout2_braid_3_32 (
output output_0,output output_1,output output_2,input input_0,input input_1,input input_2
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_1_2, output_1_0, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_0), .y(output_0_2));
wire output_2_2, output_2_0, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_0), .y(output_1_2));
wire output_3_2, output_3_0, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_0), .y(output_2_2));
wire output_1_3, output_1_1, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_1), .y(output_0_3));
wire output_2_3, output_2_1, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_1), .y(output_1_3));
wire output_3_3, output_3_1, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_1), .y(output_2_3));
wire output_1_4, output_1_2, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_2), .y(output_0_4));
wire output_2_4, output_2_2, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_2), .y(output_1_4));
wire output_3_4, output_3_2, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_2), .y(output_2_4));
wire output_1_5, output_1_0, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_0), .y(output_0_5));
wire output_2_5, output_2_0, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_0), .y(output_1_5));
wire output_3_5, output_3_0, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_0), .y(output_2_5));
wire output_1_6, output_1_1, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_1), .y(output_0_6));
wire output_2_6, output_2_1, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_1), .y(output_1_6));
wire output_3_6, output_3_1, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_1), .y(output_2_6));
wire output_1_7, output_1_2, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_2), .y(output_0_7));
wire output_2_7, output_2_2, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_2), .y(output_1_7));
wire output_3_7, output_3_2, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_2), .y(output_2_7));
wire output_1_8, output_1_0, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_0), .y(output_0_8));
wire output_2_8, output_2_0, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_0), .y(output_1_8));
wire output_3_8, output_3_0, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_0), .y(output_2_8));
wire output_1_9, output_1_1, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_1), .y(output_0_9));
wire output_2_9, output_2_1, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_1), .y(output_1_9));
wire output_3_9, output_3_1, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_1), .y(output_2_9));
wire output_1_10, output_1_2, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_2), .y(output_0_10));
wire output_2_10, output_2_2, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_2), .y(output_1_10));
wire output_3_10, output_3_2, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_2), .y(output_2_10));
wire output_1_11, output_1_0, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_0), .y(output_0_11));
wire output_2_11, output_2_0, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_0), .y(output_1_11));
wire output_3_11, output_3_0, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_0), .y(output_2_11));
wire output_1_12, output_1_1, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_1), .y(output_0_12));
wire output_2_12, output_2_1, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_1), .y(output_1_12));
wire output_3_12, output_3_1, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_1), .y(output_2_12));
wire output_1_13, output_1_2, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_2), .y(output_0_13));
wire output_2_13, output_2_2, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_2), .y(output_1_13));
wire output_3_13, output_3_2, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_2), .y(output_2_13));
wire output_1_14, output_1_0, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_0), .y(output_0_14));
wire output_2_14, output_2_0, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_0), .y(output_1_14));
wire output_3_14, output_3_0, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_0), .y(output_2_14));
wire output_1_15, output_1_1, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_1), .y(output_0_15));
wire output_2_15, output_2_1, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_1), .y(output_1_15));
wire output_3_15, output_3_1, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_1), .y(output_2_15));
wire output_1_16, output_1_2, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_2), .y(output_0_16));
wire output_2_16, output_2_2, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_2), .y(output_1_16));
wire output_3_16, output_3_2, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_2), .y(output_2_16));
wire output_1_17, output_1_0, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_0), .y(output_0_17));
wire output_2_17, output_2_0, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_0), .y(output_1_17));
wire output_3_17, output_3_0, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_0), .y(output_2_17));
wire output_1_18, output_1_1, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_1), .y(output_0_18));
wire output_2_18, output_2_1, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_1), .y(output_1_18));
wire output_3_18, output_3_1, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_1), .y(output_2_18));
wire output_1_19, output_1_2, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_2), .y(output_0_19));
wire output_2_19, output_2_2, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_2), .y(output_1_19));
wire output_3_19, output_3_2, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_2), .y(output_2_19));
wire output_1_20, output_1_0, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_0), .y(output_0_20));
wire output_2_20, output_2_0, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_0), .y(output_1_20));
wire output_3_20, output_3_0, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_0), .y(output_2_20));
wire output_1_21, output_1_1, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_1), .y(output_0_21));
wire output_2_21, output_2_1, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_1), .y(output_1_21));
wire output_3_21, output_3_1, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_1), .y(output_2_21));
wire output_1_22, output_1_2, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_2), .y(output_0_22));
wire output_2_22, output_2_2, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_2), .y(output_1_22));
wire output_3_22, output_3_2, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_2), .y(output_2_22));
wire output_1_23, output_1_0, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_0), .y(output_0_23));
wire output_2_23, output_2_0, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_0), .y(output_1_23));
wire output_3_23, output_3_0, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_0), .y(output_2_23));
wire output_1_24, output_1_1, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_1), .y(output_0_24));
wire output_2_24, output_2_1, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_1), .y(output_1_24));
wire output_3_24, output_3_1, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_1), .y(output_2_24));
wire output_1_25, output_1_2, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_2), .y(output_0_25));
wire output_2_25, output_2_2, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_2), .y(output_1_25));
wire output_3_25, output_3_2, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_2), .y(output_2_25));
wire output_1_26, output_1_0, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_0), .y(output_0_26));
wire output_2_26, output_2_0, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_0), .y(output_1_26));
wire output_3_26, output_3_0, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_0), .y(output_2_26));
wire output_1_27, output_1_1, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_1), .y(output_0_27));
wire output_2_27, output_2_1, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_1), .y(output_1_27));
wire output_3_27, output_3_1, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_1), .y(output_2_27));
wire output_1_28, output_1_2, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_2), .y(output_0_28));
wire output_2_28, output_2_2, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_2), .y(output_1_28));
wire output_3_28, output_3_2, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_2), .y(output_2_28));
wire output_1_29, output_1_0, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_0), .y(output_0_29));
wire output_2_29, output_2_0, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_0), .y(output_1_29));
wire output_3_29, output_3_0, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_0), .y(output_2_29));
wire output_1_30, output_1_1, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_1), .y(output_0_30));
wire output_2_30, output_2_1, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_1), .y(output_1_30));
wire output_3_30, output_3_1, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_1), .y(output_2_30));
wire output_1_31, output_1_2, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_2), .y(output_0_31));
wire output_2_31, output_2_2, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_2), .y(output_1_31));
wire output_3_31, output_3_2, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_2), .y(output_2_31));
assign output_0 = output_0_0;
wire output_0_32;
assign output_0_32 = input_0;
assign output_1 = output_1_0;
wire output_1_32;
assign output_1_32 = input_1;
assign output_2 = output_2_0;
wire output_2_32;
assign output_2_32 = input_2;
endmodule
