module Planar_Synthetic_5(
input Source1,
input Source2,
output Out1
);
wire flow_switch4_1_Source1;
wire flow_switch4_1_Mixer1;
wire flow_switch4_1_Mixer2;
wire flow_switch4_2_flow_switch4_1;
wire flow_switch4_2_Mixer3;
wire flow_switch4_2_Mixer4;
wire flow_switch4_3_flow_switch4_2;
wire flow_switch4_3_Mixer5;
wire flow_switch4_3_Mixer6;
wire flow_switch4_4_flow_switch4_3;
wire flow_switch4_4_Mixer7;
wire flow_switch4_4_Mixer8;
wire flow_switch4_5_flow_switch4_4;
wire flow_switch4_5_Heater1;
wire flow_switch4_5_Heater2;
wire flow_switch4_6_flow_switch4_5;
wire flow_switch4_6_Filter1;
wire flow_switch4_6_Filter2;
wire flow_switch4_7_Source2;
wire flow_switch4_7_Mixer9;
wire flow_switch4_7_Mixer10;
wire flow_switch4_8_flow_switch4_7;
wire flow_switch4_8_Mixer11;
wire flow_switch4_8_Mixer12;
wire flow_switch4_9_flow_switch4_8;
wire flow_switch4_9_Mixer13;
wire flow_switch4_9_Mixer14;
wire flow_switch4_10_flow_switch4_9;
wire flow_switch4_10_Mixer15;
wire flow_switch4_10_Mixer16;
wire flow_switch4_11_flow_switch4_10;
wire flow_switch4_11_Heater3;
wire flow_switch4_11_Heater4;
wire flow_switch4_12_flow_switch4_11;
wire flow_switch4_12_Filter3;
wire flow_switch4_12_Filter4;
wire Heater5_flow_switch4_6;
wire Heater6_flow_switch4_12;
wire Filter5_Heater5;
wire Filter6_Heater6;
wire flow_switch3_1_Filter5;
wire flow_switch3_1_Filter6;
wire Mixer17_flow_switch3_1;
wire Filter7_Mixer17;
wire Out1_Filter7;
assign flow_switch4_1_Source1 = Source1;
assign flow_switch4_7_Source2 = Source2;
chamber Mixer1(.port0(flow_switch4_1_Mixer1));
chamber Mixer2(.port1(flow_switch4_1_Mixer2));
chamber Mixer3(.port1(flow_switch4_2_Mixer3));
chamber Mixer4(.port1(flow_switch4_2_Mixer4));
chamber Mixer5(.port1(flow_switch4_3_Mixer5));
chamber Mixer6(.port1(flow_switch4_3_Mixer6));
chamber Mixer7(.port1(flow_switch4_4_Mixer7));
chamber Mixer8(.port1(flow_switch4_4_Mixer8));
chamber Mixer9(.port0(flow_switch4_7_Mixer9));
chamber Mixer10(.port1(flow_switch4_7_Mixer10));
chamber Mixer11(.port1(flow_switch4_8_Mixer11));
chamber Mixer12(.port1(flow_switch4_8_Mixer12));
chamber Mixer13(.port1(flow_switch4_9_Mixer13));
chamber Mixer14(.port1(flow_switch4_9_Mixer14));
chamber Mixer15(.port1(flow_switch4_10_Mixer15));
chamber Mixer16(.port1(flow_switch4_10_Mixer16));
chamber Mixer17(.port0(Filter7_Mixer17),.port1(Mixer17_flow_switch3_1));
heater Heater1(.port0(flow_switch4_5_Heater1));
heater Heater2(.port0(flow_switch4_5_Heater2));
heater Heater3(.port0(flow_switch4_11_Heater3));
heater Heater4(.port0(flow_switch4_11_Heater4));
heater Heater5(.port0(Filter5_Heater5),.port1(Heater5_flow_switch4_6));
heater Heater6(.port0(Heater6_flow_switch4_12),.port1(Filter6_Heater6));
filter Filter1(.port0(flow_switch4_6_Filter1));
filter Filter2(.port0(flow_switch4_6_Filter2));
filter Filter3(.port0(flow_switch4_12_Filter3));
filter Filter4(.port0(flow_switch4_12_Filter4));
filter Filter5(.port0(flow_switch3_1_Filter5),.port1(Filter5_Heater5));
filter Filter6(.port0(flow_switch3_1_Filter6),.port1(Filter6_Heater6));
filter Filter7(.port0(Filter7_Mixer17),.port1(Out1_Filter7));
assign Out1 = Out1_Filter7;
junction4 flow_switch4_1(.port0(flow_switch4_2_flow_switch4_1),.port1(flow_switch4_1_Source1),.port2(flow_switch4_1_Mixer1),.port3(flow_switch4_1_Mixer2));
junction4 flow_switch4_2(.port0(flow_switch4_2_Mixer4),.port1(flow_switch4_3_flow_switch4_2),.port2(flow_switch4_2_flow_switch4_1),.port3(flow_switch4_2_Mixer3));
junction4 flow_switch4_3(.port0(flow_switch4_3_Mixer6),.port1(flow_switch4_3_flow_switch4_2),.port2(flow_switch4_4_flow_switch4_3),.port3(flow_switch4_3_Mixer5));
junction4 flow_switch4_4(.port0(flow_switch4_4_Mixer8),.port1(flow_switch4_5_flow_switch4_4),.port2(flow_switch4_4_flow_switch4_3),.port3(flow_switch4_4_Mixer7));
junction4 flow_switch4_5(.port0(flow_switch4_5_Heater2),.port1(flow_switch4_5_flow_switch4_4),.port2(flow_switch4_6_flow_switch4_5),.port3(flow_switch4_5_Heater1));
junction4 flow_switch4_6(.port0(flow_switch4_6_Filter2),.port1(flow_switch4_6_flow_switch4_5),.port2(Heater5_flow_switch4_6),.port3(flow_switch4_6_Filter1));
junction4 flow_switch4_7(.port0(flow_switch4_7_Source2),.port1(flow_switch4_8_flow_switch4_7),.port2(flow_switch4_7_Mixer9),.port3(flow_switch4_7_Mixer10));
junction4 flow_switch4_8(.port0(flow_switch4_8_Mixer12),.port1(flow_switch4_9_flow_switch4_8),.port2(flow_switch4_8_flow_switch4_7),.port3(flow_switch4_8_Mixer11));
junction4 flow_switch4_9(.port0(flow_switch4_9_Mixer14),.port1(flow_switch4_9_flow_switch4_8),.port2(flow_switch4_10_flow_switch4_9),.port3(flow_switch4_9_Mixer13));
junction4 flow_switch4_10(.port0(flow_switch4_10_Mixer16),.port1(flow_switch4_10_flow_switch4_9),.port2(flow_switch4_11_flow_switch4_10),.port3(flow_switch4_10_Mixer15));
junction4 flow_switch4_11(.port0(flow_switch4_11_Heater4),.port1(flow_switch4_11_flow_switch4_10),.port2(flow_switch4_12_flow_switch4_11),.port3(flow_switch4_11_Heater3));
junction4 flow_switch4_12(.port0(flow_switch4_12_Filter3),.port1(Heater6_flow_switch4_12),.port2(flow_switch4_12_Filter4),.port3(flow_switch4_12_flow_switch4_11));
junction4 flow_switch3_1(.port1(Mixer17_flow_switch3_1),.port2(flow_switch3_1_Filter6),.port3(flow_switch3_1_Filter5));
endmodule
