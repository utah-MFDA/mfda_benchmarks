module fanout2_braid_8_96 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_1_7, output_1_0, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_0), .y(output_0_7));
wire output_2_7, output_2_0, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_0), .y(output_1_7));
wire output_3_7, output_3_0, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_0), .y(output_2_7));
wire output_4_7, output_4_0, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_0), .y(output_3_7));
wire output_5_7, output_5_0, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_0), .y(output_4_7));
wire output_6_7, output_6_0, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_0), .y(output_5_7));
wire output_7_7, output_7_0, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_0), .y(output_6_7));
wire output_8_7, output_8_0, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_0), .y(output_7_7));
wire output_1_8, output_1_1, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_1), .y(output_0_8));
wire output_2_8, output_2_1, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_1), .y(output_1_8));
wire output_3_8, output_3_1, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_1), .y(output_2_8));
wire output_4_8, output_4_1, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_1), .y(output_3_8));
wire output_5_8, output_5_1, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_1), .y(output_4_8));
wire output_6_8, output_6_1, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_1), .y(output_5_8));
wire output_7_8, output_7_1, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_1), .y(output_6_8));
wire output_8_8, output_8_1, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_1), .y(output_7_8));
wire output_1_9, output_1_2, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_2), .y(output_0_9));
wire output_2_9, output_2_2, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_2), .y(output_1_9));
wire output_3_9, output_3_2, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_2), .y(output_2_9));
wire output_4_9, output_4_2, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_2), .y(output_3_9));
wire output_5_9, output_5_2, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_2), .y(output_4_9));
wire output_6_9, output_6_2, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_2), .y(output_5_9));
wire output_7_9, output_7_2, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_2), .y(output_6_9));
wire output_8_9, output_8_2, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_2), .y(output_7_9));
wire output_1_10, output_1_3, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_3), .y(output_0_10));
wire output_2_10, output_2_3, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_3), .y(output_1_10));
wire output_3_10, output_3_3, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_3), .y(output_2_10));
wire output_4_10, output_4_3, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_3), .y(output_3_10));
wire output_5_10, output_5_3, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_3), .y(output_4_10));
wire output_6_10, output_6_3, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_3), .y(output_5_10));
wire output_7_10, output_7_3, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_3), .y(output_6_10));
wire output_8_10, output_8_3, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_3), .y(output_7_10));
wire output_1_11, output_1_4, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_4), .y(output_0_11));
wire output_2_11, output_2_4, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_4), .y(output_1_11));
wire output_3_11, output_3_4, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_4), .y(output_2_11));
wire output_4_11, output_4_4, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_4), .y(output_3_11));
wire output_5_11, output_5_4, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_4), .y(output_4_11));
wire output_6_11, output_6_4, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_4), .y(output_5_11));
wire output_7_11, output_7_4, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_4), .y(output_6_11));
wire output_8_11, output_8_4, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_4), .y(output_7_11));
wire output_1_12, output_1_5, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_5), .y(output_0_12));
wire output_2_12, output_2_5, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_5), .y(output_1_12));
wire output_3_12, output_3_5, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_5), .y(output_2_12));
wire output_4_12, output_4_5, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_5), .y(output_3_12));
wire output_5_12, output_5_5, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_5), .y(output_4_12));
wire output_6_12, output_6_5, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_5), .y(output_5_12));
wire output_7_12, output_7_5, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_5), .y(output_6_12));
wire output_8_12, output_8_5, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_5), .y(output_7_12));
wire output_1_13, output_1_6, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_6), .y(output_0_13));
wire output_2_13, output_2_6, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_6), .y(output_1_13));
wire output_3_13, output_3_6, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_6), .y(output_2_13));
wire output_4_13, output_4_6, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_6), .y(output_3_13));
wire output_5_13, output_5_6, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_6), .y(output_4_13));
wire output_6_13, output_6_6, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_6), .y(output_5_13));
wire output_7_13, output_7_6, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_6), .y(output_6_13));
wire output_8_13, output_8_6, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_6), .y(output_7_13));
wire output_1_14, output_1_7, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_7), .y(output_0_14));
wire output_2_14, output_2_7, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_7), .y(output_1_14));
wire output_3_14, output_3_7, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_7), .y(output_2_14));
wire output_4_14, output_4_7, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_7), .y(output_3_14));
wire output_5_14, output_5_7, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_7), .y(output_4_14));
wire output_6_14, output_6_7, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_7), .y(output_5_14));
wire output_7_14, output_7_7, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_7), .y(output_6_14));
wire output_8_14, output_8_7, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_7), .y(output_7_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
wire output_1_16, output_1_1, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_1), .y(output_0_16));
wire output_2_16, output_2_1, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_1), .y(output_1_16));
wire output_3_16, output_3_1, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_1), .y(output_2_16));
wire output_4_16, output_4_1, output_3_16;
mixer gate_output_3_16(.a(output_4_16), .b(output_4_1), .y(output_3_16));
wire output_5_16, output_5_1, output_4_16;
mixer gate_output_4_16(.a(output_5_16), .b(output_5_1), .y(output_4_16));
wire output_6_16, output_6_1, output_5_16;
mixer gate_output_5_16(.a(output_6_16), .b(output_6_1), .y(output_5_16));
wire output_7_16, output_7_1, output_6_16;
mixer gate_output_6_16(.a(output_7_16), .b(output_7_1), .y(output_6_16));
wire output_8_16, output_8_1, output_7_16;
mixer gate_output_7_16(.a(output_8_16), .b(output_8_1), .y(output_7_16));
wire output_1_17, output_1_2, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_2), .y(output_0_17));
wire output_2_17, output_2_2, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_2), .y(output_1_17));
wire output_3_17, output_3_2, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_2), .y(output_2_17));
wire output_4_17, output_4_2, output_3_17;
mixer gate_output_3_17(.a(output_4_17), .b(output_4_2), .y(output_3_17));
wire output_5_17, output_5_2, output_4_17;
mixer gate_output_4_17(.a(output_5_17), .b(output_5_2), .y(output_4_17));
wire output_6_17, output_6_2, output_5_17;
mixer gate_output_5_17(.a(output_6_17), .b(output_6_2), .y(output_5_17));
wire output_7_17, output_7_2, output_6_17;
mixer gate_output_6_17(.a(output_7_17), .b(output_7_2), .y(output_6_17));
wire output_8_17, output_8_2, output_7_17;
mixer gate_output_7_17(.a(output_8_17), .b(output_8_2), .y(output_7_17));
wire output_1_18, output_1_3, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_3), .y(output_0_18));
wire output_2_18, output_2_3, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_3), .y(output_1_18));
wire output_3_18, output_3_3, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_3), .y(output_2_18));
wire output_4_18, output_4_3, output_3_18;
mixer gate_output_3_18(.a(output_4_18), .b(output_4_3), .y(output_3_18));
wire output_5_18, output_5_3, output_4_18;
mixer gate_output_4_18(.a(output_5_18), .b(output_5_3), .y(output_4_18));
wire output_6_18, output_6_3, output_5_18;
mixer gate_output_5_18(.a(output_6_18), .b(output_6_3), .y(output_5_18));
wire output_7_18, output_7_3, output_6_18;
mixer gate_output_6_18(.a(output_7_18), .b(output_7_3), .y(output_6_18));
wire output_8_18, output_8_3, output_7_18;
mixer gate_output_7_18(.a(output_8_18), .b(output_8_3), .y(output_7_18));
wire output_1_19, output_1_4, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_4), .y(output_0_19));
wire output_2_19, output_2_4, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_4), .y(output_1_19));
wire output_3_19, output_3_4, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_4), .y(output_2_19));
wire output_4_19, output_4_4, output_3_19;
mixer gate_output_3_19(.a(output_4_19), .b(output_4_4), .y(output_3_19));
wire output_5_19, output_5_4, output_4_19;
mixer gate_output_4_19(.a(output_5_19), .b(output_5_4), .y(output_4_19));
wire output_6_19, output_6_4, output_5_19;
mixer gate_output_5_19(.a(output_6_19), .b(output_6_4), .y(output_5_19));
wire output_7_19, output_7_4, output_6_19;
mixer gate_output_6_19(.a(output_7_19), .b(output_7_4), .y(output_6_19));
wire output_8_19, output_8_4, output_7_19;
mixer gate_output_7_19(.a(output_8_19), .b(output_8_4), .y(output_7_19));
wire output_1_20, output_1_5, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_5), .y(output_0_20));
wire output_2_20, output_2_5, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_5), .y(output_1_20));
wire output_3_20, output_3_5, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_5), .y(output_2_20));
wire output_4_20, output_4_5, output_3_20;
mixer gate_output_3_20(.a(output_4_20), .b(output_4_5), .y(output_3_20));
wire output_5_20, output_5_5, output_4_20;
mixer gate_output_4_20(.a(output_5_20), .b(output_5_5), .y(output_4_20));
wire output_6_20, output_6_5, output_5_20;
mixer gate_output_5_20(.a(output_6_20), .b(output_6_5), .y(output_5_20));
wire output_7_20, output_7_5, output_6_20;
mixer gate_output_6_20(.a(output_7_20), .b(output_7_5), .y(output_6_20));
wire output_8_20, output_8_5, output_7_20;
mixer gate_output_7_20(.a(output_8_20), .b(output_8_5), .y(output_7_20));
wire output_1_21, output_1_6, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_6), .y(output_0_21));
wire output_2_21, output_2_6, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_6), .y(output_1_21));
wire output_3_21, output_3_6, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_6), .y(output_2_21));
wire output_4_21, output_4_6, output_3_21;
mixer gate_output_3_21(.a(output_4_21), .b(output_4_6), .y(output_3_21));
wire output_5_21, output_5_6, output_4_21;
mixer gate_output_4_21(.a(output_5_21), .b(output_5_6), .y(output_4_21));
wire output_6_21, output_6_6, output_5_21;
mixer gate_output_5_21(.a(output_6_21), .b(output_6_6), .y(output_5_21));
wire output_7_21, output_7_6, output_6_21;
mixer gate_output_6_21(.a(output_7_21), .b(output_7_6), .y(output_6_21));
wire output_8_21, output_8_6, output_7_21;
mixer gate_output_7_21(.a(output_8_21), .b(output_8_6), .y(output_7_21));
wire output_1_22, output_1_7, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_7), .y(output_0_22));
wire output_2_22, output_2_7, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_7), .y(output_1_22));
wire output_3_22, output_3_7, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_7), .y(output_2_22));
wire output_4_22, output_4_7, output_3_22;
mixer gate_output_3_22(.a(output_4_22), .b(output_4_7), .y(output_3_22));
wire output_5_22, output_5_7, output_4_22;
mixer gate_output_4_22(.a(output_5_22), .b(output_5_7), .y(output_4_22));
wire output_6_22, output_6_7, output_5_22;
mixer gate_output_5_22(.a(output_6_22), .b(output_6_7), .y(output_5_22));
wire output_7_22, output_7_7, output_6_22;
mixer gate_output_6_22(.a(output_7_22), .b(output_7_7), .y(output_6_22));
wire output_8_22, output_8_7, output_7_22;
mixer gate_output_7_22(.a(output_8_22), .b(output_8_7), .y(output_7_22));
wire output_1_23, output_1_0, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_0), .y(output_0_23));
wire output_2_23, output_2_0, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_0), .y(output_1_23));
wire output_3_23, output_3_0, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_0), .y(output_2_23));
wire output_4_23, output_4_0, output_3_23;
mixer gate_output_3_23(.a(output_4_23), .b(output_4_0), .y(output_3_23));
wire output_5_23, output_5_0, output_4_23;
mixer gate_output_4_23(.a(output_5_23), .b(output_5_0), .y(output_4_23));
wire output_6_23, output_6_0, output_5_23;
mixer gate_output_5_23(.a(output_6_23), .b(output_6_0), .y(output_5_23));
wire output_7_23, output_7_0, output_6_23;
mixer gate_output_6_23(.a(output_7_23), .b(output_7_0), .y(output_6_23));
wire output_8_23, output_8_0, output_7_23;
mixer gate_output_7_23(.a(output_8_23), .b(output_8_0), .y(output_7_23));
wire output_1_24, output_1_1, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_1), .y(output_0_24));
wire output_2_24, output_2_1, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_1), .y(output_1_24));
wire output_3_24, output_3_1, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_1), .y(output_2_24));
wire output_4_24, output_4_1, output_3_24;
mixer gate_output_3_24(.a(output_4_24), .b(output_4_1), .y(output_3_24));
wire output_5_24, output_5_1, output_4_24;
mixer gate_output_4_24(.a(output_5_24), .b(output_5_1), .y(output_4_24));
wire output_6_24, output_6_1, output_5_24;
mixer gate_output_5_24(.a(output_6_24), .b(output_6_1), .y(output_5_24));
wire output_7_24, output_7_1, output_6_24;
mixer gate_output_6_24(.a(output_7_24), .b(output_7_1), .y(output_6_24));
wire output_8_24, output_8_1, output_7_24;
mixer gate_output_7_24(.a(output_8_24), .b(output_8_1), .y(output_7_24));
wire output_1_25, output_1_2, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_2), .y(output_0_25));
wire output_2_25, output_2_2, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_2), .y(output_1_25));
wire output_3_25, output_3_2, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_2), .y(output_2_25));
wire output_4_25, output_4_2, output_3_25;
mixer gate_output_3_25(.a(output_4_25), .b(output_4_2), .y(output_3_25));
wire output_5_25, output_5_2, output_4_25;
mixer gate_output_4_25(.a(output_5_25), .b(output_5_2), .y(output_4_25));
wire output_6_25, output_6_2, output_5_25;
mixer gate_output_5_25(.a(output_6_25), .b(output_6_2), .y(output_5_25));
wire output_7_25, output_7_2, output_6_25;
mixer gate_output_6_25(.a(output_7_25), .b(output_7_2), .y(output_6_25));
wire output_8_25, output_8_2, output_7_25;
mixer gate_output_7_25(.a(output_8_25), .b(output_8_2), .y(output_7_25));
wire output_1_26, output_1_3, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_3), .y(output_0_26));
wire output_2_26, output_2_3, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_3), .y(output_1_26));
wire output_3_26, output_3_3, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_3), .y(output_2_26));
wire output_4_26, output_4_3, output_3_26;
mixer gate_output_3_26(.a(output_4_26), .b(output_4_3), .y(output_3_26));
wire output_5_26, output_5_3, output_4_26;
mixer gate_output_4_26(.a(output_5_26), .b(output_5_3), .y(output_4_26));
wire output_6_26, output_6_3, output_5_26;
mixer gate_output_5_26(.a(output_6_26), .b(output_6_3), .y(output_5_26));
wire output_7_26, output_7_3, output_6_26;
mixer gate_output_6_26(.a(output_7_26), .b(output_7_3), .y(output_6_26));
wire output_8_26, output_8_3, output_7_26;
mixer gate_output_7_26(.a(output_8_26), .b(output_8_3), .y(output_7_26));
wire output_1_27, output_1_4, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_4), .y(output_0_27));
wire output_2_27, output_2_4, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_4), .y(output_1_27));
wire output_3_27, output_3_4, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_4), .y(output_2_27));
wire output_4_27, output_4_4, output_3_27;
mixer gate_output_3_27(.a(output_4_27), .b(output_4_4), .y(output_3_27));
wire output_5_27, output_5_4, output_4_27;
mixer gate_output_4_27(.a(output_5_27), .b(output_5_4), .y(output_4_27));
wire output_6_27, output_6_4, output_5_27;
mixer gate_output_5_27(.a(output_6_27), .b(output_6_4), .y(output_5_27));
wire output_7_27, output_7_4, output_6_27;
mixer gate_output_6_27(.a(output_7_27), .b(output_7_4), .y(output_6_27));
wire output_8_27, output_8_4, output_7_27;
mixer gate_output_7_27(.a(output_8_27), .b(output_8_4), .y(output_7_27));
wire output_1_28, output_1_5, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_5), .y(output_0_28));
wire output_2_28, output_2_5, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_5), .y(output_1_28));
wire output_3_28, output_3_5, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_5), .y(output_2_28));
wire output_4_28, output_4_5, output_3_28;
mixer gate_output_3_28(.a(output_4_28), .b(output_4_5), .y(output_3_28));
wire output_5_28, output_5_5, output_4_28;
mixer gate_output_4_28(.a(output_5_28), .b(output_5_5), .y(output_4_28));
wire output_6_28, output_6_5, output_5_28;
mixer gate_output_5_28(.a(output_6_28), .b(output_6_5), .y(output_5_28));
wire output_7_28, output_7_5, output_6_28;
mixer gate_output_6_28(.a(output_7_28), .b(output_7_5), .y(output_6_28));
wire output_8_28, output_8_5, output_7_28;
mixer gate_output_7_28(.a(output_8_28), .b(output_8_5), .y(output_7_28));
wire output_1_29, output_1_6, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_6), .y(output_0_29));
wire output_2_29, output_2_6, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_6), .y(output_1_29));
wire output_3_29, output_3_6, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_6), .y(output_2_29));
wire output_4_29, output_4_6, output_3_29;
mixer gate_output_3_29(.a(output_4_29), .b(output_4_6), .y(output_3_29));
wire output_5_29, output_5_6, output_4_29;
mixer gate_output_4_29(.a(output_5_29), .b(output_5_6), .y(output_4_29));
wire output_6_29, output_6_6, output_5_29;
mixer gate_output_5_29(.a(output_6_29), .b(output_6_6), .y(output_5_29));
wire output_7_29, output_7_6, output_6_29;
mixer gate_output_6_29(.a(output_7_29), .b(output_7_6), .y(output_6_29));
wire output_8_29, output_8_6, output_7_29;
mixer gate_output_7_29(.a(output_8_29), .b(output_8_6), .y(output_7_29));
wire output_1_30, output_1_7, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_7), .y(output_0_30));
wire output_2_30, output_2_7, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_7), .y(output_1_30));
wire output_3_30, output_3_7, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_7), .y(output_2_30));
wire output_4_30, output_4_7, output_3_30;
mixer gate_output_3_30(.a(output_4_30), .b(output_4_7), .y(output_3_30));
wire output_5_30, output_5_7, output_4_30;
mixer gate_output_4_30(.a(output_5_30), .b(output_5_7), .y(output_4_30));
wire output_6_30, output_6_7, output_5_30;
mixer gate_output_5_30(.a(output_6_30), .b(output_6_7), .y(output_5_30));
wire output_7_30, output_7_7, output_6_30;
mixer gate_output_6_30(.a(output_7_30), .b(output_7_7), .y(output_6_30));
wire output_8_30, output_8_7, output_7_30;
mixer gate_output_7_30(.a(output_8_30), .b(output_8_7), .y(output_7_30));
wire output_1_31, output_1_0, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_0), .y(output_0_31));
wire output_2_31, output_2_0, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_0), .y(output_1_31));
wire output_3_31, output_3_0, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_0), .y(output_2_31));
wire output_4_31, output_4_0, output_3_31;
mixer gate_output_3_31(.a(output_4_31), .b(output_4_0), .y(output_3_31));
wire output_5_31, output_5_0, output_4_31;
mixer gate_output_4_31(.a(output_5_31), .b(output_5_0), .y(output_4_31));
wire output_6_31, output_6_0, output_5_31;
mixer gate_output_5_31(.a(output_6_31), .b(output_6_0), .y(output_5_31));
wire output_7_31, output_7_0, output_6_31;
mixer gate_output_6_31(.a(output_7_31), .b(output_7_0), .y(output_6_31));
wire output_8_31, output_8_0, output_7_31;
mixer gate_output_7_31(.a(output_8_31), .b(output_8_0), .y(output_7_31));
wire output_1_32, output_1_1, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_1), .y(output_0_32));
wire output_2_32, output_2_1, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_1), .y(output_1_32));
wire output_3_32, output_3_1, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_1), .y(output_2_32));
wire output_4_32, output_4_1, output_3_32;
mixer gate_output_3_32(.a(output_4_32), .b(output_4_1), .y(output_3_32));
wire output_5_32, output_5_1, output_4_32;
mixer gate_output_4_32(.a(output_5_32), .b(output_5_1), .y(output_4_32));
wire output_6_32, output_6_1, output_5_32;
mixer gate_output_5_32(.a(output_6_32), .b(output_6_1), .y(output_5_32));
wire output_7_32, output_7_1, output_6_32;
mixer gate_output_6_32(.a(output_7_32), .b(output_7_1), .y(output_6_32));
wire output_8_32, output_8_1, output_7_32;
mixer gate_output_7_32(.a(output_8_32), .b(output_8_1), .y(output_7_32));
wire output_1_33, output_1_2, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_2), .y(output_0_33));
wire output_2_33, output_2_2, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_2), .y(output_1_33));
wire output_3_33, output_3_2, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_2), .y(output_2_33));
wire output_4_33, output_4_2, output_3_33;
mixer gate_output_3_33(.a(output_4_33), .b(output_4_2), .y(output_3_33));
wire output_5_33, output_5_2, output_4_33;
mixer gate_output_4_33(.a(output_5_33), .b(output_5_2), .y(output_4_33));
wire output_6_33, output_6_2, output_5_33;
mixer gate_output_5_33(.a(output_6_33), .b(output_6_2), .y(output_5_33));
wire output_7_33, output_7_2, output_6_33;
mixer gate_output_6_33(.a(output_7_33), .b(output_7_2), .y(output_6_33));
wire output_8_33, output_8_2, output_7_33;
mixer gate_output_7_33(.a(output_8_33), .b(output_8_2), .y(output_7_33));
wire output_1_34, output_1_3, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_3), .y(output_0_34));
wire output_2_34, output_2_3, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_3), .y(output_1_34));
wire output_3_34, output_3_3, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_3), .y(output_2_34));
wire output_4_34, output_4_3, output_3_34;
mixer gate_output_3_34(.a(output_4_34), .b(output_4_3), .y(output_3_34));
wire output_5_34, output_5_3, output_4_34;
mixer gate_output_4_34(.a(output_5_34), .b(output_5_3), .y(output_4_34));
wire output_6_34, output_6_3, output_5_34;
mixer gate_output_5_34(.a(output_6_34), .b(output_6_3), .y(output_5_34));
wire output_7_34, output_7_3, output_6_34;
mixer gate_output_6_34(.a(output_7_34), .b(output_7_3), .y(output_6_34));
wire output_8_34, output_8_3, output_7_34;
mixer gate_output_7_34(.a(output_8_34), .b(output_8_3), .y(output_7_34));
wire output_1_35, output_1_4, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_4), .y(output_0_35));
wire output_2_35, output_2_4, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_4), .y(output_1_35));
wire output_3_35, output_3_4, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_4), .y(output_2_35));
wire output_4_35, output_4_4, output_3_35;
mixer gate_output_3_35(.a(output_4_35), .b(output_4_4), .y(output_3_35));
wire output_5_35, output_5_4, output_4_35;
mixer gate_output_4_35(.a(output_5_35), .b(output_5_4), .y(output_4_35));
wire output_6_35, output_6_4, output_5_35;
mixer gate_output_5_35(.a(output_6_35), .b(output_6_4), .y(output_5_35));
wire output_7_35, output_7_4, output_6_35;
mixer gate_output_6_35(.a(output_7_35), .b(output_7_4), .y(output_6_35));
wire output_8_35, output_8_4, output_7_35;
mixer gate_output_7_35(.a(output_8_35), .b(output_8_4), .y(output_7_35));
wire output_1_36, output_1_5, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_5), .y(output_0_36));
wire output_2_36, output_2_5, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_5), .y(output_1_36));
wire output_3_36, output_3_5, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_5), .y(output_2_36));
wire output_4_36, output_4_5, output_3_36;
mixer gate_output_3_36(.a(output_4_36), .b(output_4_5), .y(output_3_36));
wire output_5_36, output_5_5, output_4_36;
mixer gate_output_4_36(.a(output_5_36), .b(output_5_5), .y(output_4_36));
wire output_6_36, output_6_5, output_5_36;
mixer gate_output_5_36(.a(output_6_36), .b(output_6_5), .y(output_5_36));
wire output_7_36, output_7_5, output_6_36;
mixer gate_output_6_36(.a(output_7_36), .b(output_7_5), .y(output_6_36));
wire output_8_36, output_8_5, output_7_36;
mixer gate_output_7_36(.a(output_8_36), .b(output_8_5), .y(output_7_36));
wire output_1_37, output_1_6, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_6), .y(output_0_37));
wire output_2_37, output_2_6, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_6), .y(output_1_37));
wire output_3_37, output_3_6, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_6), .y(output_2_37));
wire output_4_37, output_4_6, output_3_37;
mixer gate_output_3_37(.a(output_4_37), .b(output_4_6), .y(output_3_37));
wire output_5_37, output_5_6, output_4_37;
mixer gate_output_4_37(.a(output_5_37), .b(output_5_6), .y(output_4_37));
wire output_6_37, output_6_6, output_5_37;
mixer gate_output_5_37(.a(output_6_37), .b(output_6_6), .y(output_5_37));
wire output_7_37, output_7_6, output_6_37;
mixer gate_output_6_37(.a(output_7_37), .b(output_7_6), .y(output_6_37));
wire output_8_37, output_8_6, output_7_37;
mixer gate_output_7_37(.a(output_8_37), .b(output_8_6), .y(output_7_37));
wire output_1_38, output_1_7, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_7), .y(output_0_38));
wire output_2_38, output_2_7, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_7), .y(output_1_38));
wire output_3_38, output_3_7, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_7), .y(output_2_38));
wire output_4_38, output_4_7, output_3_38;
mixer gate_output_3_38(.a(output_4_38), .b(output_4_7), .y(output_3_38));
wire output_5_38, output_5_7, output_4_38;
mixer gate_output_4_38(.a(output_5_38), .b(output_5_7), .y(output_4_38));
wire output_6_38, output_6_7, output_5_38;
mixer gate_output_5_38(.a(output_6_38), .b(output_6_7), .y(output_5_38));
wire output_7_38, output_7_7, output_6_38;
mixer gate_output_6_38(.a(output_7_38), .b(output_7_7), .y(output_6_38));
wire output_8_38, output_8_7, output_7_38;
mixer gate_output_7_38(.a(output_8_38), .b(output_8_7), .y(output_7_38));
wire output_1_39, output_1_0, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_0), .y(output_0_39));
wire output_2_39, output_2_0, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_0), .y(output_1_39));
wire output_3_39, output_3_0, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_0), .y(output_2_39));
wire output_4_39, output_4_0, output_3_39;
mixer gate_output_3_39(.a(output_4_39), .b(output_4_0), .y(output_3_39));
wire output_5_39, output_5_0, output_4_39;
mixer gate_output_4_39(.a(output_5_39), .b(output_5_0), .y(output_4_39));
wire output_6_39, output_6_0, output_5_39;
mixer gate_output_5_39(.a(output_6_39), .b(output_6_0), .y(output_5_39));
wire output_7_39, output_7_0, output_6_39;
mixer gate_output_6_39(.a(output_7_39), .b(output_7_0), .y(output_6_39));
wire output_8_39, output_8_0, output_7_39;
mixer gate_output_7_39(.a(output_8_39), .b(output_8_0), .y(output_7_39));
wire output_1_40, output_1_1, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_1), .y(output_0_40));
wire output_2_40, output_2_1, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_1), .y(output_1_40));
wire output_3_40, output_3_1, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_1), .y(output_2_40));
wire output_4_40, output_4_1, output_3_40;
mixer gate_output_3_40(.a(output_4_40), .b(output_4_1), .y(output_3_40));
wire output_5_40, output_5_1, output_4_40;
mixer gate_output_4_40(.a(output_5_40), .b(output_5_1), .y(output_4_40));
wire output_6_40, output_6_1, output_5_40;
mixer gate_output_5_40(.a(output_6_40), .b(output_6_1), .y(output_5_40));
wire output_7_40, output_7_1, output_6_40;
mixer gate_output_6_40(.a(output_7_40), .b(output_7_1), .y(output_6_40));
wire output_8_40, output_8_1, output_7_40;
mixer gate_output_7_40(.a(output_8_40), .b(output_8_1), .y(output_7_40));
wire output_1_41, output_1_2, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_2), .y(output_0_41));
wire output_2_41, output_2_2, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_2), .y(output_1_41));
wire output_3_41, output_3_2, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_2), .y(output_2_41));
wire output_4_41, output_4_2, output_3_41;
mixer gate_output_3_41(.a(output_4_41), .b(output_4_2), .y(output_3_41));
wire output_5_41, output_5_2, output_4_41;
mixer gate_output_4_41(.a(output_5_41), .b(output_5_2), .y(output_4_41));
wire output_6_41, output_6_2, output_5_41;
mixer gate_output_5_41(.a(output_6_41), .b(output_6_2), .y(output_5_41));
wire output_7_41, output_7_2, output_6_41;
mixer gate_output_6_41(.a(output_7_41), .b(output_7_2), .y(output_6_41));
wire output_8_41, output_8_2, output_7_41;
mixer gate_output_7_41(.a(output_8_41), .b(output_8_2), .y(output_7_41));
wire output_1_42, output_1_3, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_3), .y(output_0_42));
wire output_2_42, output_2_3, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_3), .y(output_1_42));
wire output_3_42, output_3_3, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_3), .y(output_2_42));
wire output_4_42, output_4_3, output_3_42;
mixer gate_output_3_42(.a(output_4_42), .b(output_4_3), .y(output_3_42));
wire output_5_42, output_5_3, output_4_42;
mixer gate_output_4_42(.a(output_5_42), .b(output_5_3), .y(output_4_42));
wire output_6_42, output_6_3, output_5_42;
mixer gate_output_5_42(.a(output_6_42), .b(output_6_3), .y(output_5_42));
wire output_7_42, output_7_3, output_6_42;
mixer gate_output_6_42(.a(output_7_42), .b(output_7_3), .y(output_6_42));
wire output_8_42, output_8_3, output_7_42;
mixer gate_output_7_42(.a(output_8_42), .b(output_8_3), .y(output_7_42));
wire output_1_43, output_1_4, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_4), .y(output_0_43));
wire output_2_43, output_2_4, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_4), .y(output_1_43));
wire output_3_43, output_3_4, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_4), .y(output_2_43));
wire output_4_43, output_4_4, output_3_43;
mixer gate_output_3_43(.a(output_4_43), .b(output_4_4), .y(output_3_43));
wire output_5_43, output_5_4, output_4_43;
mixer gate_output_4_43(.a(output_5_43), .b(output_5_4), .y(output_4_43));
wire output_6_43, output_6_4, output_5_43;
mixer gate_output_5_43(.a(output_6_43), .b(output_6_4), .y(output_5_43));
wire output_7_43, output_7_4, output_6_43;
mixer gate_output_6_43(.a(output_7_43), .b(output_7_4), .y(output_6_43));
wire output_8_43, output_8_4, output_7_43;
mixer gate_output_7_43(.a(output_8_43), .b(output_8_4), .y(output_7_43));
wire output_1_44, output_1_5, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_5), .y(output_0_44));
wire output_2_44, output_2_5, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_5), .y(output_1_44));
wire output_3_44, output_3_5, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_5), .y(output_2_44));
wire output_4_44, output_4_5, output_3_44;
mixer gate_output_3_44(.a(output_4_44), .b(output_4_5), .y(output_3_44));
wire output_5_44, output_5_5, output_4_44;
mixer gate_output_4_44(.a(output_5_44), .b(output_5_5), .y(output_4_44));
wire output_6_44, output_6_5, output_5_44;
mixer gate_output_5_44(.a(output_6_44), .b(output_6_5), .y(output_5_44));
wire output_7_44, output_7_5, output_6_44;
mixer gate_output_6_44(.a(output_7_44), .b(output_7_5), .y(output_6_44));
wire output_8_44, output_8_5, output_7_44;
mixer gate_output_7_44(.a(output_8_44), .b(output_8_5), .y(output_7_44));
wire output_1_45, output_1_6, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_6), .y(output_0_45));
wire output_2_45, output_2_6, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_6), .y(output_1_45));
wire output_3_45, output_3_6, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_6), .y(output_2_45));
wire output_4_45, output_4_6, output_3_45;
mixer gate_output_3_45(.a(output_4_45), .b(output_4_6), .y(output_3_45));
wire output_5_45, output_5_6, output_4_45;
mixer gate_output_4_45(.a(output_5_45), .b(output_5_6), .y(output_4_45));
wire output_6_45, output_6_6, output_5_45;
mixer gate_output_5_45(.a(output_6_45), .b(output_6_6), .y(output_5_45));
wire output_7_45, output_7_6, output_6_45;
mixer gate_output_6_45(.a(output_7_45), .b(output_7_6), .y(output_6_45));
wire output_8_45, output_8_6, output_7_45;
mixer gate_output_7_45(.a(output_8_45), .b(output_8_6), .y(output_7_45));
wire output_1_46, output_1_7, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_7), .y(output_0_46));
wire output_2_46, output_2_7, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_7), .y(output_1_46));
wire output_3_46, output_3_7, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_7), .y(output_2_46));
wire output_4_46, output_4_7, output_3_46;
mixer gate_output_3_46(.a(output_4_46), .b(output_4_7), .y(output_3_46));
wire output_5_46, output_5_7, output_4_46;
mixer gate_output_4_46(.a(output_5_46), .b(output_5_7), .y(output_4_46));
wire output_6_46, output_6_7, output_5_46;
mixer gate_output_5_46(.a(output_6_46), .b(output_6_7), .y(output_5_46));
wire output_7_46, output_7_7, output_6_46;
mixer gate_output_6_46(.a(output_7_46), .b(output_7_7), .y(output_6_46));
wire output_8_46, output_8_7, output_7_46;
mixer gate_output_7_46(.a(output_8_46), .b(output_8_7), .y(output_7_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_4_47, output_4_0, output_3_47;
mixer gate_output_3_47(.a(output_4_47), .b(output_4_0), .y(output_3_47));
wire output_5_47, output_5_0, output_4_47;
mixer gate_output_4_47(.a(output_5_47), .b(output_5_0), .y(output_4_47));
wire output_6_47, output_6_0, output_5_47;
mixer gate_output_5_47(.a(output_6_47), .b(output_6_0), .y(output_5_47));
wire output_7_47, output_7_0, output_6_47;
mixer gate_output_6_47(.a(output_7_47), .b(output_7_0), .y(output_6_47));
wire output_8_47, output_8_0, output_7_47;
mixer gate_output_7_47(.a(output_8_47), .b(output_8_0), .y(output_7_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_4_48, output_4_1, output_3_48;
mixer gate_output_3_48(.a(output_4_48), .b(output_4_1), .y(output_3_48));
wire output_5_48, output_5_1, output_4_48;
mixer gate_output_4_48(.a(output_5_48), .b(output_5_1), .y(output_4_48));
wire output_6_48, output_6_1, output_5_48;
mixer gate_output_5_48(.a(output_6_48), .b(output_6_1), .y(output_5_48));
wire output_7_48, output_7_1, output_6_48;
mixer gate_output_6_48(.a(output_7_48), .b(output_7_1), .y(output_6_48));
wire output_8_48, output_8_1, output_7_48;
mixer gate_output_7_48(.a(output_8_48), .b(output_8_1), .y(output_7_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_4_49, output_4_2, output_3_49;
mixer gate_output_3_49(.a(output_4_49), .b(output_4_2), .y(output_3_49));
wire output_5_49, output_5_2, output_4_49;
mixer gate_output_4_49(.a(output_5_49), .b(output_5_2), .y(output_4_49));
wire output_6_49, output_6_2, output_5_49;
mixer gate_output_5_49(.a(output_6_49), .b(output_6_2), .y(output_5_49));
wire output_7_49, output_7_2, output_6_49;
mixer gate_output_6_49(.a(output_7_49), .b(output_7_2), .y(output_6_49));
wire output_8_49, output_8_2, output_7_49;
mixer gate_output_7_49(.a(output_8_49), .b(output_8_2), .y(output_7_49));
wire output_1_50, output_1_3, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_3), .y(output_0_50));
wire output_2_50, output_2_3, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_3), .y(output_1_50));
wire output_3_50, output_3_3, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_3), .y(output_2_50));
wire output_4_50, output_4_3, output_3_50;
mixer gate_output_3_50(.a(output_4_50), .b(output_4_3), .y(output_3_50));
wire output_5_50, output_5_3, output_4_50;
mixer gate_output_4_50(.a(output_5_50), .b(output_5_3), .y(output_4_50));
wire output_6_50, output_6_3, output_5_50;
mixer gate_output_5_50(.a(output_6_50), .b(output_6_3), .y(output_5_50));
wire output_7_50, output_7_3, output_6_50;
mixer gate_output_6_50(.a(output_7_50), .b(output_7_3), .y(output_6_50));
wire output_8_50, output_8_3, output_7_50;
mixer gate_output_7_50(.a(output_8_50), .b(output_8_3), .y(output_7_50));
wire output_1_51, output_1_4, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_4), .y(output_0_51));
wire output_2_51, output_2_4, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_4), .y(output_1_51));
wire output_3_51, output_3_4, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_4), .y(output_2_51));
wire output_4_51, output_4_4, output_3_51;
mixer gate_output_3_51(.a(output_4_51), .b(output_4_4), .y(output_3_51));
wire output_5_51, output_5_4, output_4_51;
mixer gate_output_4_51(.a(output_5_51), .b(output_5_4), .y(output_4_51));
wire output_6_51, output_6_4, output_5_51;
mixer gate_output_5_51(.a(output_6_51), .b(output_6_4), .y(output_5_51));
wire output_7_51, output_7_4, output_6_51;
mixer gate_output_6_51(.a(output_7_51), .b(output_7_4), .y(output_6_51));
wire output_8_51, output_8_4, output_7_51;
mixer gate_output_7_51(.a(output_8_51), .b(output_8_4), .y(output_7_51));
wire output_1_52, output_1_5, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_5), .y(output_0_52));
wire output_2_52, output_2_5, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_5), .y(output_1_52));
wire output_3_52, output_3_5, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_5), .y(output_2_52));
wire output_4_52, output_4_5, output_3_52;
mixer gate_output_3_52(.a(output_4_52), .b(output_4_5), .y(output_3_52));
wire output_5_52, output_5_5, output_4_52;
mixer gate_output_4_52(.a(output_5_52), .b(output_5_5), .y(output_4_52));
wire output_6_52, output_6_5, output_5_52;
mixer gate_output_5_52(.a(output_6_52), .b(output_6_5), .y(output_5_52));
wire output_7_52, output_7_5, output_6_52;
mixer gate_output_6_52(.a(output_7_52), .b(output_7_5), .y(output_6_52));
wire output_8_52, output_8_5, output_7_52;
mixer gate_output_7_52(.a(output_8_52), .b(output_8_5), .y(output_7_52));
wire output_1_53, output_1_6, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_6), .y(output_0_53));
wire output_2_53, output_2_6, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_6), .y(output_1_53));
wire output_3_53, output_3_6, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_6), .y(output_2_53));
wire output_4_53, output_4_6, output_3_53;
mixer gate_output_3_53(.a(output_4_53), .b(output_4_6), .y(output_3_53));
wire output_5_53, output_5_6, output_4_53;
mixer gate_output_4_53(.a(output_5_53), .b(output_5_6), .y(output_4_53));
wire output_6_53, output_6_6, output_5_53;
mixer gate_output_5_53(.a(output_6_53), .b(output_6_6), .y(output_5_53));
wire output_7_53, output_7_6, output_6_53;
mixer gate_output_6_53(.a(output_7_53), .b(output_7_6), .y(output_6_53));
wire output_8_53, output_8_6, output_7_53;
mixer gate_output_7_53(.a(output_8_53), .b(output_8_6), .y(output_7_53));
wire output_1_54, output_1_7, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_7), .y(output_0_54));
wire output_2_54, output_2_7, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_7), .y(output_1_54));
wire output_3_54, output_3_7, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_7), .y(output_2_54));
wire output_4_54, output_4_7, output_3_54;
mixer gate_output_3_54(.a(output_4_54), .b(output_4_7), .y(output_3_54));
wire output_5_54, output_5_7, output_4_54;
mixer gate_output_4_54(.a(output_5_54), .b(output_5_7), .y(output_4_54));
wire output_6_54, output_6_7, output_5_54;
mixer gate_output_5_54(.a(output_6_54), .b(output_6_7), .y(output_5_54));
wire output_7_54, output_7_7, output_6_54;
mixer gate_output_6_54(.a(output_7_54), .b(output_7_7), .y(output_6_54));
wire output_8_54, output_8_7, output_7_54;
mixer gate_output_7_54(.a(output_8_54), .b(output_8_7), .y(output_7_54));
wire output_1_55, output_1_0, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_0), .y(output_0_55));
wire output_2_55, output_2_0, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_0), .y(output_1_55));
wire output_3_55, output_3_0, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_0), .y(output_2_55));
wire output_4_55, output_4_0, output_3_55;
mixer gate_output_3_55(.a(output_4_55), .b(output_4_0), .y(output_3_55));
wire output_5_55, output_5_0, output_4_55;
mixer gate_output_4_55(.a(output_5_55), .b(output_5_0), .y(output_4_55));
wire output_6_55, output_6_0, output_5_55;
mixer gate_output_5_55(.a(output_6_55), .b(output_6_0), .y(output_5_55));
wire output_7_55, output_7_0, output_6_55;
mixer gate_output_6_55(.a(output_7_55), .b(output_7_0), .y(output_6_55));
wire output_8_55, output_8_0, output_7_55;
mixer gate_output_7_55(.a(output_8_55), .b(output_8_0), .y(output_7_55));
wire output_1_56, output_1_1, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_1), .y(output_0_56));
wire output_2_56, output_2_1, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_1), .y(output_1_56));
wire output_3_56, output_3_1, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_1), .y(output_2_56));
wire output_4_56, output_4_1, output_3_56;
mixer gate_output_3_56(.a(output_4_56), .b(output_4_1), .y(output_3_56));
wire output_5_56, output_5_1, output_4_56;
mixer gate_output_4_56(.a(output_5_56), .b(output_5_1), .y(output_4_56));
wire output_6_56, output_6_1, output_5_56;
mixer gate_output_5_56(.a(output_6_56), .b(output_6_1), .y(output_5_56));
wire output_7_56, output_7_1, output_6_56;
mixer gate_output_6_56(.a(output_7_56), .b(output_7_1), .y(output_6_56));
wire output_8_56, output_8_1, output_7_56;
mixer gate_output_7_56(.a(output_8_56), .b(output_8_1), .y(output_7_56));
wire output_1_57, output_1_2, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_2), .y(output_0_57));
wire output_2_57, output_2_2, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_2), .y(output_1_57));
wire output_3_57, output_3_2, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_2), .y(output_2_57));
wire output_4_57, output_4_2, output_3_57;
mixer gate_output_3_57(.a(output_4_57), .b(output_4_2), .y(output_3_57));
wire output_5_57, output_5_2, output_4_57;
mixer gate_output_4_57(.a(output_5_57), .b(output_5_2), .y(output_4_57));
wire output_6_57, output_6_2, output_5_57;
mixer gate_output_5_57(.a(output_6_57), .b(output_6_2), .y(output_5_57));
wire output_7_57, output_7_2, output_6_57;
mixer gate_output_6_57(.a(output_7_57), .b(output_7_2), .y(output_6_57));
wire output_8_57, output_8_2, output_7_57;
mixer gate_output_7_57(.a(output_8_57), .b(output_8_2), .y(output_7_57));
wire output_1_58, output_1_3, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_3), .y(output_0_58));
wire output_2_58, output_2_3, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_3), .y(output_1_58));
wire output_3_58, output_3_3, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_3), .y(output_2_58));
wire output_4_58, output_4_3, output_3_58;
mixer gate_output_3_58(.a(output_4_58), .b(output_4_3), .y(output_3_58));
wire output_5_58, output_5_3, output_4_58;
mixer gate_output_4_58(.a(output_5_58), .b(output_5_3), .y(output_4_58));
wire output_6_58, output_6_3, output_5_58;
mixer gate_output_5_58(.a(output_6_58), .b(output_6_3), .y(output_5_58));
wire output_7_58, output_7_3, output_6_58;
mixer gate_output_6_58(.a(output_7_58), .b(output_7_3), .y(output_6_58));
wire output_8_58, output_8_3, output_7_58;
mixer gate_output_7_58(.a(output_8_58), .b(output_8_3), .y(output_7_58));
wire output_1_59, output_1_4, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_4), .y(output_0_59));
wire output_2_59, output_2_4, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_4), .y(output_1_59));
wire output_3_59, output_3_4, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_4), .y(output_2_59));
wire output_4_59, output_4_4, output_3_59;
mixer gate_output_3_59(.a(output_4_59), .b(output_4_4), .y(output_3_59));
wire output_5_59, output_5_4, output_4_59;
mixer gate_output_4_59(.a(output_5_59), .b(output_5_4), .y(output_4_59));
wire output_6_59, output_6_4, output_5_59;
mixer gate_output_5_59(.a(output_6_59), .b(output_6_4), .y(output_5_59));
wire output_7_59, output_7_4, output_6_59;
mixer gate_output_6_59(.a(output_7_59), .b(output_7_4), .y(output_6_59));
wire output_8_59, output_8_4, output_7_59;
mixer gate_output_7_59(.a(output_8_59), .b(output_8_4), .y(output_7_59));
wire output_1_60, output_1_5, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_5), .y(output_0_60));
wire output_2_60, output_2_5, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_5), .y(output_1_60));
wire output_3_60, output_3_5, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_5), .y(output_2_60));
wire output_4_60, output_4_5, output_3_60;
mixer gate_output_3_60(.a(output_4_60), .b(output_4_5), .y(output_3_60));
wire output_5_60, output_5_5, output_4_60;
mixer gate_output_4_60(.a(output_5_60), .b(output_5_5), .y(output_4_60));
wire output_6_60, output_6_5, output_5_60;
mixer gate_output_5_60(.a(output_6_60), .b(output_6_5), .y(output_5_60));
wire output_7_60, output_7_5, output_6_60;
mixer gate_output_6_60(.a(output_7_60), .b(output_7_5), .y(output_6_60));
wire output_8_60, output_8_5, output_7_60;
mixer gate_output_7_60(.a(output_8_60), .b(output_8_5), .y(output_7_60));
wire output_1_61, output_1_6, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_6), .y(output_0_61));
wire output_2_61, output_2_6, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_6), .y(output_1_61));
wire output_3_61, output_3_6, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_6), .y(output_2_61));
wire output_4_61, output_4_6, output_3_61;
mixer gate_output_3_61(.a(output_4_61), .b(output_4_6), .y(output_3_61));
wire output_5_61, output_5_6, output_4_61;
mixer gate_output_4_61(.a(output_5_61), .b(output_5_6), .y(output_4_61));
wire output_6_61, output_6_6, output_5_61;
mixer gate_output_5_61(.a(output_6_61), .b(output_6_6), .y(output_5_61));
wire output_7_61, output_7_6, output_6_61;
mixer gate_output_6_61(.a(output_7_61), .b(output_7_6), .y(output_6_61));
wire output_8_61, output_8_6, output_7_61;
mixer gate_output_7_61(.a(output_8_61), .b(output_8_6), .y(output_7_61));
wire output_1_62, output_1_7, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_7), .y(output_0_62));
wire output_2_62, output_2_7, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_7), .y(output_1_62));
wire output_3_62, output_3_7, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_7), .y(output_2_62));
wire output_4_62, output_4_7, output_3_62;
mixer gate_output_3_62(.a(output_4_62), .b(output_4_7), .y(output_3_62));
wire output_5_62, output_5_7, output_4_62;
mixer gate_output_4_62(.a(output_5_62), .b(output_5_7), .y(output_4_62));
wire output_6_62, output_6_7, output_5_62;
mixer gate_output_5_62(.a(output_6_62), .b(output_6_7), .y(output_5_62));
wire output_7_62, output_7_7, output_6_62;
mixer gate_output_6_62(.a(output_7_62), .b(output_7_7), .y(output_6_62));
wire output_8_62, output_8_7, output_7_62;
mixer gate_output_7_62(.a(output_8_62), .b(output_8_7), .y(output_7_62));
wire output_1_63, output_1_0, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_0), .y(output_0_63));
wire output_2_63, output_2_0, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_0), .y(output_1_63));
wire output_3_63, output_3_0, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_0), .y(output_2_63));
wire output_4_63, output_4_0, output_3_63;
mixer gate_output_3_63(.a(output_4_63), .b(output_4_0), .y(output_3_63));
wire output_5_63, output_5_0, output_4_63;
mixer gate_output_4_63(.a(output_5_63), .b(output_5_0), .y(output_4_63));
wire output_6_63, output_6_0, output_5_63;
mixer gate_output_5_63(.a(output_6_63), .b(output_6_0), .y(output_5_63));
wire output_7_63, output_7_0, output_6_63;
mixer gate_output_6_63(.a(output_7_63), .b(output_7_0), .y(output_6_63));
wire output_8_63, output_8_0, output_7_63;
mixer gate_output_7_63(.a(output_8_63), .b(output_8_0), .y(output_7_63));
wire output_1_64, output_1_1, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_1), .y(output_0_64));
wire output_2_64, output_2_1, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_1), .y(output_1_64));
wire output_3_64, output_3_1, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_1), .y(output_2_64));
wire output_4_64, output_4_1, output_3_64;
mixer gate_output_3_64(.a(output_4_64), .b(output_4_1), .y(output_3_64));
wire output_5_64, output_5_1, output_4_64;
mixer gate_output_4_64(.a(output_5_64), .b(output_5_1), .y(output_4_64));
wire output_6_64, output_6_1, output_5_64;
mixer gate_output_5_64(.a(output_6_64), .b(output_6_1), .y(output_5_64));
wire output_7_64, output_7_1, output_6_64;
mixer gate_output_6_64(.a(output_7_64), .b(output_7_1), .y(output_6_64));
wire output_8_64, output_8_1, output_7_64;
mixer gate_output_7_64(.a(output_8_64), .b(output_8_1), .y(output_7_64));
wire output_1_65, output_1_2, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_2), .y(output_0_65));
wire output_2_65, output_2_2, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_2), .y(output_1_65));
wire output_3_65, output_3_2, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_2), .y(output_2_65));
wire output_4_65, output_4_2, output_3_65;
mixer gate_output_3_65(.a(output_4_65), .b(output_4_2), .y(output_3_65));
wire output_5_65, output_5_2, output_4_65;
mixer gate_output_4_65(.a(output_5_65), .b(output_5_2), .y(output_4_65));
wire output_6_65, output_6_2, output_5_65;
mixer gate_output_5_65(.a(output_6_65), .b(output_6_2), .y(output_5_65));
wire output_7_65, output_7_2, output_6_65;
mixer gate_output_6_65(.a(output_7_65), .b(output_7_2), .y(output_6_65));
wire output_8_65, output_8_2, output_7_65;
mixer gate_output_7_65(.a(output_8_65), .b(output_8_2), .y(output_7_65));
wire output_1_66, output_1_3, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_3), .y(output_0_66));
wire output_2_66, output_2_3, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_3), .y(output_1_66));
wire output_3_66, output_3_3, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_3), .y(output_2_66));
wire output_4_66, output_4_3, output_3_66;
mixer gate_output_3_66(.a(output_4_66), .b(output_4_3), .y(output_3_66));
wire output_5_66, output_5_3, output_4_66;
mixer gate_output_4_66(.a(output_5_66), .b(output_5_3), .y(output_4_66));
wire output_6_66, output_6_3, output_5_66;
mixer gate_output_5_66(.a(output_6_66), .b(output_6_3), .y(output_5_66));
wire output_7_66, output_7_3, output_6_66;
mixer gate_output_6_66(.a(output_7_66), .b(output_7_3), .y(output_6_66));
wire output_8_66, output_8_3, output_7_66;
mixer gate_output_7_66(.a(output_8_66), .b(output_8_3), .y(output_7_66));
wire output_1_67, output_1_4, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_4), .y(output_0_67));
wire output_2_67, output_2_4, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_4), .y(output_1_67));
wire output_3_67, output_3_4, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_4), .y(output_2_67));
wire output_4_67, output_4_4, output_3_67;
mixer gate_output_3_67(.a(output_4_67), .b(output_4_4), .y(output_3_67));
wire output_5_67, output_5_4, output_4_67;
mixer gate_output_4_67(.a(output_5_67), .b(output_5_4), .y(output_4_67));
wire output_6_67, output_6_4, output_5_67;
mixer gate_output_5_67(.a(output_6_67), .b(output_6_4), .y(output_5_67));
wire output_7_67, output_7_4, output_6_67;
mixer gate_output_6_67(.a(output_7_67), .b(output_7_4), .y(output_6_67));
wire output_8_67, output_8_4, output_7_67;
mixer gate_output_7_67(.a(output_8_67), .b(output_8_4), .y(output_7_67));
wire output_1_68, output_1_5, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_5), .y(output_0_68));
wire output_2_68, output_2_5, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_5), .y(output_1_68));
wire output_3_68, output_3_5, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_5), .y(output_2_68));
wire output_4_68, output_4_5, output_3_68;
mixer gate_output_3_68(.a(output_4_68), .b(output_4_5), .y(output_3_68));
wire output_5_68, output_5_5, output_4_68;
mixer gate_output_4_68(.a(output_5_68), .b(output_5_5), .y(output_4_68));
wire output_6_68, output_6_5, output_5_68;
mixer gate_output_5_68(.a(output_6_68), .b(output_6_5), .y(output_5_68));
wire output_7_68, output_7_5, output_6_68;
mixer gate_output_6_68(.a(output_7_68), .b(output_7_5), .y(output_6_68));
wire output_8_68, output_8_5, output_7_68;
mixer gate_output_7_68(.a(output_8_68), .b(output_8_5), .y(output_7_68));
wire output_1_69, output_1_6, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_6), .y(output_0_69));
wire output_2_69, output_2_6, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_6), .y(output_1_69));
wire output_3_69, output_3_6, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_6), .y(output_2_69));
wire output_4_69, output_4_6, output_3_69;
mixer gate_output_3_69(.a(output_4_69), .b(output_4_6), .y(output_3_69));
wire output_5_69, output_5_6, output_4_69;
mixer gate_output_4_69(.a(output_5_69), .b(output_5_6), .y(output_4_69));
wire output_6_69, output_6_6, output_5_69;
mixer gate_output_5_69(.a(output_6_69), .b(output_6_6), .y(output_5_69));
wire output_7_69, output_7_6, output_6_69;
mixer gate_output_6_69(.a(output_7_69), .b(output_7_6), .y(output_6_69));
wire output_8_69, output_8_6, output_7_69;
mixer gate_output_7_69(.a(output_8_69), .b(output_8_6), .y(output_7_69));
wire output_1_70, output_1_7, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_7), .y(output_0_70));
wire output_2_70, output_2_7, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_7), .y(output_1_70));
wire output_3_70, output_3_7, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_7), .y(output_2_70));
wire output_4_70, output_4_7, output_3_70;
mixer gate_output_3_70(.a(output_4_70), .b(output_4_7), .y(output_3_70));
wire output_5_70, output_5_7, output_4_70;
mixer gate_output_4_70(.a(output_5_70), .b(output_5_7), .y(output_4_70));
wire output_6_70, output_6_7, output_5_70;
mixer gate_output_5_70(.a(output_6_70), .b(output_6_7), .y(output_5_70));
wire output_7_70, output_7_7, output_6_70;
mixer gate_output_6_70(.a(output_7_70), .b(output_7_7), .y(output_6_70));
wire output_8_70, output_8_7, output_7_70;
mixer gate_output_7_70(.a(output_8_70), .b(output_8_7), .y(output_7_70));
wire output_1_71, output_1_0, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_0), .y(output_0_71));
wire output_2_71, output_2_0, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_0), .y(output_1_71));
wire output_3_71, output_3_0, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_0), .y(output_2_71));
wire output_4_71, output_4_0, output_3_71;
mixer gate_output_3_71(.a(output_4_71), .b(output_4_0), .y(output_3_71));
wire output_5_71, output_5_0, output_4_71;
mixer gate_output_4_71(.a(output_5_71), .b(output_5_0), .y(output_4_71));
wire output_6_71, output_6_0, output_5_71;
mixer gate_output_5_71(.a(output_6_71), .b(output_6_0), .y(output_5_71));
wire output_7_71, output_7_0, output_6_71;
mixer gate_output_6_71(.a(output_7_71), .b(output_7_0), .y(output_6_71));
wire output_8_71, output_8_0, output_7_71;
mixer gate_output_7_71(.a(output_8_71), .b(output_8_0), .y(output_7_71));
wire output_1_72, output_1_1, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_1), .y(output_0_72));
wire output_2_72, output_2_1, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_1), .y(output_1_72));
wire output_3_72, output_3_1, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_1), .y(output_2_72));
wire output_4_72, output_4_1, output_3_72;
mixer gate_output_3_72(.a(output_4_72), .b(output_4_1), .y(output_3_72));
wire output_5_72, output_5_1, output_4_72;
mixer gate_output_4_72(.a(output_5_72), .b(output_5_1), .y(output_4_72));
wire output_6_72, output_6_1, output_5_72;
mixer gate_output_5_72(.a(output_6_72), .b(output_6_1), .y(output_5_72));
wire output_7_72, output_7_1, output_6_72;
mixer gate_output_6_72(.a(output_7_72), .b(output_7_1), .y(output_6_72));
wire output_8_72, output_8_1, output_7_72;
mixer gate_output_7_72(.a(output_8_72), .b(output_8_1), .y(output_7_72));
wire output_1_73, output_1_2, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_2), .y(output_0_73));
wire output_2_73, output_2_2, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_2), .y(output_1_73));
wire output_3_73, output_3_2, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_2), .y(output_2_73));
wire output_4_73, output_4_2, output_3_73;
mixer gate_output_3_73(.a(output_4_73), .b(output_4_2), .y(output_3_73));
wire output_5_73, output_5_2, output_4_73;
mixer gate_output_4_73(.a(output_5_73), .b(output_5_2), .y(output_4_73));
wire output_6_73, output_6_2, output_5_73;
mixer gate_output_5_73(.a(output_6_73), .b(output_6_2), .y(output_5_73));
wire output_7_73, output_7_2, output_6_73;
mixer gate_output_6_73(.a(output_7_73), .b(output_7_2), .y(output_6_73));
wire output_8_73, output_8_2, output_7_73;
mixer gate_output_7_73(.a(output_8_73), .b(output_8_2), .y(output_7_73));
wire output_1_74, output_1_3, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_3), .y(output_0_74));
wire output_2_74, output_2_3, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_3), .y(output_1_74));
wire output_3_74, output_3_3, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_3), .y(output_2_74));
wire output_4_74, output_4_3, output_3_74;
mixer gate_output_3_74(.a(output_4_74), .b(output_4_3), .y(output_3_74));
wire output_5_74, output_5_3, output_4_74;
mixer gate_output_4_74(.a(output_5_74), .b(output_5_3), .y(output_4_74));
wire output_6_74, output_6_3, output_5_74;
mixer gate_output_5_74(.a(output_6_74), .b(output_6_3), .y(output_5_74));
wire output_7_74, output_7_3, output_6_74;
mixer gate_output_6_74(.a(output_7_74), .b(output_7_3), .y(output_6_74));
wire output_8_74, output_8_3, output_7_74;
mixer gate_output_7_74(.a(output_8_74), .b(output_8_3), .y(output_7_74));
wire output_1_75, output_1_4, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_4), .y(output_0_75));
wire output_2_75, output_2_4, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_4), .y(output_1_75));
wire output_3_75, output_3_4, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_4), .y(output_2_75));
wire output_4_75, output_4_4, output_3_75;
mixer gate_output_3_75(.a(output_4_75), .b(output_4_4), .y(output_3_75));
wire output_5_75, output_5_4, output_4_75;
mixer gate_output_4_75(.a(output_5_75), .b(output_5_4), .y(output_4_75));
wire output_6_75, output_6_4, output_5_75;
mixer gate_output_5_75(.a(output_6_75), .b(output_6_4), .y(output_5_75));
wire output_7_75, output_7_4, output_6_75;
mixer gate_output_6_75(.a(output_7_75), .b(output_7_4), .y(output_6_75));
wire output_8_75, output_8_4, output_7_75;
mixer gate_output_7_75(.a(output_8_75), .b(output_8_4), .y(output_7_75));
wire output_1_76, output_1_5, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_5), .y(output_0_76));
wire output_2_76, output_2_5, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_5), .y(output_1_76));
wire output_3_76, output_3_5, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_5), .y(output_2_76));
wire output_4_76, output_4_5, output_3_76;
mixer gate_output_3_76(.a(output_4_76), .b(output_4_5), .y(output_3_76));
wire output_5_76, output_5_5, output_4_76;
mixer gate_output_4_76(.a(output_5_76), .b(output_5_5), .y(output_4_76));
wire output_6_76, output_6_5, output_5_76;
mixer gate_output_5_76(.a(output_6_76), .b(output_6_5), .y(output_5_76));
wire output_7_76, output_7_5, output_6_76;
mixer gate_output_6_76(.a(output_7_76), .b(output_7_5), .y(output_6_76));
wire output_8_76, output_8_5, output_7_76;
mixer gate_output_7_76(.a(output_8_76), .b(output_8_5), .y(output_7_76));
wire output_1_77, output_1_6, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_6), .y(output_0_77));
wire output_2_77, output_2_6, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_6), .y(output_1_77));
wire output_3_77, output_3_6, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_6), .y(output_2_77));
wire output_4_77, output_4_6, output_3_77;
mixer gate_output_3_77(.a(output_4_77), .b(output_4_6), .y(output_3_77));
wire output_5_77, output_5_6, output_4_77;
mixer gate_output_4_77(.a(output_5_77), .b(output_5_6), .y(output_4_77));
wire output_6_77, output_6_6, output_5_77;
mixer gate_output_5_77(.a(output_6_77), .b(output_6_6), .y(output_5_77));
wire output_7_77, output_7_6, output_6_77;
mixer gate_output_6_77(.a(output_7_77), .b(output_7_6), .y(output_6_77));
wire output_8_77, output_8_6, output_7_77;
mixer gate_output_7_77(.a(output_8_77), .b(output_8_6), .y(output_7_77));
wire output_1_78, output_1_7, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_7), .y(output_0_78));
wire output_2_78, output_2_7, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_7), .y(output_1_78));
wire output_3_78, output_3_7, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_7), .y(output_2_78));
wire output_4_78, output_4_7, output_3_78;
mixer gate_output_3_78(.a(output_4_78), .b(output_4_7), .y(output_3_78));
wire output_5_78, output_5_7, output_4_78;
mixer gate_output_4_78(.a(output_5_78), .b(output_5_7), .y(output_4_78));
wire output_6_78, output_6_7, output_5_78;
mixer gate_output_5_78(.a(output_6_78), .b(output_6_7), .y(output_5_78));
wire output_7_78, output_7_7, output_6_78;
mixer gate_output_6_78(.a(output_7_78), .b(output_7_7), .y(output_6_78));
wire output_8_78, output_8_7, output_7_78;
mixer gate_output_7_78(.a(output_8_78), .b(output_8_7), .y(output_7_78));
wire output_1_79, output_1_0, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_0), .y(output_0_79));
wire output_2_79, output_2_0, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_0), .y(output_1_79));
wire output_3_79, output_3_0, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_0), .y(output_2_79));
wire output_4_79, output_4_0, output_3_79;
mixer gate_output_3_79(.a(output_4_79), .b(output_4_0), .y(output_3_79));
wire output_5_79, output_5_0, output_4_79;
mixer gate_output_4_79(.a(output_5_79), .b(output_5_0), .y(output_4_79));
wire output_6_79, output_6_0, output_5_79;
mixer gate_output_5_79(.a(output_6_79), .b(output_6_0), .y(output_5_79));
wire output_7_79, output_7_0, output_6_79;
mixer gate_output_6_79(.a(output_7_79), .b(output_7_0), .y(output_6_79));
wire output_8_79, output_8_0, output_7_79;
mixer gate_output_7_79(.a(output_8_79), .b(output_8_0), .y(output_7_79));
wire output_1_80, output_1_1, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_1), .y(output_0_80));
wire output_2_80, output_2_1, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_1), .y(output_1_80));
wire output_3_80, output_3_1, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_1), .y(output_2_80));
wire output_4_80, output_4_1, output_3_80;
mixer gate_output_3_80(.a(output_4_80), .b(output_4_1), .y(output_3_80));
wire output_5_80, output_5_1, output_4_80;
mixer gate_output_4_80(.a(output_5_80), .b(output_5_1), .y(output_4_80));
wire output_6_80, output_6_1, output_5_80;
mixer gate_output_5_80(.a(output_6_80), .b(output_6_1), .y(output_5_80));
wire output_7_80, output_7_1, output_6_80;
mixer gate_output_6_80(.a(output_7_80), .b(output_7_1), .y(output_6_80));
wire output_8_80, output_8_1, output_7_80;
mixer gate_output_7_80(.a(output_8_80), .b(output_8_1), .y(output_7_80));
wire output_1_81, output_1_2, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_2), .y(output_0_81));
wire output_2_81, output_2_2, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_2), .y(output_1_81));
wire output_3_81, output_3_2, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_2), .y(output_2_81));
wire output_4_81, output_4_2, output_3_81;
mixer gate_output_3_81(.a(output_4_81), .b(output_4_2), .y(output_3_81));
wire output_5_81, output_5_2, output_4_81;
mixer gate_output_4_81(.a(output_5_81), .b(output_5_2), .y(output_4_81));
wire output_6_81, output_6_2, output_5_81;
mixer gate_output_5_81(.a(output_6_81), .b(output_6_2), .y(output_5_81));
wire output_7_81, output_7_2, output_6_81;
mixer gate_output_6_81(.a(output_7_81), .b(output_7_2), .y(output_6_81));
wire output_8_81, output_8_2, output_7_81;
mixer gate_output_7_81(.a(output_8_81), .b(output_8_2), .y(output_7_81));
wire output_1_82, output_1_3, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_3), .y(output_0_82));
wire output_2_82, output_2_3, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_3), .y(output_1_82));
wire output_3_82, output_3_3, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_3), .y(output_2_82));
wire output_4_82, output_4_3, output_3_82;
mixer gate_output_3_82(.a(output_4_82), .b(output_4_3), .y(output_3_82));
wire output_5_82, output_5_3, output_4_82;
mixer gate_output_4_82(.a(output_5_82), .b(output_5_3), .y(output_4_82));
wire output_6_82, output_6_3, output_5_82;
mixer gate_output_5_82(.a(output_6_82), .b(output_6_3), .y(output_5_82));
wire output_7_82, output_7_3, output_6_82;
mixer gate_output_6_82(.a(output_7_82), .b(output_7_3), .y(output_6_82));
wire output_8_82, output_8_3, output_7_82;
mixer gate_output_7_82(.a(output_8_82), .b(output_8_3), .y(output_7_82));
wire output_1_83, output_1_4, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_4), .y(output_0_83));
wire output_2_83, output_2_4, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_4), .y(output_1_83));
wire output_3_83, output_3_4, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_4), .y(output_2_83));
wire output_4_83, output_4_4, output_3_83;
mixer gate_output_3_83(.a(output_4_83), .b(output_4_4), .y(output_3_83));
wire output_5_83, output_5_4, output_4_83;
mixer gate_output_4_83(.a(output_5_83), .b(output_5_4), .y(output_4_83));
wire output_6_83, output_6_4, output_5_83;
mixer gate_output_5_83(.a(output_6_83), .b(output_6_4), .y(output_5_83));
wire output_7_83, output_7_4, output_6_83;
mixer gate_output_6_83(.a(output_7_83), .b(output_7_4), .y(output_6_83));
wire output_8_83, output_8_4, output_7_83;
mixer gate_output_7_83(.a(output_8_83), .b(output_8_4), .y(output_7_83));
wire output_1_84, output_1_5, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_5), .y(output_0_84));
wire output_2_84, output_2_5, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_5), .y(output_1_84));
wire output_3_84, output_3_5, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_5), .y(output_2_84));
wire output_4_84, output_4_5, output_3_84;
mixer gate_output_3_84(.a(output_4_84), .b(output_4_5), .y(output_3_84));
wire output_5_84, output_5_5, output_4_84;
mixer gate_output_4_84(.a(output_5_84), .b(output_5_5), .y(output_4_84));
wire output_6_84, output_6_5, output_5_84;
mixer gate_output_5_84(.a(output_6_84), .b(output_6_5), .y(output_5_84));
wire output_7_84, output_7_5, output_6_84;
mixer gate_output_6_84(.a(output_7_84), .b(output_7_5), .y(output_6_84));
wire output_8_84, output_8_5, output_7_84;
mixer gate_output_7_84(.a(output_8_84), .b(output_8_5), .y(output_7_84));
wire output_1_85, output_1_6, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_6), .y(output_0_85));
wire output_2_85, output_2_6, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_6), .y(output_1_85));
wire output_3_85, output_3_6, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_6), .y(output_2_85));
wire output_4_85, output_4_6, output_3_85;
mixer gate_output_3_85(.a(output_4_85), .b(output_4_6), .y(output_3_85));
wire output_5_85, output_5_6, output_4_85;
mixer gate_output_4_85(.a(output_5_85), .b(output_5_6), .y(output_4_85));
wire output_6_85, output_6_6, output_5_85;
mixer gate_output_5_85(.a(output_6_85), .b(output_6_6), .y(output_5_85));
wire output_7_85, output_7_6, output_6_85;
mixer gate_output_6_85(.a(output_7_85), .b(output_7_6), .y(output_6_85));
wire output_8_85, output_8_6, output_7_85;
mixer gate_output_7_85(.a(output_8_85), .b(output_8_6), .y(output_7_85));
wire output_1_86, output_1_7, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_7), .y(output_0_86));
wire output_2_86, output_2_7, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_7), .y(output_1_86));
wire output_3_86, output_3_7, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_7), .y(output_2_86));
wire output_4_86, output_4_7, output_3_86;
mixer gate_output_3_86(.a(output_4_86), .b(output_4_7), .y(output_3_86));
wire output_5_86, output_5_7, output_4_86;
mixer gate_output_4_86(.a(output_5_86), .b(output_5_7), .y(output_4_86));
wire output_6_86, output_6_7, output_5_86;
mixer gate_output_5_86(.a(output_6_86), .b(output_6_7), .y(output_5_86));
wire output_7_86, output_7_7, output_6_86;
mixer gate_output_6_86(.a(output_7_86), .b(output_7_7), .y(output_6_86));
wire output_8_86, output_8_7, output_7_86;
mixer gate_output_7_86(.a(output_8_86), .b(output_8_7), .y(output_7_86));
wire output_1_87, output_1_0, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_0), .y(output_0_87));
wire output_2_87, output_2_0, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_0), .y(output_1_87));
wire output_3_87, output_3_0, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_0), .y(output_2_87));
wire output_4_87, output_4_0, output_3_87;
mixer gate_output_3_87(.a(output_4_87), .b(output_4_0), .y(output_3_87));
wire output_5_87, output_5_0, output_4_87;
mixer gate_output_4_87(.a(output_5_87), .b(output_5_0), .y(output_4_87));
wire output_6_87, output_6_0, output_5_87;
mixer gate_output_5_87(.a(output_6_87), .b(output_6_0), .y(output_5_87));
wire output_7_87, output_7_0, output_6_87;
mixer gate_output_6_87(.a(output_7_87), .b(output_7_0), .y(output_6_87));
wire output_8_87, output_8_0, output_7_87;
mixer gate_output_7_87(.a(output_8_87), .b(output_8_0), .y(output_7_87));
wire output_1_88, output_1_1, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_1), .y(output_0_88));
wire output_2_88, output_2_1, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_1), .y(output_1_88));
wire output_3_88, output_3_1, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_1), .y(output_2_88));
wire output_4_88, output_4_1, output_3_88;
mixer gate_output_3_88(.a(output_4_88), .b(output_4_1), .y(output_3_88));
wire output_5_88, output_5_1, output_4_88;
mixer gate_output_4_88(.a(output_5_88), .b(output_5_1), .y(output_4_88));
wire output_6_88, output_6_1, output_5_88;
mixer gate_output_5_88(.a(output_6_88), .b(output_6_1), .y(output_5_88));
wire output_7_88, output_7_1, output_6_88;
mixer gate_output_6_88(.a(output_7_88), .b(output_7_1), .y(output_6_88));
wire output_8_88, output_8_1, output_7_88;
mixer gate_output_7_88(.a(output_8_88), .b(output_8_1), .y(output_7_88));
wire output_1_89, output_1_2, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_2), .y(output_0_89));
wire output_2_89, output_2_2, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_2), .y(output_1_89));
wire output_3_89, output_3_2, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_2), .y(output_2_89));
wire output_4_89, output_4_2, output_3_89;
mixer gate_output_3_89(.a(output_4_89), .b(output_4_2), .y(output_3_89));
wire output_5_89, output_5_2, output_4_89;
mixer gate_output_4_89(.a(output_5_89), .b(output_5_2), .y(output_4_89));
wire output_6_89, output_6_2, output_5_89;
mixer gate_output_5_89(.a(output_6_89), .b(output_6_2), .y(output_5_89));
wire output_7_89, output_7_2, output_6_89;
mixer gate_output_6_89(.a(output_7_89), .b(output_7_2), .y(output_6_89));
wire output_8_89, output_8_2, output_7_89;
mixer gate_output_7_89(.a(output_8_89), .b(output_8_2), .y(output_7_89));
wire output_1_90, output_1_3, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_3), .y(output_0_90));
wire output_2_90, output_2_3, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_3), .y(output_1_90));
wire output_3_90, output_3_3, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_3), .y(output_2_90));
wire output_4_90, output_4_3, output_3_90;
mixer gate_output_3_90(.a(output_4_90), .b(output_4_3), .y(output_3_90));
wire output_5_90, output_5_3, output_4_90;
mixer gate_output_4_90(.a(output_5_90), .b(output_5_3), .y(output_4_90));
wire output_6_90, output_6_3, output_5_90;
mixer gate_output_5_90(.a(output_6_90), .b(output_6_3), .y(output_5_90));
wire output_7_90, output_7_3, output_6_90;
mixer gate_output_6_90(.a(output_7_90), .b(output_7_3), .y(output_6_90));
wire output_8_90, output_8_3, output_7_90;
mixer gate_output_7_90(.a(output_8_90), .b(output_8_3), .y(output_7_90));
wire output_1_91, output_1_4, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_4), .y(output_0_91));
wire output_2_91, output_2_4, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_4), .y(output_1_91));
wire output_3_91, output_3_4, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_4), .y(output_2_91));
wire output_4_91, output_4_4, output_3_91;
mixer gate_output_3_91(.a(output_4_91), .b(output_4_4), .y(output_3_91));
wire output_5_91, output_5_4, output_4_91;
mixer gate_output_4_91(.a(output_5_91), .b(output_5_4), .y(output_4_91));
wire output_6_91, output_6_4, output_5_91;
mixer gate_output_5_91(.a(output_6_91), .b(output_6_4), .y(output_5_91));
wire output_7_91, output_7_4, output_6_91;
mixer gate_output_6_91(.a(output_7_91), .b(output_7_4), .y(output_6_91));
wire output_8_91, output_8_4, output_7_91;
mixer gate_output_7_91(.a(output_8_91), .b(output_8_4), .y(output_7_91));
wire output_1_92, output_1_5, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_5), .y(output_0_92));
wire output_2_92, output_2_5, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_5), .y(output_1_92));
wire output_3_92, output_3_5, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_5), .y(output_2_92));
wire output_4_92, output_4_5, output_3_92;
mixer gate_output_3_92(.a(output_4_92), .b(output_4_5), .y(output_3_92));
wire output_5_92, output_5_5, output_4_92;
mixer gate_output_4_92(.a(output_5_92), .b(output_5_5), .y(output_4_92));
wire output_6_92, output_6_5, output_5_92;
mixer gate_output_5_92(.a(output_6_92), .b(output_6_5), .y(output_5_92));
wire output_7_92, output_7_5, output_6_92;
mixer gate_output_6_92(.a(output_7_92), .b(output_7_5), .y(output_6_92));
wire output_8_92, output_8_5, output_7_92;
mixer gate_output_7_92(.a(output_8_92), .b(output_8_5), .y(output_7_92));
wire output_1_93, output_1_6, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_6), .y(output_0_93));
wire output_2_93, output_2_6, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_6), .y(output_1_93));
wire output_3_93, output_3_6, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_6), .y(output_2_93));
wire output_4_93, output_4_6, output_3_93;
mixer gate_output_3_93(.a(output_4_93), .b(output_4_6), .y(output_3_93));
wire output_5_93, output_5_6, output_4_93;
mixer gate_output_4_93(.a(output_5_93), .b(output_5_6), .y(output_4_93));
wire output_6_93, output_6_6, output_5_93;
mixer gate_output_5_93(.a(output_6_93), .b(output_6_6), .y(output_5_93));
wire output_7_93, output_7_6, output_6_93;
mixer gate_output_6_93(.a(output_7_93), .b(output_7_6), .y(output_6_93));
wire output_8_93, output_8_6, output_7_93;
mixer gate_output_7_93(.a(output_8_93), .b(output_8_6), .y(output_7_93));
wire output_1_94, output_1_7, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_7), .y(output_0_94));
wire output_2_94, output_2_7, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_7), .y(output_1_94));
wire output_3_94, output_3_7, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_7), .y(output_2_94));
wire output_4_94, output_4_7, output_3_94;
mixer gate_output_3_94(.a(output_4_94), .b(output_4_7), .y(output_3_94));
wire output_5_94, output_5_7, output_4_94;
mixer gate_output_4_94(.a(output_5_94), .b(output_5_7), .y(output_4_94));
wire output_6_94, output_6_7, output_5_94;
mixer gate_output_5_94(.a(output_6_94), .b(output_6_7), .y(output_5_94));
wire output_7_94, output_7_7, output_6_94;
mixer gate_output_6_94(.a(output_7_94), .b(output_7_7), .y(output_6_94));
wire output_8_94, output_8_7, output_7_94;
mixer gate_output_7_94(.a(output_8_94), .b(output_8_7), .y(output_7_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_4_95, output_4_0, output_3_95;
mixer gate_output_3_95(.a(output_4_95), .b(output_4_0), .y(output_3_95));
wire output_5_95, output_5_0, output_4_95;
mixer gate_output_4_95(.a(output_5_95), .b(output_5_0), .y(output_4_95));
wire output_6_95, output_6_0, output_5_95;
mixer gate_output_5_95(.a(output_6_95), .b(output_6_0), .y(output_5_95));
wire output_7_95, output_7_0, output_6_95;
mixer gate_output_6_95(.a(output_7_95), .b(output_7_0), .y(output_6_95));
wire output_8_95, output_8_0, output_7_95;
mixer gate_output_7_95(.a(output_8_95), .b(output_8_0), .y(output_7_95));
assign output_0 = output_0_0;
wire output_0_96;
assign output_0_96 = input_0;
assign output_1 = output_1_0;
wire output_1_96;
assign output_1_96 = input_1;
assign output_2 = output_2_0;
wire output_2_96;
assign output_2_96 = input_2;
assign output_3 = output_3_0;
wire output_3_96;
assign output_3_96 = input_3;
assign output_4 = output_4_0;
wire output_4_96;
assign output_4_96 = input_4;
assign output_5 = output_5_0;
wire output_5_96;
assign output_5_96 = input_5;
assign output_6 = output_6_0;
wire output_6_96;
assign output_6_96 = input_6;
assign output_7 = output_7_0;
wire output_7_96;
assign output_7_96 = input_7;
endmodule
