module chain_16 (
inout k0, k16
);
wire {wires};
chamber ch0 (.in(k0), .out(k1)
chamber ch1 (.in(k1), .out(k2)
chamber ch2 (.in(k2), .out(k3)
chamber ch3 (.in(k3), .out(k4)
chamber ch4 (.in(k4), .out(k5)
chamber ch5 (.in(k5), .out(k6)
chamber ch6 (.in(k6), .out(k7)
chamber ch7 (.in(k7), .out(k8)
chamber ch8 (.in(k8), .out(k9)
chamber ch9 (.in(k9), .out(k10)
chamber ch10 (.in(k10), .out(k11)
chamber ch11 (.in(k11), .out(k12)
chamber ch12 (.in(k12), .out(k13)
chamber ch13 (.in(k13), .out(k14)
chamber ch14 (.in(k14), .out(k15)
chamber ch15 (.in(k15), .out(k16)
endmodule
