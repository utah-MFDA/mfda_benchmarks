module complete_bipartite_32_32 (
inout input_0,inout input_1,inout input_2,inout input_3,inout input_4,inout input_5,inout input_6,inout input_7,inout input_8,inout input_9,inout input_10,inout input_11,inout input_12,inout input_13,inout input_14,inout input_15,inout input_16,inout input_17,inout input_18,inout input_19,inout input_20,inout input_21,inout input_22,inout input_23,inout input_24,inout input_25,inout input_26,inout input_27,inout input_28,inout input_29,inout input_30,inout input_31,inout output_0,inout output_1,inout output_2,inout output_3,inout output_4,inout output_5,inout output_6,inout output_7,inout output_8,inout output_9,inout output_10,inout output_11,inout output_12,inout output_13,inout output_14,inout output_15,inout output_16,inout output_17,inout output_18,inout output_19,inout output_20,inout output_21,inout output_22,inout output_23,inout output_24,inout output_25,inout output_26,inout output_27,inout output_28,inout output_29,inout output_30,inout output_31
);
assign output_0 = input_0;
assign output_1 = input_0;
assign output_2 = input_0;
assign output_3 = input_0;
assign output_4 = input_0;
assign output_5 = input_0;
assign output_6 = input_0;
assign output_7 = input_0;
assign output_8 = input_0;
assign output_9 = input_0;
assign output_10 = input_0;
assign output_11 = input_0;
assign output_12 = input_0;
assign output_13 = input_0;
assign output_14 = input_0;
assign output_15 = input_0;
assign output_16 = input_0;
assign output_17 = input_0;
assign output_18 = input_0;
assign output_19 = input_0;
assign output_20 = input_0;
assign output_21 = input_0;
assign output_22 = input_0;
assign output_23 = input_0;
assign output_24 = input_0;
assign output_25 = input_0;
assign output_26 = input_0;
assign output_27 = input_0;
assign output_28 = input_0;
assign output_29 = input_0;
assign output_30 = input_0;
assign output_31 = input_0;
assign output_0 = input_1;
assign output_1 = input_1;
assign output_2 = input_1;
assign output_3 = input_1;
assign output_4 = input_1;
assign output_5 = input_1;
assign output_6 = input_1;
assign output_7 = input_1;
assign output_8 = input_1;
assign output_9 = input_1;
assign output_10 = input_1;
assign output_11 = input_1;
assign output_12 = input_1;
assign output_13 = input_1;
assign output_14 = input_1;
assign output_15 = input_1;
assign output_16 = input_1;
assign output_17 = input_1;
assign output_18 = input_1;
assign output_19 = input_1;
assign output_20 = input_1;
assign output_21 = input_1;
assign output_22 = input_1;
assign output_23 = input_1;
assign output_24 = input_1;
assign output_25 = input_1;
assign output_26 = input_1;
assign output_27 = input_1;
assign output_28 = input_1;
assign output_29 = input_1;
assign output_30 = input_1;
assign output_31 = input_1;
assign output_0 = input_2;
assign output_1 = input_2;
assign output_2 = input_2;
assign output_3 = input_2;
assign output_4 = input_2;
assign output_5 = input_2;
assign output_6 = input_2;
assign output_7 = input_2;
assign output_8 = input_2;
assign output_9 = input_2;
assign output_10 = input_2;
assign output_11 = input_2;
assign output_12 = input_2;
assign output_13 = input_2;
assign output_14 = input_2;
assign output_15 = input_2;
assign output_16 = input_2;
assign output_17 = input_2;
assign output_18 = input_2;
assign output_19 = input_2;
assign output_20 = input_2;
assign output_21 = input_2;
assign output_22 = input_2;
assign output_23 = input_2;
assign output_24 = input_2;
assign output_25 = input_2;
assign output_26 = input_2;
assign output_27 = input_2;
assign output_28 = input_2;
assign output_29 = input_2;
assign output_30 = input_2;
assign output_31 = input_2;
assign output_0 = input_3;
assign output_1 = input_3;
assign output_2 = input_3;
assign output_3 = input_3;
assign output_4 = input_3;
assign output_5 = input_3;
assign output_6 = input_3;
assign output_7 = input_3;
assign output_8 = input_3;
assign output_9 = input_3;
assign output_10 = input_3;
assign output_11 = input_3;
assign output_12 = input_3;
assign output_13 = input_3;
assign output_14 = input_3;
assign output_15 = input_3;
assign output_16 = input_3;
assign output_17 = input_3;
assign output_18 = input_3;
assign output_19 = input_3;
assign output_20 = input_3;
assign output_21 = input_3;
assign output_22 = input_3;
assign output_23 = input_3;
assign output_24 = input_3;
assign output_25 = input_3;
assign output_26 = input_3;
assign output_27 = input_3;
assign output_28 = input_3;
assign output_29 = input_3;
assign output_30 = input_3;
assign output_31 = input_3;
assign output_0 = input_4;
assign output_1 = input_4;
assign output_2 = input_4;
assign output_3 = input_4;
assign output_4 = input_4;
assign output_5 = input_4;
assign output_6 = input_4;
assign output_7 = input_4;
assign output_8 = input_4;
assign output_9 = input_4;
assign output_10 = input_4;
assign output_11 = input_4;
assign output_12 = input_4;
assign output_13 = input_4;
assign output_14 = input_4;
assign output_15 = input_4;
assign output_16 = input_4;
assign output_17 = input_4;
assign output_18 = input_4;
assign output_19 = input_4;
assign output_20 = input_4;
assign output_21 = input_4;
assign output_22 = input_4;
assign output_23 = input_4;
assign output_24 = input_4;
assign output_25 = input_4;
assign output_26 = input_4;
assign output_27 = input_4;
assign output_28 = input_4;
assign output_29 = input_4;
assign output_30 = input_4;
assign output_31 = input_4;
assign output_0 = input_5;
assign output_1 = input_5;
assign output_2 = input_5;
assign output_3 = input_5;
assign output_4 = input_5;
assign output_5 = input_5;
assign output_6 = input_5;
assign output_7 = input_5;
assign output_8 = input_5;
assign output_9 = input_5;
assign output_10 = input_5;
assign output_11 = input_5;
assign output_12 = input_5;
assign output_13 = input_5;
assign output_14 = input_5;
assign output_15 = input_5;
assign output_16 = input_5;
assign output_17 = input_5;
assign output_18 = input_5;
assign output_19 = input_5;
assign output_20 = input_5;
assign output_21 = input_5;
assign output_22 = input_5;
assign output_23 = input_5;
assign output_24 = input_5;
assign output_25 = input_5;
assign output_26 = input_5;
assign output_27 = input_5;
assign output_28 = input_5;
assign output_29 = input_5;
assign output_30 = input_5;
assign output_31 = input_5;
assign output_0 = input_6;
assign output_1 = input_6;
assign output_2 = input_6;
assign output_3 = input_6;
assign output_4 = input_6;
assign output_5 = input_6;
assign output_6 = input_6;
assign output_7 = input_6;
assign output_8 = input_6;
assign output_9 = input_6;
assign output_10 = input_6;
assign output_11 = input_6;
assign output_12 = input_6;
assign output_13 = input_6;
assign output_14 = input_6;
assign output_15 = input_6;
assign output_16 = input_6;
assign output_17 = input_6;
assign output_18 = input_6;
assign output_19 = input_6;
assign output_20 = input_6;
assign output_21 = input_6;
assign output_22 = input_6;
assign output_23 = input_6;
assign output_24 = input_6;
assign output_25 = input_6;
assign output_26 = input_6;
assign output_27 = input_6;
assign output_28 = input_6;
assign output_29 = input_6;
assign output_30 = input_6;
assign output_31 = input_6;
assign output_0 = input_7;
assign output_1 = input_7;
assign output_2 = input_7;
assign output_3 = input_7;
assign output_4 = input_7;
assign output_5 = input_7;
assign output_6 = input_7;
assign output_7 = input_7;
assign output_8 = input_7;
assign output_9 = input_7;
assign output_10 = input_7;
assign output_11 = input_7;
assign output_12 = input_7;
assign output_13 = input_7;
assign output_14 = input_7;
assign output_15 = input_7;
assign output_16 = input_7;
assign output_17 = input_7;
assign output_18 = input_7;
assign output_19 = input_7;
assign output_20 = input_7;
assign output_21 = input_7;
assign output_22 = input_7;
assign output_23 = input_7;
assign output_24 = input_7;
assign output_25 = input_7;
assign output_26 = input_7;
assign output_27 = input_7;
assign output_28 = input_7;
assign output_29 = input_7;
assign output_30 = input_7;
assign output_31 = input_7;
assign output_0 = input_8;
assign output_1 = input_8;
assign output_2 = input_8;
assign output_3 = input_8;
assign output_4 = input_8;
assign output_5 = input_8;
assign output_6 = input_8;
assign output_7 = input_8;
assign output_8 = input_8;
assign output_9 = input_8;
assign output_10 = input_8;
assign output_11 = input_8;
assign output_12 = input_8;
assign output_13 = input_8;
assign output_14 = input_8;
assign output_15 = input_8;
assign output_16 = input_8;
assign output_17 = input_8;
assign output_18 = input_8;
assign output_19 = input_8;
assign output_20 = input_8;
assign output_21 = input_8;
assign output_22 = input_8;
assign output_23 = input_8;
assign output_24 = input_8;
assign output_25 = input_8;
assign output_26 = input_8;
assign output_27 = input_8;
assign output_28 = input_8;
assign output_29 = input_8;
assign output_30 = input_8;
assign output_31 = input_8;
assign output_0 = input_9;
assign output_1 = input_9;
assign output_2 = input_9;
assign output_3 = input_9;
assign output_4 = input_9;
assign output_5 = input_9;
assign output_6 = input_9;
assign output_7 = input_9;
assign output_8 = input_9;
assign output_9 = input_9;
assign output_10 = input_9;
assign output_11 = input_9;
assign output_12 = input_9;
assign output_13 = input_9;
assign output_14 = input_9;
assign output_15 = input_9;
assign output_16 = input_9;
assign output_17 = input_9;
assign output_18 = input_9;
assign output_19 = input_9;
assign output_20 = input_9;
assign output_21 = input_9;
assign output_22 = input_9;
assign output_23 = input_9;
assign output_24 = input_9;
assign output_25 = input_9;
assign output_26 = input_9;
assign output_27 = input_9;
assign output_28 = input_9;
assign output_29 = input_9;
assign output_30 = input_9;
assign output_31 = input_9;
assign output_0 = input_10;
assign output_1 = input_10;
assign output_2 = input_10;
assign output_3 = input_10;
assign output_4 = input_10;
assign output_5 = input_10;
assign output_6 = input_10;
assign output_7 = input_10;
assign output_8 = input_10;
assign output_9 = input_10;
assign output_10 = input_10;
assign output_11 = input_10;
assign output_12 = input_10;
assign output_13 = input_10;
assign output_14 = input_10;
assign output_15 = input_10;
assign output_16 = input_10;
assign output_17 = input_10;
assign output_18 = input_10;
assign output_19 = input_10;
assign output_20 = input_10;
assign output_21 = input_10;
assign output_22 = input_10;
assign output_23 = input_10;
assign output_24 = input_10;
assign output_25 = input_10;
assign output_26 = input_10;
assign output_27 = input_10;
assign output_28 = input_10;
assign output_29 = input_10;
assign output_30 = input_10;
assign output_31 = input_10;
assign output_0 = input_11;
assign output_1 = input_11;
assign output_2 = input_11;
assign output_3 = input_11;
assign output_4 = input_11;
assign output_5 = input_11;
assign output_6 = input_11;
assign output_7 = input_11;
assign output_8 = input_11;
assign output_9 = input_11;
assign output_10 = input_11;
assign output_11 = input_11;
assign output_12 = input_11;
assign output_13 = input_11;
assign output_14 = input_11;
assign output_15 = input_11;
assign output_16 = input_11;
assign output_17 = input_11;
assign output_18 = input_11;
assign output_19 = input_11;
assign output_20 = input_11;
assign output_21 = input_11;
assign output_22 = input_11;
assign output_23 = input_11;
assign output_24 = input_11;
assign output_25 = input_11;
assign output_26 = input_11;
assign output_27 = input_11;
assign output_28 = input_11;
assign output_29 = input_11;
assign output_30 = input_11;
assign output_31 = input_11;
assign output_0 = input_12;
assign output_1 = input_12;
assign output_2 = input_12;
assign output_3 = input_12;
assign output_4 = input_12;
assign output_5 = input_12;
assign output_6 = input_12;
assign output_7 = input_12;
assign output_8 = input_12;
assign output_9 = input_12;
assign output_10 = input_12;
assign output_11 = input_12;
assign output_12 = input_12;
assign output_13 = input_12;
assign output_14 = input_12;
assign output_15 = input_12;
assign output_16 = input_12;
assign output_17 = input_12;
assign output_18 = input_12;
assign output_19 = input_12;
assign output_20 = input_12;
assign output_21 = input_12;
assign output_22 = input_12;
assign output_23 = input_12;
assign output_24 = input_12;
assign output_25 = input_12;
assign output_26 = input_12;
assign output_27 = input_12;
assign output_28 = input_12;
assign output_29 = input_12;
assign output_30 = input_12;
assign output_31 = input_12;
assign output_0 = input_13;
assign output_1 = input_13;
assign output_2 = input_13;
assign output_3 = input_13;
assign output_4 = input_13;
assign output_5 = input_13;
assign output_6 = input_13;
assign output_7 = input_13;
assign output_8 = input_13;
assign output_9 = input_13;
assign output_10 = input_13;
assign output_11 = input_13;
assign output_12 = input_13;
assign output_13 = input_13;
assign output_14 = input_13;
assign output_15 = input_13;
assign output_16 = input_13;
assign output_17 = input_13;
assign output_18 = input_13;
assign output_19 = input_13;
assign output_20 = input_13;
assign output_21 = input_13;
assign output_22 = input_13;
assign output_23 = input_13;
assign output_24 = input_13;
assign output_25 = input_13;
assign output_26 = input_13;
assign output_27 = input_13;
assign output_28 = input_13;
assign output_29 = input_13;
assign output_30 = input_13;
assign output_31 = input_13;
assign output_0 = input_14;
assign output_1 = input_14;
assign output_2 = input_14;
assign output_3 = input_14;
assign output_4 = input_14;
assign output_5 = input_14;
assign output_6 = input_14;
assign output_7 = input_14;
assign output_8 = input_14;
assign output_9 = input_14;
assign output_10 = input_14;
assign output_11 = input_14;
assign output_12 = input_14;
assign output_13 = input_14;
assign output_14 = input_14;
assign output_15 = input_14;
assign output_16 = input_14;
assign output_17 = input_14;
assign output_18 = input_14;
assign output_19 = input_14;
assign output_20 = input_14;
assign output_21 = input_14;
assign output_22 = input_14;
assign output_23 = input_14;
assign output_24 = input_14;
assign output_25 = input_14;
assign output_26 = input_14;
assign output_27 = input_14;
assign output_28 = input_14;
assign output_29 = input_14;
assign output_30 = input_14;
assign output_31 = input_14;
assign output_0 = input_15;
assign output_1 = input_15;
assign output_2 = input_15;
assign output_3 = input_15;
assign output_4 = input_15;
assign output_5 = input_15;
assign output_6 = input_15;
assign output_7 = input_15;
assign output_8 = input_15;
assign output_9 = input_15;
assign output_10 = input_15;
assign output_11 = input_15;
assign output_12 = input_15;
assign output_13 = input_15;
assign output_14 = input_15;
assign output_15 = input_15;
assign output_16 = input_15;
assign output_17 = input_15;
assign output_18 = input_15;
assign output_19 = input_15;
assign output_20 = input_15;
assign output_21 = input_15;
assign output_22 = input_15;
assign output_23 = input_15;
assign output_24 = input_15;
assign output_25 = input_15;
assign output_26 = input_15;
assign output_27 = input_15;
assign output_28 = input_15;
assign output_29 = input_15;
assign output_30 = input_15;
assign output_31 = input_15;
assign output_0 = input_16;
assign output_1 = input_16;
assign output_2 = input_16;
assign output_3 = input_16;
assign output_4 = input_16;
assign output_5 = input_16;
assign output_6 = input_16;
assign output_7 = input_16;
assign output_8 = input_16;
assign output_9 = input_16;
assign output_10 = input_16;
assign output_11 = input_16;
assign output_12 = input_16;
assign output_13 = input_16;
assign output_14 = input_16;
assign output_15 = input_16;
assign output_16 = input_16;
assign output_17 = input_16;
assign output_18 = input_16;
assign output_19 = input_16;
assign output_20 = input_16;
assign output_21 = input_16;
assign output_22 = input_16;
assign output_23 = input_16;
assign output_24 = input_16;
assign output_25 = input_16;
assign output_26 = input_16;
assign output_27 = input_16;
assign output_28 = input_16;
assign output_29 = input_16;
assign output_30 = input_16;
assign output_31 = input_16;
assign output_0 = input_17;
assign output_1 = input_17;
assign output_2 = input_17;
assign output_3 = input_17;
assign output_4 = input_17;
assign output_5 = input_17;
assign output_6 = input_17;
assign output_7 = input_17;
assign output_8 = input_17;
assign output_9 = input_17;
assign output_10 = input_17;
assign output_11 = input_17;
assign output_12 = input_17;
assign output_13 = input_17;
assign output_14 = input_17;
assign output_15 = input_17;
assign output_16 = input_17;
assign output_17 = input_17;
assign output_18 = input_17;
assign output_19 = input_17;
assign output_20 = input_17;
assign output_21 = input_17;
assign output_22 = input_17;
assign output_23 = input_17;
assign output_24 = input_17;
assign output_25 = input_17;
assign output_26 = input_17;
assign output_27 = input_17;
assign output_28 = input_17;
assign output_29 = input_17;
assign output_30 = input_17;
assign output_31 = input_17;
assign output_0 = input_18;
assign output_1 = input_18;
assign output_2 = input_18;
assign output_3 = input_18;
assign output_4 = input_18;
assign output_5 = input_18;
assign output_6 = input_18;
assign output_7 = input_18;
assign output_8 = input_18;
assign output_9 = input_18;
assign output_10 = input_18;
assign output_11 = input_18;
assign output_12 = input_18;
assign output_13 = input_18;
assign output_14 = input_18;
assign output_15 = input_18;
assign output_16 = input_18;
assign output_17 = input_18;
assign output_18 = input_18;
assign output_19 = input_18;
assign output_20 = input_18;
assign output_21 = input_18;
assign output_22 = input_18;
assign output_23 = input_18;
assign output_24 = input_18;
assign output_25 = input_18;
assign output_26 = input_18;
assign output_27 = input_18;
assign output_28 = input_18;
assign output_29 = input_18;
assign output_30 = input_18;
assign output_31 = input_18;
assign output_0 = input_19;
assign output_1 = input_19;
assign output_2 = input_19;
assign output_3 = input_19;
assign output_4 = input_19;
assign output_5 = input_19;
assign output_6 = input_19;
assign output_7 = input_19;
assign output_8 = input_19;
assign output_9 = input_19;
assign output_10 = input_19;
assign output_11 = input_19;
assign output_12 = input_19;
assign output_13 = input_19;
assign output_14 = input_19;
assign output_15 = input_19;
assign output_16 = input_19;
assign output_17 = input_19;
assign output_18 = input_19;
assign output_19 = input_19;
assign output_20 = input_19;
assign output_21 = input_19;
assign output_22 = input_19;
assign output_23 = input_19;
assign output_24 = input_19;
assign output_25 = input_19;
assign output_26 = input_19;
assign output_27 = input_19;
assign output_28 = input_19;
assign output_29 = input_19;
assign output_30 = input_19;
assign output_31 = input_19;
assign output_0 = input_20;
assign output_1 = input_20;
assign output_2 = input_20;
assign output_3 = input_20;
assign output_4 = input_20;
assign output_5 = input_20;
assign output_6 = input_20;
assign output_7 = input_20;
assign output_8 = input_20;
assign output_9 = input_20;
assign output_10 = input_20;
assign output_11 = input_20;
assign output_12 = input_20;
assign output_13 = input_20;
assign output_14 = input_20;
assign output_15 = input_20;
assign output_16 = input_20;
assign output_17 = input_20;
assign output_18 = input_20;
assign output_19 = input_20;
assign output_20 = input_20;
assign output_21 = input_20;
assign output_22 = input_20;
assign output_23 = input_20;
assign output_24 = input_20;
assign output_25 = input_20;
assign output_26 = input_20;
assign output_27 = input_20;
assign output_28 = input_20;
assign output_29 = input_20;
assign output_30 = input_20;
assign output_31 = input_20;
assign output_0 = input_21;
assign output_1 = input_21;
assign output_2 = input_21;
assign output_3 = input_21;
assign output_4 = input_21;
assign output_5 = input_21;
assign output_6 = input_21;
assign output_7 = input_21;
assign output_8 = input_21;
assign output_9 = input_21;
assign output_10 = input_21;
assign output_11 = input_21;
assign output_12 = input_21;
assign output_13 = input_21;
assign output_14 = input_21;
assign output_15 = input_21;
assign output_16 = input_21;
assign output_17 = input_21;
assign output_18 = input_21;
assign output_19 = input_21;
assign output_20 = input_21;
assign output_21 = input_21;
assign output_22 = input_21;
assign output_23 = input_21;
assign output_24 = input_21;
assign output_25 = input_21;
assign output_26 = input_21;
assign output_27 = input_21;
assign output_28 = input_21;
assign output_29 = input_21;
assign output_30 = input_21;
assign output_31 = input_21;
assign output_0 = input_22;
assign output_1 = input_22;
assign output_2 = input_22;
assign output_3 = input_22;
assign output_4 = input_22;
assign output_5 = input_22;
assign output_6 = input_22;
assign output_7 = input_22;
assign output_8 = input_22;
assign output_9 = input_22;
assign output_10 = input_22;
assign output_11 = input_22;
assign output_12 = input_22;
assign output_13 = input_22;
assign output_14 = input_22;
assign output_15 = input_22;
assign output_16 = input_22;
assign output_17 = input_22;
assign output_18 = input_22;
assign output_19 = input_22;
assign output_20 = input_22;
assign output_21 = input_22;
assign output_22 = input_22;
assign output_23 = input_22;
assign output_24 = input_22;
assign output_25 = input_22;
assign output_26 = input_22;
assign output_27 = input_22;
assign output_28 = input_22;
assign output_29 = input_22;
assign output_30 = input_22;
assign output_31 = input_22;
assign output_0 = input_23;
assign output_1 = input_23;
assign output_2 = input_23;
assign output_3 = input_23;
assign output_4 = input_23;
assign output_5 = input_23;
assign output_6 = input_23;
assign output_7 = input_23;
assign output_8 = input_23;
assign output_9 = input_23;
assign output_10 = input_23;
assign output_11 = input_23;
assign output_12 = input_23;
assign output_13 = input_23;
assign output_14 = input_23;
assign output_15 = input_23;
assign output_16 = input_23;
assign output_17 = input_23;
assign output_18 = input_23;
assign output_19 = input_23;
assign output_20 = input_23;
assign output_21 = input_23;
assign output_22 = input_23;
assign output_23 = input_23;
assign output_24 = input_23;
assign output_25 = input_23;
assign output_26 = input_23;
assign output_27 = input_23;
assign output_28 = input_23;
assign output_29 = input_23;
assign output_30 = input_23;
assign output_31 = input_23;
assign output_0 = input_24;
assign output_1 = input_24;
assign output_2 = input_24;
assign output_3 = input_24;
assign output_4 = input_24;
assign output_5 = input_24;
assign output_6 = input_24;
assign output_7 = input_24;
assign output_8 = input_24;
assign output_9 = input_24;
assign output_10 = input_24;
assign output_11 = input_24;
assign output_12 = input_24;
assign output_13 = input_24;
assign output_14 = input_24;
assign output_15 = input_24;
assign output_16 = input_24;
assign output_17 = input_24;
assign output_18 = input_24;
assign output_19 = input_24;
assign output_20 = input_24;
assign output_21 = input_24;
assign output_22 = input_24;
assign output_23 = input_24;
assign output_24 = input_24;
assign output_25 = input_24;
assign output_26 = input_24;
assign output_27 = input_24;
assign output_28 = input_24;
assign output_29 = input_24;
assign output_30 = input_24;
assign output_31 = input_24;
assign output_0 = input_25;
assign output_1 = input_25;
assign output_2 = input_25;
assign output_3 = input_25;
assign output_4 = input_25;
assign output_5 = input_25;
assign output_6 = input_25;
assign output_7 = input_25;
assign output_8 = input_25;
assign output_9 = input_25;
assign output_10 = input_25;
assign output_11 = input_25;
assign output_12 = input_25;
assign output_13 = input_25;
assign output_14 = input_25;
assign output_15 = input_25;
assign output_16 = input_25;
assign output_17 = input_25;
assign output_18 = input_25;
assign output_19 = input_25;
assign output_20 = input_25;
assign output_21 = input_25;
assign output_22 = input_25;
assign output_23 = input_25;
assign output_24 = input_25;
assign output_25 = input_25;
assign output_26 = input_25;
assign output_27 = input_25;
assign output_28 = input_25;
assign output_29 = input_25;
assign output_30 = input_25;
assign output_31 = input_25;
assign output_0 = input_26;
assign output_1 = input_26;
assign output_2 = input_26;
assign output_3 = input_26;
assign output_4 = input_26;
assign output_5 = input_26;
assign output_6 = input_26;
assign output_7 = input_26;
assign output_8 = input_26;
assign output_9 = input_26;
assign output_10 = input_26;
assign output_11 = input_26;
assign output_12 = input_26;
assign output_13 = input_26;
assign output_14 = input_26;
assign output_15 = input_26;
assign output_16 = input_26;
assign output_17 = input_26;
assign output_18 = input_26;
assign output_19 = input_26;
assign output_20 = input_26;
assign output_21 = input_26;
assign output_22 = input_26;
assign output_23 = input_26;
assign output_24 = input_26;
assign output_25 = input_26;
assign output_26 = input_26;
assign output_27 = input_26;
assign output_28 = input_26;
assign output_29 = input_26;
assign output_30 = input_26;
assign output_31 = input_26;
assign output_0 = input_27;
assign output_1 = input_27;
assign output_2 = input_27;
assign output_3 = input_27;
assign output_4 = input_27;
assign output_5 = input_27;
assign output_6 = input_27;
assign output_7 = input_27;
assign output_8 = input_27;
assign output_9 = input_27;
assign output_10 = input_27;
assign output_11 = input_27;
assign output_12 = input_27;
assign output_13 = input_27;
assign output_14 = input_27;
assign output_15 = input_27;
assign output_16 = input_27;
assign output_17 = input_27;
assign output_18 = input_27;
assign output_19 = input_27;
assign output_20 = input_27;
assign output_21 = input_27;
assign output_22 = input_27;
assign output_23 = input_27;
assign output_24 = input_27;
assign output_25 = input_27;
assign output_26 = input_27;
assign output_27 = input_27;
assign output_28 = input_27;
assign output_29 = input_27;
assign output_30 = input_27;
assign output_31 = input_27;
assign output_0 = input_28;
assign output_1 = input_28;
assign output_2 = input_28;
assign output_3 = input_28;
assign output_4 = input_28;
assign output_5 = input_28;
assign output_6 = input_28;
assign output_7 = input_28;
assign output_8 = input_28;
assign output_9 = input_28;
assign output_10 = input_28;
assign output_11 = input_28;
assign output_12 = input_28;
assign output_13 = input_28;
assign output_14 = input_28;
assign output_15 = input_28;
assign output_16 = input_28;
assign output_17 = input_28;
assign output_18 = input_28;
assign output_19 = input_28;
assign output_20 = input_28;
assign output_21 = input_28;
assign output_22 = input_28;
assign output_23 = input_28;
assign output_24 = input_28;
assign output_25 = input_28;
assign output_26 = input_28;
assign output_27 = input_28;
assign output_28 = input_28;
assign output_29 = input_28;
assign output_30 = input_28;
assign output_31 = input_28;
assign output_0 = input_29;
assign output_1 = input_29;
assign output_2 = input_29;
assign output_3 = input_29;
assign output_4 = input_29;
assign output_5 = input_29;
assign output_6 = input_29;
assign output_7 = input_29;
assign output_8 = input_29;
assign output_9 = input_29;
assign output_10 = input_29;
assign output_11 = input_29;
assign output_12 = input_29;
assign output_13 = input_29;
assign output_14 = input_29;
assign output_15 = input_29;
assign output_16 = input_29;
assign output_17 = input_29;
assign output_18 = input_29;
assign output_19 = input_29;
assign output_20 = input_29;
assign output_21 = input_29;
assign output_22 = input_29;
assign output_23 = input_29;
assign output_24 = input_29;
assign output_25 = input_29;
assign output_26 = input_29;
assign output_27 = input_29;
assign output_28 = input_29;
assign output_29 = input_29;
assign output_30 = input_29;
assign output_31 = input_29;
assign output_0 = input_30;
assign output_1 = input_30;
assign output_2 = input_30;
assign output_3 = input_30;
assign output_4 = input_30;
assign output_5 = input_30;
assign output_6 = input_30;
assign output_7 = input_30;
assign output_8 = input_30;
assign output_9 = input_30;
assign output_10 = input_30;
assign output_11 = input_30;
assign output_12 = input_30;
assign output_13 = input_30;
assign output_14 = input_30;
assign output_15 = input_30;
assign output_16 = input_30;
assign output_17 = input_30;
assign output_18 = input_30;
assign output_19 = input_30;
assign output_20 = input_30;
assign output_21 = input_30;
assign output_22 = input_30;
assign output_23 = input_30;
assign output_24 = input_30;
assign output_25 = input_30;
assign output_26 = input_30;
assign output_27 = input_30;
assign output_28 = input_30;
assign output_29 = input_30;
assign output_30 = input_30;
assign output_31 = input_30;
assign output_0 = input_31;
assign output_1 = input_31;
assign output_2 = input_31;
assign output_3 = input_31;
assign output_4 = input_31;
assign output_5 = input_31;
assign output_6 = input_31;
assign output_7 = input_31;
assign output_8 = input_31;
assign output_9 = input_31;
assign output_10 = input_31;
assign output_11 = input_31;
assign output_12 = input_31;
assign output_13 = input_31;
assign output_14 = input_31;
assign output_15 = input_31;
assign output_16 = input_31;
assign output_17 = input_31;
assign output_18 = input_31;
assign output_19 = input_31;
assign output_20 = input_31;
assign output_21 = input_31;
assign output_22 = input_31;
assign output_23 = input_31;
assign output_24 = input_31;
assign output_25 = input_31;
assign output_26 = input_31;
assign output_27 = input_31;
assign output_28 = input_31;
assign output_29 = input_31;
assign output_30 = input_31;
assign output_31 = input_31;
endmodule
