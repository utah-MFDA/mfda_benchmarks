module fanout2_braid_16_1024 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,output output_8,output output_9,output output_10,output output_11,output output_12,output output_13,output output_14,output output_15,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_9_0, output_9_1, output_8_0;
mixer gate_output_8_0(.a(output_9_0), .b(output_9_1), .y(output_8_0));
wire output_10_0, output_10_1, output_9_0;
mixer gate_output_9_0(.a(output_10_0), .b(output_10_1), .y(output_9_0));
wire output_11_0, output_11_1, output_10_0;
mixer gate_output_10_0(.a(output_11_0), .b(output_11_1), .y(output_10_0));
wire output_12_0, output_12_1, output_11_0;
mixer gate_output_11_0(.a(output_12_0), .b(output_12_1), .y(output_11_0));
wire output_13_0, output_13_1, output_12_0;
mixer gate_output_12_0(.a(output_13_0), .b(output_13_1), .y(output_12_0));
wire output_14_0, output_14_1, output_13_0;
mixer gate_output_13_0(.a(output_14_0), .b(output_14_1), .y(output_13_0));
wire output_15_0, output_15_1, output_14_0;
mixer gate_output_14_0(.a(output_15_0), .b(output_15_1), .y(output_14_0));
wire output_16_0, output_16_1, output_15_0;
mixer gate_output_15_0(.a(output_16_0), .b(output_16_1), .y(output_15_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_9_1, output_9_2, output_8_1;
mixer gate_output_8_1(.a(output_9_1), .b(output_9_2), .y(output_8_1));
wire output_10_1, output_10_2, output_9_1;
mixer gate_output_9_1(.a(output_10_1), .b(output_10_2), .y(output_9_1));
wire output_11_1, output_11_2, output_10_1;
mixer gate_output_10_1(.a(output_11_1), .b(output_11_2), .y(output_10_1));
wire output_12_1, output_12_2, output_11_1;
mixer gate_output_11_1(.a(output_12_1), .b(output_12_2), .y(output_11_1));
wire output_13_1, output_13_2, output_12_1;
mixer gate_output_12_1(.a(output_13_1), .b(output_13_2), .y(output_12_1));
wire output_14_1, output_14_2, output_13_1;
mixer gate_output_13_1(.a(output_14_1), .b(output_14_2), .y(output_13_1));
wire output_15_1, output_15_2, output_14_1;
mixer gate_output_14_1(.a(output_15_1), .b(output_15_2), .y(output_14_1));
wire output_16_1, output_16_2, output_15_1;
mixer gate_output_15_1(.a(output_16_1), .b(output_16_2), .y(output_15_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_9_2, output_9_3, output_8_2;
mixer gate_output_8_2(.a(output_9_2), .b(output_9_3), .y(output_8_2));
wire output_10_2, output_10_3, output_9_2;
mixer gate_output_9_2(.a(output_10_2), .b(output_10_3), .y(output_9_2));
wire output_11_2, output_11_3, output_10_2;
mixer gate_output_10_2(.a(output_11_2), .b(output_11_3), .y(output_10_2));
wire output_12_2, output_12_3, output_11_2;
mixer gate_output_11_2(.a(output_12_2), .b(output_12_3), .y(output_11_2));
wire output_13_2, output_13_3, output_12_2;
mixer gate_output_12_2(.a(output_13_2), .b(output_13_3), .y(output_12_2));
wire output_14_2, output_14_3, output_13_2;
mixer gate_output_13_2(.a(output_14_2), .b(output_14_3), .y(output_13_2));
wire output_15_2, output_15_3, output_14_2;
mixer gate_output_14_2(.a(output_15_2), .b(output_15_3), .y(output_14_2));
wire output_16_2, output_16_3, output_15_2;
mixer gate_output_15_2(.a(output_16_2), .b(output_16_3), .y(output_15_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_9_3, output_9_4, output_8_3;
mixer gate_output_8_3(.a(output_9_3), .b(output_9_4), .y(output_8_3));
wire output_10_3, output_10_4, output_9_3;
mixer gate_output_9_3(.a(output_10_3), .b(output_10_4), .y(output_9_3));
wire output_11_3, output_11_4, output_10_3;
mixer gate_output_10_3(.a(output_11_3), .b(output_11_4), .y(output_10_3));
wire output_12_3, output_12_4, output_11_3;
mixer gate_output_11_3(.a(output_12_3), .b(output_12_4), .y(output_11_3));
wire output_13_3, output_13_4, output_12_3;
mixer gate_output_12_3(.a(output_13_3), .b(output_13_4), .y(output_12_3));
wire output_14_3, output_14_4, output_13_3;
mixer gate_output_13_3(.a(output_14_3), .b(output_14_4), .y(output_13_3));
wire output_15_3, output_15_4, output_14_3;
mixer gate_output_14_3(.a(output_15_3), .b(output_15_4), .y(output_14_3));
wire output_16_3, output_16_4, output_15_3;
mixer gate_output_15_3(.a(output_16_3), .b(output_16_4), .y(output_15_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_9_4, output_9_5, output_8_4;
mixer gate_output_8_4(.a(output_9_4), .b(output_9_5), .y(output_8_4));
wire output_10_4, output_10_5, output_9_4;
mixer gate_output_9_4(.a(output_10_4), .b(output_10_5), .y(output_9_4));
wire output_11_4, output_11_5, output_10_4;
mixer gate_output_10_4(.a(output_11_4), .b(output_11_5), .y(output_10_4));
wire output_12_4, output_12_5, output_11_4;
mixer gate_output_11_4(.a(output_12_4), .b(output_12_5), .y(output_11_4));
wire output_13_4, output_13_5, output_12_4;
mixer gate_output_12_4(.a(output_13_4), .b(output_13_5), .y(output_12_4));
wire output_14_4, output_14_5, output_13_4;
mixer gate_output_13_4(.a(output_14_4), .b(output_14_5), .y(output_13_4));
wire output_15_4, output_15_5, output_14_4;
mixer gate_output_14_4(.a(output_15_4), .b(output_15_5), .y(output_14_4));
wire output_16_4, output_16_5, output_15_4;
mixer gate_output_15_4(.a(output_16_4), .b(output_16_5), .y(output_15_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_9_5, output_9_6, output_8_5;
mixer gate_output_8_5(.a(output_9_5), .b(output_9_6), .y(output_8_5));
wire output_10_5, output_10_6, output_9_5;
mixer gate_output_9_5(.a(output_10_5), .b(output_10_6), .y(output_9_5));
wire output_11_5, output_11_6, output_10_5;
mixer gate_output_10_5(.a(output_11_5), .b(output_11_6), .y(output_10_5));
wire output_12_5, output_12_6, output_11_5;
mixer gate_output_11_5(.a(output_12_5), .b(output_12_6), .y(output_11_5));
wire output_13_5, output_13_6, output_12_5;
mixer gate_output_12_5(.a(output_13_5), .b(output_13_6), .y(output_12_5));
wire output_14_5, output_14_6, output_13_5;
mixer gate_output_13_5(.a(output_14_5), .b(output_14_6), .y(output_13_5));
wire output_15_5, output_15_6, output_14_5;
mixer gate_output_14_5(.a(output_15_5), .b(output_15_6), .y(output_14_5));
wire output_16_5, output_16_6, output_15_5;
mixer gate_output_15_5(.a(output_16_5), .b(output_16_6), .y(output_15_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_9_6, output_9_7, output_8_6;
mixer gate_output_8_6(.a(output_9_6), .b(output_9_7), .y(output_8_6));
wire output_10_6, output_10_7, output_9_6;
mixer gate_output_9_6(.a(output_10_6), .b(output_10_7), .y(output_9_6));
wire output_11_6, output_11_7, output_10_6;
mixer gate_output_10_6(.a(output_11_6), .b(output_11_7), .y(output_10_6));
wire output_12_6, output_12_7, output_11_6;
mixer gate_output_11_6(.a(output_12_6), .b(output_12_7), .y(output_11_6));
wire output_13_6, output_13_7, output_12_6;
mixer gate_output_12_6(.a(output_13_6), .b(output_13_7), .y(output_12_6));
wire output_14_6, output_14_7, output_13_6;
mixer gate_output_13_6(.a(output_14_6), .b(output_14_7), .y(output_13_6));
wire output_15_6, output_15_7, output_14_6;
mixer gate_output_14_6(.a(output_15_6), .b(output_15_7), .y(output_14_6));
wire output_16_6, output_16_7, output_15_6;
mixer gate_output_15_6(.a(output_16_6), .b(output_16_7), .y(output_15_6));
wire output_1_7, output_1_8, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_8), .y(output_0_7));
wire output_2_7, output_2_8, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_8), .y(output_1_7));
wire output_3_7, output_3_8, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_8), .y(output_2_7));
wire output_4_7, output_4_8, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_8), .y(output_3_7));
wire output_5_7, output_5_8, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_8), .y(output_4_7));
wire output_6_7, output_6_8, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_8), .y(output_5_7));
wire output_7_7, output_7_8, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_8), .y(output_6_7));
wire output_8_7, output_8_8, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_8), .y(output_7_7));
wire output_9_7, output_9_8, output_8_7;
mixer gate_output_8_7(.a(output_9_7), .b(output_9_8), .y(output_8_7));
wire output_10_7, output_10_8, output_9_7;
mixer gate_output_9_7(.a(output_10_7), .b(output_10_8), .y(output_9_7));
wire output_11_7, output_11_8, output_10_7;
mixer gate_output_10_7(.a(output_11_7), .b(output_11_8), .y(output_10_7));
wire output_12_7, output_12_8, output_11_7;
mixer gate_output_11_7(.a(output_12_7), .b(output_12_8), .y(output_11_7));
wire output_13_7, output_13_8, output_12_7;
mixer gate_output_12_7(.a(output_13_7), .b(output_13_8), .y(output_12_7));
wire output_14_7, output_14_8, output_13_7;
mixer gate_output_13_7(.a(output_14_7), .b(output_14_8), .y(output_13_7));
wire output_15_7, output_15_8, output_14_7;
mixer gate_output_14_7(.a(output_15_7), .b(output_15_8), .y(output_14_7));
wire output_16_7, output_16_8, output_15_7;
mixer gate_output_15_7(.a(output_16_7), .b(output_16_8), .y(output_15_7));
wire output_1_8, output_1_9, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_9), .y(output_0_8));
wire output_2_8, output_2_9, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_9), .y(output_1_8));
wire output_3_8, output_3_9, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_9), .y(output_2_8));
wire output_4_8, output_4_9, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_9), .y(output_3_8));
wire output_5_8, output_5_9, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_9), .y(output_4_8));
wire output_6_8, output_6_9, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_9), .y(output_5_8));
wire output_7_8, output_7_9, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_9), .y(output_6_8));
wire output_8_8, output_8_9, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_9), .y(output_7_8));
wire output_9_8, output_9_9, output_8_8;
mixer gate_output_8_8(.a(output_9_8), .b(output_9_9), .y(output_8_8));
wire output_10_8, output_10_9, output_9_8;
mixer gate_output_9_8(.a(output_10_8), .b(output_10_9), .y(output_9_8));
wire output_11_8, output_11_9, output_10_8;
mixer gate_output_10_8(.a(output_11_8), .b(output_11_9), .y(output_10_8));
wire output_12_8, output_12_9, output_11_8;
mixer gate_output_11_8(.a(output_12_8), .b(output_12_9), .y(output_11_8));
wire output_13_8, output_13_9, output_12_8;
mixer gate_output_12_8(.a(output_13_8), .b(output_13_9), .y(output_12_8));
wire output_14_8, output_14_9, output_13_8;
mixer gate_output_13_8(.a(output_14_8), .b(output_14_9), .y(output_13_8));
wire output_15_8, output_15_9, output_14_8;
mixer gate_output_14_8(.a(output_15_8), .b(output_15_9), .y(output_14_8));
wire output_16_8, output_16_9, output_15_8;
mixer gate_output_15_8(.a(output_16_8), .b(output_16_9), .y(output_15_8));
wire output_1_9, output_1_10, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_10), .y(output_0_9));
wire output_2_9, output_2_10, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_10), .y(output_1_9));
wire output_3_9, output_3_10, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_10), .y(output_2_9));
wire output_4_9, output_4_10, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_10), .y(output_3_9));
wire output_5_9, output_5_10, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_10), .y(output_4_9));
wire output_6_9, output_6_10, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_10), .y(output_5_9));
wire output_7_9, output_7_10, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_10), .y(output_6_9));
wire output_8_9, output_8_10, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_10), .y(output_7_9));
wire output_9_9, output_9_10, output_8_9;
mixer gate_output_8_9(.a(output_9_9), .b(output_9_10), .y(output_8_9));
wire output_10_9, output_10_10, output_9_9;
mixer gate_output_9_9(.a(output_10_9), .b(output_10_10), .y(output_9_9));
wire output_11_9, output_11_10, output_10_9;
mixer gate_output_10_9(.a(output_11_9), .b(output_11_10), .y(output_10_9));
wire output_12_9, output_12_10, output_11_9;
mixer gate_output_11_9(.a(output_12_9), .b(output_12_10), .y(output_11_9));
wire output_13_9, output_13_10, output_12_9;
mixer gate_output_12_9(.a(output_13_9), .b(output_13_10), .y(output_12_9));
wire output_14_9, output_14_10, output_13_9;
mixer gate_output_13_9(.a(output_14_9), .b(output_14_10), .y(output_13_9));
wire output_15_9, output_15_10, output_14_9;
mixer gate_output_14_9(.a(output_15_9), .b(output_15_10), .y(output_14_9));
wire output_16_9, output_16_10, output_15_9;
mixer gate_output_15_9(.a(output_16_9), .b(output_16_10), .y(output_15_9));
wire output_1_10, output_1_11, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_11), .y(output_0_10));
wire output_2_10, output_2_11, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_11), .y(output_1_10));
wire output_3_10, output_3_11, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_11), .y(output_2_10));
wire output_4_10, output_4_11, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_11), .y(output_3_10));
wire output_5_10, output_5_11, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_11), .y(output_4_10));
wire output_6_10, output_6_11, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_11), .y(output_5_10));
wire output_7_10, output_7_11, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_11), .y(output_6_10));
wire output_8_10, output_8_11, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_11), .y(output_7_10));
wire output_9_10, output_9_11, output_8_10;
mixer gate_output_8_10(.a(output_9_10), .b(output_9_11), .y(output_8_10));
wire output_10_10, output_10_11, output_9_10;
mixer gate_output_9_10(.a(output_10_10), .b(output_10_11), .y(output_9_10));
wire output_11_10, output_11_11, output_10_10;
mixer gate_output_10_10(.a(output_11_10), .b(output_11_11), .y(output_10_10));
wire output_12_10, output_12_11, output_11_10;
mixer gate_output_11_10(.a(output_12_10), .b(output_12_11), .y(output_11_10));
wire output_13_10, output_13_11, output_12_10;
mixer gate_output_12_10(.a(output_13_10), .b(output_13_11), .y(output_12_10));
wire output_14_10, output_14_11, output_13_10;
mixer gate_output_13_10(.a(output_14_10), .b(output_14_11), .y(output_13_10));
wire output_15_10, output_15_11, output_14_10;
mixer gate_output_14_10(.a(output_15_10), .b(output_15_11), .y(output_14_10));
wire output_16_10, output_16_11, output_15_10;
mixer gate_output_15_10(.a(output_16_10), .b(output_16_11), .y(output_15_10));
wire output_1_11, output_1_12, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_12), .y(output_0_11));
wire output_2_11, output_2_12, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_12), .y(output_1_11));
wire output_3_11, output_3_12, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_12), .y(output_2_11));
wire output_4_11, output_4_12, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_12), .y(output_3_11));
wire output_5_11, output_5_12, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_12), .y(output_4_11));
wire output_6_11, output_6_12, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_12), .y(output_5_11));
wire output_7_11, output_7_12, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_12), .y(output_6_11));
wire output_8_11, output_8_12, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_12), .y(output_7_11));
wire output_9_11, output_9_12, output_8_11;
mixer gate_output_8_11(.a(output_9_11), .b(output_9_12), .y(output_8_11));
wire output_10_11, output_10_12, output_9_11;
mixer gate_output_9_11(.a(output_10_11), .b(output_10_12), .y(output_9_11));
wire output_11_11, output_11_12, output_10_11;
mixer gate_output_10_11(.a(output_11_11), .b(output_11_12), .y(output_10_11));
wire output_12_11, output_12_12, output_11_11;
mixer gate_output_11_11(.a(output_12_11), .b(output_12_12), .y(output_11_11));
wire output_13_11, output_13_12, output_12_11;
mixer gate_output_12_11(.a(output_13_11), .b(output_13_12), .y(output_12_11));
wire output_14_11, output_14_12, output_13_11;
mixer gate_output_13_11(.a(output_14_11), .b(output_14_12), .y(output_13_11));
wire output_15_11, output_15_12, output_14_11;
mixer gate_output_14_11(.a(output_15_11), .b(output_15_12), .y(output_14_11));
wire output_16_11, output_16_12, output_15_11;
mixer gate_output_15_11(.a(output_16_11), .b(output_16_12), .y(output_15_11));
wire output_1_12, output_1_13, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_13), .y(output_0_12));
wire output_2_12, output_2_13, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_13), .y(output_1_12));
wire output_3_12, output_3_13, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_13), .y(output_2_12));
wire output_4_12, output_4_13, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_13), .y(output_3_12));
wire output_5_12, output_5_13, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_13), .y(output_4_12));
wire output_6_12, output_6_13, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_13), .y(output_5_12));
wire output_7_12, output_7_13, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_13), .y(output_6_12));
wire output_8_12, output_8_13, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_13), .y(output_7_12));
wire output_9_12, output_9_13, output_8_12;
mixer gate_output_8_12(.a(output_9_12), .b(output_9_13), .y(output_8_12));
wire output_10_12, output_10_13, output_9_12;
mixer gate_output_9_12(.a(output_10_12), .b(output_10_13), .y(output_9_12));
wire output_11_12, output_11_13, output_10_12;
mixer gate_output_10_12(.a(output_11_12), .b(output_11_13), .y(output_10_12));
wire output_12_12, output_12_13, output_11_12;
mixer gate_output_11_12(.a(output_12_12), .b(output_12_13), .y(output_11_12));
wire output_13_12, output_13_13, output_12_12;
mixer gate_output_12_12(.a(output_13_12), .b(output_13_13), .y(output_12_12));
wire output_14_12, output_14_13, output_13_12;
mixer gate_output_13_12(.a(output_14_12), .b(output_14_13), .y(output_13_12));
wire output_15_12, output_15_13, output_14_12;
mixer gate_output_14_12(.a(output_15_12), .b(output_15_13), .y(output_14_12));
wire output_16_12, output_16_13, output_15_12;
mixer gate_output_15_12(.a(output_16_12), .b(output_16_13), .y(output_15_12));
wire output_1_13, output_1_14, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_14), .y(output_0_13));
wire output_2_13, output_2_14, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_14), .y(output_1_13));
wire output_3_13, output_3_14, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_14), .y(output_2_13));
wire output_4_13, output_4_14, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_14), .y(output_3_13));
wire output_5_13, output_5_14, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_14), .y(output_4_13));
wire output_6_13, output_6_14, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_14), .y(output_5_13));
wire output_7_13, output_7_14, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_14), .y(output_6_13));
wire output_8_13, output_8_14, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_14), .y(output_7_13));
wire output_9_13, output_9_14, output_8_13;
mixer gate_output_8_13(.a(output_9_13), .b(output_9_14), .y(output_8_13));
wire output_10_13, output_10_14, output_9_13;
mixer gate_output_9_13(.a(output_10_13), .b(output_10_14), .y(output_9_13));
wire output_11_13, output_11_14, output_10_13;
mixer gate_output_10_13(.a(output_11_13), .b(output_11_14), .y(output_10_13));
wire output_12_13, output_12_14, output_11_13;
mixer gate_output_11_13(.a(output_12_13), .b(output_12_14), .y(output_11_13));
wire output_13_13, output_13_14, output_12_13;
mixer gate_output_12_13(.a(output_13_13), .b(output_13_14), .y(output_12_13));
wire output_14_13, output_14_14, output_13_13;
mixer gate_output_13_13(.a(output_14_13), .b(output_14_14), .y(output_13_13));
wire output_15_13, output_15_14, output_14_13;
mixer gate_output_14_13(.a(output_15_13), .b(output_15_14), .y(output_14_13));
wire output_16_13, output_16_14, output_15_13;
mixer gate_output_15_13(.a(output_16_13), .b(output_16_14), .y(output_15_13));
wire output_1_14, output_1_15, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_15), .y(output_0_14));
wire output_2_14, output_2_15, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_15), .y(output_1_14));
wire output_3_14, output_3_15, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_15), .y(output_2_14));
wire output_4_14, output_4_15, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_15), .y(output_3_14));
wire output_5_14, output_5_15, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_15), .y(output_4_14));
wire output_6_14, output_6_15, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_15), .y(output_5_14));
wire output_7_14, output_7_15, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_15), .y(output_6_14));
wire output_8_14, output_8_15, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_15), .y(output_7_14));
wire output_9_14, output_9_15, output_8_14;
mixer gate_output_8_14(.a(output_9_14), .b(output_9_15), .y(output_8_14));
wire output_10_14, output_10_15, output_9_14;
mixer gate_output_9_14(.a(output_10_14), .b(output_10_15), .y(output_9_14));
wire output_11_14, output_11_15, output_10_14;
mixer gate_output_10_14(.a(output_11_14), .b(output_11_15), .y(output_10_14));
wire output_12_14, output_12_15, output_11_14;
mixer gate_output_11_14(.a(output_12_14), .b(output_12_15), .y(output_11_14));
wire output_13_14, output_13_15, output_12_14;
mixer gate_output_12_14(.a(output_13_14), .b(output_13_15), .y(output_12_14));
wire output_14_14, output_14_15, output_13_14;
mixer gate_output_13_14(.a(output_14_14), .b(output_14_15), .y(output_13_14));
wire output_15_14, output_15_15, output_14_14;
mixer gate_output_14_14(.a(output_15_14), .b(output_15_15), .y(output_14_14));
wire output_16_14, output_16_15, output_15_14;
mixer gate_output_15_14(.a(output_16_14), .b(output_16_15), .y(output_15_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
wire output_9_15, output_9_0, output_8_15;
mixer gate_output_8_15(.a(output_9_15), .b(output_9_0), .y(output_8_15));
wire output_10_15, output_10_0, output_9_15;
mixer gate_output_9_15(.a(output_10_15), .b(output_10_0), .y(output_9_15));
wire output_11_15, output_11_0, output_10_15;
mixer gate_output_10_15(.a(output_11_15), .b(output_11_0), .y(output_10_15));
wire output_12_15, output_12_0, output_11_15;
mixer gate_output_11_15(.a(output_12_15), .b(output_12_0), .y(output_11_15));
wire output_13_15, output_13_0, output_12_15;
mixer gate_output_12_15(.a(output_13_15), .b(output_13_0), .y(output_12_15));
wire output_14_15, output_14_0, output_13_15;
mixer gate_output_13_15(.a(output_14_15), .b(output_14_0), .y(output_13_15));
wire output_15_15, output_15_0, output_14_15;
mixer gate_output_14_15(.a(output_15_15), .b(output_15_0), .y(output_14_15));
wire output_16_15, output_16_0, output_15_15;
mixer gate_output_15_15(.a(output_16_15), .b(output_16_0), .y(output_15_15));
wire output_1_16, output_1_1, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_1), .y(output_0_16));
wire output_2_16, output_2_1, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_1), .y(output_1_16));
wire output_3_16, output_3_1, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_1), .y(output_2_16));
wire output_4_16, output_4_1, output_3_16;
mixer gate_output_3_16(.a(output_4_16), .b(output_4_1), .y(output_3_16));
wire output_5_16, output_5_1, output_4_16;
mixer gate_output_4_16(.a(output_5_16), .b(output_5_1), .y(output_4_16));
wire output_6_16, output_6_1, output_5_16;
mixer gate_output_5_16(.a(output_6_16), .b(output_6_1), .y(output_5_16));
wire output_7_16, output_7_1, output_6_16;
mixer gate_output_6_16(.a(output_7_16), .b(output_7_1), .y(output_6_16));
wire output_8_16, output_8_1, output_7_16;
mixer gate_output_7_16(.a(output_8_16), .b(output_8_1), .y(output_7_16));
wire output_9_16, output_9_1, output_8_16;
mixer gate_output_8_16(.a(output_9_16), .b(output_9_1), .y(output_8_16));
wire output_10_16, output_10_1, output_9_16;
mixer gate_output_9_16(.a(output_10_16), .b(output_10_1), .y(output_9_16));
wire output_11_16, output_11_1, output_10_16;
mixer gate_output_10_16(.a(output_11_16), .b(output_11_1), .y(output_10_16));
wire output_12_16, output_12_1, output_11_16;
mixer gate_output_11_16(.a(output_12_16), .b(output_12_1), .y(output_11_16));
wire output_13_16, output_13_1, output_12_16;
mixer gate_output_12_16(.a(output_13_16), .b(output_13_1), .y(output_12_16));
wire output_14_16, output_14_1, output_13_16;
mixer gate_output_13_16(.a(output_14_16), .b(output_14_1), .y(output_13_16));
wire output_15_16, output_15_1, output_14_16;
mixer gate_output_14_16(.a(output_15_16), .b(output_15_1), .y(output_14_16));
wire output_16_16, output_16_1, output_15_16;
mixer gate_output_15_16(.a(output_16_16), .b(output_16_1), .y(output_15_16));
wire output_1_17, output_1_2, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_2), .y(output_0_17));
wire output_2_17, output_2_2, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_2), .y(output_1_17));
wire output_3_17, output_3_2, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_2), .y(output_2_17));
wire output_4_17, output_4_2, output_3_17;
mixer gate_output_3_17(.a(output_4_17), .b(output_4_2), .y(output_3_17));
wire output_5_17, output_5_2, output_4_17;
mixer gate_output_4_17(.a(output_5_17), .b(output_5_2), .y(output_4_17));
wire output_6_17, output_6_2, output_5_17;
mixer gate_output_5_17(.a(output_6_17), .b(output_6_2), .y(output_5_17));
wire output_7_17, output_7_2, output_6_17;
mixer gate_output_6_17(.a(output_7_17), .b(output_7_2), .y(output_6_17));
wire output_8_17, output_8_2, output_7_17;
mixer gate_output_7_17(.a(output_8_17), .b(output_8_2), .y(output_7_17));
wire output_9_17, output_9_2, output_8_17;
mixer gate_output_8_17(.a(output_9_17), .b(output_9_2), .y(output_8_17));
wire output_10_17, output_10_2, output_9_17;
mixer gate_output_9_17(.a(output_10_17), .b(output_10_2), .y(output_9_17));
wire output_11_17, output_11_2, output_10_17;
mixer gate_output_10_17(.a(output_11_17), .b(output_11_2), .y(output_10_17));
wire output_12_17, output_12_2, output_11_17;
mixer gate_output_11_17(.a(output_12_17), .b(output_12_2), .y(output_11_17));
wire output_13_17, output_13_2, output_12_17;
mixer gate_output_12_17(.a(output_13_17), .b(output_13_2), .y(output_12_17));
wire output_14_17, output_14_2, output_13_17;
mixer gate_output_13_17(.a(output_14_17), .b(output_14_2), .y(output_13_17));
wire output_15_17, output_15_2, output_14_17;
mixer gate_output_14_17(.a(output_15_17), .b(output_15_2), .y(output_14_17));
wire output_16_17, output_16_2, output_15_17;
mixer gate_output_15_17(.a(output_16_17), .b(output_16_2), .y(output_15_17));
wire output_1_18, output_1_3, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_3), .y(output_0_18));
wire output_2_18, output_2_3, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_3), .y(output_1_18));
wire output_3_18, output_3_3, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_3), .y(output_2_18));
wire output_4_18, output_4_3, output_3_18;
mixer gate_output_3_18(.a(output_4_18), .b(output_4_3), .y(output_3_18));
wire output_5_18, output_5_3, output_4_18;
mixer gate_output_4_18(.a(output_5_18), .b(output_5_3), .y(output_4_18));
wire output_6_18, output_6_3, output_5_18;
mixer gate_output_5_18(.a(output_6_18), .b(output_6_3), .y(output_5_18));
wire output_7_18, output_7_3, output_6_18;
mixer gate_output_6_18(.a(output_7_18), .b(output_7_3), .y(output_6_18));
wire output_8_18, output_8_3, output_7_18;
mixer gate_output_7_18(.a(output_8_18), .b(output_8_3), .y(output_7_18));
wire output_9_18, output_9_3, output_8_18;
mixer gate_output_8_18(.a(output_9_18), .b(output_9_3), .y(output_8_18));
wire output_10_18, output_10_3, output_9_18;
mixer gate_output_9_18(.a(output_10_18), .b(output_10_3), .y(output_9_18));
wire output_11_18, output_11_3, output_10_18;
mixer gate_output_10_18(.a(output_11_18), .b(output_11_3), .y(output_10_18));
wire output_12_18, output_12_3, output_11_18;
mixer gate_output_11_18(.a(output_12_18), .b(output_12_3), .y(output_11_18));
wire output_13_18, output_13_3, output_12_18;
mixer gate_output_12_18(.a(output_13_18), .b(output_13_3), .y(output_12_18));
wire output_14_18, output_14_3, output_13_18;
mixer gate_output_13_18(.a(output_14_18), .b(output_14_3), .y(output_13_18));
wire output_15_18, output_15_3, output_14_18;
mixer gate_output_14_18(.a(output_15_18), .b(output_15_3), .y(output_14_18));
wire output_16_18, output_16_3, output_15_18;
mixer gate_output_15_18(.a(output_16_18), .b(output_16_3), .y(output_15_18));
wire output_1_19, output_1_4, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_4), .y(output_0_19));
wire output_2_19, output_2_4, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_4), .y(output_1_19));
wire output_3_19, output_3_4, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_4), .y(output_2_19));
wire output_4_19, output_4_4, output_3_19;
mixer gate_output_3_19(.a(output_4_19), .b(output_4_4), .y(output_3_19));
wire output_5_19, output_5_4, output_4_19;
mixer gate_output_4_19(.a(output_5_19), .b(output_5_4), .y(output_4_19));
wire output_6_19, output_6_4, output_5_19;
mixer gate_output_5_19(.a(output_6_19), .b(output_6_4), .y(output_5_19));
wire output_7_19, output_7_4, output_6_19;
mixer gate_output_6_19(.a(output_7_19), .b(output_7_4), .y(output_6_19));
wire output_8_19, output_8_4, output_7_19;
mixer gate_output_7_19(.a(output_8_19), .b(output_8_4), .y(output_7_19));
wire output_9_19, output_9_4, output_8_19;
mixer gate_output_8_19(.a(output_9_19), .b(output_9_4), .y(output_8_19));
wire output_10_19, output_10_4, output_9_19;
mixer gate_output_9_19(.a(output_10_19), .b(output_10_4), .y(output_9_19));
wire output_11_19, output_11_4, output_10_19;
mixer gate_output_10_19(.a(output_11_19), .b(output_11_4), .y(output_10_19));
wire output_12_19, output_12_4, output_11_19;
mixer gate_output_11_19(.a(output_12_19), .b(output_12_4), .y(output_11_19));
wire output_13_19, output_13_4, output_12_19;
mixer gate_output_12_19(.a(output_13_19), .b(output_13_4), .y(output_12_19));
wire output_14_19, output_14_4, output_13_19;
mixer gate_output_13_19(.a(output_14_19), .b(output_14_4), .y(output_13_19));
wire output_15_19, output_15_4, output_14_19;
mixer gate_output_14_19(.a(output_15_19), .b(output_15_4), .y(output_14_19));
wire output_16_19, output_16_4, output_15_19;
mixer gate_output_15_19(.a(output_16_19), .b(output_16_4), .y(output_15_19));
wire output_1_20, output_1_5, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_5), .y(output_0_20));
wire output_2_20, output_2_5, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_5), .y(output_1_20));
wire output_3_20, output_3_5, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_5), .y(output_2_20));
wire output_4_20, output_4_5, output_3_20;
mixer gate_output_3_20(.a(output_4_20), .b(output_4_5), .y(output_3_20));
wire output_5_20, output_5_5, output_4_20;
mixer gate_output_4_20(.a(output_5_20), .b(output_5_5), .y(output_4_20));
wire output_6_20, output_6_5, output_5_20;
mixer gate_output_5_20(.a(output_6_20), .b(output_6_5), .y(output_5_20));
wire output_7_20, output_7_5, output_6_20;
mixer gate_output_6_20(.a(output_7_20), .b(output_7_5), .y(output_6_20));
wire output_8_20, output_8_5, output_7_20;
mixer gate_output_7_20(.a(output_8_20), .b(output_8_5), .y(output_7_20));
wire output_9_20, output_9_5, output_8_20;
mixer gate_output_8_20(.a(output_9_20), .b(output_9_5), .y(output_8_20));
wire output_10_20, output_10_5, output_9_20;
mixer gate_output_9_20(.a(output_10_20), .b(output_10_5), .y(output_9_20));
wire output_11_20, output_11_5, output_10_20;
mixer gate_output_10_20(.a(output_11_20), .b(output_11_5), .y(output_10_20));
wire output_12_20, output_12_5, output_11_20;
mixer gate_output_11_20(.a(output_12_20), .b(output_12_5), .y(output_11_20));
wire output_13_20, output_13_5, output_12_20;
mixer gate_output_12_20(.a(output_13_20), .b(output_13_5), .y(output_12_20));
wire output_14_20, output_14_5, output_13_20;
mixer gate_output_13_20(.a(output_14_20), .b(output_14_5), .y(output_13_20));
wire output_15_20, output_15_5, output_14_20;
mixer gate_output_14_20(.a(output_15_20), .b(output_15_5), .y(output_14_20));
wire output_16_20, output_16_5, output_15_20;
mixer gate_output_15_20(.a(output_16_20), .b(output_16_5), .y(output_15_20));
wire output_1_21, output_1_6, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_6), .y(output_0_21));
wire output_2_21, output_2_6, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_6), .y(output_1_21));
wire output_3_21, output_3_6, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_6), .y(output_2_21));
wire output_4_21, output_4_6, output_3_21;
mixer gate_output_3_21(.a(output_4_21), .b(output_4_6), .y(output_3_21));
wire output_5_21, output_5_6, output_4_21;
mixer gate_output_4_21(.a(output_5_21), .b(output_5_6), .y(output_4_21));
wire output_6_21, output_6_6, output_5_21;
mixer gate_output_5_21(.a(output_6_21), .b(output_6_6), .y(output_5_21));
wire output_7_21, output_7_6, output_6_21;
mixer gate_output_6_21(.a(output_7_21), .b(output_7_6), .y(output_6_21));
wire output_8_21, output_8_6, output_7_21;
mixer gate_output_7_21(.a(output_8_21), .b(output_8_6), .y(output_7_21));
wire output_9_21, output_9_6, output_8_21;
mixer gate_output_8_21(.a(output_9_21), .b(output_9_6), .y(output_8_21));
wire output_10_21, output_10_6, output_9_21;
mixer gate_output_9_21(.a(output_10_21), .b(output_10_6), .y(output_9_21));
wire output_11_21, output_11_6, output_10_21;
mixer gate_output_10_21(.a(output_11_21), .b(output_11_6), .y(output_10_21));
wire output_12_21, output_12_6, output_11_21;
mixer gate_output_11_21(.a(output_12_21), .b(output_12_6), .y(output_11_21));
wire output_13_21, output_13_6, output_12_21;
mixer gate_output_12_21(.a(output_13_21), .b(output_13_6), .y(output_12_21));
wire output_14_21, output_14_6, output_13_21;
mixer gate_output_13_21(.a(output_14_21), .b(output_14_6), .y(output_13_21));
wire output_15_21, output_15_6, output_14_21;
mixer gate_output_14_21(.a(output_15_21), .b(output_15_6), .y(output_14_21));
wire output_16_21, output_16_6, output_15_21;
mixer gate_output_15_21(.a(output_16_21), .b(output_16_6), .y(output_15_21));
wire output_1_22, output_1_7, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_7), .y(output_0_22));
wire output_2_22, output_2_7, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_7), .y(output_1_22));
wire output_3_22, output_3_7, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_7), .y(output_2_22));
wire output_4_22, output_4_7, output_3_22;
mixer gate_output_3_22(.a(output_4_22), .b(output_4_7), .y(output_3_22));
wire output_5_22, output_5_7, output_4_22;
mixer gate_output_4_22(.a(output_5_22), .b(output_5_7), .y(output_4_22));
wire output_6_22, output_6_7, output_5_22;
mixer gate_output_5_22(.a(output_6_22), .b(output_6_7), .y(output_5_22));
wire output_7_22, output_7_7, output_6_22;
mixer gate_output_6_22(.a(output_7_22), .b(output_7_7), .y(output_6_22));
wire output_8_22, output_8_7, output_7_22;
mixer gate_output_7_22(.a(output_8_22), .b(output_8_7), .y(output_7_22));
wire output_9_22, output_9_7, output_8_22;
mixer gate_output_8_22(.a(output_9_22), .b(output_9_7), .y(output_8_22));
wire output_10_22, output_10_7, output_9_22;
mixer gate_output_9_22(.a(output_10_22), .b(output_10_7), .y(output_9_22));
wire output_11_22, output_11_7, output_10_22;
mixer gate_output_10_22(.a(output_11_22), .b(output_11_7), .y(output_10_22));
wire output_12_22, output_12_7, output_11_22;
mixer gate_output_11_22(.a(output_12_22), .b(output_12_7), .y(output_11_22));
wire output_13_22, output_13_7, output_12_22;
mixer gate_output_12_22(.a(output_13_22), .b(output_13_7), .y(output_12_22));
wire output_14_22, output_14_7, output_13_22;
mixer gate_output_13_22(.a(output_14_22), .b(output_14_7), .y(output_13_22));
wire output_15_22, output_15_7, output_14_22;
mixer gate_output_14_22(.a(output_15_22), .b(output_15_7), .y(output_14_22));
wire output_16_22, output_16_7, output_15_22;
mixer gate_output_15_22(.a(output_16_22), .b(output_16_7), .y(output_15_22));
wire output_1_23, output_1_8, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_8), .y(output_0_23));
wire output_2_23, output_2_8, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_8), .y(output_1_23));
wire output_3_23, output_3_8, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_8), .y(output_2_23));
wire output_4_23, output_4_8, output_3_23;
mixer gate_output_3_23(.a(output_4_23), .b(output_4_8), .y(output_3_23));
wire output_5_23, output_5_8, output_4_23;
mixer gate_output_4_23(.a(output_5_23), .b(output_5_8), .y(output_4_23));
wire output_6_23, output_6_8, output_5_23;
mixer gate_output_5_23(.a(output_6_23), .b(output_6_8), .y(output_5_23));
wire output_7_23, output_7_8, output_6_23;
mixer gate_output_6_23(.a(output_7_23), .b(output_7_8), .y(output_6_23));
wire output_8_23, output_8_8, output_7_23;
mixer gate_output_7_23(.a(output_8_23), .b(output_8_8), .y(output_7_23));
wire output_9_23, output_9_8, output_8_23;
mixer gate_output_8_23(.a(output_9_23), .b(output_9_8), .y(output_8_23));
wire output_10_23, output_10_8, output_9_23;
mixer gate_output_9_23(.a(output_10_23), .b(output_10_8), .y(output_9_23));
wire output_11_23, output_11_8, output_10_23;
mixer gate_output_10_23(.a(output_11_23), .b(output_11_8), .y(output_10_23));
wire output_12_23, output_12_8, output_11_23;
mixer gate_output_11_23(.a(output_12_23), .b(output_12_8), .y(output_11_23));
wire output_13_23, output_13_8, output_12_23;
mixer gate_output_12_23(.a(output_13_23), .b(output_13_8), .y(output_12_23));
wire output_14_23, output_14_8, output_13_23;
mixer gate_output_13_23(.a(output_14_23), .b(output_14_8), .y(output_13_23));
wire output_15_23, output_15_8, output_14_23;
mixer gate_output_14_23(.a(output_15_23), .b(output_15_8), .y(output_14_23));
wire output_16_23, output_16_8, output_15_23;
mixer gate_output_15_23(.a(output_16_23), .b(output_16_8), .y(output_15_23));
wire output_1_24, output_1_9, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_9), .y(output_0_24));
wire output_2_24, output_2_9, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_9), .y(output_1_24));
wire output_3_24, output_3_9, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_9), .y(output_2_24));
wire output_4_24, output_4_9, output_3_24;
mixer gate_output_3_24(.a(output_4_24), .b(output_4_9), .y(output_3_24));
wire output_5_24, output_5_9, output_4_24;
mixer gate_output_4_24(.a(output_5_24), .b(output_5_9), .y(output_4_24));
wire output_6_24, output_6_9, output_5_24;
mixer gate_output_5_24(.a(output_6_24), .b(output_6_9), .y(output_5_24));
wire output_7_24, output_7_9, output_6_24;
mixer gate_output_6_24(.a(output_7_24), .b(output_7_9), .y(output_6_24));
wire output_8_24, output_8_9, output_7_24;
mixer gate_output_7_24(.a(output_8_24), .b(output_8_9), .y(output_7_24));
wire output_9_24, output_9_9, output_8_24;
mixer gate_output_8_24(.a(output_9_24), .b(output_9_9), .y(output_8_24));
wire output_10_24, output_10_9, output_9_24;
mixer gate_output_9_24(.a(output_10_24), .b(output_10_9), .y(output_9_24));
wire output_11_24, output_11_9, output_10_24;
mixer gate_output_10_24(.a(output_11_24), .b(output_11_9), .y(output_10_24));
wire output_12_24, output_12_9, output_11_24;
mixer gate_output_11_24(.a(output_12_24), .b(output_12_9), .y(output_11_24));
wire output_13_24, output_13_9, output_12_24;
mixer gate_output_12_24(.a(output_13_24), .b(output_13_9), .y(output_12_24));
wire output_14_24, output_14_9, output_13_24;
mixer gate_output_13_24(.a(output_14_24), .b(output_14_9), .y(output_13_24));
wire output_15_24, output_15_9, output_14_24;
mixer gate_output_14_24(.a(output_15_24), .b(output_15_9), .y(output_14_24));
wire output_16_24, output_16_9, output_15_24;
mixer gate_output_15_24(.a(output_16_24), .b(output_16_9), .y(output_15_24));
wire output_1_25, output_1_10, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_10), .y(output_0_25));
wire output_2_25, output_2_10, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_10), .y(output_1_25));
wire output_3_25, output_3_10, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_10), .y(output_2_25));
wire output_4_25, output_4_10, output_3_25;
mixer gate_output_3_25(.a(output_4_25), .b(output_4_10), .y(output_3_25));
wire output_5_25, output_5_10, output_4_25;
mixer gate_output_4_25(.a(output_5_25), .b(output_5_10), .y(output_4_25));
wire output_6_25, output_6_10, output_5_25;
mixer gate_output_5_25(.a(output_6_25), .b(output_6_10), .y(output_5_25));
wire output_7_25, output_7_10, output_6_25;
mixer gate_output_6_25(.a(output_7_25), .b(output_7_10), .y(output_6_25));
wire output_8_25, output_8_10, output_7_25;
mixer gate_output_7_25(.a(output_8_25), .b(output_8_10), .y(output_7_25));
wire output_9_25, output_9_10, output_8_25;
mixer gate_output_8_25(.a(output_9_25), .b(output_9_10), .y(output_8_25));
wire output_10_25, output_10_10, output_9_25;
mixer gate_output_9_25(.a(output_10_25), .b(output_10_10), .y(output_9_25));
wire output_11_25, output_11_10, output_10_25;
mixer gate_output_10_25(.a(output_11_25), .b(output_11_10), .y(output_10_25));
wire output_12_25, output_12_10, output_11_25;
mixer gate_output_11_25(.a(output_12_25), .b(output_12_10), .y(output_11_25));
wire output_13_25, output_13_10, output_12_25;
mixer gate_output_12_25(.a(output_13_25), .b(output_13_10), .y(output_12_25));
wire output_14_25, output_14_10, output_13_25;
mixer gate_output_13_25(.a(output_14_25), .b(output_14_10), .y(output_13_25));
wire output_15_25, output_15_10, output_14_25;
mixer gate_output_14_25(.a(output_15_25), .b(output_15_10), .y(output_14_25));
wire output_16_25, output_16_10, output_15_25;
mixer gate_output_15_25(.a(output_16_25), .b(output_16_10), .y(output_15_25));
wire output_1_26, output_1_11, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_11), .y(output_0_26));
wire output_2_26, output_2_11, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_11), .y(output_1_26));
wire output_3_26, output_3_11, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_11), .y(output_2_26));
wire output_4_26, output_4_11, output_3_26;
mixer gate_output_3_26(.a(output_4_26), .b(output_4_11), .y(output_3_26));
wire output_5_26, output_5_11, output_4_26;
mixer gate_output_4_26(.a(output_5_26), .b(output_5_11), .y(output_4_26));
wire output_6_26, output_6_11, output_5_26;
mixer gate_output_5_26(.a(output_6_26), .b(output_6_11), .y(output_5_26));
wire output_7_26, output_7_11, output_6_26;
mixer gate_output_6_26(.a(output_7_26), .b(output_7_11), .y(output_6_26));
wire output_8_26, output_8_11, output_7_26;
mixer gate_output_7_26(.a(output_8_26), .b(output_8_11), .y(output_7_26));
wire output_9_26, output_9_11, output_8_26;
mixer gate_output_8_26(.a(output_9_26), .b(output_9_11), .y(output_8_26));
wire output_10_26, output_10_11, output_9_26;
mixer gate_output_9_26(.a(output_10_26), .b(output_10_11), .y(output_9_26));
wire output_11_26, output_11_11, output_10_26;
mixer gate_output_10_26(.a(output_11_26), .b(output_11_11), .y(output_10_26));
wire output_12_26, output_12_11, output_11_26;
mixer gate_output_11_26(.a(output_12_26), .b(output_12_11), .y(output_11_26));
wire output_13_26, output_13_11, output_12_26;
mixer gate_output_12_26(.a(output_13_26), .b(output_13_11), .y(output_12_26));
wire output_14_26, output_14_11, output_13_26;
mixer gate_output_13_26(.a(output_14_26), .b(output_14_11), .y(output_13_26));
wire output_15_26, output_15_11, output_14_26;
mixer gate_output_14_26(.a(output_15_26), .b(output_15_11), .y(output_14_26));
wire output_16_26, output_16_11, output_15_26;
mixer gate_output_15_26(.a(output_16_26), .b(output_16_11), .y(output_15_26));
wire output_1_27, output_1_12, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_12), .y(output_0_27));
wire output_2_27, output_2_12, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_12), .y(output_1_27));
wire output_3_27, output_3_12, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_12), .y(output_2_27));
wire output_4_27, output_4_12, output_3_27;
mixer gate_output_3_27(.a(output_4_27), .b(output_4_12), .y(output_3_27));
wire output_5_27, output_5_12, output_4_27;
mixer gate_output_4_27(.a(output_5_27), .b(output_5_12), .y(output_4_27));
wire output_6_27, output_6_12, output_5_27;
mixer gate_output_5_27(.a(output_6_27), .b(output_6_12), .y(output_5_27));
wire output_7_27, output_7_12, output_6_27;
mixer gate_output_6_27(.a(output_7_27), .b(output_7_12), .y(output_6_27));
wire output_8_27, output_8_12, output_7_27;
mixer gate_output_7_27(.a(output_8_27), .b(output_8_12), .y(output_7_27));
wire output_9_27, output_9_12, output_8_27;
mixer gate_output_8_27(.a(output_9_27), .b(output_9_12), .y(output_8_27));
wire output_10_27, output_10_12, output_9_27;
mixer gate_output_9_27(.a(output_10_27), .b(output_10_12), .y(output_9_27));
wire output_11_27, output_11_12, output_10_27;
mixer gate_output_10_27(.a(output_11_27), .b(output_11_12), .y(output_10_27));
wire output_12_27, output_12_12, output_11_27;
mixer gate_output_11_27(.a(output_12_27), .b(output_12_12), .y(output_11_27));
wire output_13_27, output_13_12, output_12_27;
mixer gate_output_12_27(.a(output_13_27), .b(output_13_12), .y(output_12_27));
wire output_14_27, output_14_12, output_13_27;
mixer gate_output_13_27(.a(output_14_27), .b(output_14_12), .y(output_13_27));
wire output_15_27, output_15_12, output_14_27;
mixer gate_output_14_27(.a(output_15_27), .b(output_15_12), .y(output_14_27));
wire output_16_27, output_16_12, output_15_27;
mixer gate_output_15_27(.a(output_16_27), .b(output_16_12), .y(output_15_27));
wire output_1_28, output_1_13, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_13), .y(output_0_28));
wire output_2_28, output_2_13, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_13), .y(output_1_28));
wire output_3_28, output_3_13, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_13), .y(output_2_28));
wire output_4_28, output_4_13, output_3_28;
mixer gate_output_3_28(.a(output_4_28), .b(output_4_13), .y(output_3_28));
wire output_5_28, output_5_13, output_4_28;
mixer gate_output_4_28(.a(output_5_28), .b(output_5_13), .y(output_4_28));
wire output_6_28, output_6_13, output_5_28;
mixer gate_output_5_28(.a(output_6_28), .b(output_6_13), .y(output_5_28));
wire output_7_28, output_7_13, output_6_28;
mixer gate_output_6_28(.a(output_7_28), .b(output_7_13), .y(output_6_28));
wire output_8_28, output_8_13, output_7_28;
mixer gate_output_7_28(.a(output_8_28), .b(output_8_13), .y(output_7_28));
wire output_9_28, output_9_13, output_8_28;
mixer gate_output_8_28(.a(output_9_28), .b(output_9_13), .y(output_8_28));
wire output_10_28, output_10_13, output_9_28;
mixer gate_output_9_28(.a(output_10_28), .b(output_10_13), .y(output_9_28));
wire output_11_28, output_11_13, output_10_28;
mixer gate_output_10_28(.a(output_11_28), .b(output_11_13), .y(output_10_28));
wire output_12_28, output_12_13, output_11_28;
mixer gate_output_11_28(.a(output_12_28), .b(output_12_13), .y(output_11_28));
wire output_13_28, output_13_13, output_12_28;
mixer gate_output_12_28(.a(output_13_28), .b(output_13_13), .y(output_12_28));
wire output_14_28, output_14_13, output_13_28;
mixer gate_output_13_28(.a(output_14_28), .b(output_14_13), .y(output_13_28));
wire output_15_28, output_15_13, output_14_28;
mixer gate_output_14_28(.a(output_15_28), .b(output_15_13), .y(output_14_28));
wire output_16_28, output_16_13, output_15_28;
mixer gate_output_15_28(.a(output_16_28), .b(output_16_13), .y(output_15_28));
wire output_1_29, output_1_14, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_14), .y(output_0_29));
wire output_2_29, output_2_14, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_14), .y(output_1_29));
wire output_3_29, output_3_14, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_14), .y(output_2_29));
wire output_4_29, output_4_14, output_3_29;
mixer gate_output_3_29(.a(output_4_29), .b(output_4_14), .y(output_3_29));
wire output_5_29, output_5_14, output_4_29;
mixer gate_output_4_29(.a(output_5_29), .b(output_5_14), .y(output_4_29));
wire output_6_29, output_6_14, output_5_29;
mixer gate_output_5_29(.a(output_6_29), .b(output_6_14), .y(output_5_29));
wire output_7_29, output_7_14, output_6_29;
mixer gate_output_6_29(.a(output_7_29), .b(output_7_14), .y(output_6_29));
wire output_8_29, output_8_14, output_7_29;
mixer gate_output_7_29(.a(output_8_29), .b(output_8_14), .y(output_7_29));
wire output_9_29, output_9_14, output_8_29;
mixer gate_output_8_29(.a(output_9_29), .b(output_9_14), .y(output_8_29));
wire output_10_29, output_10_14, output_9_29;
mixer gate_output_9_29(.a(output_10_29), .b(output_10_14), .y(output_9_29));
wire output_11_29, output_11_14, output_10_29;
mixer gate_output_10_29(.a(output_11_29), .b(output_11_14), .y(output_10_29));
wire output_12_29, output_12_14, output_11_29;
mixer gate_output_11_29(.a(output_12_29), .b(output_12_14), .y(output_11_29));
wire output_13_29, output_13_14, output_12_29;
mixer gate_output_12_29(.a(output_13_29), .b(output_13_14), .y(output_12_29));
wire output_14_29, output_14_14, output_13_29;
mixer gate_output_13_29(.a(output_14_29), .b(output_14_14), .y(output_13_29));
wire output_15_29, output_15_14, output_14_29;
mixer gate_output_14_29(.a(output_15_29), .b(output_15_14), .y(output_14_29));
wire output_16_29, output_16_14, output_15_29;
mixer gate_output_15_29(.a(output_16_29), .b(output_16_14), .y(output_15_29));
wire output_1_30, output_1_15, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_15), .y(output_0_30));
wire output_2_30, output_2_15, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_15), .y(output_1_30));
wire output_3_30, output_3_15, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_15), .y(output_2_30));
wire output_4_30, output_4_15, output_3_30;
mixer gate_output_3_30(.a(output_4_30), .b(output_4_15), .y(output_3_30));
wire output_5_30, output_5_15, output_4_30;
mixer gate_output_4_30(.a(output_5_30), .b(output_5_15), .y(output_4_30));
wire output_6_30, output_6_15, output_5_30;
mixer gate_output_5_30(.a(output_6_30), .b(output_6_15), .y(output_5_30));
wire output_7_30, output_7_15, output_6_30;
mixer gate_output_6_30(.a(output_7_30), .b(output_7_15), .y(output_6_30));
wire output_8_30, output_8_15, output_7_30;
mixer gate_output_7_30(.a(output_8_30), .b(output_8_15), .y(output_7_30));
wire output_9_30, output_9_15, output_8_30;
mixer gate_output_8_30(.a(output_9_30), .b(output_9_15), .y(output_8_30));
wire output_10_30, output_10_15, output_9_30;
mixer gate_output_9_30(.a(output_10_30), .b(output_10_15), .y(output_9_30));
wire output_11_30, output_11_15, output_10_30;
mixer gate_output_10_30(.a(output_11_30), .b(output_11_15), .y(output_10_30));
wire output_12_30, output_12_15, output_11_30;
mixer gate_output_11_30(.a(output_12_30), .b(output_12_15), .y(output_11_30));
wire output_13_30, output_13_15, output_12_30;
mixer gate_output_12_30(.a(output_13_30), .b(output_13_15), .y(output_12_30));
wire output_14_30, output_14_15, output_13_30;
mixer gate_output_13_30(.a(output_14_30), .b(output_14_15), .y(output_13_30));
wire output_15_30, output_15_15, output_14_30;
mixer gate_output_14_30(.a(output_15_30), .b(output_15_15), .y(output_14_30));
wire output_16_30, output_16_15, output_15_30;
mixer gate_output_15_30(.a(output_16_30), .b(output_16_15), .y(output_15_30));
wire output_1_31, output_1_0, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_0), .y(output_0_31));
wire output_2_31, output_2_0, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_0), .y(output_1_31));
wire output_3_31, output_3_0, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_0), .y(output_2_31));
wire output_4_31, output_4_0, output_3_31;
mixer gate_output_3_31(.a(output_4_31), .b(output_4_0), .y(output_3_31));
wire output_5_31, output_5_0, output_4_31;
mixer gate_output_4_31(.a(output_5_31), .b(output_5_0), .y(output_4_31));
wire output_6_31, output_6_0, output_5_31;
mixer gate_output_5_31(.a(output_6_31), .b(output_6_0), .y(output_5_31));
wire output_7_31, output_7_0, output_6_31;
mixer gate_output_6_31(.a(output_7_31), .b(output_7_0), .y(output_6_31));
wire output_8_31, output_8_0, output_7_31;
mixer gate_output_7_31(.a(output_8_31), .b(output_8_0), .y(output_7_31));
wire output_9_31, output_9_0, output_8_31;
mixer gate_output_8_31(.a(output_9_31), .b(output_9_0), .y(output_8_31));
wire output_10_31, output_10_0, output_9_31;
mixer gate_output_9_31(.a(output_10_31), .b(output_10_0), .y(output_9_31));
wire output_11_31, output_11_0, output_10_31;
mixer gate_output_10_31(.a(output_11_31), .b(output_11_0), .y(output_10_31));
wire output_12_31, output_12_0, output_11_31;
mixer gate_output_11_31(.a(output_12_31), .b(output_12_0), .y(output_11_31));
wire output_13_31, output_13_0, output_12_31;
mixer gate_output_12_31(.a(output_13_31), .b(output_13_0), .y(output_12_31));
wire output_14_31, output_14_0, output_13_31;
mixer gate_output_13_31(.a(output_14_31), .b(output_14_0), .y(output_13_31));
wire output_15_31, output_15_0, output_14_31;
mixer gate_output_14_31(.a(output_15_31), .b(output_15_0), .y(output_14_31));
wire output_16_31, output_16_0, output_15_31;
mixer gate_output_15_31(.a(output_16_31), .b(output_16_0), .y(output_15_31));
wire output_1_32, output_1_1, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_1), .y(output_0_32));
wire output_2_32, output_2_1, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_1), .y(output_1_32));
wire output_3_32, output_3_1, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_1), .y(output_2_32));
wire output_4_32, output_4_1, output_3_32;
mixer gate_output_3_32(.a(output_4_32), .b(output_4_1), .y(output_3_32));
wire output_5_32, output_5_1, output_4_32;
mixer gate_output_4_32(.a(output_5_32), .b(output_5_1), .y(output_4_32));
wire output_6_32, output_6_1, output_5_32;
mixer gate_output_5_32(.a(output_6_32), .b(output_6_1), .y(output_5_32));
wire output_7_32, output_7_1, output_6_32;
mixer gate_output_6_32(.a(output_7_32), .b(output_7_1), .y(output_6_32));
wire output_8_32, output_8_1, output_7_32;
mixer gate_output_7_32(.a(output_8_32), .b(output_8_1), .y(output_7_32));
wire output_9_32, output_9_1, output_8_32;
mixer gate_output_8_32(.a(output_9_32), .b(output_9_1), .y(output_8_32));
wire output_10_32, output_10_1, output_9_32;
mixer gate_output_9_32(.a(output_10_32), .b(output_10_1), .y(output_9_32));
wire output_11_32, output_11_1, output_10_32;
mixer gate_output_10_32(.a(output_11_32), .b(output_11_1), .y(output_10_32));
wire output_12_32, output_12_1, output_11_32;
mixer gate_output_11_32(.a(output_12_32), .b(output_12_1), .y(output_11_32));
wire output_13_32, output_13_1, output_12_32;
mixer gate_output_12_32(.a(output_13_32), .b(output_13_1), .y(output_12_32));
wire output_14_32, output_14_1, output_13_32;
mixer gate_output_13_32(.a(output_14_32), .b(output_14_1), .y(output_13_32));
wire output_15_32, output_15_1, output_14_32;
mixer gate_output_14_32(.a(output_15_32), .b(output_15_1), .y(output_14_32));
wire output_16_32, output_16_1, output_15_32;
mixer gate_output_15_32(.a(output_16_32), .b(output_16_1), .y(output_15_32));
wire output_1_33, output_1_2, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_2), .y(output_0_33));
wire output_2_33, output_2_2, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_2), .y(output_1_33));
wire output_3_33, output_3_2, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_2), .y(output_2_33));
wire output_4_33, output_4_2, output_3_33;
mixer gate_output_3_33(.a(output_4_33), .b(output_4_2), .y(output_3_33));
wire output_5_33, output_5_2, output_4_33;
mixer gate_output_4_33(.a(output_5_33), .b(output_5_2), .y(output_4_33));
wire output_6_33, output_6_2, output_5_33;
mixer gate_output_5_33(.a(output_6_33), .b(output_6_2), .y(output_5_33));
wire output_7_33, output_7_2, output_6_33;
mixer gate_output_6_33(.a(output_7_33), .b(output_7_2), .y(output_6_33));
wire output_8_33, output_8_2, output_7_33;
mixer gate_output_7_33(.a(output_8_33), .b(output_8_2), .y(output_7_33));
wire output_9_33, output_9_2, output_8_33;
mixer gate_output_8_33(.a(output_9_33), .b(output_9_2), .y(output_8_33));
wire output_10_33, output_10_2, output_9_33;
mixer gate_output_9_33(.a(output_10_33), .b(output_10_2), .y(output_9_33));
wire output_11_33, output_11_2, output_10_33;
mixer gate_output_10_33(.a(output_11_33), .b(output_11_2), .y(output_10_33));
wire output_12_33, output_12_2, output_11_33;
mixer gate_output_11_33(.a(output_12_33), .b(output_12_2), .y(output_11_33));
wire output_13_33, output_13_2, output_12_33;
mixer gate_output_12_33(.a(output_13_33), .b(output_13_2), .y(output_12_33));
wire output_14_33, output_14_2, output_13_33;
mixer gate_output_13_33(.a(output_14_33), .b(output_14_2), .y(output_13_33));
wire output_15_33, output_15_2, output_14_33;
mixer gate_output_14_33(.a(output_15_33), .b(output_15_2), .y(output_14_33));
wire output_16_33, output_16_2, output_15_33;
mixer gate_output_15_33(.a(output_16_33), .b(output_16_2), .y(output_15_33));
wire output_1_34, output_1_3, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_3), .y(output_0_34));
wire output_2_34, output_2_3, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_3), .y(output_1_34));
wire output_3_34, output_3_3, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_3), .y(output_2_34));
wire output_4_34, output_4_3, output_3_34;
mixer gate_output_3_34(.a(output_4_34), .b(output_4_3), .y(output_3_34));
wire output_5_34, output_5_3, output_4_34;
mixer gate_output_4_34(.a(output_5_34), .b(output_5_3), .y(output_4_34));
wire output_6_34, output_6_3, output_5_34;
mixer gate_output_5_34(.a(output_6_34), .b(output_6_3), .y(output_5_34));
wire output_7_34, output_7_3, output_6_34;
mixer gate_output_6_34(.a(output_7_34), .b(output_7_3), .y(output_6_34));
wire output_8_34, output_8_3, output_7_34;
mixer gate_output_7_34(.a(output_8_34), .b(output_8_3), .y(output_7_34));
wire output_9_34, output_9_3, output_8_34;
mixer gate_output_8_34(.a(output_9_34), .b(output_9_3), .y(output_8_34));
wire output_10_34, output_10_3, output_9_34;
mixer gate_output_9_34(.a(output_10_34), .b(output_10_3), .y(output_9_34));
wire output_11_34, output_11_3, output_10_34;
mixer gate_output_10_34(.a(output_11_34), .b(output_11_3), .y(output_10_34));
wire output_12_34, output_12_3, output_11_34;
mixer gate_output_11_34(.a(output_12_34), .b(output_12_3), .y(output_11_34));
wire output_13_34, output_13_3, output_12_34;
mixer gate_output_12_34(.a(output_13_34), .b(output_13_3), .y(output_12_34));
wire output_14_34, output_14_3, output_13_34;
mixer gate_output_13_34(.a(output_14_34), .b(output_14_3), .y(output_13_34));
wire output_15_34, output_15_3, output_14_34;
mixer gate_output_14_34(.a(output_15_34), .b(output_15_3), .y(output_14_34));
wire output_16_34, output_16_3, output_15_34;
mixer gate_output_15_34(.a(output_16_34), .b(output_16_3), .y(output_15_34));
wire output_1_35, output_1_4, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_4), .y(output_0_35));
wire output_2_35, output_2_4, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_4), .y(output_1_35));
wire output_3_35, output_3_4, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_4), .y(output_2_35));
wire output_4_35, output_4_4, output_3_35;
mixer gate_output_3_35(.a(output_4_35), .b(output_4_4), .y(output_3_35));
wire output_5_35, output_5_4, output_4_35;
mixer gate_output_4_35(.a(output_5_35), .b(output_5_4), .y(output_4_35));
wire output_6_35, output_6_4, output_5_35;
mixer gate_output_5_35(.a(output_6_35), .b(output_6_4), .y(output_5_35));
wire output_7_35, output_7_4, output_6_35;
mixer gate_output_6_35(.a(output_7_35), .b(output_7_4), .y(output_6_35));
wire output_8_35, output_8_4, output_7_35;
mixer gate_output_7_35(.a(output_8_35), .b(output_8_4), .y(output_7_35));
wire output_9_35, output_9_4, output_8_35;
mixer gate_output_8_35(.a(output_9_35), .b(output_9_4), .y(output_8_35));
wire output_10_35, output_10_4, output_9_35;
mixer gate_output_9_35(.a(output_10_35), .b(output_10_4), .y(output_9_35));
wire output_11_35, output_11_4, output_10_35;
mixer gate_output_10_35(.a(output_11_35), .b(output_11_4), .y(output_10_35));
wire output_12_35, output_12_4, output_11_35;
mixer gate_output_11_35(.a(output_12_35), .b(output_12_4), .y(output_11_35));
wire output_13_35, output_13_4, output_12_35;
mixer gate_output_12_35(.a(output_13_35), .b(output_13_4), .y(output_12_35));
wire output_14_35, output_14_4, output_13_35;
mixer gate_output_13_35(.a(output_14_35), .b(output_14_4), .y(output_13_35));
wire output_15_35, output_15_4, output_14_35;
mixer gate_output_14_35(.a(output_15_35), .b(output_15_4), .y(output_14_35));
wire output_16_35, output_16_4, output_15_35;
mixer gate_output_15_35(.a(output_16_35), .b(output_16_4), .y(output_15_35));
wire output_1_36, output_1_5, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_5), .y(output_0_36));
wire output_2_36, output_2_5, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_5), .y(output_1_36));
wire output_3_36, output_3_5, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_5), .y(output_2_36));
wire output_4_36, output_4_5, output_3_36;
mixer gate_output_3_36(.a(output_4_36), .b(output_4_5), .y(output_3_36));
wire output_5_36, output_5_5, output_4_36;
mixer gate_output_4_36(.a(output_5_36), .b(output_5_5), .y(output_4_36));
wire output_6_36, output_6_5, output_5_36;
mixer gate_output_5_36(.a(output_6_36), .b(output_6_5), .y(output_5_36));
wire output_7_36, output_7_5, output_6_36;
mixer gate_output_6_36(.a(output_7_36), .b(output_7_5), .y(output_6_36));
wire output_8_36, output_8_5, output_7_36;
mixer gate_output_7_36(.a(output_8_36), .b(output_8_5), .y(output_7_36));
wire output_9_36, output_9_5, output_8_36;
mixer gate_output_8_36(.a(output_9_36), .b(output_9_5), .y(output_8_36));
wire output_10_36, output_10_5, output_9_36;
mixer gate_output_9_36(.a(output_10_36), .b(output_10_5), .y(output_9_36));
wire output_11_36, output_11_5, output_10_36;
mixer gate_output_10_36(.a(output_11_36), .b(output_11_5), .y(output_10_36));
wire output_12_36, output_12_5, output_11_36;
mixer gate_output_11_36(.a(output_12_36), .b(output_12_5), .y(output_11_36));
wire output_13_36, output_13_5, output_12_36;
mixer gate_output_12_36(.a(output_13_36), .b(output_13_5), .y(output_12_36));
wire output_14_36, output_14_5, output_13_36;
mixer gate_output_13_36(.a(output_14_36), .b(output_14_5), .y(output_13_36));
wire output_15_36, output_15_5, output_14_36;
mixer gate_output_14_36(.a(output_15_36), .b(output_15_5), .y(output_14_36));
wire output_16_36, output_16_5, output_15_36;
mixer gate_output_15_36(.a(output_16_36), .b(output_16_5), .y(output_15_36));
wire output_1_37, output_1_6, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_6), .y(output_0_37));
wire output_2_37, output_2_6, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_6), .y(output_1_37));
wire output_3_37, output_3_6, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_6), .y(output_2_37));
wire output_4_37, output_4_6, output_3_37;
mixer gate_output_3_37(.a(output_4_37), .b(output_4_6), .y(output_3_37));
wire output_5_37, output_5_6, output_4_37;
mixer gate_output_4_37(.a(output_5_37), .b(output_5_6), .y(output_4_37));
wire output_6_37, output_6_6, output_5_37;
mixer gate_output_5_37(.a(output_6_37), .b(output_6_6), .y(output_5_37));
wire output_7_37, output_7_6, output_6_37;
mixer gate_output_6_37(.a(output_7_37), .b(output_7_6), .y(output_6_37));
wire output_8_37, output_8_6, output_7_37;
mixer gate_output_7_37(.a(output_8_37), .b(output_8_6), .y(output_7_37));
wire output_9_37, output_9_6, output_8_37;
mixer gate_output_8_37(.a(output_9_37), .b(output_9_6), .y(output_8_37));
wire output_10_37, output_10_6, output_9_37;
mixer gate_output_9_37(.a(output_10_37), .b(output_10_6), .y(output_9_37));
wire output_11_37, output_11_6, output_10_37;
mixer gate_output_10_37(.a(output_11_37), .b(output_11_6), .y(output_10_37));
wire output_12_37, output_12_6, output_11_37;
mixer gate_output_11_37(.a(output_12_37), .b(output_12_6), .y(output_11_37));
wire output_13_37, output_13_6, output_12_37;
mixer gate_output_12_37(.a(output_13_37), .b(output_13_6), .y(output_12_37));
wire output_14_37, output_14_6, output_13_37;
mixer gate_output_13_37(.a(output_14_37), .b(output_14_6), .y(output_13_37));
wire output_15_37, output_15_6, output_14_37;
mixer gate_output_14_37(.a(output_15_37), .b(output_15_6), .y(output_14_37));
wire output_16_37, output_16_6, output_15_37;
mixer gate_output_15_37(.a(output_16_37), .b(output_16_6), .y(output_15_37));
wire output_1_38, output_1_7, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_7), .y(output_0_38));
wire output_2_38, output_2_7, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_7), .y(output_1_38));
wire output_3_38, output_3_7, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_7), .y(output_2_38));
wire output_4_38, output_4_7, output_3_38;
mixer gate_output_3_38(.a(output_4_38), .b(output_4_7), .y(output_3_38));
wire output_5_38, output_5_7, output_4_38;
mixer gate_output_4_38(.a(output_5_38), .b(output_5_7), .y(output_4_38));
wire output_6_38, output_6_7, output_5_38;
mixer gate_output_5_38(.a(output_6_38), .b(output_6_7), .y(output_5_38));
wire output_7_38, output_7_7, output_6_38;
mixer gate_output_6_38(.a(output_7_38), .b(output_7_7), .y(output_6_38));
wire output_8_38, output_8_7, output_7_38;
mixer gate_output_7_38(.a(output_8_38), .b(output_8_7), .y(output_7_38));
wire output_9_38, output_9_7, output_8_38;
mixer gate_output_8_38(.a(output_9_38), .b(output_9_7), .y(output_8_38));
wire output_10_38, output_10_7, output_9_38;
mixer gate_output_9_38(.a(output_10_38), .b(output_10_7), .y(output_9_38));
wire output_11_38, output_11_7, output_10_38;
mixer gate_output_10_38(.a(output_11_38), .b(output_11_7), .y(output_10_38));
wire output_12_38, output_12_7, output_11_38;
mixer gate_output_11_38(.a(output_12_38), .b(output_12_7), .y(output_11_38));
wire output_13_38, output_13_7, output_12_38;
mixer gate_output_12_38(.a(output_13_38), .b(output_13_7), .y(output_12_38));
wire output_14_38, output_14_7, output_13_38;
mixer gate_output_13_38(.a(output_14_38), .b(output_14_7), .y(output_13_38));
wire output_15_38, output_15_7, output_14_38;
mixer gate_output_14_38(.a(output_15_38), .b(output_15_7), .y(output_14_38));
wire output_16_38, output_16_7, output_15_38;
mixer gate_output_15_38(.a(output_16_38), .b(output_16_7), .y(output_15_38));
wire output_1_39, output_1_8, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_8), .y(output_0_39));
wire output_2_39, output_2_8, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_8), .y(output_1_39));
wire output_3_39, output_3_8, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_8), .y(output_2_39));
wire output_4_39, output_4_8, output_3_39;
mixer gate_output_3_39(.a(output_4_39), .b(output_4_8), .y(output_3_39));
wire output_5_39, output_5_8, output_4_39;
mixer gate_output_4_39(.a(output_5_39), .b(output_5_8), .y(output_4_39));
wire output_6_39, output_6_8, output_5_39;
mixer gate_output_5_39(.a(output_6_39), .b(output_6_8), .y(output_5_39));
wire output_7_39, output_7_8, output_6_39;
mixer gate_output_6_39(.a(output_7_39), .b(output_7_8), .y(output_6_39));
wire output_8_39, output_8_8, output_7_39;
mixer gate_output_7_39(.a(output_8_39), .b(output_8_8), .y(output_7_39));
wire output_9_39, output_9_8, output_8_39;
mixer gate_output_8_39(.a(output_9_39), .b(output_9_8), .y(output_8_39));
wire output_10_39, output_10_8, output_9_39;
mixer gate_output_9_39(.a(output_10_39), .b(output_10_8), .y(output_9_39));
wire output_11_39, output_11_8, output_10_39;
mixer gate_output_10_39(.a(output_11_39), .b(output_11_8), .y(output_10_39));
wire output_12_39, output_12_8, output_11_39;
mixer gate_output_11_39(.a(output_12_39), .b(output_12_8), .y(output_11_39));
wire output_13_39, output_13_8, output_12_39;
mixer gate_output_12_39(.a(output_13_39), .b(output_13_8), .y(output_12_39));
wire output_14_39, output_14_8, output_13_39;
mixer gate_output_13_39(.a(output_14_39), .b(output_14_8), .y(output_13_39));
wire output_15_39, output_15_8, output_14_39;
mixer gate_output_14_39(.a(output_15_39), .b(output_15_8), .y(output_14_39));
wire output_16_39, output_16_8, output_15_39;
mixer gate_output_15_39(.a(output_16_39), .b(output_16_8), .y(output_15_39));
wire output_1_40, output_1_9, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_9), .y(output_0_40));
wire output_2_40, output_2_9, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_9), .y(output_1_40));
wire output_3_40, output_3_9, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_9), .y(output_2_40));
wire output_4_40, output_4_9, output_3_40;
mixer gate_output_3_40(.a(output_4_40), .b(output_4_9), .y(output_3_40));
wire output_5_40, output_5_9, output_4_40;
mixer gate_output_4_40(.a(output_5_40), .b(output_5_9), .y(output_4_40));
wire output_6_40, output_6_9, output_5_40;
mixer gate_output_5_40(.a(output_6_40), .b(output_6_9), .y(output_5_40));
wire output_7_40, output_7_9, output_6_40;
mixer gate_output_6_40(.a(output_7_40), .b(output_7_9), .y(output_6_40));
wire output_8_40, output_8_9, output_7_40;
mixer gate_output_7_40(.a(output_8_40), .b(output_8_9), .y(output_7_40));
wire output_9_40, output_9_9, output_8_40;
mixer gate_output_8_40(.a(output_9_40), .b(output_9_9), .y(output_8_40));
wire output_10_40, output_10_9, output_9_40;
mixer gate_output_9_40(.a(output_10_40), .b(output_10_9), .y(output_9_40));
wire output_11_40, output_11_9, output_10_40;
mixer gate_output_10_40(.a(output_11_40), .b(output_11_9), .y(output_10_40));
wire output_12_40, output_12_9, output_11_40;
mixer gate_output_11_40(.a(output_12_40), .b(output_12_9), .y(output_11_40));
wire output_13_40, output_13_9, output_12_40;
mixer gate_output_12_40(.a(output_13_40), .b(output_13_9), .y(output_12_40));
wire output_14_40, output_14_9, output_13_40;
mixer gate_output_13_40(.a(output_14_40), .b(output_14_9), .y(output_13_40));
wire output_15_40, output_15_9, output_14_40;
mixer gate_output_14_40(.a(output_15_40), .b(output_15_9), .y(output_14_40));
wire output_16_40, output_16_9, output_15_40;
mixer gate_output_15_40(.a(output_16_40), .b(output_16_9), .y(output_15_40));
wire output_1_41, output_1_10, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_10), .y(output_0_41));
wire output_2_41, output_2_10, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_10), .y(output_1_41));
wire output_3_41, output_3_10, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_10), .y(output_2_41));
wire output_4_41, output_4_10, output_3_41;
mixer gate_output_3_41(.a(output_4_41), .b(output_4_10), .y(output_3_41));
wire output_5_41, output_5_10, output_4_41;
mixer gate_output_4_41(.a(output_5_41), .b(output_5_10), .y(output_4_41));
wire output_6_41, output_6_10, output_5_41;
mixer gate_output_5_41(.a(output_6_41), .b(output_6_10), .y(output_5_41));
wire output_7_41, output_7_10, output_6_41;
mixer gate_output_6_41(.a(output_7_41), .b(output_7_10), .y(output_6_41));
wire output_8_41, output_8_10, output_7_41;
mixer gate_output_7_41(.a(output_8_41), .b(output_8_10), .y(output_7_41));
wire output_9_41, output_9_10, output_8_41;
mixer gate_output_8_41(.a(output_9_41), .b(output_9_10), .y(output_8_41));
wire output_10_41, output_10_10, output_9_41;
mixer gate_output_9_41(.a(output_10_41), .b(output_10_10), .y(output_9_41));
wire output_11_41, output_11_10, output_10_41;
mixer gate_output_10_41(.a(output_11_41), .b(output_11_10), .y(output_10_41));
wire output_12_41, output_12_10, output_11_41;
mixer gate_output_11_41(.a(output_12_41), .b(output_12_10), .y(output_11_41));
wire output_13_41, output_13_10, output_12_41;
mixer gate_output_12_41(.a(output_13_41), .b(output_13_10), .y(output_12_41));
wire output_14_41, output_14_10, output_13_41;
mixer gate_output_13_41(.a(output_14_41), .b(output_14_10), .y(output_13_41));
wire output_15_41, output_15_10, output_14_41;
mixer gate_output_14_41(.a(output_15_41), .b(output_15_10), .y(output_14_41));
wire output_16_41, output_16_10, output_15_41;
mixer gate_output_15_41(.a(output_16_41), .b(output_16_10), .y(output_15_41));
wire output_1_42, output_1_11, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_11), .y(output_0_42));
wire output_2_42, output_2_11, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_11), .y(output_1_42));
wire output_3_42, output_3_11, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_11), .y(output_2_42));
wire output_4_42, output_4_11, output_3_42;
mixer gate_output_3_42(.a(output_4_42), .b(output_4_11), .y(output_3_42));
wire output_5_42, output_5_11, output_4_42;
mixer gate_output_4_42(.a(output_5_42), .b(output_5_11), .y(output_4_42));
wire output_6_42, output_6_11, output_5_42;
mixer gate_output_5_42(.a(output_6_42), .b(output_6_11), .y(output_5_42));
wire output_7_42, output_7_11, output_6_42;
mixer gate_output_6_42(.a(output_7_42), .b(output_7_11), .y(output_6_42));
wire output_8_42, output_8_11, output_7_42;
mixer gate_output_7_42(.a(output_8_42), .b(output_8_11), .y(output_7_42));
wire output_9_42, output_9_11, output_8_42;
mixer gate_output_8_42(.a(output_9_42), .b(output_9_11), .y(output_8_42));
wire output_10_42, output_10_11, output_9_42;
mixer gate_output_9_42(.a(output_10_42), .b(output_10_11), .y(output_9_42));
wire output_11_42, output_11_11, output_10_42;
mixer gate_output_10_42(.a(output_11_42), .b(output_11_11), .y(output_10_42));
wire output_12_42, output_12_11, output_11_42;
mixer gate_output_11_42(.a(output_12_42), .b(output_12_11), .y(output_11_42));
wire output_13_42, output_13_11, output_12_42;
mixer gate_output_12_42(.a(output_13_42), .b(output_13_11), .y(output_12_42));
wire output_14_42, output_14_11, output_13_42;
mixer gate_output_13_42(.a(output_14_42), .b(output_14_11), .y(output_13_42));
wire output_15_42, output_15_11, output_14_42;
mixer gate_output_14_42(.a(output_15_42), .b(output_15_11), .y(output_14_42));
wire output_16_42, output_16_11, output_15_42;
mixer gate_output_15_42(.a(output_16_42), .b(output_16_11), .y(output_15_42));
wire output_1_43, output_1_12, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_12), .y(output_0_43));
wire output_2_43, output_2_12, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_12), .y(output_1_43));
wire output_3_43, output_3_12, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_12), .y(output_2_43));
wire output_4_43, output_4_12, output_3_43;
mixer gate_output_3_43(.a(output_4_43), .b(output_4_12), .y(output_3_43));
wire output_5_43, output_5_12, output_4_43;
mixer gate_output_4_43(.a(output_5_43), .b(output_5_12), .y(output_4_43));
wire output_6_43, output_6_12, output_5_43;
mixer gate_output_5_43(.a(output_6_43), .b(output_6_12), .y(output_5_43));
wire output_7_43, output_7_12, output_6_43;
mixer gate_output_6_43(.a(output_7_43), .b(output_7_12), .y(output_6_43));
wire output_8_43, output_8_12, output_7_43;
mixer gate_output_7_43(.a(output_8_43), .b(output_8_12), .y(output_7_43));
wire output_9_43, output_9_12, output_8_43;
mixer gate_output_8_43(.a(output_9_43), .b(output_9_12), .y(output_8_43));
wire output_10_43, output_10_12, output_9_43;
mixer gate_output_9_43(.a(output_10_43), .b(output_10_12), .y(output_9_43));
wire output_11_43, output_11_12, output_10_43;
mixer gate_output_10_43(.a(output_11_43), .b(output_11_12), .y(output_10_43));
wire output_12_43, output_12_12, output_11_43;
mixer gate_output_11_43(.a(output_12_43), .b(output_12_12), .y(output_11_43));
wire output_13_43, output_13_12, output_12_43;
mixer gate_output_12_43(.a(output_13_43), .b(output_13_12), .y(output_12_43));
wire output_14_43, output_14_12, output_13_43;
mixer gate_output_13_43(.a(output_14_43), .b(output_14_12), .y(output_13_43));
wire output_15_43, output_15_12, output_14_43;
mixer gate_output_14_43(.a(output_15_43), .b(output_15_12), .y(output_14_43));
wire output_16_43, output_16_12, output_15_43;
mixer gate_output_15_43(.a(output_16_43), .b(output_16_12), .y(output_15_43));
wire output_1_44, output_1_13, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_13), .y(output_0_44));
wire output_2_44, output_2_13, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_13), .y(output_1_44));
wire output_3_44, output_3_13, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_13), .y(output_2_44));
wire output_4_44, output_4_13, output_3_44;
mixer gate_output_3_44(.a(output_4_44), .b(output_4_13), .y(output_3_44));
wire output_5_44, output_5_13, output_4_44;
mixer gate_output_4_44(.a(output_5_44), .b(output_5_13), .y(output_4_44));
wire output_6_44, output_6_13, output_5_44;
mixer gate_output_5_44(.a(output_6_44), .b(output_6_13), .y(output_5_44));
wire output_7_44, output_7_13, output_6_44;
mixer gate_output_6_44(.a(output_7_44), .b(output_7_13), .y(output_6_44));
wire output_8_44, output_8_13, output_7_44;
mixer gate_output_7_44(.a(output_8_44), .b(output_8_13), .y(output_7_44));
wire output_9_44, output_9_13, output_8_44;
mixer gate_output_8_44(.a(output_9_44), .b(output_9_13), .y(output_8_44));
wire output_10_44, output_10_13, output_9_44;
mixer gate_output_9_44(.a(output_10_44), .b(output_10_13), .y(output_9_44));
wire output_11_44, output_11_13, output_10_44;
mixer gate_output_10_44(.a(output_11_44), .b(output_11_13), .y(output_10_44));
wire output_12_44, output_12_13, output_11_44;
mixer gate_output_11_44(.a(output_12_44), .b(output_12_13), .y(output_11_44));
wire output_13_44, output_13_13, output_12_44;
mixer gate_output_12_44(.a(output_13_44), .b(output_13_13), .y(output_12_44));
wire output_14_44, output_14_13, output_13_44;
mixer gate_output_13_44(.a(output_14_44), .b(output_14_13), .y(output_13_44));
wire output_15_44, output_15_13, output_14_44;
mixer gate_output_14_44(.a(output_15_44), .b(output_15_13), .y(output_14_44));
wire output_16_44, output_16_13, output_15_44;
mixer gate_output_15_44(.a(output_16_44), .b(output_16_13), .y(output_15_44));
wire output_1_45, output_1_14, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_14), .y(output_0_45));
wire output_2_45, output_2_14, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_14), .y(output_1_45));
wire output_3_45, output_3_14, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_14), .y(output_2_45));
wire output_4_45, output_4_14, output_3_45;
mixer gate_output_3_45(.a(output_4_45), .b(output_4_14), .y(output_3_45));
wire output_5_45, output_5_14, output_4_45;
mixer gate_output_4_45(.a(output_5_45), .b(output_5_14), .y(output_4_45));
wire output_6_45, output_6_14, output_5_45;
mixer gate_output_5_45(.a(output_6_45), .b(output_6_14), .y(output_5_45));
wire output_7_45, output_7_14, output_6_45;
mixer gate_output_6_45(.a(output_7_45), .b(output_7_14), .y(output_6_45));
wire output_8_45, output_8_14, output_7_45;
mixer gate_output_7_45(.a(output_8_45), .b(output_8_14), .y(output_7_45));
wire output_9_45, output_9_14, output_8_45;
mixer gate_output_8_45(.a(output_9_45), .b(output_9_14), .y(output_8_45));
wire output_10_45, output_10_14, output_9_45;
mixer gate_output_9_45(.a(output_10_45), .b(output_10_14), .y(output_9_45));
wire output_11_45, output_11_14, output_10_45;
mixer gate_output_10_45(.a(output_11_45), .b(output_11_14), .y(output_10_45));
wire output_12_45, output_12_14, output_11_45;
mixer gate_output_11_45(.a(output_12_45), .b(output_12_14), .y(output_11_45));
wire output_13_45, output_13_14, output_12_45;
mixer gate_output_12_45(.a(output_13_45), .b(output_13_14), .y(output_12_45));
wire output_14_45, output_14_14, output_13_45;
mixer gate_output_13_45(.a(output_14_45), .b(output_14_14), .y(output_13_45));
wire output_15_45, output_15_14, output_14_45;
mixer gate_output_14_45(.a(output_15_45), .b(output_15_14), .y(output_14_45));
wire output_16_45, output_16_14, output_15_45;
mixer gate_output_15_45(.a(output_16_45), .b(output_16_14), .y(output_15_45));
wire output_1_46, output_1_15, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_15), .y(output_0_46));
wire output_2_46, output_2_15, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_15), .y(output_1_46));
wire output_3_46, output_3_15, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_15), .y(output_2_46));
wire output_4_46, output_4_15, output_3_46;
mixer gate_output_3_46(.a(output_4_46), .b(output_4_15), .y(output_3_46));
wire output_5_46, output_5_15, output_4_46;
mixer gate_output_4_46(.a(output_5_46), .b(output_5_15), .y(output_4_46));
wire output_6_46, output_6_15, output_5_46;
mixer gate_output_5_46(.a(output_6_46), .b(output_6_15), .y(output_5_46));
wire output_7_46, output_7_15, output_6_46;
mixer gate_output_6_46(.a(output_7_46), .b(output_7_15), .y(output_6_46));
wire output_8_46, output_8_15, output_7_46;
mixer gate_output_7_46(.a(output_8_46), .b(output_8_15), .y(output_7_46));
wire output_9_46, output_9_15, output_8_46;
mixer gate_output_8_46(.a(output_9_46), .b(output_9_15), .y(output_8_46));
wire output_10_46, output_10_15, output_9_46;
mixer gate_output_9_46(.a(output_10_46), .b(output_10_15), .y(output_9_46));
wire output_11_46, output_11_15, output_10_46;
mixer gate_output_10_46(.a(output_11_46), .b(output_11_15), .y(output_10_46));
wire output_12_46, output_12_15, output_11_46;
mixer gate_output_11_46(.a(output_12_46), .b(output_12_15), .y(output_11_46));
wire output_13_46, output_13_15, output_12_46;
mixer gate_output_12_46(.a(output_13_46), .b(output_13_15), .y(output_12_46));
wire output_14_46, output_14_15, output_13_46;
mixer gate_output_13_46(.a(output_14_46), .b(output_14_15), .y(output_13_46));
wire output_15_46, output_15_15, output_14_46;
mixer gate_output_14_46(.a(output_15_46), .b(output_15_15), .y(output_14_46));
wire output_16_46, output_16_15, output_15_46;
mixer gate_output_15_46(.a(output_16_46), .b(output_16_15), .y(output_15_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_4_47, output_4_0, output_3_47;
mixer gate_output_3_47(.a(output_4_47), .b(output_4_0), .y(output_3_47));
wire output_5_47, output_5_0, output_4_47;
mixer gate_output_4_47(.a(output_5_47), .b(output_5_0), .y(output_4_47));
wire output_6_47, output_6_0, output_5_47;
mixer gate_output_5_47(.a(output_6_47), .b(output_6_0), .y(output_5_47));
wire output_7_47, output_7_0, output_6_47;
mixer gate_output_6_47(.a(output_7_47), .b(output_7_0), .y(output_6_47));
wire output_8_47, output_8_0, output_7_47;
mixer gate_output_7_47(.a(output_8_47), .b(output_8_0), .y(output_7_47));
wire output_9_47, output_9_0, output_8_47;
mixer gate_output_8_47(.a(output_9_47), .b(output_9_0), .y(output_8_47));
wire output_10_47, output_10_0, output_9_47;
mixer gate_output_9_47(.a(output_10_47), .b(output_10_0), .y(output_9_47));
wire output_11_47, output_11_0, output_10_47;
mixer gate_output_10_47(.a(output_11_47), .b(output_11_0), .y(output_10_47));
wire output_12_47, output_12_0, output_11_47;
mixer gate_output_11_47(.a(output_12_47), .b(output_12_0), .y(output_11_47));
wire output_13_47, output_13_0, output_12_47;
mixer gate_output_12_47(.a(output_13_47), .b(output_13_0), .y(output_12_47));
wire output_14_47, output_14_0, output_13_47;
mixer gate_output_13_47(.a(output_14_47), .b(output_14_0), .y(output_13_47));
wire output_15_47, output_15_0, output_14_47;
mixer gate_output_14_47(.a(output_15_47), .b(output_15_0), .y(output_14_47));
wire output_16_47, output_16_0, output_15_47;
mixer gate_output_15_47(.a(output_16_47), .b(output_16_0), .y(output_15_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_4_48, output_4_1, output_3_48;
mixer gate_output_3_48(.a(output_4_48), .b(output_4_1), .y(output_3_48));
wire output_5_48, output_5_1, output_4_48;
mixer gate_output_4_48(.a(output_5_48), .b(output_5_1), .y(output_4_48));
wire output_6_48, output_6_1, output_5_48;
mixer gate_output_5_48(.a(output_6_48), .b(output_6_1), .y(output_5_48));
wire output_7_48, output_7_1, output_6_48;
mixer gate_output_6_48(.a(output_7_48), .b(output_7_1), .y(output_6_48));
wire output_8_48, output_8_1, output_7_48;
mixer gate_output_7_48(.a(output_8_48), .b(output_8_1), .y(output_7_48));
wire output_9_48, output_9_1, output_8_48;
mixer gate_output_8_48(.a(output_9_48), .b(output_9_1), .y(output_8_48));
wire output_10_48, output_10_1, output_9_48;
mixer gate_output_9_48(.a(output_10_48), .b(output_10_1), .y(output_9_48));
wire output_11_48, output_11_1, output_10_48;
mixer gate_output_10_48(.a(output_11_48), .b(output_11_1), .y(output_10_48));
wire output_12_48, output_12_1, output_11_48;
mixer gate_output_11_48(.a(output_12_48), .b(output_12_1), .y(output_11_48));
wire output_13_48, output_13_1, output_12_48;
mixer gate_output_12_48(.a(output_13_48), .b(output_13_1), .y(output_12_48));
wire output_14_48, output_14_1, output_13_48;
mixer gate_output_13_48(.a(output_14_48), .b(output_14_1), .y(output_13_48));
wire output_15_48, output_15_1, output_14_48;
mixer gate_output_14_48(.a(output_15_48), .b(output_15_1), .y(output_14_48));
wire output_16_48, output_16_1, output_15_48;
mixer gate_output_15_48(.a(output_16_48), .b(output_16_1), .y(output_15_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_4_49, output_4_2, output_3_49;
mixer gate_output_3_49(.a(output_4_49), .b(output_4_2), .y(output_3_49));
wire output_5_49, output_5_2, output_4_49;
mixer gate_output_4_49(.a(output_5_49), .b(output_5_2), .y(output_4_49));
wire output_6_49, output_6_2, output_5_49;
mixer gate_output_5_49(.a(output_6_49), .b(output_6_2), .y(output_5_49));
wire output_7_49, output_7_2, output_6_49;
mixer gate_output_6_49(.a(output_7_49), .b(output_7_2), .y(output_6_49));
wire output_8_49, output_8_2, output_7_49;
mixer gate_output_7_49(.a(output_8_49), .b(output_8_2), .y(output_7_49));
wire output_9_49, output_9_2, output_8_49;
mixer gate_output_8_49(.a(output_9_49), .b(output_9_2), .y(output_8_49));
wire output_10_49, output_10_2, output_9_49;
mixer gate_output_9_49(.a(output_10_49), .b(output_10_2), .y(output_9_49));
wire output_11_49, output_11_2, output_10_49;
mixer gate_output_10_49(.a(output_11_49), .b(output_11_2), .y(output_10_49));
wire output_12_49, output_12_2, output_11_49;
mixer gate_output_11_49(.a(output_12_49), .b(output_12_2), .y(output_11_49));
wire output_13_49, output_13_2, output_12_49;
mixer gate_output_12_49(.a(output_13_49), .b(output_13_2), .y(output_12_49));
wire output_14_49, output_14_2, output_13_49;
mixer gate_output_13_49(.a(output_14_49), .b(output_14_2), .y(output_13_49));
wire output_15_49, output_15_2, output_14_49;
mixer gate_output_14_49(.a(output_15_49), .b(output_15_2), .y(output_14_49));
wire output_16_49, output_16_2, output_15_49;
mixer gate_output_15_49(.a(output_16_49), .b(output_16_2), .y(output_15_49));
wire output_1_50, output_1_3, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_3), .y(output_0_50));
wire output_2_50, output_2_3, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_3), .y(output_1_50));
wire output_3_50, output_3_3, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_3), .y(output_2_50));
wire output_4_50, output_4_3, output_3_50;
mixer gate_output_3_50(.a(output_4_50), .b(output_4_3), .y(output_3_50));
wire output_5_50, output_5_3, output_4_50;
mixer gate_output_4_50(.a(output_5_50), .b(output_5_3), .y(output_4_50));
wire output_6_50, output_6_3, output_5_50;
mixer gate_output_5_50(.a(output_6_50), .b(output_6_3), .y(output_5_50));
wire output_7_50, output_7_3, output_6_50;
mixer gate_output_6_50(.a(output_7_50), .b(output_7_3), .y(output_6_50));
wire output_8_50, output_8_3, output_7_50;
mixer gate_output_7_50(.a(output_8_50), .b(output_8_3), .y(output_7_50));
wire output_9_50, output_9_3, output_8_50;
mixer gate_output_8_50(.a(output_9_50), .b(output_9_3), .y(output_8_50));
wire output_10_50, output_10_3, output_9_50;
mixer gate_output_9_50(.a(output_10_50), .b(output_10_3), .y(output_9_50));
wire output_11_50, output_11_3, output_10_50;
mixer gate_output_10_50(.a(output_11_50), .b(output_11_3), .y(output_10_50));
wire output_12_50, output_12_3, output_11_50;
mixer gate_output_11_50(.a(output_12_50), .b(output_12_3), .y(output_11_50));
wire output_13_50, output_13_3, output_12_50;
mixer gate_output_12_50(.a(output_13_50), .b(output_13_3), .y(output_12_50));
wire output_14_50, output_14_3, output_13_50;
mixer gate_output_13_50(.a(output_14_50), .b(output_14_3), .y(output_13_50));
wire output_15_50, output_15_3, output_14_50;
mixer gate_output_14_50(.a(output_15_50), .b(output_15_3), .y(output_14_50));
wire output_16_50, output_16_3, output_15_50;
mixer gate_output_15_50(.a(output_16_50), .b(output_16_3), .y(output_15_50));
wire output_1_51, output_1_4, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_4), .y(output_0_51));
wire output_2_51, output_2_4, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_4), .y(output_1_51));
wire output_3_51, output_3_4, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_4), .y(output_2_51));
wire output_4_51, output_4_4, output_3_51;
mixer gate_output_3_51(.a(output_4_51), .b(output_4_4), .y(output_3_51));
wire output_5_51, output_5_4, output_4_51;
mixer gate_output_4_51(.a(output_5_51), .b(output_5_4), .y(output_4_51));
wire output_6_51, output_6_4, output_5_51;
mixer gate_output_5_51(.a(output_6_51), .b(output_6_4), .y(output_5_51));
wire output_7_51, output_7_4, output_6_51;
mixer gate_output_6_51(.a(output_7_51), .b(output_7_4), .y(output_6_51));
wire output_8_51, output_8_4, output_7_51;
mixer gate_output_7_51(.a(output_8_51), .b(output_8_4), .y(output_7_51));
wire output_9_51, output_9_4, output_8_51;
mixer gate_output_8_51(.a(output_9_51), .b(output_9_4), .y(output_8_51));
wire output_10_51, output_10_4, output_9_51;
mixer gate_output_9_51(.a(output_10_51), .b(output_10_4), .y(output_9_51));
wire output_11_51, output_11_4, output_10_51;
mixer gate_output_10_51(.a(output_11_51), .b(output_11_4), .y(output_10_51));
wire output_12_51, output_12_4, output_11_51;
mixer gate_output_11_51(.a(output_12_51), .b(output_12_4), .y(output_11_51));
wire output_13_51, output_13_4, output_12_51;
mixer gate_output_12_51(.a(output_13_51), .b(output_13_4), .y(output_12_51));
wire output_14_51, output_14_4, output_13_51;
mixer gate_output_13_51(.a(output_14_51), .b(output_14_4), .y(output_13_51));
wire output_15_51, output_15_4, output_14_51;
mixer gate_output_14_51(.a(output_15_51), .b(output_15_4), .y(output_14_51));
wire output_16_51, output_16_4, output_15_51;
mixer gate_output_15_51(.a(output_16_51), .b(output_16_4), .y(output_15_51));
wire output_1_52, output_1_5, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_5), .y(output_0_52));
wire output_2_52, output_2_5, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_5), .y(output_1_52));
wire output_3_52, output_3_5, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_5), .y(output_2_52));
wire output_4_52, output_4_5, output_3_52;
mixer gate_output_3_52(.a(output_4_52), .b(output_4_5), .y(output_3_52));
wire output_5_52, output_5_5, output_4_52;
mixer gate_output_4_52(.a(output_5_52), .b(output_5_5), .y(output_4_52));
wire output_6_52, output_6_5, output_5_52;
mixer gate_output_5_52(.a(output_6_52), .b(output_6_5), .y(output_5_52));
wire output_7_52, output_7_5, output_6_52;
mixer gate_output_6_52(.a(output_7_52), .b(output_7_5), .y(output_6_52));
wire output_8_52, output_8_5, output_7_52;
mixer gate_output_7_52(.a(output_8_52), .b(output_8_5), .y(output_7_52));
wire output_9_52, output_9_5, output_8_52;
mixer gate_output_8_52(.a(output_9_52), .b(output_9_5), .y(output_8_52));
wire output_10_52, output_10_5, output_9_52;
mixer gate_output_9_52(.a(output_10_52), .b(output_10_5), .y(output_9_52));
wire output_11_52, output_11_5, output_10_52;
mixer gate_output_10_52(.a(output_11_52), .b(output_11_5), .y(output_10_52));
wire output_12_52, output_12_5, output_11_52;
mixer gate_output_11_52(.a(output_12_52), .b(output_12_5), .y(output_11_52));
wire output_13_52, output_13_5, output_12_52;
mixer gate_output_12_52(.a(output_13_52), .b(output_13_5), .y(output_12_52));
wire output_14_52, output_14_5, output_13_52;
mixer gate_output_13_52(.a(output_14_52), .b(output_14_5), .y(output_13_52));
wire output_15_52, output_15_5, output_14_52;
mixer gate_output_14_52(.a(output_15_52), .b(output_15_5), .y(output_14_52));
wire output_16_52, output_16_5, output_15_52;
mixer gate_output_15_52(.a(output_16_52), .b(output_16_5), .y(output_15_52));
wire output_1_53, output_1_6, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_6), .y(output_0_53));
wire output_2_53, output_2_6, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_6), .y(output_1_53));
wire output_3_53, output_3_6, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_6), .y(output_2_53));
wire output_4_53, output_4_6, output_3_53;
mixer gate_output_3_53(.a(output_4_53), .b(output_4_6), .y(output_3_53));
wire output_5_53, output_5_6, output_4_53;
mixer gate_output_4_53(.a(output_5_53), .b(output_5_6), .y(output_4_53));
wire output_6_53, output_6_6, output_5_53;
mixer gate_output_5_53(.a(output_6_53), .b(output_6_6), .y(output_5_53));
wire output_7_53, output_7_6, output_6_53;
mixer gate_output_6_53(.a(output_7_53), .b(output_7_6), .y(output_6_53));
wire output_8_53, output_8_6, output_7_53;
mixer gate_output_7_53(.a(output_8_53), .b(output_8_6), .y(output_7_53));
wire output_9_53, output_9_6, output_8_53;
mixer gate_output_8_53(.a(output_9_53), .b(output_9_6), .y(output_8_53));
wire output_10_53, output_10_6, output_9_53;
mixer gate_output_9_53(.a(output_10_53), .b(output_10_6), .y(output_9_53));
wire output_11_53, output_11_6, output_10_53;
mixer gate_output_10_53(.a(output_11_53), .b(output_11_6), .y(output_10_53));
wire output_12_53, output_12_6, output_11_53;
mixer gate_output_11_53(.a(output_12_53), .b(output_12_6), .y(output_11_53));
wire output_13_53, output_13_6, output_12_53;
mixer gate_output_12_53(.a(output_13_53), .b(output_13_6), .y(output_12_53));
wire output_14_53, output_14_6, output_13_53;
mixer gate_output_13_53(.a(output_14_53), .b(output_14_6), .y(output_13_53));
wire output_15_53, output_15_6, output_14_53;
mixer gate_output_14_53(.a(output_15_53), .b(output_15_6), .y(output_14_53));
wire output_16_53, output_16_6, output_15_53;
mixer gate_output_15_53(.a(output_16_53), .b(output_16_6), .y(output_15_53));
wire output_1_54, output_1_7, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_7), .y(output_0_54));
wire output_2_54, output_2_7, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_7), .y(output_1_54));
wire output_3_54, output_3_7, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_7), .y(output_2_54));
wire output_4_54, output_4_7, output_3_54;
mixer gate_output_3_54(.a(output_4_54), .b(output_4_7), .y(output_3_54));
wire output_5_54, output_5_7, output_4_54;
mixer gate_output_4_54(.a(output_5_54), .b(output_5_7), .y(output_4_54));
wire output_6_54, output_6_7, output_5_54;
mixer gate_output_5_54(.a(output_6_54), .b(output_6_7), .y(output_5_54));
wire output_7_54, output_7_7, output_6_54;
mixer gate_output_6_54(.a(output_7_54), .b(output_7_7), .y(output_6_54));
wire output_8_54, output_8_7, output_7_54;
mixer gate_output_7_54(.a(output_8_54), .b(output_8_7), .y(output_7_54));
wire output_9_54, output_9_7, output_8_54;
mixer gate_output_8_54(.a(output_9_54), .b(output_9_7), .y(output_8_54));
wire output_10_54, output_10_7, output_9_54;
mixer gate_output_9_54(.a(output_10_54), .b(output_10_7), .y(output_9_54));
wire output_11_54, output_11_7, output_10_54;
mixer gate_output_10_54(.a(output_11_54), .b(output_11_7), .y(output_10_54));
wire output_12_54, output_12_7, output_11_54;
mixer gate_output_11_54(.a(output_12_54), .b(output_12_7), .y(output_11_54));
wire output_13_54, output_13_7, output_12_54;
mixer gate_output_12_54(.a(output_13_54), .b(output_13_7), .y(output_12_54));
wire output_14_54, output_14_7, output_13_54;
mixer gate_output_13_54(.a(output_14_54), .b(output_14_7), .y(output_13_54));
wire output_15_54, output_15_7, output_14_54;
mixer gate_output_14_54(.a(output_15_54), .b(output_15_7), .y(output_14_54));
wire output_16_54, output_16_7, output_15_54;
mixer gate_output_15_54(.a(output_16_54), .b(output_16_7), .y(output_15_54));
wire output_1_55, output_1_8, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_8), .y(output_0_55));
wire output_2_55, output_2_8, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_8), .y(output_1_55));
wire output_3_55, output_3_8, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_8), .y(output_2_55));
wire output_4_55, output_4_8, output_3_55;
mixer gate_output_3_55(.a(output_4_55), .b(output_4_8), .y(output_3_55));
wire output_5_55, output_5_8, output_4_55;
mixer gate_output_4_55(.a(output_5_55), .b(output_5_8), .y(output_4_55));
wire output_6_55, output_6_8, output_5_55;
mixer gate_output_5_55(.a(output_6_55), .b(output_6_8), .y(output_5_55));
wire output_7_55, output_7_8, output_6_55;
mixer gate_output_6_55(.a(output_7_55), .b(output_7_8), .y(output_6_55));
wire output_8_55, output_8_8, output_7_55;
mixer gate_output_7_55(.a(output_8_55), .b(output_8_8), .y(output_7_55));
wire output_9_55, output_9_8, output_8_55;
mixer gate_output_8_55(.a(output_9_55), .b(output_9_8), .y(output_8_55));
wire output_10_55, output_10_8, output_9_55;
mixer gate_output_9_55(.a(output_10_55), .b(output_10_8), .y(output_9_55));
wire output_11_55, output_11_8, output_10_55;
mixer gate_output_10_55(.a(output_11_55), .b(output_11_8), .y(output_10_55));
wire output_12_55, output_12_8, output_11_55;
mixer gate_output_11_55(.a(output_12_55), .b(output_12_8), .y(output_11_55));
wire output_13_55, output_13_8, output_12_55;
mixer gate_output_12_55(.a(output_13_55), .b(output_13_8), .y(output_12_55));
wire output_14_55, output_14_8, output_13_55;
mixer gate_output_13_55(.a(output_14_55), .b(output_14_8), .y(output_13_55));
wire output_15_55, output_15_8, output_14_55;
mixer gate_output_14_55(.a(output_15_55), .b(output_15_8), .y(output_14_55));
wire output_16_55, output_16_8, output_15_55;
mixer gate_output_15_55(.a(output_16_55), .b(output_16_8), .y(output_15_55));
wire output_1_56, output_1_9, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_9), .y(output_0_56));
wire output_2_56, output_2_9, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_9), .y(output_1_56));
wire output_3_56, output_3_9, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_9), .y(output_2_56));
wire output_4_56, output_4_9, output_3_56;
mixer gate_output_3_56(.a(output_4_56), .b(output_4_9), .y(output_3_56));
wire output_5_56, output_5_9, output_4_56;
mixer gate_output_4_56(.a(output_5_56), .b(output_5_9), .y(output_4_56));
wire output_6_56, output_6_9, output_5_56;
mixer gate_output_5_56(.a(output_6_56), .b(output_6_9), .y(output_5_56));
wire output_7_56, output_7_9, output_6_56;
mixer gate_output_6_56(.a(output_7_56), .b(output_7_9), .y(output_6_56));
wire output_8_56, output_8_9, output_7_56;
mixer gate_output_7_56(.a(output_8_56), .b(output_8_9), .y(output_7_56));
wire output_9_56, output_9_9, output_8_56;
mixer gate_output_8_56(.a(output_9_56), .b(output_9_9), .y(output_8_56));
wire output_10_56, output_10_9, output_9_56;
mixer gate_output_9_56(.a(output_10_56), .b(output_10_9), .y(output_9_56));
wire output_11_56, output_11_9, output_10_56;
mixer gate_output_10_56(.a(output_11_56), .b(output_11_9), .y(output_10_56));
wire output_12_56, output_12_9, output_11_56;
mixer gate_output_11_56(.a(output_12_56), .b(output_12_9), .y(output_11_56));
wire output_13_56, output_13_9, output_12_56;
mixer gate_output_12_56(.a(output_13_56), .b(output_13_9), .y(output_12_56));
wire output_14_56, output_14_9, output_13_56;
mixer gate_output_13_56(.a(output_14_56), .b(output_14_9), .y(output_13_56));
wire output_15_56, output_15_9, output_14_56;
mixer gate_output_14_56(.a(output_15_56), .b(output_15_9), .y(output_14_56));
wire output_16_56, output_16_9, output_15_56;
mixer gate_output_15_56(.a(output_16_56), .b(output_16_9), .y(output_15_56));
wire output_1_57, output_1_10, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_10), .y(output_0_57));
wire output_2_57, output_2_10, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_10), .y(output_1_57));
wire output_3_57, output_3_10, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_10), .y(output_2_57));
wire output_4_57, output_4_10, output_3_57;
mixer gate_output_3_57(.a(output_4_57), .b(output_4_10), .y(output_3_57));
wire output_5_57, output_5_10, output_4_57;
mixer gate_output_4_57(.a(output_5_57), .b(output_5_10), .y(output_4_57));
wire output_6_57, output_6_10, output_5_57;
mixer gate_output_5_57(.a(output_6_57), .b(output_6_10), .y(output_5_57));
wire output_7_57, output_7_10, output_6_57;
mixer gate_output_6_57(.a(output_7_57), .b(output_7_10), .y(output_6_57));
wire output_8_57, output_8_10, output_7_57;
mixer gate_output_7_57(.a(output_8_57), .b(output_8_10), .y(output_7_57));
wire output_9_57, output_9_10, output_8_57;
mixer gate_output_8_57(.a(output_9_57), .b(output_9_10), .y(output_8_57));
wire output_10_57, output_10_10, output_9_57;
mixer gate_output_9_57(.a(output_10_57), .b(output_10_10), .y(output_9_57));
wire output_11_57, output_11_10, output_10_57;
mixer gate_output_10_57(.a(output_11_57), .b(output_11_10), .y(output_10_57));
wire output_12_57, output_12_10, output_11_57;
mixer gate_output_11_57(.a(output_12_57), .b(output_12_10), .y(output_11_57));
wire output_13_57, output_13_10, output_12_57;
mixer gate_output_12_57(.a(output_13_57), .b(output_13_10), .y(output_12_57));
wire output_14_57, output_14_10, output_13_57;
mixer gate_output_13_57(.a(output_14_57), .b(output_14_10), .y(output_13_57));
wire output_15_57, output_15_10, output_14_57;
mixer gate_output_14_57(.a(output_15_57), .b(output_15_10), .y(output_14_57));
wire output_16_57, output_16_10, output_15_57;
mixer gate_output_15_57(.a(output_16_57), .b(output_16_10), .y(output_15_57));
wire output_1_58, output_1_11, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_11), .y(output_0_58));
wire output_2_58, output_2_11, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_11), .y(output_1_58));
wire output_3_58, output_3_11, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_11), .y(output_2_58));
wire output_4_58, output_4_11, output_3_58;
mixer gate_output_3_58(.a(output_4_58), .b(output_4_11), .y(output_3_58));
wire output_5_58, output_5_11, output_4_58;
mixer gate_output_4_58(.a(output_5_58), .b(output_5_11), .y(output_4_58));
wire output_6_58, output_6_11, output_5_58;
mixer gate_output_5_58(.a(output_6_58), .b(output_6_11), .y(output_5_58));
wire output_7_58, output_7_11, output_6_58;
mixer gate_output_6_58(.a(output_7_58), .b(output_7_11), .y(output_6_58));
wire output_8_58, output_8_11, output_7_58;
mixer gate_output_7_58(.a(output_8_58), .b(output_8_11), .y(output_7_58));
wire output_9_58, output_9_11, output_8_58;
mixer gate_output_8_58(.a(output_9_58), .b(output_9_11), .y(output_8_58));
wire output_10_58, output_10_11, output_9_58;
mixer gate_output_9_58(.a(output_10_58), .b(output_10_11), .y(output_9_58));
wire output_11_58, output_11_11, output_10_58;
mixer gate_output_10_58(.a(output_11_58), .b(output_11_11), .y(output_10_58));
wire output_12_58, output_12_11, output_11_58;
mixer gate_output_11_58(.a(output_12_58), .b(output_12_11), .y(output_11_58));
wire output_13_58, output_13_11, output_12_58;
mixer gate_output_12_58(.a(output_13_58), .b(output_13_11), .y(output_12_58));
wire output_14_58, output_14_11, output_13_58;
mixer gate_output_13_58(.a(output_14_58), .b(output_14_11), .y(output_13_58));
wire output_15_58, output_15_11, output_14_58;
mixer gate_output_14_58(.a(output_15_58), .b(output_15_11), .y(output_14_58));
wire output_16_58, output_16_11, output_15_58;
mixer gate_output_15_58(.a(output_16_58), .b(output_16_11), .y(output_15_58));
wire output_1_59, output_1_12, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_12), .y(output_0_59));
wire output_2_59, output_2_12, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_12), .y(output_1_59));
wire output_3_59, output_3_12, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_12), .y(output_2_59));
wire output_4_59, output_4_12, output_3_59;
mixer gate_output_3_59(.a(output_4_59), .b(output_4_12), .y(output_3_59));
wire output_5_59, output_5_12, output_4_59;
mixer gate_output_4_59(.a(output_5_59), .b(output_5_12), .y(output_4_59));
wire output_6_59, output_6_12, output_5_59;
mixer gate_output_5_59(.a(output_6_59), .b(output_6_12), .y(output_5_59));
wire output_7_59, output_7_12, output_6_59;
mixer gate_output_6_59(.a(output_7_59), .b(output_7_12), .y(output_6_59));
wire output_8_59, output_8_12, output_7_59;
mixer gate_output_7_59(.a(output_8_59), .b(output_8_12), .y(output_7_59));
wire output_9_59, output_9_12, output_8_59;
mixer gate_output_8_59(.a(output_9_59), .b(output_9_12), .y(output_8_59));
wire output_10_59, output_10_12, output_9_59;
mixer gate_output_9_59(.a(output_10_59), .b(output_10_12), .y(output_9_59));
wire output_11_59, output_11_12, output_10_59;
mixer gate_output_10_59(.a(output_11_59), .b(output_11_12), .y(output_10_59));
wire output_12_59, output_12_12, output_11_59;
mixer gate_output_11_59(.a(output_12_59), .b(output_12_12), .y(output_11_59));
wire output_13_59, output_13_12, output_12_59;
mixer gate_output_12_59(.a(output_13_59), .b(output_13_12), .y(output_12_59));
wire output_14_59, output_14_12, output_13_59;
mixer gate_output_13_59(.a(output_14_59), .b(output_14_12), .y(output_13_59));
wire output_15_59, output_15_12, output_14_59;
mixer gate_output_14_59(.a(output_15_59), .b(output_15_12), .y(output_14_59));
wire output_16_59, output_16_12, output_15_59;
mixer gate_output_15_59(.a(output_16_59), .b(output_16_12), .y(output_15_59));
wire output_1_60, output_1_13, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_13), .y(output_0_60));
wire output_2_60, output_2_13, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_13), .y(output_1_60));
wire output_3_60, output_3_13, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_13), .y(output_2_60));
wire output_4_60, output_4_13, output_3_60;
mixer gate_output_3_60(.a(output_4_60), .b(output_4_13), .y(output_3_60));
wire output_5_60, output_5_13, output_4_60;
mixer gate_output_4_60(.a(output_5_60), .b(output_5_13), .y(output_4_60));
wire output_6_60, output_6_13, output_5_60;
mixer gate_output_5_60(.a(output_6_60), .b(output_6_13), .y(output_5_60));
wire output_7_60, output_7_13, output_6_60;
mixer gate_output_6_60(.a(output_7_60), .b(output_7_13), .y(output_6_60));
wire output_8_60, output_8_13, output_7_60;
mixer gate_output_7_60(.a(output_8_60), .b(output_8_13), .y(output_7_60));
wire output_9_60, output_9_13, output_8_60;
mixer gate_output_8_60(.a(output_9_60), .b(output_9_13), .y(output_8_60));
wire output_10_60, output_10_13, output_9_60;
mixer gate_output_9_60(.a(output_10_60), .b(output_10_13), .y(output_9_60));
wire output_11_60, output_11_13, output_10_60;
mixer gate_output_10_60(.a(output_11_60), .b(output_11_13), .y(output_10_60));
wire output_12_60, output_12_13, output_11_60;
mixer gate_output_11_60(.a(output_12_60), .b(output_12_13), .y(output_11_60));
wire output_13_60, output_13_13, output_12_60;
mixer gate_output_12_60(.a(output_13_60), .b(output_13_13), .y(output_12_60));
wire output_14_60, output_14_13, output_13_60;
mixer gate_output_13_60(.a(output_14_60), .b(output_14_13), .y(output_13_60));
wire output_15_60, output_15_13, output_14_60;
mixer gate_output_14_60(.a(output_15_60), .b(output_15_13), .y(output_14_60));
wire output_16_60, output_16_13, output_15_60;
mixer gate_output_15_60(.a(output_16_60), .b(output_16_13), .y(output_15_60));
wire output_1_61, output_1_14, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_14), .y(output_0_61));
wire output_2_61, output_2_14, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_14), .y(output_1_61));
wire output_3_61, output_3_14, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_14), .y(output_2_61));
wire output_4_61, output_4_14, output_3_61;
mixer gate_output_3_61(.a(output_4_61), .b(output_4_14), .y(output_3_61));
wire output_5_61, output_5_14, output_4_61;
mixer gate_output_4_61(.a(output_5_61), .b(output_5_14), .y(output_4_61));
wire output_6_61, output_6_14, output_5_61;
mixer gate_output_5_61(.a(output_6_61), .b(output_6_14), .y(output_5_61));
wire output_7_61, output_7_14, output_6_61;
mixer gate_output_6_61(.a(output_7_61), .b(output_7_14), .y(output_6_61));
wire output_8_61, output_8_14, output_7_61;
mixer gate_output_7_61(.a(output_8_61), .b(output_8_14), .y(output_7_61));
wire output_9_61, output_9_14, output_8_61;
mixer gate_output_8_61(.a(output_9_61), .b(output_9_14), .y(output_8_61));
wire output_10_61, output_10_14, output_9_61;
mixer gate_output_9_61(.a(output_10_61), .b(output_10_14), .y(output_9_61));
wire output_11_61, output_11_14, output_10_61;
mixer gate_output_10_61(.a(output_11_61), .b(output_11_14), .y(output_10_61));
wire output_12_61, output_12_14, output_11_61;
mixer gate_output_11_61(.a(output_12_61), .b(output_12_14), .y(output_11_61));
wire output_13_61, output_13_14, output_12_61;
mixer gate_output_12_61(.a(output_13_61), .b(output_13_14), .y(output_12_61));
wire output_14_61, output_14_14, output_13_61;
mixer gate_output_13_61(.a(output_14_61), .b(output_14_14), .y(output_13_61));
wire output_15_61, output_15_14, output_14_61;
mixer gate_output_14_61(.a(output_15_61), .b(output_15_14), .y(output_14_61));
wire output_16_61, output_16_14, output_15_61;
mixer gate_output_15_61(.a(output_16_61), .b(output_16_14), .y(output_15_61));
wire output_1_62, output_1_15, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_15), .y(output_0_62));
wire output_2_62, output_2_15, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_15), .y(output_1_62));
wire output_3_62, output_3_15, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_15), .y(output_2_62));
wire output_4_62, output_4_15, output_3_62;
mixer gate_output_3_62(.a(output_4_62), .b(output_4_15), .y(output_3_62));
wire output_5_62, output_5_15, output_4_62;
mixer gate_output_4_62(.a(output_5_62), .b(output_5_15), .y(output_4_62));
wire output_6_62, output_6_15, output_5_62;
mixer gate_output_5_62(.a(output_6_62), .b(output_6_15), .y(output_5_62));
wire output_7_62, output_7_15, output_6_62;
mixer gate_output_6_62(.a(output_7_62), .b(output_7_15), .y(output_6_62));
wire output_8_62, output_8_15, output_7_62;
mixer gate_output_7_62(.a(output_8_62), .b(output_8_15), .y(output_7_62));
wire output_9_62, output_9_15, output_8_62;
mixer gate_output_8_62(.a(output_9_62), .b(output_9_15), .y(output_8_62));
wire output_10_62, output_10_15, output_9_62;
mixer gate_output_9_62(.a(output_10_62), .b(output_10_15), .y(output_9_62));
wire output_11_62, output_11_15, output_10_62;
mixer gate_output_10_62(.a(output_11_62), .b(output_11_15), .y(output_10_62));
wire output_12_62, output_12_15, output_11_62;
mixer gate_output_11_62(.a(output_12_62), .b(output_12_15), .y(output_11_62));
wire output_13_62, output_13_15, output_12_62;
mixer gate_output_12_62(.a(output_13_62), .b(output_13_15), .y(output_12_62));
wire output_14_62, output_14_15, output_13_62;
mixer gate_output_13_62(.a(output_14_62), .b(output_14_15), .y(output_13_62));
wire output_15_62, output_15_15, output_14_62;
mixer gate_output_14_62(.a(output_15_62), .b(output_15_15), .y(output_14_62));
wire output_16_62, output_16_15, output_15_62;
mixer gate_output_15_62(.a(output_16_62), .b(output_16_15), .y(output_15_62));
wire output_1_63, output_1_0, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_0), .y(output_0_63));
wire output_2_63, output_2_0, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_0), .y(output_1_63));
wire output_3_63, output_3_0, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_0), .y(output_2_63));
wire output_4_63, output_4_0, output_3_63;
mixer gate_output_3_63(.a(output_4_63), .b(output_4_0), .y(output_3_63));
wire output_5_63, output_5_0, output_4_63;
mixer gate_output_4_63(.a(output_5_63), .b(output_5_0), .y(output_4_63));
wire output_6_63, output_6_0, output_5_63;
mixer gate_output_5_63(.a(output_6_63), .b(output_6_0), .y(output_5_63));
wire output_7_63, output_7_0, output_6_63;
mixer gate_output_6_63(.a(output_7_63), .b(output_7_0), .y(output_6_63));
wire output_8_63, output_8_0, output_7_63;
mixer gate_output_7_63(.a(output_8_63), .b(output_8_0), .y(output_7_63));
wire output_9_63, output_9_0, output_8_63;
mixer gate_output_8_63(.a(output_9_63), .b(output_9_0), .y(output_8_63));
wire output_10_63, output_10_0, output_9_63;
mixer gate_output_9_63(.a(output_10_63), .b(output_10_0), .y(output_9_63));
wire output_11_63, output_11_0, output_10_63;
mixer gate_output_10_63(.a(output_11_63), .b(output_11_0), .y(output_10_63));
wire output_12_63, output_12_0, output_11_63;
mixer gate_output_11_63(.a(output_12_63), .b(output_12_0), .y(output_11_63));
wire output_13_63, output_13_0, output_12_63;
mixer gate_output_12_63(.a(output_13_63), .b(output_13_0), .y(output_12_63));
wire output_14_63, output_14_0, output_13_63;
mixer gate_output_13_63(.a(output_14_63), .b(output_14_0), .y(output_13_63));
wire output_15_63, output_15_0, output_14_63;
mixer gate_output_14_63(.a(output_15_63), .b(output_15_0), .y(output_14_63));
wire output_16_63, output_16_0, output_15_63;
mixer gate_output_15_63(.a(output_16_63), .b(output_16_0), .y(output_15_63));
wire output_1_64, output_1_1, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_1), .y(output_0_64));
wire output_2_64, output_2_1, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_1), .y(output_1_64));
wire output_3_64, output_3_1, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_1), .y(output_2_64));
wire output_4_64, output_4_1, output_3_64;
mixer gate_output_3_64(.a(output_4_64), .b(output_4_1), .y(output_3_64));
wire output_5_64, output_5_1, output_4_64;
mixer gate_output_4_64(.a(output_5_64), .b(output_5_1), .y(output_4_64));
wire output_6_64, output_6_1, output_5_64;
mixer gate_output_5_64(.a(output_6_64), .b(output_6_1), .y(output_5_64));
wire output_7_64, output_7_1, output_6_64;
mixer gate_output_6_64(.a(output_7_64), .b(output_7_1), .y(output_6_64));
wire output_8_64, output_8_1, output_7_64;
mixer gate_output_7_64(.a(output_8_64), .b(output_8_1), .y(output_7_64));
wire output_9_64, output_9_1, output_8_64;
mixer gate_output_8_64(.a(output_9_64), .b(output_9_1), .y(output_8_64));
wire output_10_64, output_10_1, output_9_64;
mixer gate_output_9_64(.a(output_10_64), .b(output_10_1), .y(output_9_64));
wire output_11_64, output_11_1, output_10_64;
mixer gate_output_10_64(.a(output_11_64), .b(output_11_1), .y(output_10_64));
wire output_12_64, output_12_1, output_11_64;
mixer gate_output_11_64(.a(output_12_64), .b(output_12_1), .y(output_11_64));
wire output_13_64, output_13_1, output_12_64;
mixer gate_output_12_64(.a(output_13_64), .b(output_13_1), .y(output_12_64));
wire output_14_64, output_14_1, output_13_64;
mixer gate_output_13_64(.a(output_14_64), .b(output_14_1), .y(output_13_64));
wire output_15_64, output_15_1, output_14_64;
mixer gate_output_14_64(.a(output_15_64), .b(output_15_1), .y(output_14_64));
wire output_16_64, output_16_1, output_15_64;
mixer gate_output_15_64(.a(output_16_64), .b(output_16_1), .y(output_15_64));
wire output_1_65, output_1_2, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_2), .y(output_0_65));
wire output_2_65, output_2_2, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_2), .y(output_1_65));
wire output_3_65, output_3_2, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_2), .y(output_2_65));
wire output_4_65, output_4_2, output_3_65;
mixer gate_output_3_65(.a(output_4_65), .b(output_4_2), .y(output_3_65));
wire output_5_65, output_5_2, output_4_65;
mixer gate_output_4_65(.a(output_5_65), .b(output_5_2), .y(output_4_65));
wire output_6_65, output_6_2, output_5_65;
mixer gate_output_5_65(.a(output_6_65), .b(output_6_2), .y(output_5_65));
wire output_7_65, output_7_2, output_6_65;
mixer gate_output_6_65(.a(output_7_65), .b(output_7_2), .y(output_6_65));
wire output_8_65, output_8_2, output_7_65;
mixer gate_output_7_65(.a(output_8_65), .b(output_8_2), .y(output_7_65));
wire output_9_65, output_9_2, output_8_65;
mixer gate_output_8_65(.a(output_9_65), .b(output_9_2), .y(output_8_65));
wire output_10_65, output_10_2, output_9_65;
mixer gate_output_9_65(.a(output_10_65), .b(output_10_2), .y(output_9_65));
wire output_11_65, output_11_2, output_10_65;
mixer gate_output_10_65(.a(output_11_65), .b(output_11_2), .y(output_10_65));
wire output_12_65, output_12_2, output_11_65;
mixer gate_output_11_65(.a(output_12_65), .b(output_12_2), .y(output_11_65));
wire output_13_65, output_13_2, output_12_65;
mixer gate_output_12_65(.a(output_13_65), .b(output_13_2), .y(output_12_65));
wire output_14_65, output_14_2, output_13_65;
mixer gate_output_13_65(.a(output_14_65), .b(output_14_2), .y(output_13_65));
wire output_15_65, output_15_2, output_14_65;
mixer gate_output_14_65(.a(output_15_65), .b(output_15_2), .y(output_14_65));
wire output_16_65, output_16_2, output_15_65;
mixer gate_output_15_65(.a(output_16_65), .b(output_16_2), .y(output_15_65));
wire output_1_66, output_1_3, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_3), .y(output_0_66));
wire output_2_66, output_2_3, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_3), .y(output_1_66));
wire output_3_66, output_3_3, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_3), .y(output_2_66));
wire output_4_66, output_4_3, output_3_66;
mixer gate_output_3_66(.a(output_4_66), .b(output_4_3), .y(output_3_66));
wire output_5_66, output_5_3, output_4_66;
mixer gate_output_4_66(.a(output_5_66), .b(output_5_3), .y(output_4_66));
wire output_6_66, output_6_3, output_5_66;
mixer gate_output_5_66(.a(output_6_66), .b(output_6_3), .y(output_5_66));
wire output_7_66, output_7_3, output_6_66;
mixer gate_output_6_66(.a(output_7_66), .b(output_7_3), .y(output_6_66));
wire output_8_66, output_8_3, output_7_66;
mixer gate_output_7_66(.a(output_8_66), .b(output_8_3), .y(output_7_66));
wire output_9_66, output_9_3, output_8_66;
mixer gate_output_8_66(.a(output_9_66), .b(output_9_3), .y(output_8_66));
wire output_10_66, output_10_3, output_9_66;
mixer gate_output_9_66(.a(output_10_66), .b(output_10_3), .y(output_9_66));
wire output_11_66, output_11_3, output_10_66;
mixer gate_output_10_66(.a(output_11_66), .b(output_11_3), .y(output_10_66));
wire output_12_66, output_12_3, output_11_66;
mixer gate_output_11_66(.a(output_12_66), .b(output_12_3), .y(output_11_66));
wire output_13_66, output_13_3, output_12_66;
mixer gate_output_12_66(.a(output_13_66), .b(output_13_3), .y(output_12_66));
wire output_14_66, output_14_3, output_13_66;
mixer gate_output_13_66(.a(output_14_66), .b(output_14_3), .y(output_13_66));
wire output_15_66, output_15_3, output_14_66;
mixer gate_output_14_66(.a(output_15_66), .b(output_15_3), .y(output_14_66));
wire output_16_66, output_16_3, output_15_66;
mixer gate_output_15_66(.a(output_16_66), .b(output_16_3), .y(output_15_66));
wire output_1_67, output_1_4, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_4), .y(output_0_67));
wire output_2_67, output_2_4, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_4), .y(output_1_67));
wire output_3_67, output_3_4, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_4), .y(output_2_67));
wire output_4_67, output_4_4, output_3_67;
mixer gate_output_3_67(.a(output_4_67), .b(output_4_4), .y(output_3_67));
wire output_5_67, output_5_4, output_4_67;
mixer gate_output_4_67(.a(output_5_67), .b(output_5_4), .y(output_4_67));
wire output_6_67, output_6_4, output_5_67;
mixer gate_output_5_67(.a(output_6_67), .b(output_6_4), .y(output_5_67));
wire output_7_67, output_7_4, output_6_67;
mixer gate_output_6_67(.a(output_7_67), .b(output_7_4), .y(output_6_67));
wire output_8_67, output_8_4, output_7_67;
mixer gate_output_7_67(.a(output_8_67), .b(output_8_4), .y(output_7_67));
wire output_9_67, output_9_4, output_8_67;
mixer gate_output_8_67(.a(output_9_67), .b(output_9_4), .y(output_8_67));
wire output_10_67, output_10_4, output_9_67;
mixer gate_output_9_67(.a(output_10_67), .b(output_10_4), .y(output_9_67));
wire output_11_67, output_11_4, output_10_67;
mixer gate_output_10_67(.a(output_11_67), .b(output_11_4), .y(output_10_67));
wire output_12_67, output_12_4, output_11_67;
mixer gate_output_11_67(.a(output_12_67), .b(output_12_4), .y(output_11_67));
wire output_13_67, output_13_4, output_12_67;
mixer gate_output_12_67(.a(output_13_67), .b(output_13_4), .y(output_12_67));
wire output_14_67, output_14_4, output_13_67;
mixer gate_output_13_67(.a(output_14_67), .b(output_14_4), .y(output_13_67));
wire output_15_67, output_15_4, output_14_67;
mixer gate_output_14_67(.a(output_15_67), .b(output_15_4), .y(output_14_67));
wire output_16_67, output_16_4, output_15_67;
mixer gate_output_15_67(.a(output_16_67), .b(output_16_4), .y(output_15_67));
wire output_1_68, output_1_5, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_5), .y(output_0_68));
wire output_2_68, output_2_5, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_5), .y(output_1_68));
wire output_3_68, output_3_5, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_5), .y(output_2_68));
wire output_4_68, output_4_5, output_3_68;
mixer gate_output_3_68(.a(output_4_68), .b(output_4_5), .y(output_3_68));
wire output_5_68, output_5_5, output_4_68;
mixer gate_output_4_68(.a(output_5_68), .b(output_5_5), .y(output_4_68));
wire output_6_68, output_6_5, output_5_68;
mixer gate_output_5_68(.a(output_6_68), .b(output_6_5), .y(output_5_68));
wire output_7_68, output_7_5, output_6_68;
mixer gate_output_6_68(.a(output_7_68), .b(output_7_5), .y(output_6_68));
wire output_8_68, output_8_5, output_7_68;
mixer gate_output_7_68(.a(output_8_68), .b(output_8_5), .y(output_7_68));
wire output_9_68, output_9_5, output_8_68;
mixer gate_output_8_68(.a(output_9_68), .b(output_9_5), .y(output_8_68));
wire output_10_68, output_10_5, output_9_68;
mixer gate_output_9_68(.a(output_10_68), .b(output_10_5), .y(output_9_68));
wire output_11_68, output_11_5, output_10_68;
mixer gate_output_10_68(.a(output_11_68), .b(output_11_5), .y(output_10_68));
wire output_12_68, output_12_5, output_11_68;
mixer gate_output_11_68(.a(output_12_68), .b(output_12_5), .y(output_11_68));
wire output_13_68, output_13_5, output_12_68;
mixer gate_output_12_68(.a(output_13_68), .b(output_13_5), .y(output_12_68));
wire output_14_68, output_14_5, output_13_68;
mixer gate_output_13_68(.a(output_14_68), .b(output_14_5), .y(output_13_68));
wire output_15_68, output_15_5, output_14_68;
mixer gate_output_14_68(.a(output_15_68), .b(output_15_5), .y(output_14_68));
wire output_16_68, output_16_5, output_15_68;
mixer gate_output_15_68(.a(output_16_68), .b(output_16_5), .y(output_15_68));
wire output_1_69, output_1_6, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_6), .y(output_0_69));
wire output_2_69, output_2_6, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_6), .y(output_1_69));
wire output_3_69, output_3_6, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_6), .y(output_2_69));
wire output_4_69, output_4_6, output_3_69;
mixer gate_output_3_69(.a(output_4_69), .b(output_4_6), .y(output_3_69));
wire output_5_69, output_5_6, output_4_69;
mixer gate_output_4_69(.a(output_5_69), .b(output_5_6), .y(output_4_69));
wire output_6_69, output_6_6, output_5_69;
mixer gate_output_5_69(.a(output_6_69), .b(output_6_6), .y(output_5_69));
wire output_7_69, output_7_6, output_6_69;
mixer gate_output_6_69(.a(output_7_69), .b(output_7_6), .y(output_6_69));
wire output_8_69, output_8_6, output_7_69;
mixer gate_output_7_69(.a(output_8_69), .b(output_8_6), .y(output_7_69));
wire output_9_69, output_9_6, output_8_69;
mixer gate_output_8_69(.a(output_9_69), .b(output_9_6), .y(output_8_69));
wire output_10_69, output_10_6, output_9_69;
mixer gate_output_9_69(.a(output_10_69), .b(output_10_6), .y(output_9_69));
wire output_11_69, output_11_6, output_10_69;
mixer gate_output_10_69(.a(output_11_69), .b(output_11_6), .y(output_10_69));
wire output_12_69, output_12_6, output_11_69;
mixer gate_output_11_69(.a(output_12_69), .b(output_12_6), .y(output_11_69));
wire output_13_69, output_13_6, output_12_69;
mixer gate_output_12_69(.a(output_13_69), .b(output_13_6), .y(output_12_69));
wire output_14_69, output_14_6, output_13_69;
mixer gate_output_13_69(.a(output_14_69), .b(output_14_6), .y(output_13_69));
wire output_15_69, output_15_6, output_14_69;
mixer gate_output_14_69(.a(output_15_69), .b(output_15_6), .y(output_14_69));
wire output_16_69, output_16_6, output_15_69;
mixer gate_output_15_69(.a(output_16_69), .b(output_16_6), .y(output_15_69));
wire output_1_70, output_1_7, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_7), .y(output_0_70));
wire output_2_70, output_2_7, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_7), .y(output_1_70));
wire output_3_70, output_3_7, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_7), .y(output_2_70));
wire output_4_70, output_4_7, output_3_70;
mixer gate_output_3_70(.a(output_4_70), .b(output_4_7), .y(output_3_70));
wire output_5_70, output_5_7, output_4_70;
mixer gate_output_4_70(.a(output_5_70), .b(output_5_7), .y(output_4_70));
wire output_6_70, output_6_7, output_5_70;
mixer gate_output_5_70(.a(output_6_70), .b(output_6_7), .y(output_5_70));
wire output_7_70, output_7_7, output_6_70;
mixer gate_output_6_70(.a(output_7_70), .b(output_7_7), .y(output_6_70));
wire output_8_70, output_8_7, output_7_70;
mixer gate_output_7_70(.a(output_8_70), .b(output_8_7), .y(output_7_70));
wire output_9_70, output_9_7, output_8_70;
mixer gate_output_8_70(.a(output_9_70), .b(output_9_7), .y(output_8_70));
wire output_10_70, output_10_7, output_9_70;
mixer gate_output_9_70(.a(output_10_70), .b(output_10_7), .y(output_9_70));
wire output_11_70, output_11_7, output_10_70;
mixer gate_output_10_70(.a(output_11_70), .b(output_11_7), .y(output_10_70));
wire output_12_70, output_12_7, output_11_70;
mixer gate_output_11_70(.a(output_12_70), .b(output_12_7), .y(output_11_70));
wire output_13_70, output_13_7, output_12_70;
mixer gate_output_12_70(.a(output_13_70), .b(output_13_7), .y(output_12_70));
wire output_14_70, output_14_7, output_13_70;
mixer gate_output_13_70(.a(output_14_70), .b(output_14_7), .y(output_13_70));
wire output_15_70, output_15_7, output_14_70;
mixer gate_output_14_70(.a(output_15_70), .b(output_15_7), .y(output_14_70));
wire output_16_70, output_16_7, output_15_70;
mixer gate_output_15_70(.a(output_16_70), .b(output_16_7), .y(output_15_70));
wire output_1_71, output_1_8, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_8), .y(output_0_71));
wire output_2_71, output_2_8, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_8), .y(output_1_71));
wire output_3_71, output_3_8, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_8), .y(output_2_71));
wire output_4_71, output_4_8, output_3_71;
mixer gate_output_3_71(.a(output_4_71), .b(output_4_8), .y(output_3_71));
wire output_5_71, output_5_8, output_4_71;
mixer gate_output_4_71(.a(output_5_71), .b(output_5_8), .y(output_4_71));
wire output_6_71, output_6_8, output_5_71;
mixer gate_output_5_71(.a(output_6_71), .b(output_6_8), .y(output_5_71));
wire output_7_71, output_7_8, output_6_71;
mixer gate_output_6_71(.a(output_7_71), .b(output_7_8), .y(output_6_71));
wire output_8_71, output_8_8, output_7_71;
mixer gate_output_7_71(.a(output_8_71), .b(output_8_8), .y(output_7_71));
wire output_9_71, output_9_8, output_8_71;
mixer gate_output_8_71(.a(output_9_71), .b(output_9_8), .y(output_8_71));
wire output_10_71, output_10_8, output_9_71;
mixer gate_output_9_71(.a(output_10_71), .b(output_10_8), .y(output_9_71));
wire output_11_71, output_11_8, output_10_71;
mixer gate_output_10_71(.a(output_11_71), .b(output_11_8), .y(output_10_71));
wire output_12_71, output_12_8, output_11_71;
mixer gate_output_11_71(.a(output_12_71), .b(output_12_8), .y(output_11_71));
wire output_13_71, output_13_8, output_12_71;
mixer gate_output_12_71(.a(output_13_71), .b(output_13_8), .y(output_12_71));
wire output_14_71, output_14_8, output_13_71;
mixer gate_output_13_71(.a(output_14_71), .b(output_14_8), .y(output_13_71));
wire output_15_71, output_15_8, output_14_71;
mixer gate_output_14_71(.a(output_15_71), .b(output_15_8), .y(output_14_71));
wire output_16_71, output_16_8, output_15_71;
mixer gate_output_15_71(.a(output_16_71), .b(output_16_8), .y(output_15_71));
wire output_1_72, output_1_9, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_9), .y(output_0_72));
wire output_2_72, output_2_9, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_9), .y(output_1_72));
wire output_3_72, output_3_9, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_9), .y(output_2_72));
wire output_4_72, output_4_9, output_3_72;
mixer gate_output_3_72(.a(output_4_72), .b(output_4_9), .y(output_3_72));
wire output_5_72, output_5_9, output_4_72;
mixer gate_output_4_72(.a(output_5_72), .b(output_5_9), .y(output_4_72));
wire output_6_72, output_6_9, output_5_72;
mixer gate_output_5_72(.a(output_6_72), .b(output_6_9), .y(output_5_72));
wire output_7_72, output_7_9, output_6_72;
mixer gate_output_6_72(.a(output_7_72), .b(output_7_9), .y(output_6_72));
wire output_8_72, output_8_9, output_7_72;
mixer gate_output_7_72(.a(output_8_72), .b(output_8_9), .y(output_7_72));
wire output_9_72, output_9_9, output_8_72;
mixer gate_output_8_72(.a(output_9_72), .b(output_9_9), .y(output_8_72));
wire output_10_72, output_10_9, output_9_72;
mixer gate_output_9_72(.a(output_10_72), .b(output_10_9), .y(output_9_72));
wire output_11_72, output_11_9, output_10_72;
mixer gate_output_10_72(.a(output_11_72), .b(output_11_9), .y(output_10_72));
wire output_12_72, output_12_9, output_11_72;
mixer gate_output_11_72(.a(output_12_72), .b(output_12_9), .y(output_11_72));
wire output_13_72, output_13_9, output_12_72;
mixer gate_output_12_72(.a(output_13_72), .b(output_13_9), .y(output_12_72));
wire output_14_72, output_14_9, output_13_72;
mixer gate_output_13_72(.a(output_14_72), .b(output_14_9), .y(output_13_72));
wire output_15_72, output_15_9, output_14_72;
mixer gate_output_14_72(.a(output_15_72), .b(output_15_9), .y(output_14_72));
wire output_16_72, output_16_9, output_15_72;
mixer gate_output_15_72(.a(output_16_72), .b(output_16_9), .y(output_15_72));
wire output_1_73, output_1_10, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_10), .y(output_0_73));
wire output_2_73, output_2_10, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_10), .y(output_1_73));
wire output_3_73, output_3_10, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_10), .y(output_2_73));
wire output_4_73, output_4_10, output_3_73;
mixer gate_output_3_73(.a(output_4_73), .b(output_4_10), .y(output_3_73));
wire output_5_73, output_5_10, output_4_73;
mixer gate_output_4_73(.a(output_5_73), .b(output_5_10), .y(output_4_73));
wire output_6_73, output_6_10, output_5_73;
mixer gate_output_5_73(.a(output_6_73), .b(output_6_10), .y(output_5_73));
wire output_7_73, output_7_10, output_6_73;
mixer gate_output_6_73(.a(output_7_73), .b(output_7_10), .y(output_6_73));
wire output_8_73, output_8_10, output_7_73;
mixer gate_output_7_73(.a(output_8_73), .b(output_8_10), .y(output_7_73));
wire output_9_73, output_9_10, output_8_73;
mixer gate_output_8_73(.a(output_9_73), .b(output_9_10), .y(output_8_73));
wire output_10_73, output_10_10, output_9_73;
mixer gate_output_9_73(.a(output_10_73), .b(output_10_10), .y(output_9_73));
wire output_11_73, output_11_10, output_10_73;
mixer gate_output_10_73(.a(output_11_73), .b(output_11_10), .y(output_10_73));
wire output_12_73, output_12_10, output_11_73;
mixer gate_output_11_73(.a(output_12_73), .b(output_12_10), .y(output_11_73));
wire output_13_73, output_13_10, output_12_73;
mixer gate_output_12_73(.a(output_13_73), .b(output_13_10), .y(output_12_73));
wire output_14_73, output_14_10, output_13_73;
mixer gate_output_13_73(.a(output_14_73), .b(output_14_10), .y(output_13_73));
wire output_15_73, output_15_10, output_14_73;
mixer gate_output_14_73(.a(output_15_73), .b(output_15_10), .y(output_14_73));
wire output_16_73, output_16_10, output_15_73;
mixer gate_output_15_73(.a(output_16_73), .b(output_16_10), .y(output_15_73));
wire output_1_74, output_1_11, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_11), .y(output_0_74));
wire output_2_74, output_2_11, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_11), .y(output_1_74));
wire output_3_74, output_3_11, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_11), .y(output_2_74));
wire output_4_74, output_4_11, output_3_74;
mixer gate_output_3_74(.a(output_4_74), .b(output_4_11), .y(output_3_74));
wire output_5_74, output_5_11, output_4_74;
mixer gate_output_4_74(.a(output_5_74), .b(output_5_11), .y(output_4_74));
wire output_6_74, output_6_11, output_5_74;
mixer gate_output_5_74(.a(output_6_74), .b(output_6_11), .y(output_5_74));
wire output_7_74, output_7_11, output_6_74;
mixer gate_output_6_74(.a(output_7_74), .b(output_7_11), .y(output_6_74));
wire output_8_74, output_8_11, output_7_74;
mixer gate_output_7_74(.a(output_8_74), .b(output_8_11), .y(output_7_74));
wire output_9_74, output_9_11, output_8_74;
mixer gate_output_8_74(.a(output_9_74), .b(output_9_11), .y(output_8_74));
wire output_10_74, output_10_11, output_9_74;
mixer gate_output_9_74(.a(output_10_74), .b(output_10_11), .y(output_9_74));
wire output_11_74, output_11_11, output_10_74;
mixer gate_output_10_74(.a(output_11_74), .b(output_11_11), .y(output_10_74));
wire output_12_74, output_12_11, output_11_74;
mixer gate_output_11_74(.a(output_12_74), .b(output_12_11), .y(output_11_74));
wire output_13_74, output_13_11, output_12_74;
mixer gate_output_12_74(.a(output_13_74), .b(output_13_11), .y(output_12_74));
wire output_14_74, output_14_11, output_13_74;
mixer gate_output_13_74(.a(output_14_74), .b(output_14_11), .y(output_13_74));
wire output_15_74, output_15_11, output_14_74;
mixer gate_output_14_74(.a(output_15_74), .b(output_15_11), .y(output_14_74));
wire output_16_74, output_16_11, output_15_74;
mixer gate_output_15_74(.a(output_16_74), .b(output_16_11), .y(output_15_74));
wire output_1_75, output_1_12, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_12), .y(output_0_75));
wire output_2_75, output_2_12, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_12), .y(output_1_75));
wire output_3_75, output_3_12, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_12), .y(output_2_75));
wire output_4_75, output_4_12, output_3_75;
mixer gate_output_3_75(.a(output_4_75), .b(output_4_12), .y(output_3_75));
wire output_5_75, output_5_12, output_4_75;
mixer gate_output_4_75(.a(output_5_75), .b(output_5_12), .y(output_4_75));
wire output_6_75, output_6_12, output_5_75;
mixer gate_output_5_75(.a(output_6_75), .b(output_6_12), .y(output_5_75));
wire output_7_75, output_7_12, output_6_75;
mixer gate_output_6_75(.a(output_7_75), .b(output_7_12), .y(output_6_75));
wire output_8_75, output_8_12, output_7_75;
mixer gate_output_7_75(.a(output_8_75), .b(output_8_12), .y(output_7_75));
wire output_9_75, output_9_12, output_8_75;
mixer gate_output_8_75(.a(output_9_75), .b(output_9_12), .y(output_8_75));
wire output_10_75, output_10_12, output_9_75;
mixer gate_output_9_75(.a(output_10_75), .b(output_10_12), .y(output_9_75));
wire output_11_75, output_11_12, output_10_75;
mixer gate_output_10_75(.a(output_11_75), .b(output_11_12), .y(output_10_75));
wire output_12_75, output_12_12, output_11_75;
mixer gate_output_11_75(.a(output_12_75), .b(output_12_12), .y(output_11_75));
wire output_13_75, output_13_12, output_12_75;
mixer gate_output_12_75(.a(output_13_75), .b(output_13_12), .y(output_12_75));
wire output_14_75, output_14_12, output_13_75;
mixer gate_output_13_75(.a(output_14_75), .b(output_14_12), .y(output_13_75));
wire output_15_75, output_15_12, output_14_75;
mixer gate_output_14_75(.a(output_15_75), .b(output_15_12), .y(output_14_75));
wire output_16_75, output_16_12, output_15_75;
mixer gate_output_15_75(.a(output_16_75), .b(output_16_12), .y(output_15_75));
wire output_1_76, output_1_13, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_13), .y(output_0_76));
wire output_2_76, output_2_13, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_13), .y(output_1_76));
wire output_3_76, output_3_13, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_13), .y(output_2_76));
wire output_4_76, output_4_13, output_3_76;
mixer gate_output_3_76(.a(output_4_76), .b(output_4_13), .y(output_3_76));
wire output_5_76, output_5_13, output_4_76;
mixer gate_output_4_76(.a(output_5_76), .b(output_5_13), .y(output_4_76));
wire output_6_76, output_6_13, output_5_76;
mixer gate_output_5_76(.a(output_6_76), .b(output_6_13), .y(output_5_76));
wire output_7_76, output_7_13, output_6_76;
mixer gate_output_6_76(.a(output_7_76), .b(output_7_13), .y(output_6_76));
wire output_8_76, output_8_13, output_7_76;
mixer gate_output_7_76(.a(output_8_76), .b(output_8_13), .y(output_7_76));
wire output_9_76, output_9_13, output_8_76;
mixer gate_output_8_76(.a(output_9_76), .b(output_9_13), .y(output_8_76));
wire output_10_76, output_10_13, output_9_76;
mixer gate_output_9_76(.a(output_10_76), .b(output_10_13), .y(output_9_76));
wire output_11_76, output_11_13, output_10_76;
mixer gate_output_10_76(.a(output_11_76), .b(output_11_13), .y(output_10_76));
wire output_12_76, output_12_13, output_11_76;
mixer gate_output_11_76(.a(output_12_76), .b(output_12_13), .y(output_11_76));
wire output_13_76, output_13_13, output_12_76;
mixer gate_output_12_76(.a(output_13_76), .b(output_13_13), .y(output_12_76));
wire output_14_76, output_14_13, output_13_76;
mixer gate_output_13_76(.a(output_14_76), .b(output_14_13), .y(output_13_76));
wire output_15_76, output_15_13, output_14_76;
mixer gate_output_14_76(.a(output_15_76), .b(output_15_13), .y(output_14_76));
wire output_16_76, output_16_13, output_15_76;
mixer gate_output_15_76(.a(output_16_76), .b(output_16_13), .y(output_15_76));
wire output_1_77, output_1_14, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_14), .y(output_0_77));
wire output_2_77, output_2_14, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_14), .y(output_1_77));
wire output_3_77, output_3_14, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_14), .y(output_2_77));
wire output_4_77, output_4_14, output_3_77;
mixer gate_output_3_77(.a(output_4_77), .b(output_4_14), .y(output_3_77));
wire output_5_77, output_5_14, output_4_77;
mixer gate_output_4_77(.a(output_5_77), .b(output_5_14), .y(output_4_77));
wire output_6_77, output_6_14, output_5_77;
mixer gate_output_5_77(.a(output_6_77), .b(output_6_14), .y(output_5_77));
wire output_7_77, output_7_14, output_6_77;
mixer gate_output_6_77(.a(output_7_77), .b(output_7_14), .y(output_6_77));
wire output_8_77, output_8_14, output_7_77;
mixer gate_output_7_77(.a(output_8_77), .b(output_8_14), .y(output_7_77));
wire output_9_77, output_9_14, output_8_77;
mixer gate_output_8_77(.a(output_9_77), .b(output_9_14), .y(output_8_77));
wire output_10_77, output_10_14, output_9_77;
mixer gate_output_9_77(.a(output_10_77), .b(output_10_14), .y(output_9_77));
wire output_11_77, output_11_14, output_10_77;
mixer gate_output_10_77(.a(output_11_77), .b(output_11_14), .y(output_10_77));
wire output_12_77, output_12_14, output_11_77;
mixer gate_output_11_77(.a(output_12_77), .b(output_12_14), .y(output_11_77));
wire output_13_77, output_13_14, output_12_77;
mixer gate_output_12_77(.a(output_13_77), .b(output_13_14), .y(output_12_77));
wire output_14_77, output_14_14, output_13_77;
mixer gate_output_13_77(.a(output_14_77), .b(output_14_14), .y(output_13_77));
wire output_15_77, output_15_14, output_14_77;
mixer gate_output_14_77(.a(output_15_77), .b(output_15_14), .y(output_14_77));
wire output_16_77, output_16_14, output_15_77;
mixer gate_output_15_77(.a(output_16_77), .b(output_16_14), .y(output_15_77));
wire output_1_78, output_1_15, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_15), .y(output_0_78));
wire output_2_78, output_2_15, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_15), .y(output_1_78));
wire output_3_78, output_3_15, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_15), .y(output_2_78));
wire output_4_78, output_4_15, output_3_78;
mixer gate_output_3_78(.a(output_4_78), .b(output_4_15), .y(output_3_78));
wire output_5_78, output_5_15, output_4_78;
mixer gate_output_4_78(.a(output_5_78), .b(output_5_15), .y(output_4_78));
wire output_6_78, output_6_15, output_5_78;
mixer gate_output_5_78(.a(output_6_78), .b(output_6_15), .y(output_5_78));
wire output_7_78, output_7_15, output_6_78;
mixer gate_output_6_78(.a(output_7_78), .b(output_7_15), .y(output_6_78));
wire output_8_78, output_8_15, output_7_78;
mixer gate_output_7_78(.a(output_8_78), .b(output_8_15), .y(output_7_78));
wire output_9_78, output_9_15, output_8_78;
mixer gate_output_8_78(.a(output_9_78), .b(output_9_15), .y(output_8_78));
wire output_10_78, output_10_15, output_9_78;
mixer gate_output_9_78(.a(output_10_78), .b(output_10_15), .y(output_9_78));
wire output_11_78, output_11_15, output_10_78;
mixer gate_output_10_78(.a(output_11_78), .b(output_11_15), .y(output_10_78));
wire output_12_78, output_12_15, output_11_78;
mixer gate_output_11_78(.a(output_12_78), .b(output_12_15), .y(output_11_78));
wire output_13_78, output_13_15, output_12_78;
mixer gate_output_12_78(.a(output_13_78), .b(output_13_15), .y(output_12_78));
wire output_14_78, output_14_15, output_13_78;
mixer gate_output_13_78(.a(output_14_78), .b(output_14_15), .y(output_13_78));
wire output_15_78, output_15_15, output_14_78;
mixer gate_output_14_78(.a(output_15_78), .b(output_15_15), .y(output_14_78));
wire output_16_78, output_16_15, output_15_78;
mixer gate_output_15_78(.a(output_16_78), .b(output_16_15), .y(output_15_78));
wire output_1_79, output_1_0, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_0), .y(output_0_79));
wire output_2_79, output_2_0, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_0), .y(output_1_79));
wire output_3_79, output_3_0, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_0), .y(output_2_79));
wire output_4_79, output_4_0, output_3_79;
mixer gate_output_3_79(.a(output_4_79), .b(output_4_0), .y(output_3_79));
wire output_5_79, output_5_0, output_4_79;
mixer gate_output_4_79(.a(output_5_79), .b(output_5_0), .y(output_4_79));
wire output_6_79, output_6_0, output_5_79;
mixer gate_output_5_79(.a(output_6_79), .b(output_6_0), .y(output_5_79));
wire output_7_79, output_7_0, output_6_79;
mixer gate_output_6_79(.a(output_7_79), .b(output_7_0), .y(output_6_79));
wire output_8_79, output_8_0, output_7_79;
mixer gate_output_7_79(.a(output_8_79), .b(output_8_0), .y(output_7_79));
wire output_9_79, output_9_0, output_8_79;
mixer gate_output_8_79(.a(output_9_79), .b(output_9_0), .y(output_8_79));
wire output_10_79, output_10_0, output_9_79;
mixer gate_output_9_79(.a(output_10_79), .b(output_10_0), .y(output_9_79));
wire output_11_79, output_11_0, output_10_79;
mixer gate_output_10_79(.a(output_11_79), .b(output_11_0), .y(output_10_79));
wire output_12_79, output_12_0, output_11_79;
mixer gate_output_11_79(.a(output_12_79), .b(output_12_0), .y(output_11_79));
wire output_13_79, output_13_0, output_12_79;
mixer gate_output_12_79(.a(output_13_79), .b(output_13_0), .y(output_12_79));
wire output_14_79, output_14_0, output_13_79;
mixer gate_output_13_79(.a(output_14_79), .b(output_14_0), .y(output_13_79));
wire output_15_79, output_15_0, output_14_79;
mixer gate_output_14_79(.a(output_15_79), .b(output_15_0), .y(output_14_79));
wire output_16_79, output_16_0, output_15_79;
mixer gate_output_15_79(.a(output_16_79), .b(output_16_0), .y(output_15_79));
wire output_1_80, output_1_1, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_1), .y(output_0_80));
wire output_2_80, output_2_1, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_1), .y(output_1_80));
wire output_3_80, output_3_1, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_1), .y(output_2_80));
wire output_4_80, output_4_1, output_3_80;
mixer gate_output_3_80(.a(output_4_80), .b(output_4_1), .y(output_3_80));
wire output_5_80, output_5_1, output_4_80;
mixer gate_output_4_80(.a(output_5_80), .b(output_5_1), .y(output_4_80));
wire output_6_80, output_6_1, output_5_80;
mixer gate_output_5_80(.a(output_6_80), .b(output_6_1), .y(output_5_80));
wire output_7_80, output_7_1, output_6_80;
mixer gate_output_6_80(.a(output_7_80), .b(output_7_1), .y(output_6_80));
wire output_8_80, output_8_1, output_7_80;
mixer gate_output_7_80(.a(output_8_80), .b(output_8_1), .y(output_7_80));
wire output_9_80, output_9_1, output_8_80;
mixer gate_output_8_80(.a(output_9_80), .b(output_9_1), .y(output_8_80));
wire output_10_80, output_10_1, output_9_80;
mixer gate_output_9_80(.a(output_10_80), .b(output_10_1), .y(output_9_80));
wire output_11_80, output_11_1, output_10_80;
mixer gate_output_10_80(.a(output_11_80), .b(output_11_1), .y(output_10_80));
wire output_12_80, output_12_1, output_11_80;
mixer gate_output_11_80(.a(output_12_80), .b(output_12_1), .y(output_11_80));
wire output_13_80, output_13_1, output_12_80;
mixer gate_output_12_80(.a(output_13_80), .b(output_13_1), .y(output_12_80));
wire output_14_80, output_14_1, output_13_80;
mixer gate_output_13_80(.a(output_14_80), .b(output_14_1), .y(output_13_80));
wire output_15_80, output_15_1, output_14_80;
mixer gate_output_14_80(.a(output_15_80), .b(output_15_1), .y(output_14_80));
wire output_16_80, output_16_1, output_15_80;
mixer gate_output_15_80(.a(output_16_80), .b(output_16_1), .y(output_15_80));
wire output_1_81, output_1_2, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_2), .y(output_0_81));
wire output_2_81, output_2_2, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_2), .y(output_1_81));
wire output_3_81, output_3_2, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_2), .y(output_2_81));
wire output_4_81, output_4_2, output_3_81;
mixer gate_output_3_81(.a(output_4_81), .b(output_4_2), .y(output_3_81));
wire output_5_81, output_5_2, output_4_81;
mixer gate_output_4_81(.a(output_5_81), .b(output_5_2), .y(output_4_81));
wire output_6_81, output_6_2, output_5_81;
mixer gate_output_5_81(.a(output_6_81), .b(output_6_2), .y(output_5_81));
wire output_7_81, output_7_2, output_6_81;
mixer gate_output_6_81(.a(output_7_81), .b(output_7_2), .y(output_6_81));
wire output_8_81, output_8_2, output_7_81;
mixer gate_output_7_81(.a(output_8_81), .b(output_8_2), .y(output_7_81));
wire output_9_81, output_9_2, output_8_81;
mixer gate_output_8_81(.a(output_9_81), .b(output_9_2), .y(output_8_81));
wire output_10_81, output_10_2, output_9_81;
mixer gate_output_9_81(.a(output_10_81), .b(output_10_2), .y(output_9_81));
wire output_11_81, output_11_2, output_10_81;
mixer gate_output_10_81(.a(output_11_81), .b(output_11_2), .y(output_10_81));
wire output_12_81, output_12_2, output_11_81;
mixer gate_output_11_81(.a(output_12_81), .b(output_12_2), .y(output_11_81));
wire output_13_81, output_13_2, output_12_81;
mixer gate_output_12_81(.a(output_13_81), .b(output_13_2), .y(output_12_81));
wire output_14_81, output_14_2, output_13_81;
mixer gate_output_13_81(.a(output_14_81), .b(output_14_2), .y(output_13_81));
wire output_15_81, output_15_2, output_14_81;
mixer gate_output_14_81(.a(output_15_81), .b(output_15_2), .y(output_14_81));
wire output_16_81, output_16_2, output_15_81;
mixer gate_output_15_81(.a(output_16_81), .b(output_16_2), .y(output_15_81));
wire output_1_82, output_1_3, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_3), .y(output_0_82));
wire output_2_82, output_2_3, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_3), .y(output_1_82));
wire output_3_82, output_3_3, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_3), .y(output_2_82));
wire output_4_82, output_4_3, output_3_82;
mixer gate_output_3_82(.a(output_4_82), .b(output_4_3), .y(output_3_82));
wire output_5_82, output_5_3, output_4_82;
mixer gate_output_4_82(.a(output_5_82), .b(output_5_3), .y(output_4_82));
wire output_6_82, output_6_3, output_5_82;
mixer gate_output_5_82(.a(output_6_82), .b(output_6_3), .y(output_5_82));
wire output_7_82, output_7_3, output_6_82;
mixer gate_output_6_82(.a(output_7_82), .b(output_7_3), .y(output_6_82));
wire output_8_82, output_8_3, output_7_82;
mixer gate_output_7_82(.a(output_8_82), .b(output_8_3), .y(output_7_82));
wire output_9_82, output_9_3, output_8_82;
mixer gate_output_8_82(.a(output_9_82), .b(output_9_3), .y(output_8_82));
wire output_10_82, output_10_3, output_9_82;
mixer gate_output_9_82(.a(output_10_82), .b(output_10_3), .y(output_9_82));
wire output_11_82, output_11_3, output_10_82;
mixer gate_output_10_82(.a(output_11_82), .b(output_11_3), .y(output_10_82));
wire output_12_82, output_12_3, output_11_82;
mixer gate_output_11_82(.a(output_12_82), .b(output_12_3), .y(output_11_82));
wire output_13_82, output_13_3, output_12_82;
mixer gate_output_12_82(.a(output_13_82), .b(output_13_3), .y(output_12_82));
wire output_14_82, output_14_3, output_13_82;
mixer gate_output_13_82(.a(output_14_82), .b(output_14_3), .y(output_13_82));
wire output_15_82, output_15_3, output_14_82;
mixer gate_output_14_82(.a(output_15_82), .b(output_15_3), .y(output_14_82));
wire output_16_82, output_16_3, output_15_82;
mixer gate_output_15_82(.a(output_16_82), .b(output_16_3), .y(output_15_82));
wire output_1_83, output_1_4, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_4), .y(output_0_83));
wire output_2_83, output_2_4, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_4), .y(output_1_83));
wire output_3_83, output_3_4, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_4), .y(output_2_83));
wire output_4_83, output_4_4, output_3_83;
mixer gate_output_3_83(.a(output_4_83), .b(output_4_4), .y(output_3_83));
wire output_5_83, output_5_4, output_4_83;
mixer gate_output_4_83(.a(output_5_83), .b(output_5_4), .y(output_4_83));
wire output_6_83, output_6_4, output_5_83;
mixer gate_output_5_83(.a(output_6_83), .b(output_6_4), .y(output_5_83));
wire output_7_83, output_7_4, output_6_83;
mixer gate_output_6_83(.a(output_7_83), .b(output_7_4), .y(output_6_83));
wire output_8_83, output_8_4, output_7_83;
mixer gate_output_7_83(.a(output_8_83), .b(output_8_4), .y(output_7_83));
wire output_9_83, output_9_4, output_8_83;
mixer gate_output_8_83(.a(output_9_83), .b(output_9_4), .y(output_8_83));
wire output_10_83, output_10_4, output_9_83;
mixer gate_output_9_83(.a(output_10_83), .b(output_10_4), .y(output_9_83));
wire output_11_83, output_11_4, output_10_83;
mixer gate_output_10_83(.a(output_11_83), .b(output_11_4), .y(output_10_83));
wire output_12_83, output_12_4, output_11_83;
mixer gate_output_11_83(.a(output_12_83), .b(output_12_4), .y(output_11_83));
wire output_13_83, output_13_4, output_12_83;
mixer gate_output_12_83(.a(output_13_83), .b(output_13_4), .y(output_12_83));
wire output_14_83, output_14_4, output_13_83;
mixer gate_output_13_83(.a(output_14_83), .b(output_14_4), .y(output_13_83));
wire output_15_83, output_15_4, output_14_83;
mixer gate_output_14_83(.a(output_15_83), .b(output_15_4), .y(output_14_83));
wire output_16_83, output_16_4, output_15_83;
mixer gate_output_15_83(.a(output_16_83), .b(output_16_4), .y(output_15_83));
wire output_1_84, output_1_5, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_5), .y(output_0_84));
wire output_2_84, output_2_5, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_5), .y(output_1_84));
wire output_3_84, output_3_5, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_5), .y(output_2_84));
wire output_4_84, output_4_5, output_3_84;
mixer gate_output_3_84(.a(output_4_84), .b(output_4_5), .y(output_3_84));
wire output_5_84, output_5_5, output_4_84;
mixer gate_output_4_84(.a(output_5_84), .b(output_5_5), .y(output_4_84));
wire output_6_84, output_6_5, output_5_84;
mixer gate_output_5_84(.a(output_6_84), .b(output_6_5), .y(output_5_84));
wire output_7_84, output_7_5, output_6_84;
mixer gate_output_6_84(.a(output_7_84), .b(output_7_5), .y(output_6_84));
wire output_8_84, output_8_5, output_7_84;
mixer gate_output_7_84(.a(output_8_84), .b(output_8_5), .y(output_7_84));
wire output_9_84, output_9_5, output_8_84;
mixer gate_output_8_84(.a(output_9_84), .b(output_9_5), .y(output_8_84));
wire output_10_84, output_10_5, output_9_84;
mixer gate_output_9_84(.a(output_10_84), .b(output_10_5), .y(output_9_84));
wire output_11_84, output_11_5, output_10_84;
mixer gate_output_10_84(.a(output_11_84), .b(output_11_5), .y(output_10_84));
wire output_12_84, output_12_5, output_11_84;
mixer gate_output_11_84(.a(output_12_84), .b(output_12_5), .y(output_11_84));
wire output_13_84, output_13_5, output_12_84;
mixer gate_output_12_84(.a(output_13_84), .b(output_13_5), .y(output_12_84));
wire output_14_84, output_14_5, output_13_84;
mixer gate_output_13_84(.a(output_14_84), .b(output_14_5), .y(output_13_84));
wire output_15_84, output_15_5, output_14_84;
mixer gate_output_14_84(.a(output_15_84), .b(output_15_5), .y(output_14_84));
wire output_16_84, output_16_5, output_15_84;
mixer gate_output_15_84(.a(output_16_84), .b(output_16_5), .y(output_15_84));
wire output_1_85, output_1_6, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_6), .y(output_0_85));
wire output_2_85, output_2_6, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_6), .y(output_1_85));
wire output_3_85, output_3_6, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_6), .y(output_2_85));
wire output_4_85, output_4_6, output_3_85;
mixer gate_output_3_85(.a(output_4_85), .b(output_4_6), .y(output_3_85));
wire output_5_85, output_5_6, output_4_85;
mixer gate_output_4_85(.a(output_5_85), .b(output_5_6), .y(output_4_85));
wire output_6_85, output_6_6, output_5_85;
mixer gate_output_5_85(.a(output_6_85), .b(output_6_6), .y(output_5_85));
wire output_7_85, output_7_6, output_6_85;
mixer gate_output_6_85(.a(output_7_85), .b(output_7_6), .y(output_6_85));
wire output_8_85, output_8_6, output_7_85;
mixer gate_output_7_85(.a(output_8_85), .b(output_8_6), .y(output_7_85));
wire output_9_85, output_9_6, output_8_85;
mixer gate_output_8_85(.a(output_9_85), .b(output_9_6), .y(output_8_85));
wire output_10_85, output_10_6, output_9_85;
mixer gate_output_9_85(.a(output_10_85), .b(output_10_6), .y(output_9_85));
wire output_11_85, output_11_6, output_10_85;
mixer gate_output_10_85(.a(output_11_85), .b(output_11_6), .y(output_10_85));
wire output_12_85, output_12_6, output_11_85;
mixer gate_output_11_85(.a(output_12_85), .b(output_12_6), .y(output_11_85));
wire output_13_85, output_13_6, output_12_85;
mixer gate_output_12_85(.a(output_13_85), .b(output_13_6), .y(output_12_85));
wire output_14_85, output_14_6, output_13_85;
mixer gate_output_13_85(.a(output_14_85), .b(output_14_6), .y(output_13_85));
wire output_15_85, output_15_6, output_14_85;
mixer gate_output_14_85(.a(output_15_85), .b(output_15_6), .y(output_14_85));
wire output_16_85, output_16_6, output_15_85;
mixer gate_output_15_85(.a(output_16_85), .b(output_16_6), .y(output_15_85));
wire output_1_86, output_1_7, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_7), .y(output_0_86));
wire output_2_86, output_2_7, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_7), .y(output_1_86));
wire output_3_86, output_3_7, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_7), .y(output_2_86));
wire output_4_86, output_4_7, output_3_86;
mixer gate_output_3_86(.a(output_4_86), .b(output_4_7), .y(output_3_86));
wire output_5_86, output_5_7, output_4_86;
mixer gate_output_4_86(.a(output_5_86), .b(output_5_7), .y(output_4_86));
wire output_6_86, output_6_7, output_5_86;
mixer gate_output_5_86(.a(output_6_86), .b(output_6_7), .y(output_5_86));
wire output_7_86, output_7_7, output_6_86;
mixer gate_output_6_86(.a(output_7_86), .b(output_7_7), .y(output_6_86));
wire output_8_86, output_8_7, output_7_86;
mixer gate_output_7_86(.a(output_8_86), .b(output_8_7), .y(output_7_86));
wire output_9_86, output_9_7, output_8_86;
mixer gate_output_8_86(.a(output_9_86), .b(output_9_7), .y(output_8_86));
wire output_10_86, output_10_7, output_9_86;
mixer gate_output_9_86(.a(output_10_86), .b(output_10_7), .y(output_9_86));
wire output_11_86, output_11_7, output_10_86;
mixer gate_output_10_86(.a(output_11_86), .b(output_11_7), .y(output_10_86));
wire output_12_86, output_12_7, output_11_86;
mixer gate_output_11_86(.a(output_12_86), .b(output_12_7), .y(output_11_86));
wire output_13_86, output_13_7, output_12_86;
mixer gate_output_12_86(.a(output_13_86), .b(output_13_7), .y(output_12_86));
wire output_14_86, output_14_7, output_13_86;
mixer gate_output_13_86(.a(output_14_86), .b(output_14_7), .y(output_13_86));
wire output_15_86, output_15_7, output_14_86;
mixer gate_output_14_86(.a(output_15_86), .b(output_15_7), .y(output_14_86));
wire output_16_86, output_16_7, output_15_86;
mixer gate_output_15_86(.a(output_16_86), .b(output_16_7), .y(output_15_86));
wire output_1_87, output_1_8, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_8), .y(output_0_87));
wire output_2_87, output_2_8, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_8), .y(output_1_87));
wire output_3_87, output_3_8, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_8), .y(output_2_87));
wire output_4_87, output_4_8, output_3_87;
mixer gate_output_3_87(.a(output_4_87), .b(output_4_8), .y(output_3_87));
wire output_5_87, output_5_8, output_4_87;
mixer gate_output_4_87(.a(output_5_87), .b(output_5_8), .y(output_4_87));
wire output_6_87, output_6_8, output_5_87;
mixer gate_output_5_87(.a(output_6_87), .b(output_6_8), .y(output_5_87));
wire output_7_87, output_7_8, output_6_87;
mixer gate_output_6_87(.a(output_7_87), .b(output_7_8), .y(output_6_87));
wire output_8_87, output_8_8, output_7_87;
mixer gate_output_7_87(.a(output_8_87), .b(output_8_8), .y(output_7_87));
wire output_9_87, output_9_8, output_8_87;
mixer gate_output_8_87(.a(output_9_87), .b(output_9_8), .y(output_8_87));
wire output_10_87, output_10_8, output_9_87;
mixer gate_output_9_87(.a(output_10_87), .b(output_10_8), .y(output_9_87));
wire output_11_87, output_11_8, output_10_87;
mixer gate_output_10_87(.a(output_11_87), .b(output_11_8), .y(output_10_87));
wire output_12_87, output_12_8, output_11_87;
mixer gate_output_11_87(.a(output_12_87), .b(output_12_8), .y(output_11_87));
wire output_13_87, output_13_8, output_12_87;
mixer gate_output_12_87(.a(output_13_87), .b(output_13_8), .y(output_12_87));
wire output_14_87, output_14_8, output_13_87;
mixer gate_output_13_87(.a(output_14_87), .b(output_14_8), .y(output_13_87));
wire output_15_87, output_15_8, output_14_87;
mixer gate_output_14_87(.a(output_15_87), .b(output_15_8), .y(output_14_87));
wire output_16_87, output_16_8, output_15_87;
mixer gate_output_15_87(.a(output_16_87), .b(output_16_8), .y(output_15_87));
wire output_1_88, output_1_9, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_9), .y(output_0_88));
wire output_2_88, output_2_9, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_9), .y(output_1_88));
wire output_3_88, output_3_9, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_9), .y(output_2_88));
wire output_4_88, output_4_9, output_3_88;
mixer gate_output_3_88(.a(output_4_88), .b(output_4_9), .y(output_3_88));
wire output_5_88, output_5_9, output_4_88;
mixer gate_output_4_88(.a(output_5_88), .b(output_5_9), .y(output_4_88));
wire output_6_88, output_6_9, output_5_88;
mixer gate_output_5_88(.a(output_6_88), .b(output_6_9), .y(output_5_88));
wire output_7_88, output_7_9, output_6_88;
mixer gate_output_6_88(.a(output_7_88), .b(output_7_9), .y(output_6_88));
wire output_8_88, output_8_9, output_7_88;
mixer gate_output_7_88(.a(output_8_88), .b(output_8_9), .y(output_7_88));
wire output_9_88, output_9_9, output_8_88;
mixer gate_output_8_88(.a(output_9_88), .b(output_9_9), .y(output_8_88));
wire output_10_88, output_10_9, output_9_88;
mixer gate_output_9_88(.a(output_10_88), .b(output_10_9), .y(output_9_88));
wire output_11_88, output_11_9, output_10_88;
mixer gate_output_10_88(.a(output_11_88), .b(output_11_9), .y(output_10_88));
wire output_12_88, output_12_9, output_11_88;
mixer gate_output_11_88(.a(output_12_88), .b(output_12_9), .y(output_11_88));
wire output_13_88, output_13_9, output_12_88;
mixer gate_output_12_88(.a(output_13_88), .b(output_13_9), .y(output_12_88));
wire output_14_88, output_14_9, output_13_88;
mixer gate_output_13_88(.a(output_14_88), .b(output_14_9), .y(output_13_88));
wire output_15_88, output_15_9, output_14_88;
mixer gate_output_14_88(.a(output_15_88), .b(output_15_9), .y(output_14_88));
wire output_16_88, output_16_9, output_15_88;
mixer gate_output_15_88(.a(output_16_88), .b(output_16_9), .y(output_15_88));
wire output_1_89, output_1_10, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_10), .y(output_0_89));
wire output_2_89, output_2_10, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_10), .y(output_1_89));
wire output_3_89, output_3_10, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_10), .y(output_2_89));
wire output_4_89, output_4_10, output_3_89;
mixer gate_output_3_89(.a(output_4_89), .b(output_4_10), .y(output_3_89));
wire output_5_89, output_5_10, output_4_89;
mixer gate_output_4_89(.a(output_5_89), .b(output_5_10), .y(output_4_89));
wire output_6_89, output_6_10, output_5_89;
mixer gate_output_5_89(.a(output_6_89), .b(output_6_10), .y(output_5_89));
wire output_7_89, output_7_10, output_6_89;
mixer gate_output_6_89(.a(output_7_89), .b(output_7_10), .y(output_6_89));
wire output_8_89, output_8_10, output_7_89;
mixer gate_output_7_89(.a(output_8_89), .b(output_8_10), .y(output_7_89));
wire output_9_89, output_9_10, output_8_89;
mixer gate_output_8_89(.a(output_9_89), .b(output_9_10), .y(output_8_89));
wire output_10_89, output_10_10, output_9_89;
mixer gate_output_9_89(.a(output_10_89), .b(output_10_10), .y(output_9_89));
wire output_11_89, output_11_10, output_10_89;
mixer gate_output_10_89(.a(output_11_89), .b(output_11_10), .y(output_10_89));
wire output_12_89, output_12_10, output_11_89;
mixer gate_output_11_89(.a(output_12_89), .b(output_12_10), .y(output_11_89));
wire output_13_89, output_13_10, output_12_89;
mixer gate_output_12_89(.a(output_13_89), .b(output_13_10), .y(output_12_89));
wire output_14_89, output_14_10, output_13_89;
mixer gate_output_13_89(.a(output_14_89), .b(output_14_10), .y(output_13_89));
wire output_15_89, output_15_10, output_14_89;
mixer gate_output_14_89(.a(output_15_89), .b(output_15_10), .y(output_14_89));
wire output_16_89, output_16_10, output_15_89;
mixer gate_output_15_89(.a(output_16_89), .b(output_16_10), .y(output_15_89));
wire output_1_90, output_1_11, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_11), .y(output_0_90));
wire output_2_90, output_2_11, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_11), .y(output_1_90));
wire output_3_90, output_3_11, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_11), .y(output_2_90));
wire output_4_90, output_4_11, output_3_90;
mixer gate_output_3_90(.a(output_4_90), .b(output_4_11), .y(output_3_90));
wire output_5_90, output_5_11, output_4_90;
mixer gate_output_4_90(.a(output_5_90), .b(output_5_11), .y(output_4_90));
wire output_6_90, output_6_11, output_5_90;
mixer gate_output_5_90(.a(output_6_90), .b(output_6_11), .y(output_5_90));
wire output_7_90, output_7_11, output_6_90;
mixer gate_output_6_90(.a(output_7_90), .b(output_7_11), .y(output_6_90));
wire output_8_90, output_8_11, output_7_90;
mixer gate_output_7_90(.a(output_8_90), .b(output_8_11), .y(output_7_90));
wire output_9_90, output_9_11, output_8_90;
mixer gate_output_8_90(.a(output_9_90), .b(output_9_11), .y(output_8_90));
wire output_10_90, output_10_11, output_9_90;
mixer gate_output_9_90(.a(output_10_90), .b(output_10_11), .y(output_9_90));
wire output_11_90, output_11_11, output_10_90;
mixer gate_output_10_90(.a(output_11_90), .b(output_11_11), .y(output_10_90));
wire output_12_90, output_12_11, output_11_90;
mixer gate_output_11_90(.a(output_12_90), .b(output_12_11), .y(output_11_90));
wire output_13_90, output_13_11, output_12_90;
mixer gate_output_12_90(.a(output_13_90), .b(output_13_11), .y(output_12_90));
wire output_14_90, output_14_11, output_13_90;
mixer gate_output_13_90(.a(output_14_90), .b(output_14_11), .y(output_13_90));
wire output_15_90, output_15_11, output_14_90;
mixer gate_output_14_90(.a(output_15_90), .b(output_15_11), .y(output_14_90));
wire output_16_90, output_16_11, output_15_90;
mixer gate_output_15_90(.a(output_16_90), .b(output_16_11), .y(output_15_90));
wire output_1_91, output_1_12, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_12), .y(output_0_91));
wire output_2_91, output_2_12, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_12), .y(output_1_91));
wire output_3_91, output_3_12, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_12), .y(output_2_91));
wire output_4_91, output_4_12, output_3_91;
mixer gate_output_3_91(.a(output_4_91), .b(output_4_12), .y(output_3_91));
wire output_5_91, output_5_12, output_4_91;
mixer gate_output_4_91(.a(output_5_91), .b(output_5_12), .y(output_4_91));
wire output_6_91, output_6_12, output_5_91;
mixer gate_output_5_91(.a(output_6_91), .b(output_6_12), .y(output_5_91));
wire output_7_91, output_7_12, output_6_91;
mixer gate_output_6_91(.a(output_7_91), .b(output_7_12), .y(output_6_91));
wire output_8_91, output_8_12, output_7_91;
mixer gate_output_7_91(.a(output_8_91), .b(output_8_12), .y(output_7_91));
wire output_9_91, output_9_12, output_8_91;
mixer gate_output_8_91(.a(output_9_91), .b(output_9_12), .y(output_8_91));
wire output_10_91, output_10_12, output_9_91;
mixer gate_output_9_91(.a(output_10_91), .b(output_10_12), .y(output_9_91));
wire output_11_91, output_11_12, output_10_91;
mixer gate_output_10_91(.a(output_11_91), .b(output_11_12), .y(output_10_91));
wire output_12_91, output_12_12, output_11_91;
mixer gate_output_11_91(.a(output_12_91), .b(output_12_12), .y(output_11_91));
wire output_13_91, output_13_12, output_12_91;
mixer gate_output_12_91(.a(output_13_91), .b(output_13_12), .y(output_12_91));
wire output_14_91, output_14_12, output_13_91;
mixer gate_output_13_91(.a(output_14_91), .b(output_14_12), .y(output_13_91));
wire output_15_91, output_15_12, output_14_91;
mixer gate_output_14_91(.a(output_15_91), .b(output_15_12), .y(output_14_91));
wire output_16_91, output_16_12, output_15_91;
mixer gate_output_15_91(.a(output_16_91), .b(output_16_12), .y(output_15_91));
wire output_1_92, output_1_13, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_13), .y(output_0_92));
wire output_2_92, output_2_13, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_13), .y(output_1_92));
wire output_3_92, output_3_13, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_13), .y(output_2_92));
wire output_4_92, output_4_13, output_3_92;
mixer gate_output_3_92(.a(output_4_92), .b(output_4_13), .y(output_3_92));
wire output_5_92, output_5_13, output_4_92;
mixer gate_output_4_92(.a(output_5_92), .b(output_5_13), .y(output_4_92));
wire output_6_92, output_6_13, output_5_92;
mixer gate_output_5_92(.a(output_6_92), .b(output_6_13), .y(output_5_92));
wire output_7_92, output_7_13, output_6_92;
mixer gate_output_6_92(.a(output_7_92), .b(output_7_13), .y(output_6_92));
wire output_8_92, output_8_13, output_7_92;
mixer gate_output_7_92(.a(output_8_92), .b(output_8_13), .y(output_7_92));
wire output_9_92, output_9_13, output_8_92;
mixer gate_output_8_92(.a(output_9_92), .b(output_9_13), .y(output_8_92));
wire output_10_92, output_10_13, output_9_92;
mixer gate_output_9_92(.a(output_10_92), .b(output_10_13), .y(output_9_92));
wire output_11_92, output_11_13, output_10_92;
mixer gate_output_10_92(.a(output_11_92), .b(output_11_13), .y(output_10_92));
wire output_12_92, output_12_13, output_11_92;
mixer gate_output_11_92(.a(output_12_92), .b(output_12_13), .y(output_11_92));
wire output_13_92, output_13_13, output_12_92;
mixer gate_output_12_92(.a(output_13_92), .b(output_13_13), .y(output_12_92));
wire output_14_92, output_14_13, output_13_92;
mixer gate_output_13_92(.a(output_14_92), .b(output_14_13), .y(output_13_92));
wire output_15_92, output_15_13, output_14_92;
mixer gate_output_14_92(.a(output_15_92), .b(output_15_13), .y(output_14_92));
wire output_16_92, output_16_13, output_15_92;
mixer gate_output_15_92(.a(output_16_92), .b(output_16_13), .y(output_15_92));
wire output_1_93, output_1_14, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_14), .y(output_0_93));
wire output_2_93, output_2_14, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_14), .y(output_1_93));
wire output_3_93, output_3_14, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_14), .y(output_2_93));
wire output_4_93, output_4_14, output_3_93;
mixer gate_output_3_93(.a(output_4_93), .b(output_4_14), .y(output_3_93));
wire output_5_93, output_5_14, output_4_93;
mixer gate_output_4_93(.a(output_5_93), .b(output_5_14), .y(output_4_93));
wire output_6_93, output_6_14, output_5_93;
mixer gate_output_5_93(.a(output_6_93), .b(output_6_14), .y(output_5_93));
wire output_7_93, output_7_14, output_6_93;
mixer gate_output_6_93(.a(output_7_93), .b(output_7_14), .y(output_6_93));
wire output_8_93, output_8_14, output_7_93;
mixer gate_output_7_93(.a(output_8_93), .b(output_8_14), .y(output_7_93));
wire output_9_93, output_9_14, output_8_93;
mixer gate_output_8_93(.a(output_9_93), .b(output_9_14), .y(output_8_93));
wire output_10_93, output_10_14, output_9_93;
mixer gate_output_9_93(.a(output_10_93), .b(output_10_14), .y(output_9_93));
wire output_11_93, output_11_14, output_10_93;
mixer gate_output_10_93(.a(output_11_93), .b(output_11_14), .y(output_10_93));
wire output_12_93, output_12_14, output_11_93;
mixer gate_output_11_93(.a(output_12_93), .b(output_12_14), .y(output_11_93));
wire output_13_93, output_13_14, output_12_93;
mixer gate_output_12_93(.a(output_13_93), .b(output_13_14), .y(output_12_93));
wire output_14_93, output_14_14, output_13_93;
mixer gate_output_13_93(.a(output_14_93), .b(output_14_14), .y(output_13_93));
wire output_15_93, output_15_14, output_14_93;
mixer gate_output_14_93(.a(output_15_93), .b(output_15_14), .y(output_14_93));
wire output_16_93, output_16_14, output_15_93;
mixer gate_output_15_93(.a(output_16_93), .b(output_16_14), .y(output_15_93));
wire output_1_94, output_1_15, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_15), .y(output_0_94));
wire output_2_94, output_2_15, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_15), .y(output_1_94));
wire output_3_94, output_3_15, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_15), .y(output_2_94));
wire output_4_94, output_4_15, output_3_94;
mixer gate_output_3_94(.a(output_4_94), .b(output_4_15), .y(output_3_94));
wire output_5_94, output_5_15, output_4_94;
mixer gate_output_4_94(.a(output_5_94), .b(output_5_15), .y(output_4_94));
wire output_6_94, output_6_15, output_5_94;
mixer gate_output_5_94(.a(output_6_94), .b(output_6_15), .y(output_5_94));
wire output_7_94, output_7_15, output_6_94;
mixer gate_output_6_94(.a(output_7_94), .b(output_7_15), .y(output_6_94));
wire output_8_94, output_8_15, output_7_94;
mixer gate_output_7_94(.a(output_8_94), .b(output_8_15), .y(output_7_94));
wire output_9_94, output_9_15, output_8_94;
mixer gate_output_8_94(.a(output_9_94), .b(output_9_15), .y(output_8_94));
wire output_10_94, output_10_15, output_9_94;
mixer gate_output_9_94(.a(output_10_94), .b(output_10_15), .y(output_9_94));
wire output_11_94, output_11_15, output_10_94;
mixer gate_output_10_94(.a(output_11_94), .b(output_11_15), .y(output_10_94));
wire output_12_94, output_12_15, output_11_94;
mixer gate_output_11_94(.a(output_12_94), .b(output_12_15), .y(output_11_94));
wire output_13_94, output_13_15, output_12_94;
mixer gate_output_12_94(.a(output_13_94), .b(output_13_15), .y(output_12_94));
wire output_14_94, output_14_15, output_13_94;
mixer gate_output_13_94(.a(output_14_94), .b(output_14_15), .y(output_13_94));
wire output_15_94, output_15_15, output_14_94;
mixer gate_output_14_94(.a(output_15_94), .b(output_15_15), .y(output_14_94));
wire output_16_94, output_16_15, output_15_94;
mixer gate_output_15_94(.a(output_16_94), .b(output_16_15), .y(output_15_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_4_95, output_4_0, output_3_95;
mixer gate_output_3_95(.a(output_4_95), .b(output_4_0), .y(output_3_95));
wire output_5_95, output_5_0, output_4_95;
mixer gate_output_4_95(.a(output_5_95), .b(output_5_0), .y(output_4_95));
wire output_6_95, output_6_0, output_5_95;
mixer gate_output_5_95(.a(output_6_95), .b(output_6_0), .y(output_5_95));
wire output_7_95, output_7_0, output_6_95;
mixer gate_output_6_95(.a(output_7_95), .b(output_7_0), .y(output_6_95));
wire output_8_95, output_8_0, output_7_95;
mixer gate_output_7_95(.a(output_8_95), .b(output_8_0), .y(output_7_95));
wire output_9_95, output_9_0, output_8_95;
mixer gate_output_8_95(.a(output_9_95), .b(output_9_0), .y(output_8_95));
wire output_10_95, output_10_0, output_9_95;
mixer gate_output_9_95(.a(output_10_95), .b(output_10_0), .y(output_9_95));
wire output_11_95, output_11_0, output_10_95;
mixer gate_output_10_95(.a(output_11_95), .b(output_11_0), .y(output_10_95));
wire output_12_95, output_12_0, output_11_95;
mixer gate_output_11_95(.a(output_12_95), .b(output_12_0), .y(output_11_95));
wire output_13_95, output_13_0, output_12_95;
mixer gate_output_12_95(.a(output_13_95), .b(output_13_0), .y(output_12_95));
wire output_14_95, output_14_0, output_13_95;
mixer gate_output_13_95(.a(output_14_95), .b(output_14_0), .y(output_13_95));
wire output_15_95, output_15_0, output_14_95;
mixer gate_output_14_95(.a(output_15_95), .b(output_15_0), .y(output_14_95));
wire output_16_95, output_16_0, output_15_95;
mixer gate_output_15_95(.a(output_16_95), .b(output_16_0), .y(output_15_95));
wire output_1_96, output_1_1, output_0_96;
mixer gate_output_0_96(.a(output_1_96), .b(output_1_1), .y(output_0_96));
wire output_2_96, output_2_1, output_1_96;
mixer gate_output_1_96(.a(output_2_96), .b(output_2_1), .y(output_1_96));
wire output_3_96, output_3_1, output_2_96;
mixer gate_output_2_96(.a(output_3_96), .b(output_3_1), .y(output_2_96));
wire output_4_96, output_4_1, output_3_96;
mixer gate_output_3_96(.a(output_4_96), .b(output_4_1), .y(output_3_96));
wire output_5_96, output_5_1, output_4_96;
mixer gate_output_4_96(.a(output_5_96), .b(output_5_1), .y(output_4_96));
wire output_6_96, output_6_1, output_5_96;
mixer gate_output_5_96(.a(output_6_96), .b(output_6_1), .y(output_5_96));
wire output_7_96, output_7_1, output_6_96;
mixer gate_output_6_96(.a(output_7_96), .b(output_7_1), .y(output_6_96));
wire output_8_96, output_8_1, output_7_96;
mixer gate_output_7_96(.a(output_8_96), .b(output_8_1), .y(output_7_96));
wire output_9_96, output_9_1, output_8_96;
mixer gate_output_8_96(.a(output_9_96), .b(output_9_1), .y(output_8_96));
wire output_10_96, output_10_1, output_9_96;
mixer gate_output_9_96(.a(output_10_96), .b(output_10_1), .y(output_9_96));
wire output_11_96, output_11_1, output_10_96;
mixer gate_output_10_96(.a(output_11_96), .b(output_11_1), .y(output_10_96));
wire output_12_96, output_12_1, output_11_96;
mixer gate_output_11_96(.a(output_12_96), .b(output_12_1), .y(output_11_96));
wire output_13_96, output_13_1, output_12_96;
mixer gate_output_12_96(.a(output_13_96), .b(output_13_1), .y(output_12_96));
wire output_14_96, output_14_1, output_13_96;
mixer gate_output_13_96(.a(output_14_96), .b(output_14_1), .y(output_13_96));
wire output_15_96, output_15_1, output_14_96;
mixer gate_output_14_96(.a(output_15_96), .b(output_15_1), .y(output_14_96));
wire output_16_96, output_16_1, output_15_96;
mixer gate_output_15_96(.a(output_16_96), .b(output_16_1), .y(output_15_96));
wire output_1_97, output_1_2, output_0_97;
mixer gate_output_0_97(.a(output_1_97), .b(output_1_2), .y(output_0_97));
wire output_2_97, output_2_2, output_1_97;
mixer gate_output_1_97(.a(output_2_97), .b(output_2_2), .y(output_1_97));
wire output_3_97, output_3_2, output_2_97;
mixer gate_output_2_97(.a(output_3_97), .b(output_3_2), .y(output_2_97));
wire output_4_97, output_4_2, output_3_97;
mixer gate_output_3_97(.a(output_4_97), .b(output_4_2), .y(output_3_97));
wire output_5_97, output_5_2, output_4_97;
mixer gate_output_4_97(.a(output_5_97), .b(output_5_2), .y(output_4_97));
wire output_6_97, output_6_2, output_5_97;
mixer gate_output_5_97(.a(output_6_97), .b(output_6_2), .y(output_5_97));
wire output_7_97, output_7_2, output_6_97;
mixer gate_output_6_97(.a(output_7_97), .b(output_7_2), .y(output_6_97));
wire output_8_97, output_8_2, output_7_97;
mixer gate_output_7_97(.a(output_8_97), .b(output_8_2), .y(output_7_97));
wire output_9_97, output_9_2, output_8_97;
mixer gate_output_8_97(.a(output_9_97), .b(output_9_2), .y(output_8_97));
wire output_10_97, output_10_2, output_9_97;
mixer gate_output_9_97(.a(output_10_97), .b(output_10_2), .y(output_9_97));
wire output_11_97, output_11_2, output_10_97;
mixer gate_output_10_97(.a(output_11_97), .b(output_11_2), .y(output_10_97));
wire output_12_97, output_12_2, output_11_97;
mixer gate_output_11_97(.a(output_12_97), .b(output_12_2), .y(output_11_97));
wire output_13_97, output_13_2, output_12_97;
mixer gate_output_12_97(.a(output_13_97), .b(output_13_2), .y(output_12_97));
wire output_14_97, output_14_2, output_13_97;
mixer gate_output_13_97(.a(output_14_97), .b(output_14_2), .y(output_13_97));
wire output_15_97, output_15_2, output_14_97;
mixer gate_output_14_97(.a(output_15_97), .b(output_15_2), .y(output_14_97));
wire output_16_97, output_16_2, output_15_97;
mixer gate_output_15_97(.a(output_16_97), .b(output_16_2), .y(output_15_97));
wire output_1_98, output_1_3, output_0_98;
mixer gate_output_0_98(.a(output_1_98), .b(output_1_3), .y(output_0_98));
wire output_2_98, output_2_3, output_1_98;
mixer gate_output_1_98(.a(output_2_98), .b(output_2_3), .y(output_1_98));
wire output_3_98, output_3_3, output_2_98;
mixer gate_output_2_98(.a(output_3_98), .b(output_3_3), .y(output_2_98));
wire output_4_98, output_4_3, output_3_98;
mixer gate_output_3_98(.a(output_4_98), .b(output_4_3), .y(output_3_98));
wire output_5_98, output_5_3, output_4_98;
mixer gate_output_4_98(.a(output_5_98), .b(output_5_3), .y(output_4_98));
wire output_6_98, output_6_3, output_5_98;
mixer gate_output_5_98(.a(output_6_98), .b(output_6_3), .y(output_5_98));
wire output_7_98, output_7_3, output_6_98;
mixer gate_output_6_98(.a(output_7_98), .b(output_7_3), .y(output_6_98));
wire output_8_98, output_8_3, output_7_98;
mixer gate_output_7_98(.a(output_8_98), .b(output_8_3), .y(output_7_98));
wire output_9_98, output_9_3, output_8_98;
mixer gate_output_8_98(.a(output_9_98), .b(output_9_3), .y(output_8_98));
wire output_10_98, output_10_3, output_9_98;
mixer gate_output_9_98(.a(output_10_98), .b(output_10_3), .y(output_9_98));
wire output_11_98, output_11_3, output_10_98;
mixer gate_output_10_98(.a(output_11_98), .b(output_11_3), .y(output_10_98));
wire output_12_98, output_12_3, output_11_98;
mixer gate_output_11_98(.a(output_12_98), .b(output_12_3), .y(output_11_98));
wire output_13_98, output_13_3, output_12_98;
mixer gate_output_12_98(.a(output_13_98), .b(output_13_3), .y(output_12_98));
wire output_14_98, output_14_3, output_13_98;
mixer gate_output_13_98(.a(output_14_98), .b(output_14_3), .y(output_13_98));
wire output_15_98, output_15_3, output_14_98;
mixer gate_output_14_98(.a(output_15_98), .b(output_15_3), .y(output_14_98));
wire output_16_98, output_16_3, output_15_98;
mixer gate_output_15_98(.a(output_16_98), .b(output_16_3), .y(output_15_98));
wire output_1_99, output_1_4, output_0_99;
mixer gate_output_0_99(.a(output_1_99), .b(output_1_4), .y(output_0_99));
wire output_2_99, output_2_4, output_1_99;
mixer gate_output_1_99(.a(output_2_99), .b(output_2_4), .y(output_1_99));
wire output_3_99, output_3_4, output_2_99;
mixer gate_output_2_99(.a(output_3_99), .b(output_3_4), .y(output_2_99));
wire output_4_99, output_4_4, output_3_99;
mixer gate_output_3_99(.a(output_4_99), .b(output_4_4), .y(output_3_99));
wire output_5_99, output_5_4, output_4_99;
mixer gate_output_4_99(.a(output_5_99), .b(output_5_4), .y(output_4_99));
wire output_6_99, output_6_4, output_5_99;
mixer gate_output_5_99(.a(output_6_99), .b(output_6_4), .y(output_5_99));
wire output_7_99, output_7_4, output_6_99;
mixer gate_output_6_99(.a(output_7_99), .b(output_7_4), .y(output_6_99));
wire output_8_99, output_8_4, output_7_99;
mixer gate_output_7_99(.a(output_8_99), .b(output_8_4), .y(output_7_99));
wire output_9_99, output_9_4, output_8_99;
mixer gate_output_8_99(.a(output_9_99), .b(output_9_4), .y(output_8_99));
wire output_10_99, output_10_4, output_9_99;
mixer gate_output_9_99(.a(output_10_99), .b(output_10_4), .y(output_9_99));
wire output_11_99, output_11_4, output_10_99;
mixer gate_output_10_99(.a(output_11_99), .b(output_11_4), .y(output_10_99));
wire output_12_99, output_12_4, output_11_99;
mixer gate_output_11_99(.a(output_12_99), .b(output_12_4), .y(output_11_99));
wire output_13_99, output_13_4, output_12_99;
mixer gate_output_12_99(.a(output_13_99), .b(output_13_4), .y(output_12_99));
wire output_14_99, output_14_4, output_13_99;
mixer gate_output_13_99(.a(output_14_99), .b(output_14_4), .y(output_13_99));
wire output_15_99, output_15_4, output_14_99;
mixer gate_output_14_99(.a(output_15_99), .b(output_15_4), .y(output_14_99));
wire output_16_99, output_16_4, output_15_99;
mixer gate_output_15_99(.a(output_16_99), .b(output_16_4), .y(output_15_99));
wire output_1_100, output_1_5, output_0_100;
mixer gate_output_0_100(.a(output_1_100), .b(output_1_5), .y(output_0_100));
wire output_2_100, output_2_5, output_1_100;
mixer gate_output_1_100(.a(output_2_100), .b(output_2_5), .y(output_1_100));
wire output_3_100, output_3_5, output_2_100;
mixer gate_output_2_100(.a(output_3_100), .b(output_3_5), .y(output_2_100));
wire output_4_100, output_4_5, output_3_100;
mixer gate_output_3_100(.a(output_4_100), .b(output_4_5), .y(output_3_100));
wire output_5_100, output_5_5, output_4_100;
mixer gate_output_4_100(.a(output_5_100), .b(output_5_5), .y(output_4_100));
wire output_6_100, output_6_5, output_5_100;
mixer gate_output_5_100(.a(output_6_100), .b(output_6_5), .y(output_5_100));
wire output_7_100, output_7_5, output_6_100;
mixer gate_output_6_100(.a(output_7_100), .b(output_7_5), .y(output_6_100));
wire output_8_100, output_8_5, output_7_100;
mixer gate_output_7_100(.a(output_8_100), .b(output_8_5), .y(output_7_100));
wire output_9_100, output_9_5, output_8_100;
mixer gate_output_8_100(.a(output_9_100), .b(output_9_5), .y(output_8_100));
wire output_10_100, output_10_5, output_9_100;
mixer gate_output_9_100(.a(output_10_100), .b(output_10_5), .y(output_9_100));
wire output_11_100, output_11_5, output_10_100;
mixer gate_output_10_100(.a(output_11_100), .b(output_11_5), .y(output_10_100));
wire output_12_100, output_12_5, output_11_100;
mixer gate_output_11_100(.a(output_12_100), .b(output_12_5), .y(output_11_100));
wire output_13_100, output_13_5, output_12_100;
mixer gate_output_12_100(.a(output_13_100), .b(output_13_5), .y(output_12_100));
wire output_14_100, output_14_5, output_13_100;
mixer gate_output_13_100(.a(output_14_100), .b(output_14_5), .y(output_13_100));
wire output_15_100, output_15_5, output_14_100;
mixer gate_output_14_100(.a(output_15_100), .b(output_15_5), .y(output_14_100));
wire output_16_100, output_16_5, output_15_100;
mixer gate_output_15_100(.a(output_16_100), .b(output_16_5), .y(output_15_100));
wire output_1_101, output_1_6, output_0_101;
mixer gate_output_0_101(.a(output_1_101), .b(output_1_6), .y(output_0_101));
wire output_2_101, output_2_6, output_1_101;
mixer gate_output_1_101(.a(output_2_101), .b(output_2_6), .y(output_1_101));
wire output_3_101, output_3_6, output_2_101;
mixer gate_output_2_101(.a(output_3_101), .b(output_3_6), .y(output_2_101));
wire output_4_101, output_4_6, output_3_101;
mixer gate_output_3_101(.a(output_4_101), .b(output_4_6), .y(output_3_101));
wire output_5_101, output_5_6, output_4_101;
mixer gate_output_4_101(.a(output_5_101), .b(output_5_6), .y(output_4_101));
wire output_6_101, output_6_6, output_5_101;
mixer gate_output_5_101(.a(output_6_101), .b(output_6_6), .y(output_5_101));
wire output_7_101, output_7_6, output_6_101;
mixer gate_output_6_101(.a(output_7_101), .b(output_7_6), .y(output_6_101));
wire output_8_101, output_8_6, output_7_101;
mixer gate_output_7_101(.a(output_8_101), .b(output_8_6), .y(output_7_101));
wire output_9_101, output_9_6, output_8_101;
mixer gate_output_8_101(.a(output_9_101), .b(output_9_6), .y(output_8_101));
wire output_10_101, output_10_6, output_9_101;
mixer gate_output_9_101(.a(output_10_101), .b(output_10_6), .y(output_9_101));
wire output_11_101, output_11_6, output_10_101;
mixer gate_output_10_101(.a(output_11_101), .b(output_11_6), .y(output_10_101));
wire output_12_101, output_12_6, output_11_101;
mixer gate_output_11_101(.a(output_12_101), .b(output_12_6), .y(output_11_101));
wire output_13_101, output_13_6, output_12_101;
mixer gate_output_12_101(.a(output_13_101), .b(output_13_6), .y(output_12_101));
wire output_14_101, output_14_6, output_13_101;
mixer gate_output_13_101(.a(output_14_101), .b(output_14_6), .y(output_13_101));
wire output_15_101, output_15_6, output_14_101;
mixer gate_output_14_101(.a(output_15_101), .b(output_15_6), .y(output_14_101));
wire output_16_101, output_16_6, output_15_101;
mixer gate_output_15_101(.a(output_16_101), .b(output_16_6), .y(output_15_101));
wire output_1_102, output_1_7, output_0_102;
mixer gate_output_0_102(.a(output_1_102), .b(output_1_7), .y(output_0_102));
wire output_2_102, output_2_7, output_1_102;
mixer gate_output_1_102(.a(output_2_102), .b(output_2_7), .y(output_1_102));
wire output_3_102, output_3_7, output_2_102;
mixer gate_output_2_102(.a(output_3_102), .b(output_3_7), .y(output_2_102));
wire output_4_102, output_4_7, output_3_102;
mixer gate_output_3_102(.a(output_4_102), .b(output_4_7), .y(output_3_102));
wire output_5_102, output_5_7, output_4_102;
mixer gate_output_4_102(.a(output_5_102), .b(output_5_7), .y(output_4_102));
wire output_6_102, output_6_7, output_5_102;
mixer gate_output_5_102(.a(output_6_102), .b(output_6_7), .y(output_5_102));
wire output_7_102, output_7_7, output_6_102;
mixer gate_output_6_102(.a(output_7_102), .b(output_7_7), .y(output_6_102));
wire output_8_102, output_8_7, output_7_102;
mixer gate_output_7_102(.a(output_8_102), .b(output_8_7), .y(output_7_102));
wire output_9_102, output_9_7, output_8_102;
mixer gate_output_8_102(.a(output_9_102), .b(output_9_7), .y(output_8_102));
wire output_10_102, output_10_7, output_9_102;
mixer gate_output_9_102(.a(output_10_102), .b(output_10_7), .y(output_9_102));
wire output_11_102, output_11_7, output_10_102;
mixer gate_output_10_102(.a(output_11_102), .b(output_11_7), .y(output_10_102));
wire output_12_102, output_12_7, output_11_102;
mixer gate_output_11_102(.a(output_12_102), .b(output_12_7), .y(output_11_102));
wire output_13_102, output_13_7, output_12_102;
mixer gate_output_12_102(.a(output_13_102), .b(output_13_7), .y(output_12_102));
wire output_14_102, output_14_7, output_13_102;
mixer gate_output_13_102(.a(output_14_102), .b(output_14_7), .y(output_13_102));
wire output_15_102, output_15_7, output_14_102;
mixer gate_output_14_102(.a(output_15_102), .b(output_15_7), .y(output_14_102));
wire output_16_102, output_16_7, output_15_102;
mixer gate_output_15_102(.a(output_16_102), .b(output_16_7), .y(output_15_102));
wire output_1_103, output_1_8, output_0_103;
mixer gate_output_0_103(.a(output_1_103), .b(output_1_8), .y(output_0_103));
wire output_2_103, output_2_8, output_1_103;
mixer gate_output_1_103(.a(output_2_103), .b(output_2_8), .y(output_1_103));
wire output_3_103, output_3_8, output_2_103;
mixer gate_output_2_103(.a(output_3_103), .b(output_3_8), .y(output_2_103));
wire output_4_103, output_4_8, output_3_103;
mixer gate_output_3_103(.a(output_4_103), .b(output_4_8), .y(output_3_103));
wire output_5_103, output_5_8, output_4_103;
mixer gate_output_4_103(.a(output_5_103), .b(output_5_8), .y(output_4_103));
wire output_6_103, output_6_8, output_5_103;
mixer gate_output_5_103(.a(output_6_103), .b(output_6_8), .y(output_5_103));
wire output_7_103, output_7_8, output_6_103;
mixer gate_output_6_103(.a(output_7_103), .b(output_7_8), .y(output_6_103));
wire output_8_103, output_8_8, output_7_103;
mixer gate_output_7_103(.a(output_8_103), .b(output_8_8), .y(output_7_103));
wire output_9_103, output_9_8, output_8_103;
mixer gate_output_8_103(.a(output_9_103), .b(output_9_8), .y(output_8_103));
wire output_10_103, output_10_8, output_9_103;
mixer gate_output_9_103(.a(output_10_103), .b(output_10_8), .y(output_9_103));
wire output_11_103, output_11_8, output_10_103;
mixer gate_output_10_103(.a(output_11_103), .b(output_11_8), .y(output_10_103));
wire output_12_103, output_12_8, output_11_103;
mixer gate_output_11_103(.a(output_12_103), .b(output_12_8), .y(output_11_103));
wire output_13_103, output_13_8, output_12_103;
mixer gate_output_12_103(.a(output_13_103), .b(output_13_8), .y(output_12_103));
wire output_14_103, output_14_8, output_13_103;
mixer gate_output_13_103(.a(output_14_103), .b(output_14_8), .y(output_13_103));
wire output_15_103, output_15_8, output_14_103;
mixer gate_output_14_103(.a(output_15_103), .b(output_15_8), .y(output_14_103));
wire output_16_103, output_16_8, output_15_103;
mixer gate_output_15_103(.a(output_16_103), .b(output_16_8), .y(output_15_103));
wire output_1_104, output_1_9, output_0_104;
mixer gate_output_0_104(.a(output_1_104), .b(output_1_9), .y(output_0_104));
wire output_2_104, output_2_9, output_1_104;
mixer gate_output_1_104(.a(output_2_104), .b(output_2_9), .y(output_1_104));
wire output_3_104, output_3_9, output_2_104;
mixer gate_output_2_104(.a(output_3_104), .b(output_3_9), .y(output_2_104));
wire output_4_104, output_4_9, output_3_104;
mixer gate_output_3_104(.a(output_4_104), .b(output_4_9), .y(output_3_104));
wire output_5_104, output_5_9, output_4_104;
mixer gate_output_4_104(.a(output_5_104), .b(output_5_9), .y(output_4_104));
wire output_6_104, output_6_9, output_5_104;
mixer gate_output_5_104(.a(output_6_104), .b(output_6_9), .y(output_5_104));
wire output_7_104, output_7_9, output_6_104;
mixer gate_output_6_104(.a(output_7_104), .b(output_7_9), .y(output_6_104));
wire output_8_104, output_8_9, output_7_104;
mixer gate_output_7_104(.a(output_8_104), .b(output_8_9), .y(output_7_104));
wire output_9_104, output_9_9, output_8_104;
mixer gate_output_8_104(.a(output_9_104), .b(output_9_9), .y(output_8_104));
wire output_10_104, output_10_9, output_9_104;
mixer gate_output_9_104(.a(output_10_104), .b(output_10_9), .y(output_9_104));
wire output_11_104, output_11_9, output_10_104;
mixer gate_output_10_104(.a(output_11_104), .b(output_11_9), .y(output_10_104));
wire output_12_104, output_12_9, output_11_104;
mixer gate_output_11_104(.a(output_12_104), .b(output_12_9), .y(output_11_104));
wire output_13_104, output_13_9, output_12_104;
mixer gate_output_12_104(.a(output_13_104), .b(output_13_9), .y(output_12_104));
wire output_14_104, output_14_9, output_13_104;
mixer gate_output_13_104(.a(output_14_104), .b(output_14_9), .y(output_13_104));
wire output_15_104, output_15_9, output_14_104;
mixer gate_output_14_104(.a(output_15_104), .b(output_15_9), .y(output_14_104));
wire output_16_104, output_16_9, output_15_104;
mixer gate_output_15_104(.a(output_16_104), .b(output_16_9), .y(output_15_104));
wire output_1_105, output_1_10, output_0_105;
mixer gate_output_0_105(.a(output_1_105), .b(output_1_10), .y(output_0_105));
wire output_2_105, output_2_10, output_1_105;
mixer gate_output_1_105(.a(output_2_105), .b(output_2_10), .y(output_1_105));
wire output_3_105, output_3_10, output_2_105;
mixer gate_output_2_105(.a(output_3_105), .b(output_3_10), .y(output_2_105));
wire output_4_105, output_4_10, output_3_105;
mixer gate_output_3_105(.a(output_4_105), .b(output_4_10), .y(output_3_105));
wire output_5_105, output_5_10, output_4_105;
mixer gate_output_4_105(.a(output_5_105), .b(output_5_10), .y(output_4_105));
wire output_6_105, output_6_10, output_5_105;
mixer gate_output_5_105(.a(output_6_105), .b(output_6_10), .y(output_5_105));
wire output_7_105, output_7_10, output_6_105;
mixer gate_output_6_105(.a(output_7_105), .b(output_7_10), .y(output_6_105));
wire output_8_105, output_8_10, output_7_105;
mixer gate_output_7_105(.a(output_8_105), .b(output_8_10), .y(output_7_105));
wire output_9_105, output_9_10, output_8_105;
mixer gate_output_8_105(.a(output_9_105), .b(output_9_10), .y(output_8_105));
wire output_10_105, output_10_10, output_9_105;
mixer gate_output_9_105(.a(output_10_105), .b(output_10_10), .y(output_9_105));
wire output_11_105, output_11_10, output_10_105;
mixer gate_output_10_105(.a(output_11_105), .b(output_11_10), .y(output_10_105));
wire output_12_105, output_12_10, output_11_105;
mixer gate_output_11_105(.a(output_12_105), .b(output_12_10), .y(output_11_105));
wire output_13_105, output_13_10, output_12_105;
mixer gate_output_12_105(.a(output_13_105), .b(output_13_10), .y(output_12_105));
wire output_14_105, output_14_10, output_13_105;
mixer gate_output_13_105(.a(output_14_105), .b(output_14_10), .y(output_13_105));
wire output_15_105, output_15_10, output_14_105;
mixer gate_output_14_105(.a(output_15_105), .b(output_15_10), .y(output_14_105));
wire output_16_105, output_16_10, output_15_105;
mixer gate_output_15_105(.a(output_16_105), .b(output_16_10), .y(output_15_105));
wire output_1_106, output_1_11, output_0_106;
mixer gate_output_0_106(.a(output_1_106), .b(output_1_11), .y(output_0_106));
wire output_2_106, output_2_11, output_1_106;
mixer gate_output_1_106(.a(output_2_106), .b(output_2_11), .y(output_1_106));
wire output_3_106, output_3_11, output_2_106;
mixer gate_output_2_106(.a(output_3_106), .b(output_3_11), .y(output_2_106));
wire output_4_106, output_4_11, output_3_106;
mixer gate_output_3_106(.a(output_4_106), .b(output_4_11), .y(output_3_106));
wire output_5_106, output_5_11, output_4_106;
mixer gate_output_4_106(.a(output_5_106), .b(output_5_11), .y(output_4_106));
wire output_6_106, output_6_11, output_5_106;
mixer gate_output_5_106(.a(output_6_106), .b(output_6_11), .y(output_5_106));
wire output_7_106, output_7_11, output_6_106;
mixer gate_output_6_106(.a(output_7_106), .b(output_7_11), .y(output_6_106));
wire output_8_106, output_8_11, output_7_106;
mixer gate_output_7_106(.a(output_8_106), .b(output_8_11), .y(output_7_106));
wire output_9_106, output_9_11, output_8_106;
mixer gate_output_8_106(.a(output_9_106), .b(output_9_11), .y(output_8_106));
wire output_10_106, output_10_11, output_9_106;
mixer gate_output_9_106(.a(output_10_106), .b(output_10_11), .y(output_9_106));
wire output_11_106, output_11_11, output_10_106;
mixer gate_output_10_106(.a(output_11_106), .b(output_11_11), .y(output_10_106));
wire output_12_106, output_12_11, output_11_106;
mixer gate_output_11_106(.a(output_12_106), .b(output_12_11), .y(output_11_106));
wire output_13_106, output_13_11, output_12_106;
mixer gate_output_12_106(.a(output_13_106), .b(output_13_11), .y(output_12_106));
wire output_14_106, output_14_11, output_13_106;
mixer gate_output_13_106(.a(output_14_106), .b(output_14_11), .y(output_13_106));
wire output_15_106, output_15_11, output_14_106;
mixer gate_output_14_106(.a(output_15_106), .b(output_15_11), .y(output_14_106));
wire output_16_106, output_16_11, output_15_106;
mixer gate_output_15_106(.a(output_16_106), .b(output_16_11), .y(output_15_106));
wire output_1_107, output_1_12, output_0_107;
mixer gate_output_0_107(.a(output_1_107), .b(output_1_12), .y(output_0_107));
wire output_2_107, output_2_12, output_1_107;
mixer gate_output_1_107(.a(output_2_107), .b(output_2_12), .y(output_1_107));
wire output_3_107, output_3_12, output_2_107;
mixer gate_output_2_107(.a(output_3_107), .b(output_3_12), .y(output_2_107));
wire output_4_107, output_4_12, output_3_107;
mixer gate_output_3_107(.a(output_4_107), .b(output_4_12), .y(output_3_107));
wire output_5_107, output_5_12, output_4_107;
mixer gate_output_4_107(.a(output_5_107), .b(output_5_12), .y(output_4_107));
wire output_6_107, output_6_12, output_5_107;
mixer gate_output_5_107(.a(output_6_107), .b(output_6_12), .y(output_5_107));
wire output_7_107, output_7_12, output_6_107;
mixer gate_output_6_107(.a(output_7_107), .b(output_7_12), .y(output_6_107));
wire output_8_107, output_8_12, output_7_107;
mixer gate_output_7_107(.a(output_8_107), .b(output_8_12), .y(output_7_107));
wire output_9_107, output_9_12, output_8_107;
mixer gate_output_8_107(.a(output_9_107), .b(output_9_12), .y(output_8_107));
wire output_10_107, output_10_12, output_9_107;
mixer gate_output_9_107(.a(output_10_107), .b(output_10_12), .y(output_9_107));
wire output_11_107, output_11_12, output_10_107;
mixer gate_output_10_107(.a(output_11_107), .b(output_11_12), .y(output_10_107));
wire output_12_107, output_12_12, output_11_107;
mixer gate_output_11_107(.a(output_12_107), .b(output_12_12), .y(output_11_107));
wire output_13_107, output_13_12, output_12_107;
mixer gate_output_12_107(.a(output_13_107), .b(output_13_12), .y(output_12_107));
wire output_14_107, output_14_12, output_13_107;
mixer gate_output_13_107(.a(output_14_107), .b(output_14_12), .y(output_13_107));
wire output_15_107, output_15_12, output_14_107;
mixer gate_output_14_107(.a(output_15_107), .b(output_15_12), .y(output_14_107));
wire output_16_107, output_16_12, output_15_107;
mixer gate_output_15_107(.a(output_16_107), .b(output_16_12), .y(output_15_107));
wire output_1_108, output_1_13, output_0_108;
mixer gate_output_0_108(.a(output_1_108), .b(output_1_13), .y(output_0_108));
wire output_2_108, output_2_13, output_1_108;
mixer gate_output_1_108(.a(output_2_108), .b(output_2_13), .y(output_1_108));
wire output_3_108, output_3_13, output_2_108;
mixer gate_output_2_108(.a(output_3_108), .b(output_3_13), .y(output_2_108));
wire output_4_108, output_4_13, output_3_108;
mixer gate_output_3_108(.a(output_4_108), .b(output_4_13), .y(output_3_108));
wire output_5_108, output_5_13, output_4_108;
mixer gate_output_4_108(.a(output_5_108), .b(output_5_13), .y(output_4_108));
wire output_6_108, output_6_13, output_5_108;
mixer gate_output_5_108(.a(output_6_108), .b(output_6_13), .y(output_5_108));
wire output_7_108, output_7_13, output_6_108;
mixer gate_output_6_108(.a(output_7_108), .b(output_7_13), .y(output_6_108));
wire output_8_108, output_8_13, output_7_108;
mixer gate_output_7_108(.a(output_8_108), .b(output_8_13), .y(output_7_108));
wire output_9_108, output_9_13, output_8_108;
mixer gate_output_8_108(.a(output_9_108), .b(output_9_13), .y(output_8_108));
wire output_10_108, output_10_13, output_9_108;
mixer gate_output_9_108(.a(output_10_108), .b(output_10_13), .y(output_9_108));
wire output_11_108, output_11_13, output_10_108;
mixer gate_output_10_108(.a(output_11_108), .b(output_11_13), .y(output_10_108));
wire output_12_108, output_12_13, output_11_108;
mixer gate_output_11_108(.a(output_12_108), .b(output_12_13), .y(output_11_108));
wire output_13_108, output_13_13, output_12_108;
mixer gate_output_12_108(.a(output_13_108), .b(output_13_13), .y(output_12_108));
wire output_14_108, output_14_13, output_13_108;
mixer gate_output_13_108(.a(output_14_108), .b(output_14_13), .y(output_13_108));
wire output_15_108, output_15_13, output_14_108;
mixer gate_output_14_108(.a(output_15_108), .b(output_15_13), .y(output_14_108));
wire output_16_108, output_16_13, output_15_108;
mixer gate_output_15_108(.a(output_16_108), .b(output_16_13), .y(output_15_108));
wire output_1_109, output_1_14, output_0_109;
mixer gate_output_0_109(.a(output_1_109), .b(output_1_14), .y(output_0_109));
wire output_2_109, output_2_14, output_1_109;
mixer gate_output_1_109(.a(output_2_109), .b(output_2_14), .y(output_1_109));
wire output_3_109, output_3_14, output_2_109;
mixer gate_output_2_109(.a(output_3_109), .b(output_3_14), .y(output_2_109));
wire output_4_109, output_4_14, output_3_109;
mixer gate_output_3_109(.a(output_4_109), .b(output_4_14), .y(output_3_109));
wire output_5_109, output_5_14, output_4_109;
mixer gate_output_4_109(.a(output_5_109), .b(output_5_14), .y(output_4_109));
wire output_6_109, output_6_14, output_5_109;
mixer gate_output_5_109(.a(output_6_109), .b(output_6_14), .y(output_5_109));
wire output_7_109, output_7_14, output_6_109;
mixer gate_output_6_109(.a(output_7_109), .b(output_7_14), .y(output_6_109));
wire output_8_109, output_8_14, output_7_109;
mixer gate_output_7_109(.a(output_8_109), .b(output_8_14), .y(output_7_109));
wire output_9_109, output_9_14, output_8_109;
mixer gate_output_8_109(.a(output_9_109), .b(output_9_14), .y(output_8_109));
wire output_10_109, output_10_14, output_9_109;
mixer gate_output_9_109(.a(output_10_109), .b(output_10_14), .y(output_9_109));
wire output_11_109, output_11_14, output_10_109;
mixer gate_output_10_109(.a(output_11_109), .b(output_11_14), .y(output_10_109));
wire output_12_109, output_12_14, output_11_109;
mixer gate_output_11_109(.a(output_12_109), .b(output_12_14), .y(output_11_109));
wire output_13_109, output_13_14, output_12_109;
mixer gate_output_12_109(.a(output_13_109), .b(output_13_14), .y(output_12_109));
wire output_14_109, output_14_14, output_13_109;
mixer gate_output_13_109(.a(output_14_109), .b(output_14_14), .y(output_13_109));
wire output_15_109, output_15_14, output_14_109;
mixer gate_output_14_109(.a(output_15_109), .b(output_15_14), .y(output_14_109));
wire output_16_109, output_16_14, output_15_109;
mixer gate_output_15_109(.a(output_16_109), .b(output_16_14), .y(output_15_109));
wire output_1_110, output_1_15, output_0_110;
mixer gate_output_0_110(.a(output_1_110), .b(output_1_15), .y(output_0_110));
wire output_2_110, output_2_15, output_1_110;
mixer gate_output_1_110(.a(output_2_110), .b(output_2_15), .y(output_1_110));
wire output_3_110, output_3_15, output_2_110;
mixer gate_output_2_110(.a(output_3_110), .b(output_3_15), .y(output_2_110));
wire output_4_110, output_4_15, output_3_110;
mixer gate_output_3_110(.a(output_4_110), .b(output_4_15), .y(output_3_110));
wire output_5_110, output_5_15, output_4_110;
mixer gate_output_4_110(.a(output_5_110), .b(output_5_15), .y(output_4_110));
wire output_6_110, output_6_15, output_5_110;
mixer gate_output_5_110(.a(output_6_110), .b(output_6_15), .y(output_5_110));
wire output_7_110, output_7_15, output_6_110;
mixer gate_output_6_110(.a(output_7_110), .b(output_7_15), .y(output_6_110));
wire output_8_110, output_8_15, output_7_110;
mixer gate_output_7_110(.a(output_8_110), .b(output_8_15), .y(output_7_110));
wire output_9_110, output_9_15, output_8_110;
mixer gate_output_8_110(.a(output_9_110), .b(output_9_15), .y(output_8_110));
wire output_10_110, output_10_15, output_9_110;
mixer gate_output_9_110(.a(output_10_110), .b(output_10_15), .y(output_9_110));
wire output_11_110, output_11_15, output_10_110;
mixer gate_output_10_110(.a(output_11_110), .b(output_11_15), .y(output_10_110));
wire output_12_110, output_12_15, output_11_110;
mixer gate_output_11_110(.a(output_12_110), .b(output_12_15), .y(output_11_110));
wire output_13_110, output_13_15, output_12_110;
mixer gate_output_12_110(.a(output_13_110), .b(output_13_15), .y(output_12_110));
wire output_14_110, output_14_15, output_13_110;
mixer gate_output_13_110(.a(output_14_110), .b(output_14_15), .y(output_13_110));
wire output_15_110, output_15_15, output_14_110;
mixer gate_output_14_110(.a(output_15_110), .b(output_15_15), .y(output_14_110));
wire output_16_110, output_16_15, output_15_110;
mixer gate_output_15_110(.a(output_16_110), .b(output_16_15), .y(output_15_110));
wire output_1_111, output_1_0, output_0_111;
mixer gate_output_0_111(.a(output_1_111), .b(output_1_0), .y(output_0_111));
wire output_2_111, output_2_0, output_1_111;
mixer gate_output_1_111(.a(output_2_111), .b(output_2_0), .y(output_1_111));
wire output_3_111, output_3_0, output_2_111;
mixer gate_output_2_111(.a(output_3_111), .b(output_3_0), .y(output_2_111));
wire output_4_111, output_4_0, output_3_111;
mixer gate_output_3_111(.a(output_4_111), .b(output_4_0), .y(output_3_111));
wire output_5_111, output_5_0, output_4_111;
mixer gate_output_4_111(.a(output_5_111), .b(output_5_0), .y(output_4_111));
wire output_6_111, output_6_0, output_5_111;
mixer gate_output_5_111(.a(output_6_111), .b(output_6_0), .y(output_5_111));
wire output_7_111, output_7_0, output_6_111;
mixer gate_output_6_111(.a(output_7_111), .b(output_7_0), .y(output_6_111));
wire output_8_111, output_8_0, output_7_111;
mixer gate_output_7_111(.a(output_8_111), .b(output_8_0), .y(output_7_111));
wire output_9_111, output_9_0, output_8_111;
mixer gate_output_8_111(.a(output_9_111), .b(output_9_0), .y(output_8_111));
wire output_10_111, output_10_0, output_9_111;
mixer gate_output_9_111(.a(output_10_111), .b(output_10_0), .y(output_9_111));
wire output_11_111, output_11_0, output_10_111;
mixer gate_output_10_111(.a(output_11_111), .b(output_11_0), .y(output_10_111));
wire output_12_111, output_12_0, output_11_111;
mixer gate_output_11_111(.a(output_12_111), .b(output_12_0), .y(output_11_111));
wire output_13_111, output_13_0, output_12_111;
mixer gate_output_12_111(.a(output_13_111), .b(output_13_0), .y(output_12_111));
wire output_14_111, output_14_0, output_13_111;
mixer gate_output_13_111(.a(output_14_111), .b(output_14_0), .y(output_13_111));
wire output_15_111, output_15_0, output_14_111;
mixer gate_output_14_111(.a(output_15_111), .b(output_15_0), .y(output_14_111));
wire output_16_111, output_16_0, output_15_111;
mixer gate_output_15_111(.a(output_16_111), .b(output_16_0), .y(output_15_111));
wire output_1_112, output_1_1, output_0_112;
mixer gate_output_0_112(.a(output_1_112), .b(output_1_1), .y(output_0_112));
wire output_2_112, output_2_1, output_1_112;
mixer gate_output_1_112(.a(output_2_112), .b(output_2_1), .y(output_1_112));
wire output_3_112, output_3_1, output_2_112;
mixer gate_output_2_112(.a(output_3_112), .b(output_3_1), .y(output_2_112));
wire output_4_112, output_4_1, output_3_112;
mixer gate_output_3_112(.a(output_4_112), .b(output_4_1), .y(output_3_112));
wire output_5_112, output_5_1, output_4_112;
mixer gate_output_4_112(.a(output_5_112), .b(output_5_1), .y(output_4_112));
wire output_6_112, output_6_1, output_5_112;
mixer gate_output_5_112(.a(output_6_112), .b(output_6_1), .y(output_5_112));
wire output_7_112, output_7_1, output_6_112;
mixer gate_output_6_112(.a(output_7_112), .b(output_7_1), .y(output_6_112));
wire output_8_112, output_8_1, output_7_112;
mixer gate_output_7_112(.a(output_8_112), .b(output_8_1), .y(output_7_112));
wire output_9_112, output_9_1, output_8_112;
mixer gate_output_8_112(.a(output_9_112), .b(output_9_1), .y(output_8_112));
wire output_10_112, output_10_1, output_9_112;
mixer gate_output_9_112(.a(output_10_112), .b(output_10_1), .y(output_9_112));
wire output_11_112, output_11_1, output_10_112;
mixer gate_output_10_112(.a(output_11_112), .b(output_11_1), .y(output_10_112));
wire output_12_112, output_12_1, output_11_112;
mixer gate_output_11_112(.a(output_12_112), .b(output_12_1), .y(output_11_112));
wire output_13_112, output_13_1, output_12_112;
mixer gate_output_12_112(.a(output_13_112), .b(output_13_1), .y(output_12_112));
wire output_14_112, output_14_1, output_13_112;
mixer gate_output_13_112(.a(output_14_112), .b(output_14_1), .y(output_13_112));
wire output_15_112, output_15_1, output_14_112;
mixer gate_output_14_112(.a(output_15_112), .b(output_15_1), .y(output_14_112));
wire output_16_112, output_16_1, output_15_112;
mixer gate_output_15_112(.a(output_16_112), .b(output_16_1), .y(output_15_112));
wire output_1_113, output_1_2, output_0_113;
mixer gate_output_0_113(.a(output_1_113), .b(output_1_2), .y(output_0_113));
wire output_2_113, output_2_2, output_1_113;
mixer gate_output_1_113(.a(output_2_113), .b(output_2_2), .y(output_1_113));
wire output_3_113, output_3_2, output_2_113;
mixer gate_output_2_113(.a(output_3_113), .b(output_3_2), .y(output_2_113));
wire output_4_113, output_4_2, output_3_113;
mixer gate_output_3_113(.a(output_4_113), .b(output_4_2), .y(output_3_113));
wire output_5_113, output_5_2, output_4_113;
mixer gate_output_4_113(.a(output_5_113), .b(output_5_2), .y(output_4_113));
wire output_6_113, output_6_2, output_5_113;
mixer gate_output_5_113(.a(output_6_113), .b(output_6_2), .y(output_5_113));
wire output_7_113, output_7_2, output_6_113;
mixer gate_output_6_113(.a(output_7_113), .b(output_7_2), .y(output_6_113));
wire output_8_113, output_8_2, output_7_113;
mixer gate_output_7_113(.a(output_8_113), .b(output_8_2), .y(output_7_113));
wire output_9_113, output_9_2, output_8_113;
mixer gate_output_8_113(.a(output_9_113), .b(output_9_2), .y(output_8_113));
wire output_10_113, output_10_2, output_9_113;
mixer gate_output_9_113(.a(output_10_113), .b(output_10_2), .y(output_9_113));
wire output_11_113, output_11_2, output_10_113;
mixer gate_output_10_113(.a(output_11_113), .b(output_11_2), .y(output_10_113));
wire output_12_113, output_12_2, output_11_113;
mixer gate_output_11_113(.a(output_12_113), .b(output_12_2), .y(output_11_113));
wire output_13_113, output_13_2, output_12_113;
mixer gate_output_12_113(.a(output_13_113), .b(output_13_2), .y(output_12_113));
wire output_14_113, output_14_2, output_13_113;
mixer gate_output_13_113(.a(output_14_113), .b(output_14_2), .y(output_13_113));
wire output_15_113, output_15_2, output_14_113;
mixer gate_output_14_113(.a(output_15_113), .b(output_15_2), .y(output_14_113));
wire output_16_113, output_16_2, output_15_113;
mixer gate_output_15_113(.a(output_16_113), .b(output_16_2), .y(output_15_113));
wire output_1_114, output_1_3, output_0_114;
mixer gate_output_0_114(.a(output_1_114), .b(output_1_3), .y(output_0_114));
wire output_2_114, output_2_3, output_1_114;
mixer gate_output_1_114(.a(output_2_114), .b(output_2_3), .y(output_1_114));
wire output_3_114, output_3_3, output_2_114;
mixer gate_output_2_114(.a(output_3_114), .b(output_3_3), .y(output_2_114));
wire output_4_114, output_4_3, output_3_114;
mixer gate_output_3_114(.a(output_4_114), .b(output_4_3), .y(output_3_114));
wire output_5_114, output_5_3, output_4_114;
mixer gate_output_4_114(.a(output_5_114), .b(output_5_3), .y(output_4_114));
wire output_6_114, output_6_3, output_5_114;
mixer gate_output_5_114(.a(output_6_114), .b(output_6_3), .y(output_5_114));
wire output_7_114, output_7_3, output_6_114;
mixer gate_output_6_114(.a(output_7_114), .b(output_7_3), .y(output_6_114));
wire output_8_114, output_8_3, output_7_114;
mixer gate_output_7_114(.a(output_8_114), .b(output_8_3), .y(output_7_114));
wire output_9_114, output_9_3, output_8_114;
mixer gate_output_8_114(.a(output_9_114), .b(output_9_3), .y(output_8_114));
wire output_10_114, output_10_3, output_9_114;
mixer gate_output_9_114(.a(output_10_114), .b(output_10_3), .y(output_9_114));
wire output_11_114, output_11_3, output_10_114;
mixer gate_output_10_114(.a(output_11_114), .b(output_11_3), .y(output_10_114));
wire output_12_114, output_12_3, output_11_114;
mixer gate_output_11_114(.a(output_12_114), .b(output_12_3), .y(output_11_114));
wire output_13_114, output_13_3, output_12_114;
mixer gate_output_12_114(.a(output_13_114), .b(output_13_3), .y(output_12_114));
wire output_14_114, output_14_3, output_13_114;
mixer gate_output_13_114(.a(output_14_114), .b(output_14_3), .y(output_13_114));
wire output_15_114, output_15_3, output_14_114;
mixer gate_output_14_114(.a(output_15_114), .b(output_15_3), .y(output_14_114));
wire output_16_114, output_16_3, output_15_114;
mixer gate_output_15_114(.a(output_16_114), .b(output_16_3), .y(output_15_114));
wire output_1_115, output_1_4, output_0_115;
mixer gate_output_0_115(.a(output_1_115), .b(output_1_4), .y(output_0_115));
wire output_2_115, output_2_4, output_1_115;
mixer gate_output_1_115(.a(output_2_115), .b(output_2_4), .y(output_1_115));
wire output_3_115, output_3_4, output_2_115;
mixer gate_output_2_115(.a(output_3_115), .b(output_3_4), .y(output_2_115));
wire output_4_115, output_4_4, output_3_115;
mixer gate_output_3_115(.a(output_4_115), .b(output_4_4), .y(output_3_115));
wire output_5_115, output_5_4, output_4_115;
mixer gate_output_4_115(.a(output_5_115), .b(output_5_4), .y(output_4_115));
wire output_6_115, output_6_4, output_5_115;
mixer gate_output_5_115(.a(output_6_115), .b(output_6_4), .y(output_5_115));
wire output_7_115, output_7_4, output_6_115;
mixer gate_output_6_115(.a(output_7_115), .b(output_7_4), .y(output_6_115));
wire output_8_115, output_8_4, output_7_115;
mixer gate_output_7_115(.a(output_8_115), .b(output_8_4), .y(output_7_115));
wire output_9_115, output_9_4, output_8_115;
mixer gate_output_8_115(.a(output_9_115), .b(output_9_4), .y(output_8_115));
wire output_10_115, output_10_4, output_9_115;
mixer gate_output_9_115(.a(output_10_115), .b(output_10_4), .y(output_9_115));
wire output_11_115, output_11_4, output_10_115;
mixer gate_output_10_115(.a(output_11_115), .b(output_11_4), .y(output_10_115));
wire output_12_115, output_12_4, output_11_115;
mixer gate_output_11_115(.a(output_12_115), .b(output_12_4), .y(output_11_115));
wire output_13_115, output_13_4, output_12_115;
mixer gate_output_12_115(.a(output_13_115), .b(output_13_4), .y(output_12_115));
wire output_14_115, output_14_4, output_13_115;
mixer gate_output_13_115(.a(output_14_115), .b(output_14_4), .y(output_13_115));
wire output_15_115, output_15_4, output_14_115;
mixer gate_output_14_115(.a(output_15_115), .b(output_15_4), .y(output_14_115));
wire output_16_115, output_16_4, output_15_115;
mixer gate_output_15_115(.a(output_16_115), .b(output_16_4), .y(output_15_115));
wire output_1_116, output_1_5, output_0_116;
mixer gate_output_0_116(.a(output_1_116), .b(output_1_5), .y(output_0_116));
wire output_2_116, output_2_5, output_1_116;
mixer gate_output_1_116(.a(output_2_116), .b(output_2_5), .y(output_1_116));
wire output_3_116, output_3_5, output_2_116;
mixer gate_output_2_116(.a(output_3_116), .b(output_3_5), .y(output_2_116));
wire output_4_116, output_4_5, output_3_116;
mixer gate_output_3_116(.a(output_4_116), .b(output_4_5), .y(output_3_116));
wire output_5_116, output_5_5, output_4_116;
mixer gate_output_4_116(.a(output_5_116), .b(output_5_5), .y(output_4_116));
wire output_6_116, output_6_5, output_5_116;
mixer gate_output_5_116(.a(output_6_116), .b(output_6_5), .y(output_5_116));
wire output_7_116, output_7_5, output_6_116;
mixer gate_output_6_116(.a(output_7_116), .b(output_7_5), .y(output_6_116));
wire output_8_116, output_8_5, output_7_116;
mixer gate_output_7_116(.a(output_8_116), .b(output_8_5), .y(output_7_116));
wire output_9_116, output_9_5, output_8_116;
mixer gate_output_8_116(.a(output_9_116), .b(output_9_5), .y(output_8_116));
wire output_10_116, output_10_5, output_9_116;
mixer gate_output_9_116(.a(output_10_116), .b(output_10_5), .y(output_9_116));
wire output_11_116, output_11_5, output_10_116;
mixer gate_output_10_116(.a(output_11_116), .b(output_11_5), .y(output_10_116));
wire output_12_116, output_12_5, output_11_116;
mixer gate_output_11_116(.a(output_12_116), .b(output_12_5), .y(output_11_116));
wire output_13_116, output_13_5, output_12_116;
mixer gate_output_12_116(.a(output_13_116), .b(output_13_5), .y(output_12_116));
wire output_14_116, output_14_5, output_13_116;
mixer gate_output_13_116(.a(output_14_116), .b(output_14_5), .y(output_13_116));
wire output_15_116, output_15_5, output_14_116;
mixer gate_output_14_116(.a(output_15_116), .b(output_15_5), .y(output_14_116));
wire output_16_116, output_16_5, output_15_116;
mixer gate_output_15_116(.a(output_16_116), .b(output_16_5), .y(output_15_116));
wire output_1_117, output_1_6, output_0_117;
mixer gate_output_0_117(.a(output_1_117), .b(output_1_6), .y(output_0_117));
wire output_2_117, output_2_6, output_1_117;
mixer gate_output_1_117(.a(output_2_117), .b(output_2_6), .y(output_1_117));
wire output_3_117, output_3_6, output_2_117;
mixer gate_output_2_117(.a(output_3_117), .b(output_3_6), .y(output_2_117));
wire output_4_117, output_4_6, output_3_117;
mixer gate_output_3_117(.a(output_4_117), .b(output_4_6), .y(output_3_117));
wire output_5_117, output_5_6, output_4_117;
mixer gate_output_4_117(.a(output_5_117), .b(output_5_6), .y(output_4_117));
wire output_6_117, output_6_6, output_5_117;
mixer gate_output_5_117(.a(output_6_117), .b(output_6_6), .y(output_5_117));
wire output_7_117, output_7_6, output_6_117;
mixer gate_output_6_117(.a(output_7_117), .b(output_7_6), .y(output_6_117));
wire output_8_117, output_8_6, output_7_117;
mixer gate_output_7_117(.a(output_8_117), .b(output_8_6), .y(output_7_117));
wire output_9_117, output_9_6, output_8_117;
mixer gate_output_8_117(.a(output_9_117), .b(output_9_6), .y(output_8_117));
wire output_10_117, output_10_6, output_9_117;
mixer gate_output_9_117(.a(output_10_117), .b(output_10_6), .y(output_9_117));
wire output_11_117, output_11_6, output_10_117;
mixer gate_output_10_117(.a(output_11_117), .b(output_11_6), .y(output_10_117));
wire output_12_117, output_12_6, output_11_117;
mixer gate_output_11_117(.a(output_12_117), .b(output_12_6), .y(output_11_117));
wire output_13_117, output_13_6, output_12_117;
mixer gate_output_12_117(.a(output_13_117), .b(output_13_6), .y(output_12_117));
wire output_14_117, output_14_6, output_13_117;
mixer gate_output_13_117(.a(output_14_117), .b(output_14_6), .y(output_13_117));
wire output_15_117, output_15_6, output_14_117;
mixer gate_output_14_117(.a(output_15_117), .b(output_15_6), .y(output_14_117));
wire output_16_117, output_16_6, output_15_117;
mixer gate_output_15_117(.a(output_16_117), .b(output_16_6), .y(output_15_117));
wire output_1_118, output_1_7, output_0_118;
mixer gate_output_0_118(.a(output_1_118), .b(output_1_7), .y(output_0_118));
wire output_2_118, output_2_7, output_1_118;
mixer gate_output_1_118(.a(output_2_118), .b(output_2_7), .y(output_1_118));
wire output_3_118, output_3_7, output_2_118;
mixer gate_output_2_118(.a(output_3_118), .b(output_3_7), .y(output_2_118));
wire output_4_118, output_4_7, output_3_118;
mixer gate_output_3_118(.a(output_4_118), .b(output_4_7), .y(output_3_118));
wire output_5_118, output_5_7, output_4_118;
mixer gate_output_4_118(.a(output_5_118), .b(output_5_7), .y(output_4_118));
wire output_6_118, output_6_7, output_5_118;
mixer gate_output_5_118(.a(output_6_118), .b(output_6_7), .y(output_5_118));
wire output_7_118, output_7_7, output_6_118;
mixer gate_output_6_118(.a(output_7_118), .b(output_7_7), .y(output_6_118));
wire output_8_118, output_8_7, output_7_118;
mixer gate_output_7_118(.a(output_8_118), .b(output_8_7), .y(output_7_118));
wire output_9_118, output_9_7, output_8_118;
mixer gate_output_8_118(.a(output_9_118), .b(output_9_7), .y(output_8_118));
wire output_10_118, output_10_7, output_9_118;
mixer gate_output_9_118(.a(output_10_118), .b(output_10_7), .y(output_9_118));
wire output_11_118, output_11_7, output_10_118;
mixer gate_output_10_118(.a(output_11_118), .b(output_11_7), .y(output_10_118));
wire output_12_118, output_12_7, output_11_118;
mixer gate_output_11_118(.a(output_12_118), .b(output_12_7), .y(output_11_118));
wire output_13_118, output_13_7, output_12_118;
mixer gate_output_12_118(.a(output_13_118), .b(output_13_7), .y(output_12_118));
wire output_14_118, output_14_7, output_13_118;
mixer gate_output_13_118(.a(output_14_118), .b(output_14_7), .y(output_13_118));
wire output_15_118, output_15_7, output_14_118;
mixer gate_output_14_118(.a(output_15_118), .b(output_15_7), .y(output_14_118));
wire output_16_118, output_16_7, output_15_118;
mixer gate_output_15_118(.a(output_16_118), .b(output_16_7), .y(output_15_118));
wire output_1_119, output_1_8, output_0_119;
mixer gate_output_0_119(.a(output_1_119), .b(output_1_8), .y(output_0_119));
wire output_2_119, output_2_8, output_1_119;
mixer gate_output_1_119(.a(output_2_119), .b(output_2_8), .y(output_1_119));
wire output_3_119, output_3_8, output_2_119;
mixer gate_output_2_119(.a(output_3_119), .b(output_3_8), .y(output_2_119));
wire output_4_119, output_4_8, output_3_119;
mixer gate_output_3_119(.a(output_4_119), .b(output_4_8), .y(output_3_119));
wire output_5_119, output_5_8, output_4_119;
mixer gate_output_4_119(.a(output_5_119), .b(output_5_8), .y(output_4_119));
wire output_6_119, output_6_8, output_5_119;
mixer gate_output_5_119(.a(output_6_119), .b(output_6_8), .y(output_5_119));
wire output_7_119, output_7_8, output_6_119;
mixer gate_output_6_119(.a(output_7_119), .b(output_7_8), .y(output_6_119));
wire output_8_119, output_8_8, output_7_119;
mixer gate_output_7_119(.a(output_8_119), .b(output_8_8), .y(output_7_119));
wire output_9_119, output_9_8, output_8_119;
mixer gate_output_8_119(.a(output_9_119), .b(output_9_8), .y(output_8_119));
wire output_10_119, output_10_8, output_9_119;
mixer gate_output_9_119(.a(output_10_119), .b(output_10_8), .y(output_9_119));
wire output_11_119, output_11_8, output_10_119;
mixer gate_output_10_119(.a(output_11_119), .b(output_11_8), .y(output_10_119));
wire output_12_119, output_12_8, output_11_119;
mixer gate_output_11_119(.a(output_12_119), .b(output_12_8), .y(output_11_119));
wire output_13_119, output_13_8, output_12_119;
mixer gate_output_12_119(.a(output_13_119), .b(output_13_8), .y(output_12_119));
wire output_14_119, output_14_8, output_13_119;
mixer gate_output_13_119(.a(output_14_119), .b(output_14_8), .y(output_13_119));
wire output_15_119, output_15_8, output_14_119;
mixer gate_output_14_119(.a(output_15_119), .b(output_15_8), .y(output_14_119));
wire output_16_119, output_16_8, output_15_119;
mixer gate_output_15_119(.a(output_16_119), .b(output_16_8), .y(output_15_119));
wire output_1_120, output_1_9, output_0_120;
mixer gate_output_0_120(.a(output_1_120), .b(output_1_9), .y(output_0_120));
wire output_2_120, output_2_9, output_1_120;
mixer gate_output_1_120(.a(output_2_120), .b(output_2_9), .y(output_1_120));
wire output_3_120, output_3_9, output_2_120;
mixer gate_output_2_120(.a(output_3_120), .b(output_3_9), .y(output_2_120));
wire output_4_120, output_4_9, output_3_120;
mixer gate_output_3_120(.a(output_4_120), .b(output_4_9), .y(output_3_120));
wire output_5_120, output_5_9, output_4_120;
mixer gate_output_4_120(.a(output_5_120), .b(output_5_9), .y(output_4_120));
wire output_6_120, output_6_9, output_5_120;
mixer gate_output_5_120(.a(output_6_120), .b(output_6_9), .y(output_5_120));
wire output_7_120, output_7_9, output_6_120;
mixer gate_output_6_120(.a(output_7_120), .b(output_7_9), .y(output_6_120));
wire output_8_120, output_8_9, output_7_120;
mixer gate_output_7_120(.a(output_8_120), .b(output_8_9), .y(output_7_120));
wire output_9_120, output_9_9, output_8_120;
mixer gate_output_8_120(.a(output_9_120), .b(output_9_9), .y(output_8_120));
wire output_10_120, output_10_9, output_9_120;
mixer gate_output_9_120(.a(output_10_120), .b(output_10_9), .y(output_9_120));
wire output_11_120, output_11_9, output_10_120;
mixer gate_output_10_120(.a(output_11_120), .b(output_11_9), .y(output_10_120));
wire output_12_120, output_12_9, output_11_120;
mixer gate_output_11_120(.a(output_12_120), .b(output_12_9), .y(output_11_120));
wire output_13_120, output_13_9, output_12_120;
mixer gate_output_12_120(.a(output_13_120), .b(output_13_9), .y(output_12_120));
wire output_14_120, output_14_9, output_13_120;
mixer gate_output_13_120(.a(output_14_120), .b(output_14_9), .y(output_13_120));
wire output_15_120, output_15_9, output_14_120;
mixer gate_output_14_120(.a(output_15_120), .b(output_15_9), .y(output_14_120));
wire output_16_120, output_16_9, output_15_120;
mixer gate_output_15_120(.a(output_16_120), .b(output_16_9), .y(output_15_120));
wire output_1_121, output_1_10, output_0_121;
mixer gate_output_0_121(.a(output_1_121), .b(output_1_10), .y(output_0_121));
wire output_2_121, output_2_10, output_1_121;
mixer gate_output_1_121(.a(output_2_121), .b(output_2_10), .y(output_1_121));
wire output_3_121, output_3_10, output_2_121;
mixer gate_output_2_121(.a(output_3_121), .b(output_3_10), .y(output_2_121));
wire output_4_121, output_4_10, output_3_121;
mixer gate_output_3_121(.a(output_4_121), .b(output_4_10), .y(output_3_121));
wire output_5_121, output_5_10, output_4_121;
mixer gate_output_4_121(.a(output_5_121), .b(output_5_10), .y(output_4_121));
wire output_6_121, output_6_10, output_5_121;
mixer gate_output_5_121(.a(output_6_121), .b(output_6_10), .y(output_5_121));
wire output_7_121, output_7_10, output_6_121;
mixer gate_output_6_121(.a(output_7_121), .b(output_7_10), .y(output_6_121));
wire output_8_121, output_8_10, output_7_121;
mixer gate_output_7_121(.a(output_8_121), .b(output_8_10), .y(output_7_121));
wire output_9_121, output_9_10, output_8_121;
mixer gate_output_8_121(.a(output_9_121), .b(output_9_10), .y(output_8_121));
wire output_10_121, output_10_10, output_9_121;
mixer gate_output_9_121(.a(output_10_121), .b(output_10_10), .y(output_9_121));
wire output_11_121, output_11_10, output_10_121;
mixer gate_output_10_121(.a(output_11_121), .b(output_11_10), .y(output_10_121));
wire output_12_121, output_12_10, output_11_121;
mixer gate_output_11_121(.a(output_12_121), .b(output_12_10), .y(output_11_121));
wire output_13_121, output_13_10, output_12_121;
mixer gate_output_12_121(.a(output_13_121), .b(output_13_10), .y(output_12_121));
wire output_14_121, output_14_10, output_13_121;
mixer gate_output_13_121(.a(output_14_121), .b(output_14_10), .y(output_13_121));
wire output_15_121, output_15_10, output_14_121;
mixer gate_output_14_121(.a(output_15_121), .b(output_15_10), .y(output_14_121));
wire output_16_121, output_16_10, output_15_121;
mixer gate_output_15_121(.a(output_16_121), .b(output_16_10), .y(output_15_121));
wire output_1_122, output_1_11, output_0_122;
mixer gate_output_0_122(.a(output_1_122), .b(output_1_11), .y(output_0_122));
wire output_2_122, output_2_11, output_1_122;
mixer gate_output_1_122(.a(output_2_122), .b(output_2_11), .y(output_1_122));
wire output_3_122, output_3_11, output_2_122;
mixer gate_output_2_122(.a(output_3_122), .b(output_3_11), .y(output_2_122));
wire output_4_122, output_4_11, output_3_122;
mixer gate_output_3_122(.a(output_4_122), .b(output_4_11), .y(output_3_122));
wire output_5_122, output_5_11, output_4_122;
mixer gate_output_4_122(.a(output_5_122), .b(output_5_11), .y(output_4_122));
wire output_6_122, output_6_11, output_5_122;
mixer gate_output_5_122(.a(output_6_122), .b(output_6_11), .y(output_5_122));
wire output_7_122, output_7_11, output_6_122;
mixer gate_output_6_122(.a(output_7_122), .b(output_7_11), .y(output_6_122));
wire output_8_122, output_8_11, output_7_122;
mixer gate_output_7_122(.a(output_8_122), .b(output_8_11), .y(output_7_122));
wire output_9_122, output_9_11, output_8_122;
mixer gate_output_8_122(.a(output_9_122), .b(output_9_11), .y(output_8_122));
wire output_10_122, output_10_11, output_9_122;
mixer gate_output_9_122(.a(output_10_122), .b(output_10_11), .y(output_9_122));
wire output_11_122, output_11_11, output_10_122;
mixer gate_output_10_122(.a(output_11_122), .b(output_11_11), .y(output_10_122));
wire output_12_122, output_12_11, output_11_122;
mixer gate_output_11_122(.a(output_12_122), .b(output_12_11), .y(output_11_122));
wire output_13_122, output_13_11, output_12_122;
mixer gate_output_12_122(.a(output_13_122), .b(output_13_11), .y(output_12_122));
wire output_14_122, output_14_11, output_13_122;
mixer gate_output_13_122(.a(output_14_122), .b(output_14_11), .y(output_13_122));
wire output_15_122, output_15_11, output_14_122;
mixer gate_output_14_122(.a(output_15_122), .b(output_15_11), .y(output_14_122));
wire output_16_122, output_16_11, output_15_122;
mixer gate_output_15_122(.a(output_16_122), .b(output_16_11), .y(output_15_122));
wire output_1_123, output_1_12, output_0_123;
mixer gate_output_0_123(.a(output_1_123), .b(output_1_12), .y(output_0_123));
wire output_2_123, output_2_12, output_1_123;
mixer gate_output_1_123(.a(output_2_123), .b(output_2_12), .y(output_1_123));
wire output_3_123, output_3_12, output_2_123;
mixer gate_output_2_123(.a(output_3_123), .b(output_3_12), .y(output_2_123));
wire output_4_123, output_4_12, output_3_123;
mixer gate_output_3_123(.a(output_4_123), .b(output_4_12), .y(output_3_123));
wire output_5_123, output_5_12, output_4_123;
mixer gate_output_4_123(.a(output_5_123), .b(output_5_12), .y(output_4_123));
wire output_6_123, output_6_12, output_5_123;
mixer gate_output_5_123(.a(output_6_123), .b(output_6_12), .y(output_5_123));
wire output_7_123, output_7_12, output_6_123;
mixer gate_output_6_123(.a(output_7_123), .b(output_7_12), .y(output_6_123));
wire output_8_123, output_8_12, output_7_123;
mixer gate_output_7_123(.a(output_8_123), .b(output_8_12), .y(output_7_123));
wire output_9_123, output_9_12, output_8_123;
mixer gate_output_8_123(.a(output_9_123), .b(output_9_12), .y(output_8_123));
wire output_10_123, output_10_12, output_9_123;
mixer gate_output_9_123(.a(output_10_123), .b(output_10_12), .y(output_9_123));
wire output_11_123, output_11_12, output_10_123;
mixer gate_output_10_123(.a(output_11_123), .b(output_11_12), .y(output_10_123));
wire output_12_123, output_12_12, output_11_123;
mixer gate_output_11_123(.a(output_12_123), .b(output_12_12), .y(output_11_123));
wire output_13_123, output_13_12, output_12_123;
mixer gate_output_12_123(.a(output_13_123), .b(output_13_12), .y(output_12_123));
wire output_14_123, output_14_12, output_13_123;
mixer gate_output_13_123(.a(output_14_123), .b(output_14_12), .y(output_13_123));
wire output_15_123, output_15_12, output_14_123;
mixer gate_output_14_123(.a(output_15_123), .b(output_15_12), .y(output_14_123));
wire output_16_123, output_16_12, output_15_123;
mixer gate_output_15_123(.a(output_16_123), .b(output_16_12), .y(output_15_123));
wire output_1_124, output_1_13, output_0_124;
mixer gate_output_0_124(.a(output_1_124), .b(output_1_13), .y(output_0_124));
wire output_2_124, output_2_13, output_1_124;
mixer gate_output_1_124(.a(output_2_124), .b(output_2_13), .y(output_1_124));
wire output_3_124, output_3_13, output_2_124;
mixer gate_output_2_124(.a(output_3_124), .b(output_3_13), .y(output_2_124));
wire output_4_124, output_4_13, output_3_124;
mixer gate_output_3_124(.a(output_4_124), .b(output_4_13), .y(output_3_124));
wire output_5_124, output_5_13, output_4_124;
mixer gate_output_4_124(.a(output_5_124), .b(output_5_13), .y(output_4_124));
wire output_6_124, output_6_13, output_5_124;
mixer gate_output_5_124(.a(output_6_124), .b(output_6_13), .y(output_5_124));
wire output_7_124, output_7_13, output_6_124;
mixer gate_output_6_124(.a(output_7_124), .b(output_7_13), .y(output_6_124));
wire output_8_124, output_8_13, output_7_124;
mixer gate_output_7_124(.a(output_8_124), .b(output_8_13), .y(output_7_124));
wire output_9_124, output_9_13, output_8_124;
mixer gate_output_8_124(.a(output_9_124), .b(output_9_13), .y(output_8_124));
wire output_10_124, output_10_13, output_9_124;
mixer gate_output_9_124(.a(output_10_124), .b(output_10_13), .y(output_9_124));
wire output_11_124, output_11_13, output_10_124;
mixer gate_output_10_124(.a(output_11_124), .b(output_11_13), .y(output_10_124));
wire output_12_124, output_12_13, output_11_124;
mixer gate_output_11_124(.a(output_12_124), .b(output_12_13), .y(output_11_124));
wire output_13_124, output_13_13, output_12_124;
mixer gate_output_12_124(.a(output_13_124), .b(output_13_13), .y(output_12_124));
wire output_14_124, output_14_13, output_13_124;
mixer gate_output_13_124(.a(output_14_124), .b(output_14_13), .y(output_13_124));
wire output_15_124, output_15_13, output_14_124;
mixer gate_output_14_124(.a(output_15_124), .b(output_15_13), .y(output_14_124));
wire output_16_124, output_16_13, output_15_124;
mixer gate_output_15_124(.a(output_16_124), .b(output_16_13), .y(output_15_124));
wire output_1_125, output_1_14, output_0_125;
mixer gate_output_0_125(.a(output_1_125), .b(output_1_14), .y(output_0_125));
wire output_2_125, output_2_14, output_1_125;
mixer gate_output_1_125(.a(output_2_125), .b(output_2_14), .y(output_1_125));
wire output_3_125, output_3_14, output_2_125;
mixer gate_output_2_125(.a(output_3_125), .b(output_3_14), .y(output_2_125));
wire output_4_125, output_4_14, output_3_125;
mixer gate_output_3_125(.a(output_4_125), .b(output_4_14), .y(output_3_125));
wire output_5_125, output_5_14, output_4_125;
mixer gate_output_4_125(.a(output_5_125), .b(output_5_14), .y(output_4_125));
wire output_6_125, output_6_14, output_5_125;
mixer gate_output_5_125(.a(output_6_125), .b(output_6_14), .y(output_5_125));
wire output_7_125, output_7_14, output_6_125;
mixer gate_output_6_125(.a(output_7_125), .b(output_7_14), .y(output_6_125));
wire output_8_125, output_8_14, output_7_125;
mixer gate_output_7_125(.a(output_8_125), .b(output_8_14), .y(output_7_125));
wire output_9_125, output_9_14, output_8_125;
mixer gate_output_8_125(.a(output_9_125), .b(output_9_14), .y(output_8_125));
wire output_10_125, output_10_14, output_9_125;
mixer gate_output_9_125(.a(output_10_125), .b(output_10_14), .y(output_9_125));
wire output_11_125, output_11_14, output_10_125;
mixer gate_output_10_125(.a(output_11_125), .b(output_11_14), .y(output_10_125));
wire output_12_125, output_12_14, output_11_125;
mixer gate_output_11_125(.a(output_12_125), .b(output_12_14), .y(output_11_125));
wire output_13_125, output_13_14, output_12_125;
mixer gate_output_12_125(.a(output_13_125), .b(output_13_14), .y(output_12_125));
wire output_14_125, output_14_14, output_13_125;
mixer gate_output_13_125(.a(output_14_125), .b(output_14_14), .y(output_13_125));
wire output_15_125, output_15_14, output_14_125;
mixer gate_output_14_125(.a(output_15_125), .b(output_15_14), .y(output_14_125));
wire output_16_125, output_16_14, output_15_125;
mixer gate_output_15_125(.a(output_16_125), .b(output_16_14), .y(output_15_125));
wire output_1_126, output_1_15, output_0_126;
mixer gate_output_0_126(.a(output_1_126), .b(output_1_15), .y(output_0_126));
wire output_2_126, output_2_15, output_1_126;
mixer gate_output_1_126(.a(output_2_126), .b(output_2_15), .y(output_1_126));
wire output_3_126, output_3_15, output_2_126;
mixer gate_output_2_126(.a(output_3_126), .b(output_3_15), .y(output_2_126));
wire output_4_126, output_4_15, output_3_126;
mixer gate_output_3_126(.a(output_4_126), .b(output_4_15), .y(output_3_126));
wire output_5_126, output_5_15, output_4_126;
mixer gate_output_4_126(.a(output_5_126), .b(output_5_15), .y(output_4_126));
wire output_6_126, output_6_15, output_5_126;
mixer gate_output_5_126(.a(output_6_126), .b(output_6_15), .y(output_5_126));
wire output_7_126, output_7_15, output_6_126;
mixer gate_output_6_126(.a(output_7_126), .b(output_7_15), .y(output_6_126));
wire output_8_126, output_8_15, output_7_126;
mixer gate_output_7_126(.a(output_8_126), .b(output_8_15), .y(output_7_126));
wire output_9_126, output_9_15, output_8_126;
mixer gate_output_8_126(.a(output_9_126), .b(output_9_15), .y(output_8_126));
wire output_10_126, output_10_15, output_9_126;
mixer gate_output_9_126(.a(output_10_126), .b(output_10_15), .y(output_9_126));
wire output_11_126, output_11_15, output_10_126;
mixer gate_output_10_126(.a(output_11_126), .b(output_11_15), .y(output_10_126));
wire output_12_126, output_12_15, output_11_126;
mixer gate_output_11_126(.a(output_12_126), .b(output_12_15), .y(output_11_126));
wire output_13_126, output_13_15, output_12_126;
mixer gate_output_12_126(.a(output_13_126), .b(output_13_15), .y(output_12_126));
wire output_14_126, output_14_15, output_13_126;
mixer gate_output_13_126(.a(output_14_126), .b(output_14_15), .y(output_13_126));
wire output_15_126, output_15_15, output_14_126;
mixer gate_output_14_126(.a(output_15_126), .b(output_15_15), .y(output_14_126));
wire output_16_126, output_16_15, output_15_126;
mixer gate_output_15_126(.a(output_16_126), .b(output_16_15), .y(output_15_126));
wire output_1_127, output_1_0, output_0_127;
mixer gate_output_0_127(.a(output_1_127), .b(output_1_0), .y(output_0_127));
wire output_2_127, output_2_0, output_1_127;
mixer gate_output_1_127(.a(output_2_127), .b(output_2_0), .y(output_1_127));
wire output_3_127, output_3_0, output_2_127;
mixer gate_output_2_127(.a(output_3_127), .b(output_3_0), .y(output_2_127));
wire output_4_127, output_4_0, output_3_127;
mixer gate_output_3_127(.a(output_4_127), .b(output_4_0), .y(output_3_127));
wire output_5_127, output_5_0, output_4_127;
mixer gate_output_4_127(.a(output_5_127), .b(output_5_0), .y(output_4_127));
wire output_6_127, output_6_0, output_5_127;
mixer gate_output_5_127(.a(output_6_127), .b(output_6_0), .y(output_5_127));
wire output_7_127, output_7_0, output_6_127;
mixer gate_output_6_127(.a(output_7_127), .b(output_7_0), .y(output_6_127));
wire output_8_127, output_8_0, output_7_127;
mixer gate_output_7_127(.a(output_8_127), .b(output_8_0), .y(output_7_127));
wire output_9_127, output_9_0, output_8_127;
mixer gate_output_8_127(.a(output_9_127), .b(output_9_0), .y(output_8_127));
wire output_10_127, output_10_0, output_9_127;
mixer gate_output_9_127(.a(output_10_127), .b(output_10_0), .y(output_9_127));
wire output_11_127, output_11_0, output_10_127;
mixer gate_output_10_127(.a(output_11_127), .b(output_11_0), .y(output_10_127));
wire output_12_127, output_12_0, output_11_127;
mixer gate_output_11_127(.a(output_12_127), .b(output_12_0), .y(output_11_127));
wire output_13_127, output_13_0, output_12_127;
mixer gate_output_12_127(.a(output_13_127), .b(output_13_0), .y(output_12_127));
wire output_14_127, output_14_0, output_13_127;
mixer gate_output_13_127(.a(output_14_127), .b(output_14_0), .y(output_13_127));
wire output_15_127, output_15_0, output_14_127;
mixer gate_output_14_127(.a(output_15_127), .b(output_15_0), .y(output_14_127));
wire output_16_127, output_16_0, output_15_127;
mixer gate_output_15_127(.a(output_16_127), .b(output_16_0), .y(output_15_127));
wire output_1_128, output_1_1, output_0_128;
mixer gate_output_0_128(.a(output_1_128), .b(output_1_1), .y(output_0_128));
wire output_2_128, output_2_1, output_1_128;
mixer gate_output_1_128(.a(output_2_128), .b(output_2_1), .y(output_1_128));
wire output_3_128, output_3_1, output_2_128;
mixer gate_output_2_128(.a(output_3_128), .b(output_3_1), .y(output_2_128));
wire output_4_128, output_4_1, output_3_128;
mixer gate_output_3_128(.a(output_4_128), .b(output_4_1), .y(output_3_128));
wire output_5_128, output_5_1, output_4_128;
mixer gate_output_4_128(.a(output_5_128), .b(output_5_1), .y(output_4_128));
wire output_6_128, output_6_1, output_5_128;
mixer gate_output_5_128(.a(output_6_128), .b(output_6_1), .y(output_5_128));
wire output_7_128, output_7_1, output_6_128;
mixer gate_output_6_128(.a(output_7_128), .b(output_7_1), .y(output_6_128));
wire output_8_128, output_8_1, output_7_128;
mixer gate_output_7_128(.a(output_8_128), .b(output_8_1), .y(output_7_128));
wire output_9_128, output_9_1, output_8_128;
mixer gate_output_8_128(.a(output_9_128), .b(output_9_1), .y(output_8_128));
wire output_10_128, output_10_1, output_9_128;
mixer gate_output_9_128(.a(output_10_128), .b(output_10_1), .y(output_9_128));
wire output_11_128, output_11_1, output_10_128;
mixer gate_output_10_128(.a(output_11_128), .b(output_11_1), .y(output_10_128));
wire output_12_128, output_12_1, output_11_128;
mixer gate_output_11_128(.a(output_12_128), .b(output_12_1), .y(output_11_128));
wire output_13_128, output_13_1, output_12_128;
mixer gate_output_12_128(.a(output_13_128), .b(output_13_1), .y(output_12_128));
wire output_14_128, output_14_1, output_13_128;
mixer gate_output_13_128(.a(output_14_128), .b(output_14_1), .y(output_13_128));
wire output_15_128, output_15_1, output_14_128;
mixer gate_output_14_128(.a(output_15_128), .b(output_15_1), .y(output_14_128));
wire output_16_128, output_16_1, output_15_128;
mixer gate_output_15_128(.a(output_16_128), .b(output_16_1), .y(output_15_128));
wire output_1_129, output_1_2, output_0_129;
mixer gate_output_0_129(.a(output_1_129), .b(output_1_2), .y(output_0_129));
wire output_2_129, output_2_2, output_1_129;
mixer gate_output_1_129(.a(output_2_129), .b(output_2_2), .y(output_1_129));
wire output_3_129, output_3_2, output_2_129;
mixer gate_output_2_129(.a(output_3_129), .b(output_3_2), .y(output_2_129));
wire output_4_129, output_4_2, output_3_129;
mixer gate_output_3_129(.a(output_4_129), .b(output_4_2), .y(output_3_129));
wire output_5_129, output_5_2, output_4_129;
mixer gate_output_4_129(.a(output_5_129), .b(output_5_2), .y(output_4_129));
wire output_6_129, output_6_2, output_5_129;
mixer gate_output_5_129(.a(output_6_129), .b(output_6_2), .y(output_5_129));
wire output_7_129, output_7_2, output_6_129;
mixer gate_output_6_129(.a(output_7_129), .b(output_7_2), .y(output_6_129));
wire output_8_129, output_8_2, output_7_129;
mixer gate_output_7_129(.a(output_8_129), .b(output_8_2), .y(output_7_129));
wire output_9_129, output_9_2, output_8_129;
mixer gate_output_8_129(.a(output_9_129), .b(output_9_2), .y(output_8_129));
wire output_10_129, output_10_2, output_9_129;
mixer gate_output_9_129(.a(output_10_129), .b(output_10_2), .y(output_9_129));
wire output_11_129, output_11_2, output_10_129;
mixer gate_output_10_129(.a(output_11_129), .b(output_11_2), .y(output_10_129));
wire output_12_129, output_12_2, output_11_129;
mixer gate_output_11_129(.a(output_12_129), .b(output_12_2), .y(output_11_129));
wire output_13_129, output_13_2, output_12_129;
mixer gate_output_12_129(.a(output_13_129), .b(output_13_2), .y(output_12_129));
wire output_14_129, output_14_2, output_13_129;
mixer gate_output_13_129(.a(output_14_129), .b(output_14_2), .y(output_13_129));
wire output_15_129, output_15_2, output_14_129;
mixer gate_output_14_129(.a(output_15_129), .b(output_15_2), .y(output_14_129));
wire output_16_129, output_16_2, output_15_129;
mixer gate_output_15_129(.a(output_16_129), .b(output_16_2), .y(output_15_129));
wire output_1_130, output_1_3, output_0_130;
mixer gate_output_0_130(.a(output_1_130), .b(output_1_3), .y(output_0_130));
wire output_2_130, output_2_3, output_1_130;
mixer gate_output_1_130(.a(output_2_130), .b(output_2_3), .y(output_1_130));
wire output_3_130, output_3_3, output_2_130;
mixer gate_output_2_130(.a(output_3_130), .b(output_3_3), .y(output_2_130));
wire output_4_130, output_4_3, output_3_130;
mixer gate_output_3_130(.a(output_4_130), .b(output_4_3), .y(output_3_130));
wire output_5_130, output_5_3, output_4_130;
mixer gate_output_4_130(.a(output_5_130), .b(output_5_3), .y(output_4_130));
wire output_6_130, output_6_3, output_5_130;
mixer gate_output_5_130(.a(output_6_130), .b(output_6_3), .y(output_5_130));
wire output_7_130, output_7_3, output_6_130;
mixer gate_output_6_130(.a(output_7_130), .b(output_7_3), .y(output_6_130));
wire output_8_130, output_8_3, output_7_130;
mixer gate_output_7_130(.a(output_8_130), .b(output_8_3), .y(output_7_130));
wire output_9_130, output_9_3, output_8_130;
mixer gate_output_8_130(.a(output_9_130), .b(output_9_3), .y(output_8_130));
wire output_10_130, output_10_3, output_9_130;
mixer gate_output_9_130(.a(output_10_130), .b(output_10_3), .y(output_9_130));
wire output_11_130, output_11_3, output_10_130;
mixer gate_output_10_130(.a(output_11_130), .b(output_11_3), .y(output_10_130));
wire output_12_130, output_12_3, output_11_130;
mixer gate_output_11_130(.a(output_12_130), .b(output_12_3), .y(output_11_130));
wire output_13_130, output_13_3, output_12_130;
mixer gate_output_12_130(.a(output_13_130), .b(output_13_3), .y(output_12_130));
wire output_14_130, output_14_3, output_13_130;
mixer gate_output_13_130(.a(output_14_130), .b(output_14_3), .y(output_13_130));
wire output_15_130, output_15_3, output_14_130;
mixer gate_output_14_130(.a(output_15_130), .b(output_15_3), .y(output_14_130));
wire output_16_130, output_16_3, output_15_130;
mixer gate_output_15_130(.a(output_16_130), .b(output_16_3), .y(output_15_130));
wire output_1_131, output_1_4, output_0_131;
mixer gate_output_0_131(.a(output_1_131), .b(output_1_4), .y(output_0_131));
wire output_2_131, output_2_4, output_1_131;
mixer gate_output_1_131(.a(output_2_131), .b(output_2_4), .y(output_1_131));
wire output_3_131, output_3_4, output_2_131;
mixer gate_output_2_131(.a(output_3_131), .b(output_3_4), .y(output_2_131));
wire output_4_131, output_4_4, output_3_131;
mixer gate_output_3_131(.a(output_4_131), .b(output_4_4), .y(output_3_131));
wire output_5_131, output_5_4, output_4_131;
mixer gate_output_4_131(.a(output_5_131), .b(output_5_4), .y(output_4_131));
wire output_6_131, output_6_4, output_5_131;
mixer gate_output_5_131(.a(output_6_131), .b(output_6_4), .y(output_5_131));
wire output_7_131, output_7_4, output_6_131;
mixer gate_output_6_131(.a(output_7_131), .b(output_7_4), .y(output_6_131));
wire output_8_131, output_8_4, output_7_131;
mixer gate_output_7_131(.a(output_8_131), .b(output_8_4), .y(output_7_131));
wire output_9_131, output_9_4, output_8_131;
mixer gate_output_8_131(.a(output_9_131), .b(output_9_4), .y(output_8_131));
wire output_10_131, output_10_4, output_9_131;
mixer gate_output_9_131(.a(output_10_131), .b(output_10_4), .y(output_9_131));
wire output_11_131, output_11_4, output_10_131;
mixer gate_output_10_131(.a(output_11_131), .b(output_11_4), .y(output_10_131));
wire output_12_131, output_12_4, output_11_131;
mixer gate_output_11_131(.a(output_12_131), .b(output_12_4), .y(output_11_131));
wire output_13_131, output_13_4, output_12_131;
mixer gate_output_12_131(.a(output_13_131), .b(output_13_4), .y(output_12_131));
wire output_14_131, output_14_4, output_13_131;
mixer gate_output_13_131(.a(output_14_131), .b(output_14_4), .y(output_13_131));
wire output_15_131, output_15_4, output_14_131;
mixer gate_output_14_131(.a(output_15_131), .b(output_15_4), .y(output_14_131));
wire output_16_131, output_16_4, output_15_131;
mixer gate_output_15_131(.a(output_16_131), .b(output_16_4), .y(output_15_131));
wire output_1_132, output_1_5, output_0_132;
mixer gate_output_0_132(.a(output_1_132), .b(output_1_5), .y(output_0_132));
wire output_2_132, output_2_5, output_1_132;
mixer gate_output_1_132(.a(output_2_132), .b(output_2_5), .y(output_1_132));
wire output_3_132, output_3_5, output_2_132;
mixer gate_output_2_132(.a(output_3_132), .b(output_3_5), .y(output_2_132));
wire output_4_132, output_4_5, output_3_132;
mixer gate_output_3_132(.a(output_4_132), .b(output_4_5), .y(output_3_132));
wire output_5_132, output_5_5, output_4_132;
mixer gate_output_4_132(.a(output_5_132), .b(output_5_5), .y(output_4_132));
wire output_6_132, output_6_5, output_5_132;
mixer gate_output_5_132(.a(output_6_132), .b(output_6_5), .y(output_5_132));
wire output_7_132, output_7_5, output_6_132;
mixer gate_output_6_132(.a(output_7_132), .b(output_7_5), .y(output_6_132));
wire output_8_132, output_8_5, output_7_132;
mixer gate_output_7_132(.a(output_8_132), .b(output_8_5), .y(output_7_132));
wire output_9_132, output_9_5, output_8_132;
mixer gate_output_8_132(.a(output_9_132), .b(output_9_5), .y(output_8_132));
wire output_10_132, output_10_5, output_9_132;
mixer gate_output_9_132(.a(output_10_132), .b(output_10_5), .y(output_9_132));
wire output_11_132, output_11_5, output_10_132;
mixer gate_output_10_132(.a(output_11_132), .b(output_11_5), .y(output_10_132));
wire output_12_132, output_12_5, output_11_132;
mixer gate_output_11_132(.a(output_12_132), .b(output_12_5), .y(output_11_132));
wire output_13_132, output_13_5, output_12_132;
mixer gate_output_12_132(.a(output_13_132), .b(output_13_5), .y(output_12_132));
wire output_14_132, output_14_5, output_13_132;
mixer gate_output_13_132(.a(output_14_132), .b(output_14_5), .y(output_13_132));
wire output_15_132, output_15_5, output_14_132;
mixer gate_output_14_132(.a(output_15_132), .b(output_15_5), .y(output_14_132));
wire output_16_132, output_16_5, output_15_132;
mixer gate_output_15_132(.a(output_16_132), .b(output_16_5), .y(output_15_132));
wire output_1_133, output_1_6, output_0_133;
mixer gate_output_0_133(.a(output_1_133), .b(output_1_6), .y(output_0_133));
wire output_2_133, output_2_6, output_1_133;
mixer gate_output_1_133(.a(output_2_133), .b(output_2_6), .y(output_1_133));
wire output_3_133, output_3_6, output_2_133;
mixer gate_output_2_133(.a(output_3_133), .b(output_3_6), .y(output_2_133));
wire output_4_133, output_4_6, output_3_133;
mixer gate_output_3_133(.a(output_4_133), .b(output_4_6), .y(output_3_133));
wire output_5_133, output_5_6, output_4_133;
mixer gate_output_4_133(.a(output_5_133), .b(output_5_6), .y(output_4_133));
wire output_6_133, output_6_6, output_5_133;
mixer gate_output_5_133(.a(output_6_133), .b(output_6_6), .y(output_5_133));
wire output_7_133, output_7_6, output_6_133;
mixer gate_output_6_133(.a(output_7_133), .b(output_7_6), .y(output_6_133));
wire output_8_133, output_8_6, output_7_133;
mixer gate_output_7_133(.a(output_8_133), .b(output_8_6), .y(output_7_133));
wire output_9_133, output_9_6, output_8_133;
mixer gate_output_8_133(.a(output_9_133), .b(output_9_6), .y(output_8_133));
wire output_10_133, output_10_6, output_9_133;
mixer gate_output_9_133(.a(output_10_133), .b(output_10_6), .y(output_9_133));
wire output_11_133, output_11_6, output_10_133;
mixer gate_output_10_133(.a(output_11_133), .b(output_11_6), .y(output_10_133));
wire output_12_133, output_12_6, output_11_133;
mixer gate_output_11_133(.a(output_12_133), .b(output_12_6), .y(output_11_133));
wire output_13_133, output_13_6, output_12_133;
mixer gate_output_12_133(.a(output_13_133), .b(output_13_6), .y(output_12_133));
wire output_14_133, output_14_6, output_13_133;
mixer gate_output_13_133(.a(output_14_133), .b(output_14_6), .y(output_13_133));
wire output_15_133, output_15_6, output_14_133;
mixer gate_output_14_133(.a(output_15_133), .b(output_15_6), .y(output_14_133));
wire output_16_133, output_16_6, output_15_133;
mixer gate_output_15_133(.a(output_16_133), .b(output_16_6), .y(output_15_133));
wire output_1_134, output_1_7, output_0_134;
mixer gate_output_0_134(.a(output_1_134), .b(output_1_7), .y(output_0_134));
wire output_2_134, output_2_7, output_1_134;
mixer gate_output_1_134(.a(output_2_134), .b(output_2_7), .y(output_1_134));
wire output_3_134, output_3_7, output_2_134;
mixer gate_output_2_134(.a(output_3_134), .b(output_3_7), .y(output_2_134));
wire output_4_134, output_4_7, output_3_134;
mixer gate_output_3_134(.a(output_4_134), .b(output_4_7), .y(output_3_134));
wire output_5_134, output_5_7, output_4_134;
mixer gate_output_4_134(.a(output_5_134), .b(output_5_7), .y(output_4_134));
wire output_6_134, output_6_7, output_5_134;
mixer gate_output_5_134(.a(output_6_134), .b(output_6_7), .y(output_5_134));
wire output_7_134, output_7_7, output_6_134;
mixer gate_output_6_134(.a(output_7_134), .b(output_7_7), .y(output_6_134));
wire output_8_134, output_8_7, output_7_134;
mixer gate_output_7_134(.a(output_8_134), .b(output_8_7), .y(output_7_134));
wire output_9_134, output_9_7, output_8_134;
mixer gate_output_8_134(.a(output_9_134), .b(output_9_7), .y(output_8_134));
wire output_10_134, output_10_7, output_9_134;
mixer gate_output_9_134(.a(output_10_134), .b(output_10_7), .y(output_9_134));
wire output_11_134, output_11_7, output_10_134;
mixer gate_output_10_134(.a(output_11_134), .b(output_11_7), .y(output_10_134));
wire output_12_134, output_12_7, output_11_134;
mixer gate_output_11_134(.a(output_12_134), .b(output_12_7), .y(output_11_134));
wire output_13_134, output_13_7, output_12_134;
mixer gate_output_12_134(.a(output_13_134), .b(output_13_7), .y(output_12_134));
wire output_14_134, output_14_7, output_13_134;
mixer gate_output_13_134(.a(output_14_134), .b(output_14_7), .y(output_13_134));
wire output_15_134, output_15_7, output_14_134;
mixer gate_output_14_134(.a(output_15_134), .b(output_15_7), .y(output_14_134));
wire output_16_134, output_16_7, output_15_134;
mixer gate_output_15_134(.a(output_16_134), .b(output_16_7), .y(output_15_134));
wire output_1_135, output_1_8, output_0_135;
mixer gate_output_0_135(.a(output_1_135), .b(output_1_8), .y(output_0_135));
wire output_2_135, output_2_8, output_1_135;
mixer gate_output_1_135(.a(output_2_135), .b(output_2_8), .y(output_1_135));
wire output_3_135, output_3_8, output_2_135;
mixer gate_output_2_135(.a(output_3_135), .b(output_3_8), .y(output_2_135));
wire output_4_135, output_4_8, output_3_135;
mixer gate_output_3_135(.a(output_4_135), .b(output_4_8), .y(output_3_135));
wire output_5_135, output_5_8, output_4_135;
mixer gate_output_4_135(.a(output_5_135), .b(output_5_8), .y(output_4_135));
wire output_6_135, output_6_8, output_5_135;
mixer gate_output_5_135(.a(output_6_135), .b(output_6_8), .y(output_5_135));
wire output_7_135, output_7_8, output_6_135;
mixer gate_output_6_135(.a(output_7_135), .b(output_7_8), .y(output_6_135));
wire output_8_135, output_8_8, output_7_135;
mixer gate_output_7_135(.a(output_8_135), .b(output_8_8), .y(output_7_135));
wire output_9_135, output_9_8, output_8_135;
mixer gate_output_8_135(.a(output_9_135), .b(output_9_8), .y(output_8_135));
wire output_10_135, output_10_8, output_9_135;
mixer gate_output_9_135(.a(output_10_135), .b(output_10_8), .y(output_9_135));
wire output_11_135, output_11_8, output_10_135;
mixer gate_output_10_135(.a(output_11_135), .b(output_11_8), .y(output_10_135));
wire output_12_135, output_12_8, output_11_135;
mixer gate_output_11_135(.a(output_12_135), .b(output_12_8), .y(output_11_135));
wire output_13_135, output_13_8, output_12_135;
mixer gate_output_12_135(.a(output_13_135), .b(output_13_8), .y(output_12_135));
wire output_14_135, output_14_8, output_13_135;
mixer gate_output_13_135(.a(output_14_135), .b(output_14_8), .y(output_13_135));
wire output_15_135, output_15_8, output_14_135;
mixer gate_output_14_135(.a(output_15_135), .b(output_15_8), .y(output_14_135));
wire output_16_135, output_16_8, output_15_135;
mixer gate_output_15_135(.a(output_16_135), .b(output_16_8), .y(output_15_135));
wire output_1_136, output_1_9, output_0_136;
mixer gate_output_0_136(.a(output_1_136), .b(output_1_9), .y(output_0_136));
wire output_2_136, output_2_9, output_1_136;
mixer gate_output_1_136(.a(output_2_136), .b(output_2_9), .y(output_1_136));
wire output_3_136, output_3_9, output_2_136;
mixer gate_output_2_136(.a(output_3_136), .b(output_3_9), .y(output_2_136));
wire output_4_136, output_4_9, output_3_136;
mixer gate_output_3_136(.a(output_4_136), .b(output_4_9), .y(output_3_136));
wire output_5_136, output_5_9, output_4_136;
mixer gate_output_4_136(.a(output_5_136), .b(output_5_9), .y(output_4_136));
wire output_6_136, output_6_9, output_5_136;
mixer gate_output_5_136(.a(output_6_136), .b(output_6_9), .y(output_5_136));
wire output_7_136, output_7_9, output_6_136;
mixer gate_output_6_136(.a(output_7_136), .b(output_7_9), .y(output_6_136));
wire output_8_136, output_8_9, output_7_136;
mixer gate_output_7_136(.a(output_8_136), .b(output_8_9), .y(output_7_136));
wire output_9_136, output_9_9, output_8_136;
mixer gate_output_8_136(.a(output_9_136), .b(output_9_9), .y(output_8_136));
wire output_10_136, output_10_9, output_9_136;
mixer gate_output_9_136(.a(output_10_136), .b(output_10_9), .y(output_9_136));
wire output_11_136, output_11_9, output_10_136;
mixer gate_output_10_136(.a(output_11_136), .b(output_11_9), .y(output_10_136));
wire output_12_136, output_12_9, output_11_136;
mixer gate_output_11_136(.a(output_12_136), .b(output_12_9), .y(output_11_136));
wire output_13_136, output_13_9, output_12_136;
mixer gate_output_12_136(.a(output_13_136), .b(output_13_9), .y(output_12_136));
wire output_14_136, output_14_9, output_13_136;
mixer gate_output_13_136(.a(output_14_136), .b(output_14_9), .y(output_13_136));
wire output_15_136, output_15_9, output_14_136;
mixer gate_output_14_136(.a(output_15_136), .b(output_15_9), .y(output_14_136));
wire output_16_136, output_16_9, output_15_136;
mixer gate_output_15_136(.a(output_16_136), .b(output_16_9), .y(output_15_136));
wire output_1_137, output_1_10, output_0_137;
mixer gate_output_0_137(.a(output_1_137), .b(output_1_10), .y(output_0_137));
wire output_2_137, output_2_10, output_1_137;
mixer gate_output_1_137(.a(output_2_137), .b(output_2_10), .y(output_1_137));
wire output_3_137, output_3_10, output_2_137;
mixer gate_output_2_137(.a(output_3_137), .b(output_3_10), .y(output_2_137));
wire output_4_137, output_4_10, output_3_137;
mixer gate_output_3_137(.a(output_4_137), .b(output_4_10), .y(output_3_137));
wire output_5_137, output_5_10, output_4_137;
mixer gate_output_4_137(.a(output_5_137), .b(output_5_10), .y(output_4_137));
wire output_6_137, output_6_10, output_5_137;
mixer gate_output_5_137(.a(output_6_137), .b(output_6_10), .y(output_5_137));
wire output_7_137, output_7_10, output_6_137;
mixer gate_output_6_137(.a(output_7_137), .b(output_7_10), .y(output_6_137));
wire output_8_137, output_8_10, output_7_137;
mixer gate_output_7_137(.a(output_8_137), .b(output_8_10), .y(output_7_137));
wire output_9_137, output_9_10, output_8_137;
mixer gate_output_8_137(.a(output_9_137), .b(output_9_10), .y(output_8_137));
wire output_10_137, output_10_10, output_9_137;
mixer gate_output_9_137(.a(output_10_137), .b(output_10_10), .y(output_9_137));
wire output_11_137, output_11_10, output_10_137;
mixer gate_output_10_137(.a(output_11_137), .b(output_11_10), .y(output_10_137));
wire output_12_137, output_12_10, output_11_137;
mixer gate_output_11_137(.a(output_12_137), .b(output_12_10), .y(output_11_137));
wire output_13_137, output_13_10, output_12_137;
mixer gate_output_12_137(.a(output_13_137), .b(output_13_10), .y(output_12_137));
wire output_14_137, output_14_10, output_13_137;
mixer gate_output_13_137(.a(output_14_137), .b(output_14_10), .y(output_13_137));
wire output_15_137, output_15_10, output_14_137;
mixer gate_output_14_137(.a(output_15_137), .b(output_15_10), .y(output_14_137));
wire output_16_137, output_16_10, output_15_137;
mixer gate_output_15_137(.a(output_16_137), .b(output_16_10), .y(output_15_137));
wire output_1_138, output_1_11, output_0_138;
mixer gate_output_0_138(.a(output_1_138), .b(output_1_11), .y(output_0_138));
wire output_2_138, output_2_11, output_1_138;
mixer gate_output_1_138(.a(output_2_138), .b(output_2_11), .y(output_1_138));
wire output_3_138, output_3_11, output_2_138;
mixer gate_output_2_138(.a(output_3_138), .b(output_3_11), .y(output_2_138));
wire output_4_138, output_4_11, output_3_138;
mixer gate_output_3_138(.a(output_4_138), .b(output_4_11), .y(output_3_138));
wire output_5_138, output_5_11, output_4_138;
mixer gate_output_4_138(.a(output_5_138), .b(output_5_11), .y(output_4_138));
wire output_6_138, output_6_11, output_5_138;
mixer gate_output_5_138(.a(output_6_138), .b(output_6_11), .y(output_5_138));
wire output_7_138, output_7_11, output_6_138;
mixer gate_output_6_138(.a(output_7_138), .b(output_7_11), .y(output_6_138));
wire output_8_138, output_8_11, output_7_138;
mixer gate_output_7_138(.a(output_8_138), .b(output_8_11), .y(output_7_138));
wire output_9_138, output_9_11, output_8_138;
mixer gate_output_8_138(.a(output_9_138), .b(output_9_11), .y(output_8_138));
wire output_10_138, output_10_11, output_9_138;
mixer gate_output_9_138(.a(output_10_138), .b(output_10_11), .y(output_9_138));
wire output_11_138, output_11_11, output_10_138;
mixer gate_output_10_138(.a(output_11_138), .b(output_11_11), .y(output_10_138));
wire output_12_138, output_12_11, output_11_138;
mixer gate_output_11_138(.a(output_12_138), .b(output_12_11), .y(output_11_138));
wire output_13_138, output_13_11, output_12_138;
mixer gate_output_12_138(.a(output_13_138), .b(output_13_11), .y(output_12_138));
wire output_14_138, output_14_11, output_13_138;
mixer gate_output_13_138(.a(output_14_138), .b(output_14_11), .y(output_13_138));
wire output_15_138, output_15_11, output_14_138;
mixer gate_output_14_138(.a(output_15_138), .b(output_15_11), .y(output_14_138));
wire output_16_138, output_16_11, output_15_138;
mixer gate_output_15_138(.a(output_16_138), .b(output_16_11), .y(output_15_138));
wire output_1_139, output_1_12, output_0_139;
mixer gate_output_0_139(.a(output_1_139), .b(output_1_12), .y(output_0_139));
wire output_2_139, output_2_12, output_1_139;
mixer gate_output_1_139(.a(output_2_139), .b(output_2_12), .y(output_1_139));
wire output_3_139, output_3_12, output_2_139;
mixer gate_output_2_139(.a(output_3_139), .b(output_3_12), .y(output_2_139));
wire output_4_139, output_4_12, output_3_139;
mixer gate_output_3_139(.a(output_4_139), .b(output_4_12), .y(output_3_139));
wire output_5_139, output_5_12, output_4_139;
mixer gate_output_4_139(.a(output_5_139), .b(output_5_12), .y(output_4_139));
wire output_6_139, output_6_12, output_5_139;
mixer gate_output_5_139(.a(output_6_139), .b(output_6_12), .y(output_5_139));
wire output_7_139, output_7_12, output_6_139;
mixer gate_output_6_139(.a(output_7_139), .b(output_7_12), .y(output_6_139));
wire output_8_139, output_8_12, output_7_139;
mixer gate_output_7_139(.a(output_8_139), .b(output_8_12), .y(output_7_139));
wire output_9_139, output_9_12, output_8_139;
mixer gate_output_8_139(.a(output_9_139), .b(output_9_12), .y(output_8_139));
wire output_10_139, output_10_12, output_9_139;
mixer gate_output_9_139(.a(output_10_139), .b(output_10_12), .y(output_9_139));
wire output_11_139, output_11_12, output_10_139;
mixer gate_output_10_139(.a(output_11_139), .b(output_11_12), .y(output_10_139));
wire output_12_139, output_12_12, output_11_139;
mixer gate_output_11_139(.a(output_12_139), .b(output_12_12), .y(output_11_139));
wire output_13_139, output_13_12, output_12_139;
mixer gate_output_12_139(.a(output_13_139), .b(output_13_12), .y(output_12_139));
wire output_14_139, output_14_12, output_13_139;
mixer gate_output_13_139(.a(output_14_139), .b(output_14_12), .y(output_13_139));
wire output_15_139, output_15_12, output_14_139;
mixer gate_output_14_139(.a(output_15_139), .b(output_15_12), .y(output_14_139));
wire output_16_139, output_16_12, output_15_139;
mixer gate_output_15_139(.a(output_16_139), .b(output_16_12), .y(output_15_139));
wire output_1_140, output_1_13, output_0_140;
mixer gate_output_0_140(.a(output_1_140), .b(output_1_13), .y(output_0_140));
wire output_2_140, output_2_13, output_1_140;
mixer gate_output_1_140(.a(output_2_140), .b(output_2_13), .y(output_1_140));
wire output_3_140, output_3_13, output_2_140;
mixer gate_output_2_140(.a(output_3_140), .b(output_3_13), .y(output_2_140));
wire output_4_140, output_4_13, output_3_140;
mixer gate_output_3_140(.a(output_4_140), .b(output_4_13), .y(output_3_140));
wire output_5_140, output_5_13, output_4_140;
mixer gate_output_4_140(.a(output_5_140), .b(output_5_13), .y(output_4_140));
wire output_6_140, output_6_13, output_5_140;
mixer gate_output_5_140(.a(output_6_140), .b(output_6_13), .y(output_5_140));
wire output_7_140, output_7_13, output_6_140;
mixer gate_output_6_140(.a(output_7_140), .b(output_7_13), .y(output_6_140));
wire output_8_140, output_8_13, output_7_140;
mixer gate_output_7_140(.a(output_8_140), .b(output_8_13), .y(output_7_140));
wire output_9_140, output_9_13, output_8_140;
mixer gate_output_8_140(.a(output_9_140), .b(output_9_13), .y(output_8_140));
wire output_10_140, output_10_13, output_9_140;
mixer gate_output_9_140(.a(output_10_140), .b(output_10_13), .y(output_9_140));
wire output_11_140, output_11_13, output_10_140;
mixer gate_output_10_140(.a(output_11_140), .b(output_11_13), .y(output_10_140));
wire output_12_140, output_12_13, output_11_140;
mixer gate_output_11_140(.a(output_12_140), .b(output_12_13), .y(output_11_140));
wire output_13_140, output_13_13, output_12_140;
mixer gate_output_12_140(.a(output_13_140), .b(output_13_13), .y(output_12_140));
wire output_14_140, output_14_13, output_13_140;
mixer gate_output_13_140(.a(output_14_140), .b(output_14_13), .y(output_13_140));
wire output_15_140, output_15_13, output_14_140;
mixer gate_output_14_140(.a(output_15_140), .b(output_15_13), .y(output_14_140));
wire output_16_140, output_16_13, output_15_140;
mixer gate_output_15_140(.a(output_16_140), .b(output_16_13), .y(output_15_140));
wire output_1_141, output_1_14, output_0_141;
mixer gate_output_0_141(.a(output_1_141), .b(output_1_14), .y(output_0_141));
wire output_2_141, output_2_14, output_1_141;
mixer gate_output_1_141(.a(output_2_141), .b(output_2_14), .y(output_1_141));
wire output_3_141, output_3_14, output_2_141;
mixer gate_output_2_141(.a(output_3_141), .b(output_3_14), .y(output_2_141));
wire output_4_141, output_4_14, output_3_141;
mixer gate_output_3_141(.a(output_4_141), .b(output_4_14), .y(output_3_141));
wire output_5_141, output_5_14, output_4_141;
mixer gate_output_4_141(.a(output_5_141), .b(output_5_14), .y(output_4_141));
wire output_6_141, output_6_14, output_5_141;
mixer gate_output_5_141(.a(output_6_141), .b(output_6_14), .y(output_5_141));
wire output_7_141, output_7_14, output_6_141;
mixer gate_output_6_141(.a(output_7_141), .b(output_7_14), .y(output_6_141));
wire output_8_141, output_8_14, output_7_141;
mixer gate_output_7_141(.a(output_8_141), .b(output_8_14), .y(output_7_141));
wire output_9_141, output_9_14, output_8_141;
mixer gate_output_8_141(.a(output_9_141), .b(output_9_14), .y(output_8_141));
wire output_10_141, output_10_14, output_9_141;
mixer gate_output_9_141(.a(output_10_141), .b(output_10_14), .y(output_9_141));
wire output_11_141, output_11_14, output_10_141;
mixer gate_output_10_141(.a(output_11_141), .b(output_11_14), .y(output_10_141));
wire output_12_141, output_12_14, output_11_141;
mixer gate_output_11_141(.a(output_12_141), .b(output_12_14), .y(output_11_141));
wire output_13_141, output_13_14, output_12_141;
mixer gate_output_12_141(.a(output_13_141), .b(output_13_14), .y(output_12_141));
wire output_14_141, output_14_14, output_13_141;
mixer gate_output_13_141(.a(output_14_141), .b(output_14_14), .y(output_13_141));
wire output_15_141, output_15_14, output_14_141;
mixer gate_output_14_141(.a(output_15_141), .b(output_15_14), .y(output_14_141));
wire output_16_141, output_16_14, output_15_141;
mixer gate_output_15_141(.a(output_16_141), .b(output_16_14), .y(output_15_141));
wire output_1_142, output_1_15, output_0_142;
mixer gate_output_0_142(.a(output_1_142), .b(output_1_15), .y(output_0_142));
wire output_2_142, output_2_15, output_1_142;
mixer gate_output_1_142(.a(output_2_142), .b(output_2_15), .y(output_1_142));
wire output_3_142, output_3_15, output_2_142;
mixer gate_output_2_142(.a(output_3_142), .b(output_3_15), .y(output_2_142));
wire output_4_142, output_4_15, output_3_142;
mixer gate_output_3_142(.a(output_4_142), .b(output_4_15), .y(output_3_142));
wire output_5_142, output_5_15, output_4_142;
mixer gate_output_4_142(.a(output_5_142), .b(output_5_15), .y(output_4_142));
wire output_6_142, output_6_15, output_5_142;
mixer gate_output_5_142(.a(output_6_142), .b(output_6_15), .y(output_5_142));
wire output_7_142, output_7_15, output_6_142;
mixer gate_output_6_142(.a(output_7_142), .b(output_7_15), .y(output_6_142));
wire output_8_142, output_8_15, output_7_142;
mixer gate_output_7_142(.a(output_8_142), .b(output_8_15), .y(output_7_142));
wire output_9_142, output_9_15, output_8_142;
mixer gate_output_8_142(.a(output_9_142), .b(output_9_15), .y(output_8_142));
wire output_10_142, output_10_15, output_9_142;
mixer gate_output_9_142(.a(output_10_142), .b(output_10_15), .y(output_9_142));
wire output_11_142, output_11_15, output_10_142;
mixer gate_output_10_142(.a(output_11_142), .b(output_11_15), .y(output_10_142));
wire output_12_142, output_12_15, output_11_142;
mixer gate_output_11_142(.a(output_12_142), .b(output_12_15), .y(output_11_142));
wire output_13_142, output_13_15, output_12_142;
mixer gate_output_12_142(.a(output_13_142), .b(output_13_15), .y(output_12_142));
wire output_14_142, output_14_15, output_13_142;
mixer gate_output_13_142(.a(output_14_142), .b(output_14_15), .y(output_13_142));
wire output_15_142, output_15_15, output_14_142;
mixer gate_output_14_142(.a(output_15_142), .b(output_15_15), .y(output_14_142));
wire output_16_142, output_16_15, output_15_142;
mixer gate_output_15_142(.a(output_16_142), .b(output_16_15), .y(output_15_142));
wire output_1_143, output_1_0, output_0_143;
mixer gate_output_0_143(.a(output_1_143), .b(output_1_0), .y(output_0_143));
wire output_2_143, output_2_0, output_1_143;
mixer gate_output_1_143(.a(output_2_143), .b(output_2_0), .y(output_1_143));
wire output_3_143, output_3_0, output_2_143;
mixer gate_output_2_143(.a(output_3_143), .b(output_3_0), .y(output_2_143));
wire output_4_143, output_4_0, output_3_143;
mixer gate_output_3_143(.a(output_4_143), .b(output_4_0), .y(output_3_143));
wire output_5_143, output_5_0, output_4_143;
mixer gate_output_4_143(.a(output_5_143), .b(output_5_0), .y(output_4_143));
wire output_6_143, output_6_0, output_5_143;
mixer gate_output_5_143(.a(output_6_143), .b(output_6_0), .y(output_5_143));
wire output_7_143, output_7_0, output_6_143;
mixer gate_output_6_143(.a(output_7_143), .b(output_7_0), .y(output_6_143));
wire output_8_143, output_8_0, output_7_143;
mixer gate_output_7_143(.a(output_8_143), .b(output_8_0), .y(output_7_143));
wire output_9_143, output_9_0, output_8_143;
mixer gate_output_8_143(.a(output_9_143), .b(output_9_0), .y(output_8_143));
wire output_10_143, output_10_0, output_9_143;
mixer gate_output_9_143(.a(output_10_143), .b(output_10_0), .y(output_9_143));
wire output_11_143, output_11_0, output_10_143;
mixer gate_output_10_143(.a(output_11_143), .b(output_11_0), .y(output_10_143));
wire output_12_143, output_12_0, output_11_143;
mixer gate_output_11_143(.a(output_12_143), .b(output_12_0), .y(output_11_143));
wire output_13_143, output_13_0, output_12_143;
mixer gate_output_12_143(.a(output_13_143), .b(output_13_0), .y(output_12_143));
wire output_14_143, output_14_0, output_13_143;
mixer gate_output_13_143(.a(output_14_143), .b(output_14_0), .y(output_13_143));
wire output_15_143, output_15_0, output_14_143;
mixer gate_output_14_143(.a(output_15_143), .b(output_15_0), .y(output_14_143));
wire output_16_143, output_16_0, output_15_143;
mixer gate_output_15_143(.a(output_16_143), .b(output_16_0), .y(output_15_143));
wire output_1_144, output_1_1, output_0_144;
mixer gate_output_0_144(.a(output_1_144), .b(output_1_1), .y(output_0_144));
wire output_2_144, output_2_1, output_1_144;
mixer gate_output_1_144(.a(output_2_144), .b(output_2_1), .y(output_1_144));
wire output_3_144, output_3_1, output_2_144;
mixer gate_output_2_144(.a(output_3_144), .b(output_3_1), .y(output_2_144));
wire output_4_144, output_4_1, output_3_144;
mixer gate_output_3_144(.a(output_4_144), .b(output_4_1), .y(output_3_144));
wire output_5_144, output_5_1, output_4_144;
mixer gate_output_4_144(.a(output_5_144), .b(output_5_1), .y(output_4_144));
wire output_6_144, output_6_1, output_5_144;
mixer gate_output_5_144(.a(output_6_144), .b(output_6_1), .y(output_5_144));
wire output_7_144, output_7_1, output_6_144;
mixer gate_output_6_144(.a(output_7_144), .b(output_7_1), .y(output_6_144));
wire output_8_144, output_8_1, output_7_144;
mixer gate_output_7_144(.a(output_8_144), .b(output_8_1), .y(output_7_144));
wire output_9_144, output_9_1, output_8_144;
mixer gate_output_8_144(.a(output_9_144), .b(output_9_1), .y(output_8_144));
wire output_10_144, output_10_1, output_9_144;
mixer gate_output_9_144(.a(output_10_144), .b(output_10_1), .y(output_9_144));
wire output_11_144, output_11_1, output_10_144;
mixer gate_output_10_144(.a(output_11_144), .b(output_11_1), .y(output_10_144));
wire output_12_144, output_12_1, output_11_144;
mixer gate_output_11_144(.a(output_12_144), .b(output_12_1), .y(output_11_144));
wire output_13_144, output_13_1, output_12_144;
mixer gate_output_12_144(.a(output_13_144), .b(output_13_1), .y(output_12_144));
wire output_14_144, output_14_1, output_13_144;
mixer gate_output_13_144(.a(output_14_144), .b(output_14_1), .y(output_13_144));
wire output_15_144, output_15_1, output_14_144;
mixer gate_output_14_144(.a(output_15_144), .b(output_15_1), .y(output_14_144));
wire output_16_144, output_16_1, output_15_144;
mixer gate_output_15_144(.a(output_16_144), .b(output_16_1), .y(output_15_144));
wire output_1_145, output_1_2, output_0_145;
mixer gate_output_0_145(.a(output_1_145), .b(output_1_2), .y(output_0_145));
wire output_2_145, output_2_2, output_1_145;
mixer gate_output_1_145(.a(output_2_145), .b(output_2_2), .y(output_1_145));
wire output_3_145, output_3_2, output_2_145;
mixer gate_output_2_145(.a(output_3_145), .b(output_3_2), .y(output_2_145));
wire output_4_145, output_4_2, output_3_145;
mixer gate_output_3_145(.a(output_4_145), .b(output_4_2), .y(output_3_145));
wire output_5_145, output_5_2, output_4_145;
mixer gate_output_4_145(.a(output_5_145), .b(output_5_2), .y(output_4_145));
wire output_6_145, output_6_2, output_5_145;
mixer gate_output_5_145(.a(output_6_145), .b(output_6_2), .y(output_5_145));
wire output_7_145, output_7_2, output_6_145;
mixer gate_output_6_145(.a(output_7_145), .b(output_7_2), .y(output_6_145));
wire output_8_145, output_8_2, output_7_145;
mixer gate_output_7_145(.a(output_8_145), .b(output_8_2), .y(output_7_145));
wire output_9_145, output_9_2, output_8_145;
mixer gate_output_8_145(.a(output_9_145), .b(output_9_2), .y(output_8_145));
wire output_10_145, output_10_2, output_9_145;
mixer gate_output_9_145(.a(output_10_145), .b(output_10_2), .y(output_9_145));
wire output_11_145, output_11_2, output_10_145;
mixer gate_output_10_145(.a(output_11_145), .b(output_11_2), .y(output_10_145));
wire output_12_145, output_12_2, output_11_145;
mixer gate_output_11_145(.a(output_12_145), .b(output_12_2), .y(output_11_145));
wire output_13_145, output_13_2, output_12_145;
mixer gate_output_12_145(.a(output_13_145), .b(output_13_2), .y(output_12_145));
wire output_14_145, output_14_2, output_13_145;
mixer gate_output_13_145(.a(output_14_145), .b(output_14_2), .y(output_13_145));
wire output_15_145, output_15_2, output_14_145;
mixer gate_output_14_145(.a(output_15_145), .b(output_15_2), .y(output_14_145));
wire output_16_145, output_16_2, output_15_145;
mixer gate_output_15_145(.a(output_16_145), .b(output_16_2), .y(output_15_145));
wire output_1_146, output_1_3, output_0_146;
mixer gate_output_0_146(.a(output_1_146), .b(output_1_3), .y(output_0_146));
wire output_2_146, output_2_3, output_1_146;
mixer gate_output_1_146(.a(output_2_146), .b(output_2_3), .y(output_1_146));
wire output_3_146, output_3_3, output_2_146;
mixer gate_output_2_146(.a(output_3_146), .b(output_3_3), .y(output_2_146));
wire output_4_146, output_4_3, output_3_146;
mixer gate_output_3_146(.a(output_4_146), .b(output_4_3), .y(output_3_146));
wire output_5_146, output_5_3, output_4_146;
mixer gate_output_4_146(.a(output_5_146), .b(output_5_3), .y(output_4_146));
wire output_6_146, output_6_3, output_5_146;
mixer gate_output_5_146(.a(output_6_146), .b(output_6_3), .y(output_5_146));
wire output_7_146, output_7_3, output_6_146;
mixer gate_output_6_146(.a(output_7_146), .b(output_7_3), .y(output_6_146));
wire output_8_146, output_8_3, output_7_146;
mixer gate_output_7_146(.a(output_8_146), .b(output_8_3), .y(output_7_146));
wire output_9_146, output_9_3, output_8_146;
mixer gate_output_8_146(.a(output_9_146), .b(output_9_3), .y(output_8_146));
wire output_10_146, output_10_3, output_9_146;
mixer gate_output_9_146(.a(output_10_146), .b(output_10_3), .y(output_9_146));
wire output_11_146, output_11_3, output_10_146;
mixer gate_output_10_146(.a(output_11_146), .b(output_11_3), .y(output_10_146));
wire output_12_146, output_12_3, output_11_146;
mixer gate_output_11_146(.a(output_12_146), .b(output_12_3), .y(output_11_146));
wire output_13_146, output_13_3, output_12_146;
mixer gate_output_12_146(.a(output_13_146), .b(output_13_3), .y(output_12_146));
wire output_14_146, output_14_3, output_13_146;
mixer gate_output_13_146(.a(output_14_146), .b(output_14_3), .y(output_13_146));
wire output_15_146, output_15_3, output_14_146;
mixer gate_output_14_146(.a(output_15_146), .b(output_15_3), .y(output_14_146));
wire output_16_146, output_16_3, output_15_146;
mixer gate_output_15_146(.a(output_16_146), .b(output_16_3), .y(output_15_146));
wire output_1_147, output_1_4, output_0_147;
mixer gate_output_0_147(.a(output_1_147), .b(output_1_4), .y(output_0_147));
wire output_2_147, output_2_4, output_1_147;
mixer gate_output_1_147(.a(output_2_147), .b(output_2_4), .y(output_1_147));
wire output_3_147, output_3_4, output_2_147;
mixer gate_output_2_147(.a(output_3_147), .b(output_3_4), .y(output_2_147));
wire output_4_147, output_4_4, output_3_147;
mixer gate_output_3_147(.a(output_4_147), .b(output_4_4), .y(output_3_147));
wire output_5_147, output_5_4, output_4_147;
mixer gate_output_4_147(.a(output_5_147), .b(output_5_4), .y(output_4_147));
wire output_6_147, output_6_4, output_5_147;
mixer gate_output_5_147(.a(output_6_147), .b(output_6_4), .y(output_5_147));
wire output_7_147, output_7_4, output_6_147;
mixer gate_output_6_147(.a(output_7_147), .b(output_7_4), .y(output_6_147));
wire output_8_147, output_8_4, output_7_147;
mixer gate_output_7_147(.a(output_8_147), .b(output_8_4), .y(output_7_147));
wire output_9_147, output_9_4, output_8_147;
mixer gate_output_8_147(.a(output_9_147), .b(output_9_4), .y(output_8_147));
wire output_10_147, output_10_4, output_9_147;
mixer gate_output_9_147(.a(output_10_147), .b(output_10_4), .y(output_9_147));
wire output_11_147, output_11_4, output_10_147;
mixer gate_output_10_147(.a(output_11_147), .b(output_11_4), .y(output_10_147));
wire output_12_147, output_12_4, output_11_147;
mixer gate_output_11_147(.a(output_12_147), .b(output_12_4), .y(output_11_147));
wire output_13_147, output_13_4, output_12_147;
mixer gate_output_12_147(.a(output_13_147), .b(output_13_4), .y(output_12_147));
wire output_14_147, output_14_4, output_13_147;
mixer gate_output_13_147(.a(output_14_147), .b(output_14_4), .y(output_13_147));
wire output_15_147, output_15_4, output_14_147;
mixer gate_output_14_147(.a(output_15_147), .b(output_15_4), .y(output_14_147));
wire output_16_147, output_16_4, output_15_147;
mixer gate_output_15_147(.a(output_16_147), .b(output_16_4), .y(output_15_147));
wire output_1_148, output_1_5, output_0_148;
mixer gate_output_0_148(.a(output_1_148), .b(output_1_5), .y(output_0_148));
wire output_2_148, output_2_5, output_1_148;
mixer gate_output_1_148(.a(output_2_148), .b(output_2_5), .y(output_1_148));
wire output_3_148, output_3_5, output_2_148;
mixer gate_output_2_148(.a(output_3_148), .b(output_3_5), .y(output_2_148));
wire output_4_148, output_4_5, output_3_148;
mixer gate_output_3_148(.a(output_4_148), .b(output_4_5), .y(output_3_148));
wire output_5_148, output_5_5, output_4_148;
mixer gate_output_4_148(.a(output_5_148), .b(output_5_5), .y(output_4_148));
wire output_6_148, output_6_5, output_5_148;
mixer gate_output_5_148(.a(output_6_148), .b(output_6_5), .y(output_5_148));
wire output_7_148, output_7_5, output_6_148;
mixer gate_output_6_148(.a(output_7_148), .b(output_7_5), .y(output_6_148));
wire output_8_148, output_8_5, output_7_148;
mixer gate_output_7_148(.a(output_8_148), .b(output_8_5), .y(output_7_148));
wire output_9_148, output_9_5, output_8_148;
mixer gate_output_8_148(.a(output_9_148), .b(output_9_5), .y(output_8_148));
wire output_10_148, output_10_5, output_9_148;
mixer gate_output_9_148(.a(output_10_148), .b(output_10_5), .y(output_9_148));
wire output_11_148, output_11_5, output_10_148;
mixer gate_output_10_148(.a(output_11_148), .b(output_11_5), .y(output_10_148));
wire output_12_148, output_12_5, output_11_148;
mixer gate_output_11_148(.a(output_12_148), .b(output_12_5), .y(output_11_148));
wire output_13_148, output_13_5, output_12_148;
mixer gate_output_12_148(.a(output_13_148), .b(output_13_5), .y(output_12_148));
wire output_14_148, output_14_5, output_13_148;
mixer gate_output_13_148(.a(output_14_148), .b(output_14_5), .y(output_13_148));
wire output_15_148, output_15_5, output_14_148;
mixer gate_output_14_148(.a(output_15_148), .b(output_15_5), .y(output_14_148));
wire output_16_148, output_16_5, output_15_148;
mixer gate_output_15_148(.a(output_16_148), .b(output_16_5), .y(output_15_148));
wire output_1_149, output_1_6, output_0_149;
mixer gate_output_0_149(.a(output_1_149), .b(output_1_6), .y(output_0_149));
wire output_2_149, output_2_6, output_1_149;
mixer gate_output_1_149(.a(output_2_149), .b(output_2_6), .y(output_1_149));
wire output_3_149, output_3_6, output_2_149;
mixer gate_output_2_149(.a(output_3_149), .b(output_3_6), .y(output_2_149));
wire output_4_149, output_4_6, output_3_149;
mixer gate_output_3_149(.a(output_4_149), .b(output_4_6), .y(output_3_149));
wire output_5_149, output_5_6, output_4_149;
mixer gate_output_4_149(.a(output_5_149), .b(output_5_6), .y(output_4_149));
wire output_6_149, output_6_6, output_5_149;
mixer gate_output_5_149(.a(output_6_149), .b(output_6_6), .y(output_5_149));
wire output_7_149, output_7_6, output_6_149;
mixer gate_output_6_149(.a(output_7_149), .b(output_7_6), .y(output_6_149));
wire output_8_149, output_8_6, output_7_149;
mixer gate_output_7_149(.a(output_8_149), .b(output_8_6), .y(output_7_149));
wire output_9_149, output_9_6, output_8_149;
mixer gate_output_8_149(.a(output_9_149), .b(output_9_6), .y(output_8_149));
wire output_10_149, output_10_6, output_9_149;
mixer gate_output_9_149(.a(output_10_149), .b(output_10_6), .y(output_9_149));
wire output_11_149, output_11_6, output_10_149;
mixer gate_output_10_149(.a(output_11_149), .b(output_11_6), .y(output_10_149));
wire output_12_149, output_12_6, output_11_149;
mixer gate_output_11_149(.a(output_12_149), .b(output_12_6), .y(output_11_149));
wire output_13_149, output_13_6, output_12_149;
mixer gate_output_12_149(.a(output_13_149), .b(output_13_6), .y(output_12_149));
wire output_14_149, output_14_6, output_13_149;
mixer gate_output_13_149(.a(output_14_149), .b(output_14_6), .y(output_13_149));
wire output_15_149, output_15_6, output_14_149;
mixer gate_output_14_149(.a(output_15_149), .b(output_15_6), .y(output_14_149));
wire output_16_149, output_16_6, output_15_149;
mixer gate_output_15_149(.a(output_16_149), .b(output_16_6), .y(output_15_149));
wire output_1_150, output_1_7, output_0_150;
mixer gate_output_0_150(.a(output_1_150), .b(output_1_7), .y(output_0_150));
wire output_2_150, output_2_7, output_1_150;
mixer gate_output_1_150(.a(output_2_150), .b(output_2_7), .y(output_1_150));
wire output_3_150, output_3_7, output_2_150;
mixer gate_output_2_150(.a(output_3_150), .b(output_3_7), .y(output_2_150));
wire output_4_150, output_4_7, output_3_150;
mixer gate_output_3_150(.a(output_4_150), .b(output_4_7), .y(output_3_150));
wire output_5_150, output_5_7, output_4_150;
mixer gate_output_4_150(.a(output_5_150), .b(output_5_7), .y(output_4_150));
wire output_6_150, output_6_7, output_5_150;
mixer gate_output_5_150(.a(output_6_150), .b(output_6_7), .y(output_5_150));
wire output_7_150, output_7_7, output_6_150;
mixer gate_output_6_150(.a(output_7_150), .b(output_7_7), .y(output_6_150));
wire output_8_150, output_8_7, output_7_150;
mixer gate_output_7_150(.a(output_8_150), .b(output_8_7), .y(output_7_150));
wire output_9_150, output_9_7, output_8_150;
mixer gate_output_8_150(.a(output_9_150), .b(output_9_7), .y(output_8_150));
wire output_10_150, output_10_7, output_9_150;
mixer gate_output_9_150(.a(output_10_150), .b(output_10_7), .y(output_9_150));
wire output_11_150, output_11_7, output_10_150;
mixer gate_output_10_150(.a(output_11_150), .b(output_11_7), .y(output_10_150));
wire output_12_150, output_12_7, output_11_150;
mixer gate_output_11_150(.a(output_12_150), .b(output_12_7), .y(output_11_150));
wire output_13_150, output_13_7, output_12_150;
mixer gate_output_12_150(.a(output_13_150), .b(output_13_7), .y(output_12_150));
wire output_14_150, output_14_7, output_13_150;
mixer gate_output_13_150(.a(output_14_150), .b(output_14_7), .y(output_13_150));
wire output_15_150, output_15_7, output_14_150;
mixer gate_output_14_150(.a(output_15_150), .b(output_15_7), .y(output_14_150));
wire output_16_150, output_16_7, output_15_150;
mixer gate_output_15_150(.a(output_16_150), .b(output_16_7), .y(output_15_150));
wire output_1_151, output_1_8, output_0_151;
mixer gate_output_0_151(.a(output_1_151), .b(output_1_8), .y(output_0_151));
wire output_2_151, output_2_8, output_1_151;
mixer gate_output_1_151(.a(output_2_151), .b(output_2_8), .y(output_1_151));
wire output_3_151, output_3_8, output_2_151;
mixer gate_output_2_151(.a(output_3_151), .b(output_3_8), .y(output_2_151));
wire output_4_151, output_4_8, output_3_151;
mixer gate_output_3_151(.a(output_4_151), .b(output_4_8), .y(output_3_151));
wire output_5_151, output_5_8, output_4_151;
mixer gate_output_4_151(.a(output_5_151), .b(output_5_8), .y(output_4_151));
wire output_6_151, output_6_8, output_5_151;
mixer gate_output_5_151(.a(output_6_151), .b(output_6_8), .y(output_5_151));
wire output_7_151, output_7_8, output_6_151;
mixer gate_output_6_151(.a(output_7_151), .b(output_7_8), .y(output_6_151));
wire output_8_151, output_8_8, output_7_151;
mixer gate_output_7_151(.a(output_8_151), .b(output_8_8), .y(output_7_151));
wire output_9_151, output_9_8, output_8_151;
mixer gate_output_8_151(.a(output_9_151), .b(output_9_8), .y(output_8_151));
wire output_10_151, output_10_8, output_9_151;
mixer gate_output_9_151(.a(output_10_151), .b(output_10_8), .y(output_9_151));
wire output_11_151, output_11_8, output_10_151;
mixer gate_output_10_151(.a(output_11_151), .b(output_11_8), .y(output_10_151));
wire output_12_151, output_12_8, output_11_151;
mixer gate_output_11_151(.a(output_12_151), .b(output_12_8), .y(output_11_151));
wire output_13_151, output_13_8, output_12_151;
mixer gate_output_12_151(.a(output_13_151), .b(output_13_8), .y(output_12_151));
wire output_14_151, output_14_8, output_13_151;
mixer gate_output_13_151(.a(output_14_151), .b(output_14_8), .y(output_13_151));
wire output_15_151, output_15_8, output_14_151;
mixer gate_output_14_151(.a(output_15_151), .b(output_15_8), .y(output_14_151));
wire output_16_151, output_16_8, output_15_151;
mixer gate_output_15_151(.a(output_16_151), .b(output_16_8), .y(output_15_151));
wire output_1_152, output_1_9, output_0_152;
mixer gate_output_0_152(.a(output_1_152), .b(output_1_9), .y(output_0_152));
wire output_2_152, output_2_9, output_1_152;
mixer gate_output_1_152(.a(output_2_152), .b(output_2_9), .y(output_1_152));
wire output_3_152, output_3_9, output_2_152;
mixer gate_output_2_152(.a(output_3_152), .b(output_3_9), .y(output_2_152));
wire output_4_152, output_4_9, output_3_152;
mixer gate_output_3_152(.a(output_4_152), .b(output_4_9), .y(output_3_152));
wire output_5_152, output_5_9, output_4_152;
mixer gate_output_4_152(.a(output_5_152), .b(output_5_9), .y(output_4_152));
wire output_6_152, output_6_9, output_5_152;
mixer gate_output_5_152(.a(output_6_152), .b(output_6_9), .y(output_5_152));
wire output_7_152, output_7_9, output_6_152;
mixer gate_output_6_152(.a(output_7_152), .b(output_7_9), .y(output_6_152));
wire output_8_152, output_8_9, output_7_152;
mixer gate_output_7_152(.a(output_8_152), .b(output_8_9), .y(output_7_152));
wire output_9_152, output_9_9, output_8_152;
mixer gate_output_8_152(.a(output_9_152), .b(output_9_9), .y(output_8_152));
wire output_10_152, output_10_9, output_9_152;
mixer gate_output_9_152(.a(output_10_152), .b(output_10_9), .y(output_9_152));
wire output_11_152, output_11_9, output_10_152;
mixer gate_output_10_152(.a(output_11_152), .b(output_11_9), .y(output_10_152));
wire output_12_152, output_12_9, output_11_152;
mixer gate_output_11_152(.a(output_12_152), .b(output_12_9), .y(output_11_152));
wire output_13_152, output_13_9, output_12_152;
mixer gate_output_12_152(.a(output_13_152), .b(output_13_9), .y(output_12_152));
wire output_14_152, output_14_9, output_13_152;
mixer gate_output_13_152(.a(output_14_152), .b(output_14_9), .y(output_13_152));
wire output_15_152, output_15_9, output_14_152;
mixer gate_output_14_152(.a(output_15_152), .b(output_15_9), .y(output_14_152));
wire output_16_152, output_16_9, output_15_152;
mixer gate_output_15_152(.a(output_16_152), .b(output_16_9), .y(output_15_152));
wire output_1_153, output_1_10, output_0_153;
mixer gate_output_0_153(.a(output_1_153), .b(output_1_10), .y(output_0_153));
wire output_2_153, output_2_10, output_1_153;
mixer gate_output_1_153(.a(output_2_153), .b(output_2_10), .y(output_1_153));
wire output_3_153, output_3_10, output_2_153;
mixer gate_output_2_153(.a(output_3_153), .b(output_3_10), .y(output_2_153));
wire output_4_153, output_4_10, output_3_153;
mixer gate_output_3_153(.a(output_4_153), .b(output_4_10), .y(output_3_153));
wire output_5_153, output_5_10, output_4_153;
mixer gate_output_4_153(.a(output_5_153), .b(output_5_10), .y(output_4_153));
wire output_6_153, output_6_10, output_5_153;
mixer gate_output_5_153(.a(output_6_153), .b(output_6_10), .y(output_5_153));
wire output_7_153, output_7_10, output_6_153;
mixer gate_output_6_153(.a(output_7_153), .b(output_7_10), .y(output_6_153));
wire output_8_153, output_8_10, output_7_153;
mixer gate_output_7_153(.a(output_8_153), .b(output_8_10), .y(output_7_153));
wire output_9_153, output_9_10, output_8_153;
mixer gate_output_8_153(.a(output_9_153), .b(output_9_10), .y(output_8_153));
wire output_10_153, output_10_10, output_9_153;
mixer gate_output_9_153(.a(output_10_153), .b(output_10_10), .y(output_9_153));
wire output_11_153, output_11_10, output_10_153;
mixer gate_output_10_153(.a(output_11_153), .b(output_11_10), .y(output_10_153));
wire output_12_153, output_12_10, output_11_153;
mixer gate_output_11_153(.a(output_12_153), .b(output_12_10), .y(output_11_153));
wire output_13_153, output_13_10, output_12_153;
mixer gate_output_12_153(.a(output_13_153), .b(output_13_10), .y(output_12_153));
wire output_14_153, output_14_10, output_13_153;
mixer gate_output_13_153(.a(output_14_153), .b(output_14_10), .y(output_13_153));
wire output_15_153, output_15_10, output_14_153;
mixer gate_output_14_153(.a(output_15_153), .b(output_15_10), .y(output_14_153));
wire output_16_153, output_16_10, output_15_153;
mixer gate_output_15_153(.a(output_16_153), .b(output_16_10), .y(output_15_153));
wire output_1_154, output_1_11, output_0_154;
mixer gate_output_0_154(.a(output_1_154), .b(output_1_11), .y(output_0_154));
wire output_2_154, output_2_11, output_1_154;
mixer gate_output_1_154(.a(output_2_154), .b(output_2_11), .y(output_1_154));
wire output_3_154, output_3_11, output_2_154;
mixer gate_output_2_154(.a(output_3_154), .b(output_3_11), .y(output_2_154));
wire output_4_154, output_4_11, output_3_154;
mixer gate_output_3_154(.a(output_4_154), .b(output_4_11), .y(output_3_154));
wire output_5_154, output_5_11, output_4_154;
mixer gate_output_4_154(.a(output_5_154), .b(output_5_11), .y(output_4_154));
wire output_6_154, output_6_11, output_5_154;
mixer gate_output_5_154(.a(output_6_154), .b(output_6_11), .y(output_5_154));
wire output_7_154, output_7_11, output_6_154;
mixer gate_output_6_154(.a(output_7_154), .b(output_7_11), .y(output_6_154));
wire output_8_154, output_8_11, output_7_154;
mixer gate_output_7_154(.a(output_8_154), .b(output_8_11), .y(output_7_154));
wire output_9_154, output_9_11, output_8_154;
mixer gate_output_8_154(.a(output_9_154), .b(output_9_11), .y(output_8_154));
wire output_10_154, output_10_11, output_9_154;
mixer gate_output_9_154(.a(output_10_154), .b(output_10_11), .y(output_9_154));
wire output_11_154, output_11_11, output_10_154;
mixer gate_output_10_154(.a(output_11_154), .b(output_11_11), .y(output_10_154));
wire output_12_154, output_12_11, output_11_154;
mixer gate_output_11_154(.a(output_12_154), .b(output_12_11), .y(output_11_154));
wire output_13_154, output_13_11, output_12_154;
mixer gate_output_12_154(.a(output_13_154), .b(output_13_11), .y(output_12_154));
wire output_14_154, output_14_11, output_13_154;
mixer gate_output_13_154(.a(output_14_154), .b(output_14_11), .y(output_13_154));
wire output_15_154, output_15_11, output_14_154;
mixer gate_output_14_154(.a(output_15_154), .b(output_15_11), .y(output_14_154));
wire output_16_154, output_16_11, output_15_154;
mixer gate_output_15_154(.a(output_16_154), .b(output_16_11), .y(output_15_154));
wire output_1_155, output_1_12, output_0_155;
mixer gate_output_0_155(.a(output_1_155), .b(output_1_12), .y(output_0_155));
wire output_2_155, output_2_12, output_1_155;
mixer gate_output_1_155(.a(output_2_155), .b(output_2_12), .y(output_1_155));
wire output_3_155, output_3_12, output_2_155;
mixer gate_output_2_155(.a(output_3_155), .b(output_3_12), .y(output_2_155));
wire output_4_155, output_4_12, output_3_155;
mixer gate_output_3_155(.a(output_4_155), .b(output_4_12), .y(output_3_155));
wire output_5_155, output_5_12, output_4_155;
mixer gate_output_4_155(.a(output_5_155), .b(output_5_12), .y(output_4_155));
wire output_6_155, output_6_12, output_5_155;
mixer gate_output_5_155(.a(output_6_155), .b(output_6_12), .y(output_5_155));
wire output_7_155, output_7_12, output_6_155;
mixer gate_output_6_155(.a(output_7_155), .b(output_7_12), .y(output_6_155));
wire output_8_155, output_8_12, output_7_155;
mixer gate_output_7_155(.a(output_8_155), .b(output_8_12), .y(output_7_155));
wire output_9_155, output_9_12, output_8_155;
mixer gate_output_8_155(.a(output_9_155), .b(output_9_12), .y(output_8_155));
wire output_10_155, output_10_12, output_9_155;
mixer gate_output_9_155(.a(output_10_155), .b(output_10_12), .y(output_9_155));
wire output_11_155, output_11_12, output_10_155;
mixer gate_output_10_155(.a(output_11_155), .b(output_11_12), .y(output_10_155));
wire output_12_155, output_12_12, output_11_155;
mixer gate_output_11_155(.a(output_12_155), .b(output_12_12), .y(output_11_155));
wire output_13_155, output_13_12, output_12_155;
mixer gate_output_12_155(.a(output_13_155), .b(output_13_12), .y(output_12_155));
wire output_14_155, output_14_12, output_13_155;
mixer gate_output_13_155(.a(output_14_155), .b(output_14_12), .y(output_13_155));
wire output_15_155, output_15_12, output_14_155;
mixer gate_output_14_155(.a(output_15_155), .b(output_15_12), .y(output_14_155));
wire output_16_155, output_16_12, output_15_155;
mixer gate_output_15_155(.a(output_16_155), .b(output_16_12), .y(output_15_155));
wire output_1_156, output_1_13, output_0_156;
mixer gate_output_0_156(.a(output_1_156), .b(output_1_13), .y(output_0_156));
wire output_2_156, output_2_13, output_1_156;
mixer gate_output_1_156(.a(output_2_156), .b(output_2_13), .y(output_1_156));
wire output_3_156, output_3_13, output_2_156;
mixer gate_output_2_156(.a(output_3_156), .b(output_3_13), .y(output_2_156));
wire output_4_156, output_4_13, output_3_156;
mixer gate_output_3_156(.a(output_4_156), .b(output_4_13), .y(output_3_156));
wire output_5_156, output_5_13, output_4_156;
mixer gate_output_4_156(.a(output_5_156), .b(output_5_13), .y(output_4_156));
wire output_6_156, output_6_13, output_5_156;
mixer gate_output_5_156(.a(output_6_156), .b(output_6_13), .y(output_5_156));
wire output_7_156, output_7_13, output_6_156;
mixer gate_output_6_156(.a(output_7_156), .b(output_7_13), .y(output_6_156));
wire output_8_156, output_8_13, output_7_156;
mixer gate_output_7_156(.a(output_8_156), .b(output_8_13), .y(output_7_156));
wire output_9_156, output_9_13, output_8_156;
mixer gate_output_8_156(.a(output_9_156), .b(output_9_13), .y(output_8_156));
wire output_10_156, output_10_13, output_9_156;
mixer gate_output_9_156(.a(output_10_156), .b(output_10_13), .y(output_9_156));
wire output_11_156, output_11_13, output_10_156;
mixer gate_output_10_156(.a(output_11_156), .b(output_11_13), .y(output_10_156));
wire output_12_156, output_12_13, output_11_156;
mixer gate_output_11_156(.a(output_12_156), .b(output_12_13), .y(output_11_156));
wire output_13_156, output_13_13, output_12_156;
mixer gate_output_12_156(.a(output_13_156), .b(output_13_13), .y(output_12_156));
wire output_14_156, output_14_13, output_13_156;
mixer gate_output_13_156(.a(output_14_156), .b(output_14_13), .y(output_13_156));
wire output_15_156, output_15_13, output_14_156;
mixer gate_output_14_156(.a(output_15_156), .b(output_15_13), .y(output_14_156));
wire output_16_156, output_16_13, output_15_156;
mixer gate_output_15_156(.a(output_16_156), .b(output_16_13), .y(output_15_156));
wire output_1_157, output_1_14, output_0_157;
mixer gate_output_0_157(.a(output_1_157), .b(output_1_14), .y(output_0_157));
wire output_2_157, output_2_14, output_1_157;
mixer gate_output_1_157(.a(output_2_157), .b(output_2_14), .y(output_1_157));
wire output_3_157, output_3_14, output_2_157;
mixer gate_output_2_157(.a(output_3_157), .b(output_3_14), .y(output_2_157));
wire output_4_157, output_4_14, output_3_157;
mixer gate_output_3_157(.a(output_4_157), .b(output_4_14), .y(output_3_157));
wire output_5_157, output_5_14, output_4_157;
mixer gate_output_4_157(.a(output_5_157), .b(output_5_14), .y(output_4_157));
wire output_6_157, output_6_14, output_5_157;
mixer gate_output_5_157(.a(output_6_157), .b(output_6_14), .y(output_5_157));
wire output_7_157, output_7_14, output_6_157;
mixer gate_output_6_157(.a(output_7_157), .b(output_7_14), .y(output_6_157));
wire output_8_157, output_8_14, output_7_157;
mixer gate_output_7_157(.a(output_8_157), .b(output_8_14), .y(output_7_157));
wire output_9_157, output_9_14, output_8_157;
mixer gate_output_8_157(.a(output_9_157), .b(output_9_14), .y(output_8_157));
wire output_10_157, output_10_14, output_9_157;
mixer gate_output_9_157(.a(output_10_157), .b(output_10_14), .y(output_9_157));
wire output_11_157, output_11_14, output_10_157;
mixer gate_output_10_157(.a(output_11_157), .b(output_11_14), .y(output_10_157));
wire output_12_157, output_12_14, output_11_157;
mixer gate_output_11_157(.a(output_12_157), .b(output_12_14), .y(output_11_157));
wire output_13_157, output_13_14, output_12_157;
mixer gate_output_12_157(.a(output_13_157), .b(output_13_14), .y(output_12_157));
wire output_14_157, output_14_14, output_13_157;
mixer gate_output_13_157(.a(output_14_157), .b(output_14_14), .y(output_13_157));
wire output_15_157, output_15_14, output_14_157;
mixer gate_output_14_157(.a(output_15_157), .b(output_15_14), .y(output_14_157));
wire output_16_157, output_16_14, output_15_157;
mixer gate_output_15_157(.a(output_16_157), .b(output_16_14), .y(output_15_157));
wire output_1_158, output_1_15, output_0_158;
mixer gate_output_0_158(.a(output_1_158), .b(output_1_15), .y(output_0_158));
wire output_2_158, output_2_15, output_1_158;
mixer gate_output_1_158(.a(output_2_158), .b(output_2_15), .y(output_1_158));
wire output_3_158, output_3_15, output_2_158;
mixer gate_output_2_158(.a(output_3_158), .b(output_3_15), .y(output_2_158));
wire output_4_158, output_4_15, output_3_158;
mixer gate_output_3_158(.a(output_4_158), .b(output_4_15), .y(output_3_158));
wire output_5_158, output_5_15, output_4_158;
mixer gate_output_4_158(.a(output_5_158), .b(output_5_15), .y(output_4_158));
wire output_6_158, output_6_15, output_5_158;
mixer gate_output_5_158(.a(output_6_158), .b(output_6_15), .y(output_5_158));
wire output_7_158, output_7_15, output_6_158;
mixer gate_output_6_158(.a(output_7_158), .b(output_7_15), .y(output_6_158));
wire output_8_158, output_8_15, output_7_158;
mixer gate_output_7_158(.a(output_8_158), .b(output_8_15), .y(output_7_158));
wire output_9_158, output_9_15, output_8_158;
mixer gate_output_8_158(.a(output_9_158), .b(output_9_15), .y(output_8_158));
wire output_10_158, output_10_15, output_9_158;
mixer gate_output_9_158(.a(output_10_158), .b(output_10_15), .y(output_9_158));
wire output_11_158, output_11_15, output_10_158;
mixer gate_output_10_158(.a(output_11_158), .b(output_11_15), .y(output_10_158));
wire output_12_158, output_12_15, output_11_158;
mixer gate_output_11_158(.a(output_12_158), .b(output_12_15), .y(output_11_158));
wire output_13_158, output_13_15, output_12_158;
mixer gate_output_12_158(.a(output_13_158), .b(output_13_15), .y(output_12_158));
wire output_14_158, output_14_15, output_13_158;
mixer gate_output_13_158(.a(output_14_158), .b(output_14_15), .y(output_13_158));
wire output_15_158, output_15_15, output_14_158;
mixer gate_output_14_158(.a(output_15_158), .b(output_15_15), .y(output_14_158));
wire output_16_158, output_16_15, output_15_158;
mixer gate_output_15_158(.a(output_16_158), .b(output_16_15), .y(output_15_158));
wire output_1_159, output_1_0, output_0_159;
mixer gate_output_0_159(.a(output_1_159), .b(output_1_0), .y(output_0_159));
wire output_2_159, output_2_0, output_1_159;
mixer gate_output_1_159(.a(output_2_159), .b(output_2_0), .y(output_1_159));
wire output_3_159, output_3_0, output_2_159;
mixer gate_output_2_159(.a(output_3_159), .b(output_3_0), .y(output_2_159));
wire output_4_159, output_4_0, output_3_159;
mixer gate_output_3_159(.a(output_4_159), .b(output_4_0), .y(output_3_159));
wire output_5_159, output_5_0, output_4_159;
mixer gate_output_4_159(.a(output_5_159), .b(output_5_0), .y(output_4_159));
wire output_6_159, output_6_0, output_5_159;
mixer gate_output_5_159(.a(output_6_159), .b(output_6_0), .y(output_5_159));
wire output_7_159, output_7_0, output_6_159;
mixer gate_output_6_159(.a(output_7_159), .b(output_7_0), .y(output_6_159));
wire output_8_159, output_8_0, output_7_159;
mixer gate_output_7_159(.a(output_8_159), .b(output_8_0), .y(output_7_159));
wire output_9_159, output_9_0, output_8_159;
mixer gate_output_8_159(.a(output_9_159), .b(output_9_0), .y(output_8_159));
wire output_10_159, output_10_0, output_9_159;
mixer gate_output_9_159(.a(output_10_159), .b(output_10_0), .y(output_9_159));
wire output_11_159, output_11_0, output_10_159;
mixer gate_output_10_159(.a(output_11_159), .b(output_11_0), .y(output_10_159));
wire output_12_159, output_12_0, output_11_159;
mixer gate_output_11_159(.a(output_12_159), .b(output_12_0), .y(output_11_159));
wire output_13_159, output_13_0, output_12_159;
mixer gate_output_12_159(.a(output_13_159), .b(output_13_0), .y(output_12_159));
wire output_14_159, output_14_0, output_13_159;
mixer gate_output_13_159(.a(output_14_159), .b(output_14_0), .y(output_13_159));
wire output_15_159, output_15_0, output_14_159;
mixer gate_output_14_159(.a(output_15_159), .b(output_15_0), .y(output_14_159));
wire output_16_159, output_16_0, output_15_159;
mixer gate_output_15_159(.a(output_16_159), .b(output_16_0), .y(output_15_159));
wire output_1_160, output_1_1, output_0_160;
mixer gate_output_0_160(.a(output_1_160), .b(output_1_1), .y(output_0_160));
wire output_2_160, output_2_1, output_1_160;
mixer gate_output_1_160(.a(output_2_160), .b(output_2_1), .y(output_1_160));
wire output_3_160, output_3_1, output_2_160;
mixer gate_output_2_160(.a(output_3_160), .b(output_3_1), .y(output_2_160));
wire output_4_160, output_4_1, output_3_160;
mixer gate_output_3_160(.a(output_4_160), .b(output_4_1), .y(output_3_160));
wire output_5_160, output_5_1, output_4_160;
mixer gate_output_4_160(.a(output_5_160), .b(output_5_1), .y(output_4_160));
wire output_6_160, output_6_1, output_5_160;
mixer gate_output_5_160(.a(output_6_160), .b(output_6_1), .y(output_5_160));
wire output_7_160, output_7_1, output_6_160;
mixer gate_output_6_160(.a(output_7_160), .b(output_7_1), .y(output_6_160));
wire output_8_160, output_8_1, output_7_160;
mixer gate_output_7_160(.a(output_8_160), .b(output_8_1), .y(output_7_160));
wire output_9_160, output_9_1, output_8_160;
mixer gate_output_8_160(.a(output_9_160), .b(output_9_1), .y(output_8_160));
wire output_10_160, output_10_1, output_9_160;
mixer gate_output_9_160(.a(output_10_160), .b(output_10_1), .y(output_9_160));
wire output_11_160, output_11_1, output_10_160;
mixer gate_output_10_160(.a(output_11_160), .b(output_11_1), .y(output_10_160));
wire output_12_160, output_12_1, output_11_160;
mixer gate_output_11_160(.a(output_12_160), .b(output_12_1), .y(output_11_160));
wire output_13_160, output_13_1, output_12_160;
mixer gate_output_12_160(.a(output_13_160), .b(output_13_1), .y(output_12_160));
wire output_14_160, output_14_1, output_13_160;
mixer gate_output_13_160(.a(output_14_160), .b(output_14_1), .y(output_13_160));
wire output_15_160, output_15_1, output_14_160;
mixer gate_output_14_160(.a(output_15_160), .b(output_15_1), .y(output_14_160));
wire output_16_160, output_16_1, output_15_160;
mixer gate_output_15_160(.a(output_16_160), .b(output_16_1), .y(output_15_160));
wire output_1_161, output_1_2, output_0_161;
mixer gate_output_0_161(.a(output_1_161), .b(output_1_2), .y(output_0_161));
wire output_2_161, output_2_2, output_1_161;
mixer gate_output_1_161(.a(output_2_161), .b(output_2_2), .y(output_1_161));
wire output_3_161, output_3_2, output_2_161;
mixer gate_output_2_161(.a(output_3_161), .b(output_3_2), .y(output_2_161));
wire output_4_161, output_4_2, output_3_161;
mixer gate_output_3_161(.a(output_4_161), .b(output_4_2), .y(output_3_161));
wire output_5_161, output_5_2, output_4_161;
mixer gate_output_4_161(.a(output_5_161), .b(output_5_2), .y(output_4_161));
wire output_6_161, output_6_2, output_5_161;
mixer gate_output_5_161(.a(output_6_161), .b(output_6_2), .y(output_5_161));
wire output_7_161, output_7_2, output_6_161;
mixer gate_output_6_161(.a(output_7_161), .b(output_7_2), .y(output_6_161));
wire output_8_161, output_8_2, output_7_161;
mixer gate_output_7_161(.a(output_8_161), .b(output_8_2), .y(output_7_161));
wire output_9_161, output_9_2, output_8_161;
mixer gate_output_8_161(.a(output_9_161), .b(output_9_2), .y(output_8_161));
wire output_10_161, output_10_2, output_9_161;
mixer gate_output_9_161(.a(output_10_161), .b(output_10_2), .y(output_9_161));
wire output_11_161, output_11_2, output_10_161;
mixer gate_output_10_161(.a(output_11_161), .b(output_11_2), .y(output_10_161));
wire output_12_161, output_12_2, output_11_161;
mixer gate_output_11_161(.a(output_12_161), .b(output_12_2), .y(output_11_161));
wire output_13_161, output_13_2, output_12_161;
mixer gate_output_12_161(.a(output_13_161), .b(output_13_2), .y(output_12_161));
wire output_14_161, output_14_2, output_13_161;
mixer gate_output_13_161(.a(output_14_161), .b(output_14_2), .y(output_13_161));
wire output_15_161, output_15_2, output_14_161;
mixer gate_output_14_161(.a(output_15_161), .b(output_15_2), .y(output_14_161));
wire output_16_161, output_16_2, output_15_161;
mixer gate_output_15_161(.a(output_16_161), .b(output_16_2), .y(output_15_161));
wire output_1_162, output_1_3, output_0_162;
mixer gate_output_0_162(.a(output_1_162), .b(output_1_3), .y(output_0_162));
wire output_2_162, output_2_3, output_1_162;
mixer gate_output_1_162(.a(output_2_162), .b(output_2_3), .y(output_1_162));
wire output_3_162, output_3_3, output_2_162;
mixer gate_output_2_162(.a(output_3_162), .b(output_3_3), .y(output_2_162));
wire output_4_162, output_4_3, output_3_162;
mixer gate_output_3_162(.a(output_4_162), .b(output_4_3), .y(output_3_162));
wire output_5_162, output_5_3, output_4_162;
mixer gate_output_4_162(.a(output_5_162), .b(output_5_3), .y(output_4_162));
wire output_6_162, output_6_3, output_5_162;
mixer gate_output_5_162(.a(output_6_162), .b(output_6_3), .y(output_5_162));
wire output_7_162, output_7_3, output_6_162;
mixer gate_output_6_162(.a(output_7_162), .b(output_7_3), .y(output_6_162));
wire output_8_162, output_8_3, output_7_162;
mixer gate_output_7_162(.a(output_8_162), .b(output_8_3), .y(output_7_162));
wire output_9_162, output_9_3, output_8_162;
mixer gate_output_8_162(.a(output_9_162), .b(output_9_3), .y(output_8_162));
wire output_10_162, output_10_3, output_9_162;
mixer gate_output_9_162(.a(output_10_162), .b(output_10_3), .y(output_9_162));
wire output_11_162, output_11_3, output_10_162;
mixer gate_output_10_162(.a(output_11_162), .b(output_11_3), .y(output_10_162));
wire output_12_162, output_12_3, output_11_162;
mixer gate_output_11_162(.a(output_12_162), .b(output_12_3), .y(output_11_162));
wire output_13_162, output_13_3, output_12_162;
mixer gate_output_12_162(.a(output_13_162), .b(output_13_3), .y(output_12_162));
wire output_14_162, output_14_3, output_13_162;
mixer gate_output_13_162(.a(output_14_162), .b(output_14_3), .y(output_13_162));
wire output_15_162, output_15_3, output_14_162;
mixer gate_output_14_162(.a(output_15_162), .b(output_15_3), .y(output_14_162));
wire output_16_162, output_16_3, output_15_162;
mixer gate_output_15_162(.a(output_16_162), .b(output_16_3), .y(output_15_162));
wire output_1_163, output_1_4, output_0_163;
mixer gate_output_0_163(.a(output_1_163), .b(output_1_4), .y(output_0_163));
wire output_2_163, output_2_4, output_1_163;
mixer gate_output_1_163(.a(output_2_163), .b(output_2_4), .y(output_1_163));
wire output_3_163, output_3_4, output_2_163;
mixer gate_output_2_163(.a(output_3_163), .b(output_3_4), .y(output_2_163));
wire output_4_163, output_4_4, output_3_163;
mixer gate_output_3_163(.a(output_4_163), .b(output_4_4), .y(output_3_163));
wire output_5_163, output_5_4, output_4_163;
mixer gate_output_4_163(.a(output_5_163), .b(output_5_4), .y(output_4_163));
wire output_6_163, output_6_4, output_5_163;
mixer gate_output_5_163(.a(output_6_163), .b(output_6_4), .y(output_5_163));
wire output_7_163, output_7_4, output_6_163;
mixer gate_output_6_163(.a(output_7_163), .b(output_7_4), .y(output_6_163));
wire output_8_163, output_8_4, output_7_163;
mixer gate_output_7_163(.a(output_8_163), .b(output_8_4), .y(output_7_163));
wire output_9_163, output_9_4, output_8_163;
mixer gate_output_8_163(.a(output_9_163), .b(output_9_4), .y(output_8_163));
wire output_10_163, output_10_4, output_9_163;
mixer gate_output_9_163(.a(output_10_163), .b(output_10_4), .y(output_9_163));
wire output_11_163, output_11_4, output_10_163;
mixer gate_output_10_163(.a(output_11_163), .b(output_11_4), .y(output_10_163));
wire output_12_163, output_12_4, output_11_163;
mixer gate_output_11_163(.a(output_12_163), .b(output_12_4), .y(output_11_163));
wire output_13_163, output_13_4, output_12_163;
mixer gate_output_12_163(.a(output_13_163), .b(output_13_4), .y(output_12_163));
wire output_14_163, output_14_4, output_13_163;
mixer gate_output_13_163(.a(output_14_163), .b(output_14_4), .y(output_13_163));
wire output_15_163, output_15_4, output_14_163;
mixer gate_output_14_163(.a(output_15_163), .b(output_15_4), .y(output_14_163));
wire output_16_163, output_16_4, output_15_163;
mixer gate_output_15_163(.a(output_16_163), .b(output_16_4), .y(output_15_163));
wire output_1_164, output_1_5, output_0_164;
mixer gate_output_0_164(.a(output_1_164), .b(output_1_5), .y(output_0_164));
wire output_2_164, output_2_5, output_1_164;
mixer gate_output_1_164(.a(output_2_164), .b(output_2_5), .y(output_1_164));
wire output_3_164, output_3_5, output_2_164;
mixer gate_output_2_164(.a(output_3_164), .b(output_3_5), .y(output_2_164));
wire output_4_164, output_4_5, output_3_164;
mixer gate_output_3_164(.a(output_4_164), .b(output_4_5), .y(output_3_164));
wire output_5_164, output_5_5, output_4_164;
mixer gate_output_4_164(.a(output_5_164), .b(output_5_5), .y(output_4_164));
wire output_6_164, output_6_5, output_5_164;
mixer gate_output_5_164(.a(output_6_164), .b(output_6_5), .y(output_5_164));
wire output_7_164, output_7_5, output_6_164;
mixer gate_output_6_164(.a(output_7_164), .b(output_7_5), .y(output_6_164));
wire output_8_164, output_8_5, output_7_164;
mixer gate_output_7_164(.a(output_8_164), .b(output_8_5), .y(output_7_164));
wire output_9_164, output_9_5, output_8_164;
mixer gate_output_8_164(.a(output_9_164), .b(output_9_5), .y(output_8_164));
wire output_10_164, output_10_5, output_9_164;
mixer gate_output_9_164(.a(output_10_164), .b(output_10_5), .y(output_9_164));
wire output_11_164, output_11_5, output_10_164;
mixer gate_output_10_164(.a(output_11_164), .b(output_11_5), .y(output_10_164));
wire output_12_164, output_12_5, output_11_164;
mixer gate_output_11_164(.a(output_12_164), .b(output_12_5), .y(output_11_164));
wire output_13_164, output_13_5, output_12_164;
mixer gate_output_12_164(.a(output_13_164), .b(output_13_5), .y(output_12_164));
wire output_14_164, output_14_5, output_13_164;
mixer gate_output_13_164(.a(output_14_164), .b(output_14_5), .y(output_13_164));
wire output_15_164, output_15_5, output_14_164;
mixer gate_output_14_164(.a(output_15_164), .b(output_15_5), .y(output_14_164));
wire output_16_164, output_16_5, output_15_164;
mixer gate_output_15_164(.a(output_16_164), .b(output_16_5), .y(output_15_164));
wire output_1_165, output_1_6, output_0_165;
mixer gate_output_0_165(.a(output_1_165), .b(output_1_6), .y(output_0_165));
wire output_2_165, output_2_6, output_1_165;
mixer gate_output_1_165(.a(output_2_165), .b(output_2_6), .y(output_1_165));
wire output_3_165, output_3_6, output_2_165;
mixer gate_output_2_165(.a(output_3_165), .b(output_3_6), .y(output_2_165));
wire output_4_165, output_4_6, output_3_165;
mixer gate_output_3_165(.a(output_4_165), .b(output_4_6), .y(output_3_165));
wire output_5_165, output_5_6, output_4_165;
mixer gate_output_4_165(.a(output_5_165), .b(output_5_6), .y(output_4_165));
wire output_6_165, output_6_6, output_5_165;
mixer gate_output_5_165(.a(output_6_165), .b(output_6_6), .y(output_5_165));
wire output_7_165, output_7_6, output_6_165;
mixer gate_output_6_165(.a(output_7_165), .b(output_7_6), .y(output_6_165));
wire output_8_165, output_8_6, output_7_165;
mixer gate_output_7_165(.a(output_8_165), .b(output_8_6), .y(output_7_165));
wire output_9_165, output_9_6, output_8_165;
mixer gate_output_8_165(.a(output_9_165), .b(output_9_6), .y(output_8_165));
wire output_10_165, output_10_6, output_9_165;
mixer gate_output_9_165(.a(output_10_165), .b(output_10_6), .y(output_9_165));
wire output_11_165, output_11_6, output_10_165;
mixer gate_output_10_165(.a(output_11_165), .b(output_11_6), .y(output_10_165));
wire output_12_165, output_12_6, output_11_165;
mixer gate_output_11_165(.a(output_12_165), .b(output_12_6), .y(output_11_165));
wire output_13_165, output_13_6, output_12_165;
mixer gate_output_12_165(.a(output_13_165), .b(output_13_6), .y(output_12_165));
wire output_14_165, output_14_6, output_13_165;
mixer gate_output_13_165(.a(output_14_165), .b(output_14_6), .y(output_13_165));
wire output_15_165, output_15_6, output_14_165;
mixer gate_output_14_165(.a(output_15_165), .b(output_15_6), .y(output_14_165));
wire output_16_165, output_16_6, output_15_165;
mixer gate_output_15_165(.a(output_16_165), .b(output_16_6), .y(output_15_165));
wire output_1_166, output_1_7, output_0_166;
mixer gate_output_0_166(.a(output_1_166), .b(output_1_7), .y(output_0_166));
wire output_2_166, output_2_7, output_1_166;
mixer gate_output_1_166(.a(output_2_166), .b(output_2_7), .y(output_1_166));
wire output_3_166, output_3_7, output_2_166;
mixer gate_output_2_166(.a(output_3_166), .b(output_3_7), .y(output_2_166));
wire output_4_166, output_4_7, output_3_166;
mixer gate_output_3_166(.a(output_4_166), .b(output_4_7), .y(output_3_166));
wire output_5_166, output_5_7, output_4_166;
mixer gate_output_4_166(.a(output_5_166), .b(output_5_7), .y(output_4_166));
wire output_6_166, output_6_7, output_5_166;
mixer gate_output_5_166(.a(output_6_166), .b(output_6_7), .y(output_5_166));
wire output_7_166, output_7_7, output_6_166;
mixer gate_output_6_166(.a(output_7_166), .b(output_7_7), .y(output_6_166));
wire output_8_166, output_8_7, output_7_166;
mixer gate_output_7_166(.a(output_8_166), .b(output_8_7), .y(output_7_166));
wire output_9_166, output_9_7, output_8_166;
mixer gate_output_8_166(.a(output_9_166), .b(output_9_7), .y(output_8_166));
wire output_10_166, output_10_7, output_9_166;
mixer gate_output_9_166(.a(output_10_166), .b(output_10_7), .y(output_9_166));
wire output_11_166, output_11_7, output_10_166;
mixer gate_output_10_166(.a(output_11_166), .b(output_11_7), .y(output_10_166));
wire output_12_166, output_12_7, output_11_166;
mixer gate_output_11_166(.a(output_12_166), .b(output_12_7), .y(output_11_166));
wire output_13_166, output_13_7, output_12_166;
mixer gate_output_12_166(.a(output_13_166), .b(output_13_7), .y(output_12_166));
wire output_14_166, output_14_7, output_13_166;
mixer gate_output_13_166(.a(output_14_166), .b(output_14_7), .y(output_13_166));
wire output_15_166, output_15_7, output_14_166;
mixer gate_output_14_166(.a(output_15_166), .b(output_15_7), .y(output_14_166));
wire output_16_166, output_16_7, output_15_166;
mixer gate_output_15_166(.a(output_16_166), .b(output_16_7), .y(output_15_166));
wire output_1_167, output_1_8, output_0_167;
mixer gate_output_0_167(.a(output_1_167), .b(output_1_8), .y(output_0_167));
wire output_2_167, output_2_8, output_1_167;
mixer gate_output_1_167(.a(output_2_167), .b(output_2_8), .y(output_1_167));
wire output_3_167, output_3_8, output_2_167;
mixer gate_output_2_167(.a(output_3_167), .b(output_3_8), .y(output_2_167));
wire output_4_167, output_4_8, output_3_167;
mixer gate_output_3_167(.a(output_4_167), .b(output_4_8), .y(output_3_167));
wire output_5_167, output_5_8, output_4_167;
mixer gate_output_4_167(.a(output_5_167), .b(output_5_8), .y(output_4_167));
wire output_6_167, output_6_8, output_5_167;
mixer gate_output_5_167(.a(output_6_167), .b(output_6_8), .y(output_5_167));
wire output_7_167, output_7_8, output_6_167;
mixer gate_output_6_167(.a(output_7_167), .b(output_7_8), .y(output_6_167));
wire output_8_167, output_8_8, output_7_167;
mixer gate_output_7_167(.a(output_8_167), .b(output_8_8), .y(output_7_167));
wire output_9_167, output_9_8, output_8_167;
mixer gate_output_8_167(.a(output_9_167), .b(output_9_8), .y(output_8_167));
wire output_10_167, output_10_8, output_9_167;
mixer gate_output_9_167(.a(output_10_167), .b(output_10_8), .y(output_9_167));
wire output_11_167, output_11_8, output_10_167;
mixer gate_output_10_167(.a(output_11_167), .b(output_11_8), .y(output_10_167));
wire output_12_167, output_12_8, output_11_167;
mixer gate_output_11_167(.a(output_12_167), .b(output_12_8), .y(output_11_167));
wire output_13_167, output_13_8, output_12_167;
mixer gate_output_12_167(.a(output_13_167), .b(output_13_8), .y(output_12_167));
wire output_14_167, output_14_8, output_13_167;
mixer gate_output_13_167(.a(output_14_167), .b(output_14_8), .y(output_13_167));
wire output_15_167, output_15_8, output_14_167;
mixer gate_output_14_167(.a(output_15_167), .b(output_15_8), .y(output_14_167));
wire output_16_167, output_16_8, output_15_167;
mixer gate_output_15_167(.a(output_16_167), .b(output_16_8), .y(output_15_167));
wire output_1_168, output_1_9, output_0_168;
mixer gate_output_0_168(.a(output_1_168), .b(output_1_9), .y(output_0_168));
wire output_2_168, output_2_9, output_1_168;
mixer gate_output_1_168(.a(output_2_168), .b(output_2_9), .y(output_1_168));
wire output_3_168, output_3_9, output_2_168;
mixer gate_output_2_168(.a(output_3_168), .b(output_3_9), .y(output_2_168));
wire output_4_168, output_4_9, output_3_168;
mixer gate_output_3_168(.a(output_4_168), .b(output_4_9), .y(output_3_168));
wire output_5_168, output_5_9, output_4_168;
mixer gate_output_4_168(.a(output_5_168), .b(output_5_9), .y(output_4_168));
wire output_6_168, output_6_9, output_5_168;
mixer gate_output_5_168(.a(output_6_168), .b(output_6_9), .y(output_5_168));
wire output_7_168, output_7_9, output_6_168;
mixer gate_output_6_168(.a(output_7_168), .b(output_7_9), .y(output_6_168));
wire output_8_168, output_8_9, output_7_168;
mixer gate_output_7_168(.a(output_8_168), .b(output_8_9), .y(output_7_168));
wire output_9_168, output_9_9, output_8_168;
mixer gate_output_8_168(.a(output_9_168), .b(output_9_9), .y(output_8_168));
wire output_10_168, output_10_9, output_9_168;
mixer gate_output_9_168(.a(output_10_168), .b(output_10_9), .y(output_9_168));
wire output_11_168, output_11_9, output_10_168;
mixer gate_output_10_168(.a(output_11_168), .b(output_11_9), .y(output_10_168));
wire output_12_168, output_12_9, output_11_168;
mixer gate_output_11_168(.a(output_12_168), .b(output_12_9), .y(output_11_168));
wire output_13_168, output_13_9, output_12_168;
mixer gate_output_12_168(.a(output_13_168), .b(output_13_9), .y(output_12_168));
wire output_14_168, output_14_9, output_13_168;
mixer gate_output_13_168(.a(output_14_168), .b(output_14_9), .y(output_13_168));
wire output_15_168, output_15_9, output_14_168;
mixer gate_output_14_168(.a(output_15_168), .b(output_15_9), .y(output_14_168));
wire output_16_168, output_16_9, output_15_168;
mixer gate_output_15_168(.a(output_16_168), .b(output_16_9), .y(output_15_168));
wire output_1_169, output_1_10, output_0_169;
mixer gate_output_0_169(.a(output_1_169), .b(output_1_10), .y(output_0_169));
wire output_2_169, output_2_10, output_1_169;
mixer gate_output_1_169(.a(output_2_169), .b(output_2_10), .y(output_1_169));
wire output_3_169, output_3_10, output_2_169;
mixer gate_output_2_169(.a(output_3_169), .b(output_3_10), .y(output_2_169));
wire output_4_169, output_4_10, output_3_169;
mixer gate_output_3_169(.a(output_4_169), .b(output_4_10), .y(output_3_169));
wire output_5_169, output_5_10, output_4_169;
mixer gate_output_4_169(.a(output_5_169), .b(output_5_10), .y(output_4_169));
wire output_6_169, output_6_10, output_5_169;
mixer gate_output_5_169(.a(output_6_169), .b(output_6_10), .y(output_5_169));
wire output_7_169, output_7_10, output_6_169;
mixer gate_output_6_169(.a(output_7_169), .b(output_7_10), .y(output_6_169));
wire output_8_169, output_8_10, output_7_169;
mixer gate_output_7_169(.a(output_8_169), .b(output_8_10), .y(output_7_169));
wire output_9_169, output_9_10, output_8_169;
mixer gate_output_8_169(.a(output_9_169), .b(output_9_10), .y(output_8_169));
wire output_10_169, output_10_10, output_9_169;
mixer gate_output_9_169(.a(output_10_169), .b(output_10_10), .y(output_9_169));
wire output_11_169, output_11_10, output_10_169;
mixer gate_output_10_169(.a(output_11_169), .b(output_11_10), .y(output_10_169));
wire output_12_169, output_12_10, output_11_169;
mixer gate_output_11_169(.a(output_12_169), .b(output_12_10), .y(output_11_169));
wire output_13_169, output_13_10, output_12_169;
mixer gate_output_12_169(.a(output_13_169), .b(output_13_10), .y(output_12_169));
wire output_14_169, output_14_10, output_13_169;
mixer gate_output_13_169(.a(output_14_169), .b(output_14_10), .y(output_13_169));
wire output_15_169, output_15_10, output_14_169;
mixer gate_output_14_169(.a(output_15_169), .b(output_15_10), .y(output_14_169));
wire output_16_169, output_16_10, output_15_169;
mixer gate_output_15_169(.a(output_16_169), .b(output_16_10), .y(output_15_169));
wire output_1_170, output_1_11, output_0_170;
mixer gate_output_0_170(.a(output_1_170), .b(output_1_11), .y(output_0_170));
wire output_2_170, output_2_11, output_1_170;
mixer gate_output_1_170(.a(output_2_170), .b(output_2_11), .y(output_1_170));
wire output_3_170, output_3_11, output_2_170;
mixer gate_output_2_170(.a(output_3_170), .b(output_3_11), .y(output_2_170));
wire output_4_170, output_4_11, output_3_170;
mixer gate_output_3_170(.a(output_4_170), .b(output_4_11), .y(output_3_170));
wire output_5_170, output_5_11, output_4_170;
mixer gate_output_4_170(.a(output_5_170), .b(output_5_11), .y(output_4_170));
wire output_6_170, output_6_11, output_5_170;
mixer gate_output_5_170(.a(output_6_170), .b(output_6_11), .y(output_5_170));
wire output_7_170, output_7_11, output_6_170;
mixer gate_output_6_170(.a(output_7_170), .b(output_7_11), .y(output_6_170));
wire output_8_170, output_8_11, output_7_170;
mixer gate_output_7_170(.a(output_8_170), .b(output_8_11), .y(output_7_170));
wire output_9_170, output_9_11, output_8_170;
mixer gate_output_8_170(.a(output_9_170), .b(output_9_11), .y(output_8_170));
wire output_10_170, output_10_11, output_9_170;
mixer gate_output_9_170(.a(output_10_170), .b(output_10_11), .y(output_9_170));
wire output_11_170, output_11_11, output_10_170;
mixer gate_output_10_170(.a(output_11_170), .b(output_11_11), .y(output_10_170));
wire output_12_170, output_12_11, output_11_170;
mixer gate_output_11_170(.a(output_12_170), .b(output_12_11), .y(output_11_170));
wire output_13_170, output_13_11, output_12_170;
mixer gate_output_12_170(.a(output_13_170), .b(output_13_11), .y(output_12_170));
wire output_14_170, output_14_11, output_13_170;
mixer gate_output_13_170(.a(output_14_170), .b(output_14_11), .y(output_13_170));
wire output_15_170, output_15_11, output_14_170;
mixer gate_output_14_170(.a(output_15_170), .b(output_15_11), .y(output_14_170));
wire output_16_170, output_16_11, output_15_170;
mixer gate_output_15_170(.a(output_16_170), .b(output_16_11), .y(output_15_170));
wire output_1_171, output_1_12, output_0_171;
mixer gate_output_0_171(.a(output_1_171), .b(output_1_12), .y(output_0_171));
wire output_2_171, output_2_12, output_1_171;
mixer gate_output_1_171(.a(output_2_171), .b(output_2_12), .y(output_1_171));
wire output_3_171, output_3_12, output_2_171;
mixer gate_output_2_171(.a(output_3_171), .b(output_3_12), .y(output_2_171));
wire output_4_171, output_4_12, output_3_171;
mixer gate_output_3_171(.a(output_4_171), .b(output_4_12), .y(output_3_171));
wire output_5_171, output_5_12, output_4_171;
mixer gate_output_4_171(.a(output_5_171), .b(output_5_12), .y(output_4_171));
wire output_6_171, output_6_12, output_5_171;
mixer gate_output_5_171(.a(output_6_171), .b(output_6_12), .y(output_5_171));
wire output_7_171, output_7_12, output_6_171;
mixer gate_output_6_171(.a(output_7_171), .b(output_7_12), .y(output_6_171));
wire output_8_171, output_8_12, output_7_171;
mixer gate_output_7_171(.a(output_8_171), .b(output_8_12), .y(output_7_171));
wire output_9_171, output_9_12, output_8_171;
mixer gate_output_8_171(.a(output_9_171), .b(output_9_12), .y(output_8_171));
wire output_10_171, output_10_12, output_9_171;
mixer gate_output_9_171(.a(output_10_171), .b(output_10_12), .y(output_9_171));
wire output_11_171, output_11_12, output_10_171;
mixer gate_output_10_171(.a(output_11_171), .b(output_11_12), .y(output_10_171));
wire output_12_171, output_12_12, output_11_171;
mixer gate_output_11_171(.a(output_12_171), .b(output_12_12), .y(output_11_171));
wire output_13_171, output_13_12, output_12_171;
mixer gate_output_12_171(.a(output_13_171), .b(output_13_12), .y(output_12_171));
wire output_14_171, output_14_12, output_13_171;
mixer gate_output_13_171(.a(output_14_171), .b(output_14_12), .y(output_13_171));
wire output_15_171, output_15_12, output_14_171;
mixer gate_output_14_171(.a(output_15_171), .b(output_15_12), .y(output_14_171));
wire output_16_171, output_16_12, output_15_171;
mixer gate_output_15_171(.a(output_16_171), .b(output_16_12), .y(output_15_171));
wire output_1_172, output_1_13, output_0_172;
mixer gate_output_0_172(.a(output_1_172), .b(output_1_13), .y(output_0_172));
wire output_2_172, output_2_13, output_1_172;
mixer gate_output_1_172(.a(output_2_172), .b(output_2_13), .y(output_1_172));
wire output_3_172, output_3_13, output_2_172;
mixer gate_output_2_172(.a(output_3_172), .b(output_3_13), .y(output_2_172));
wire output_4_172, output_4_13, output_3_172;
mixer gate_output_3_172(.a(output_4_172), .b(output_4_13), .y(output_3_172));
wire output_5_172, output_5_13, output_4_172;
mixer gate_output_4_172(.a(output_5_172), .b(output_5_13), .y(output_4_172));
wire output_6_172, output_6_13, output_5_172;
mixer gate_output_5_172(.a(output_6_172), .b(output_6_13), .y(output_5_172));
wire output_7_172, output_7_13, output_6_172;
mixer gate_output_6_172(.a(output_7_172), .b(output_7_13), .y(output_6_172));
wire output_8_172, output_8_13, output_7_172;
mixer gate_output_7_172(.a(output_8_172), .b(output_8_13), .y(output_7_172));
wire output_9_172, output_9_13, output_8_172;
mixer gate_output_8_172(.a(output_9_172), .b(output_9_13), .y(output_8_172));
wire output_10_172, output_10_13, output_9_172;
mixer gate_output_9_172(.a(output_10_172), .b(output_10_13), .y(output_9_172));
wire output_11_172, output_11_13, output_10_172;
mixer gate_output_10_172(.a(output_11_172), .b(output_11_13), .y(output_10_172));
wire output_12_172, output_12_13, output_11_172;
mixer gate_output_11_172(.a(output_12_172), .b(output_12_13), .y(output_11_172));
wire output_13_172, output_13_13, output_12_172;
mixer gate_output_12_172(.a(output_13_172), .b(output_13_13), .y(output_12_172));
wire output_14_172, output_14_13, output_13_172;
mixer gate_output_13_172(.a(output_14_172), .b(output_14_13), .y(output_13_172));
wire output_15_172, output_15_13, output_14_172;
mixer gate_output_14_172(.a(output_15_172), .b(output_15_13), .y(output_14_172));
wire output_16_172, output_16_13, output_15_172;
mixer gate_output_15_172(.a(output_16_172), .b(output_16_13), .y(output_15_172));
wire output_1_173, output_1_14, output_0_173;
mixer gate_output_0_173(.a(output_1_173), .b(output_1_14), .y(output_0_173));
wire output_2_173, output_2_14, output_1_173;
mixer gate_output_1_173(.a(output_2_173), .b(output_2_14), .y(output_1_173));
wire output_3_173, output_3_14, output_2_173;
mixer gate_output_2_173(.a(output_3_173), .b(output_3_14), .y(output_2_173));
wire output_4_173, output_4_14, output_3_173;
mixer gate_output_3_173(.a(output_4_173), .b(output_4_14), .y(output_3_173));
wire output_5_173, output_5_14, output_4_173;
mixer gate_output_4_173(.a(output_5_173), .b(output_5_14), .y(output_4_173));
wire output_6_173, output_6_14, output_5_173;
mixer gate_output_5_173(.a(output_6_173), .b(output_6_14), .y(output_5_173));
wire output_7_173, output_7_14, output_6_173;
mixer gate_output_6_173(.a(output_7_173), .b(output_7_14), .y(output_6_173));
wire output_8_173, output_8_14, output_7_173;
mixer gate_output_7_173(.a(output_8_173), .b(output_8_14), .y(output_7_173));
wire output_9_173, output_9_14, output_8_173;
mixer gate_output_8_173(.a(output_9_173), .b(output_9_14), .y(output_8_173));
wire output_10_173, output_10_14, output_9_173;
mixer gate_output_9_173(.a(output_10_173), .b(output_10_14), .y(output_9_173));
wire output_11_173, output_11_14, output_10_173;
mixer gate_output_10_173(.a(output_11_173), .b(output_11_14), .y(output_10_173));
wire output_12_173, output_12_14, output_11_173;
mixer gate_output_11_173(.a(output_12_173), .b(output_12_14), .y(output_11_173));
wire output_13_173, output_13_14, output_12_173;
mixer gate_output_12_173(.a(output_13_173), .b(output_13_14), .y(output_12_173));
wire output_14_173, output_14_14, output_13_173;
mixer gate_output_13_173(.a(output_14_173), .b(output_14_14), .y(output_13_173));
wire output_15_173, output_15_14, output_14_173;
mixer gate_output_14_173(.a(output_15_173), .b(output_15_14), .y(output_14_173));
wire output_16_173, output_16_14, output_15_173;
mixer gate_output_15_173(.a(output_16_173), .b(output_16_14), .y(output_15_173));
wire output_1_174, output_1_15, output_0_174;
mixer gate_output_0_174(.a(output_1_174), .b(output_1_15), .y(output_0_174));
wire output_2_174, output_2_15, output_1_174;
mixer gate_output_1_174(.a(output_2_174), .b(output_2_15), .y(output_1_174));
wire output_3_174, output_3_15, output_2_174;
mixer gate_output_2_174(.a(output_3_174), .b(output_3_15), .y(output_2_174));
wire output_4_174, output_4_15, output_3_174;
mixer gate_output_3_174(.a(output_4_174), .b(output_4_15), .y(output_3_174));
wire output_5_174, output_5_15, output_4_174;
mixer gate_output_4_174(.a(output_5_174), .b(output_5_15), .y(output_4_174));
wire output_6_174, output_6_15, output_5_174;
mixer gate_output_5_174(.a(output_6_174), .b(output_6_15), .y(output_5_174));
wire output_7_174, output_7_15, output_6_174;
mixer gate_output_6_174(.a(output_7_174), .b(output_7_15), .y(output_6_174));
wire output_8_174, output_8_15, output_7_174;
mixer gate_output_7_174(.a(output_8_174), .b(output_8_15), .y(output_7_174));
wire output_9_174, output_9_15, output_8_174;
mixer gate_output_8_174(.a(output_9_174), .b(output_9_15), .y(output_8_174));
wire output_10_174, output_10_15, output_9_174;
mixer gate_output_9_174(.a(output_10_174), .b(output_10_15), .y(output_9_174));
wire output_11_174, output_11_15, output_10_174;
mixer gate_output_10_174(.a(output_11_174), .b(output_11_15), .y(output_10_174));
wire output_12_174, output_12_15, output_11_174;
mixer gate_output_11_174(.a(output_12_174), .b(output_12_15), .y(output_11_174));
wire output_13_174, output_13_15, output_12_174;
mixer gate_output_12_174(.a(output_13_174), .b(output_13_15), .y(output_12_174));
wire output_14_174, output_14_15, output_13_174;
mixer gate_output_13_174(.a(output_14_174), .b(output_14_15), .y(output_13_174));
wire output_15_174, output_15_15, output_14_174;
mixer gate_output_14_174(.a(output_15_174), .b(output_15_15), .y(output_14_174));
wire output_16_174, output_16_15, output_15_174;
mixer gate_output_15_174(.a(output_16_174), .b(output_16_15), .y(output_15_174));
wire output_1_175, output_1_0, output_0_175;
mixer gate_output_0_175(.a(output_1_175), .b(output_1_0), .y(output_0_175));
wire output_2_175, output_2_0, output_1_175;
mixer gate_output_1_175(.a(output_2_175), .b(output_2_0), .y(output_1_175));
wire output_3_175, output_3_0, output_2_175;
mixer gate_output_2_175(.a(output_3_175), .b(output_3_0), .y(output_2_175));
wire output_4_175, output_4_0, output_3_175;
mixer gate_output_3_175(.a(output_4_175), .b(output_4_0), .y(output_3_175));
wire output_5_175, output_5_0, output_4_175;
mixer gate_output_4_175(.a(output_5_175), .b(output_5_0), .y(output_4_175));
wire output_6_175, output_6_0, output_5_175;
mixer gate_output_5_175(.a(output_6_175), .b(output_6_0), .y(output_5_175));
wire output_7_175, output_7_0, output_6_175;
mixer gate_output_6_175(.a(output_7_175), .b(output_7_0), .y(output_6_175));
wire output_8_175, output_8_0, output_7_175;
mixer gate_output_7_175(.a(output_8_175), .b(output_8_0), .y(output_7_175));
wire output_9_175, output_9_0, output_8_175;
mixer gate_output_8_175(.a(output_9_175), .b(output_9_0), .y(output_8_175));
wire output_10_175, output_10_0, output_9_175;
mixer gate_output_9_175(.a(output_10_175), .b(output_10_0), .y(output_9_175));
wire output_11_175, output_11_0, output_10_175;
mixer gate_output_10_175(.a(output_11_175), .b(output_11_0), .y(output_10_175));
wire output_12_175, output_12_0, output_11_175;
mixer gate_output_11_175(.a(output_12_175), .b(output_12_0), .y(output_11_175));
wire output_13_175, output_13_0, output_12_175;
mixer gate_output_12_175(.a(output_13_175), .b(output_13_0), .y(output_12_175));
wire output_14_175, output_14_0, output_13_175;
mixer gate_output_13_175(.a(output_14_175), .b(output_14_0), .y(output_13_175));
wire output_15_175, output_15_0, output_14_175;
mixer gate_output_14_175(.a(output_15_175), .b(output_15_0), .y(output_14_175));
wire output_16_175, output_16_0, output_15_175;
mixer gate_output_15_175(.a(output_16_175), .b(output_16_0), .y(output_15_175));
wire output_1_176, output_1_1, output_0_176;
mixer gate_output_0_176(.a(output_1_176), .b(output_1_1), .y(output_0_176));
wire output_2_176, output_2_1, output_1_176;
mixer gate_output_1_176(.a(output_2_176), .b(output_2_1), .y(output_1_176));
wire output_3_176, output_3_1, output_2_176;
mixer gate_output_2_176(.a(output_3_176), .b(output_3_1), .y(output_2_176));
wire output_4_176, output_4_1, output_3_176;
mixer gate_output_3_176(.a(output_4_176), .b(output_4_1), .y(output_3_176));
wire output_5_176, output_5_1, output_4_176;
mixer gate_output_4_176(.a(output_5_176), .b(output_5_1), .y(output_4_176));
wire output_6_176, output_6_1, output_5_176;
mixer gate_output_5_176(.a(output_6_176), .b(output_6_1), .y(output_5_176));
wire output_7_176, output_7_1, output_6_176;
mixer gate_output_6_176(.a(output_7_176), .b(output_7_1), .y(output_6_176));
wire output_8_176, output_8_1, output_7_176;
mixer gate_output_7_176(.a(output_8_176), .b(output_8_1), .y(output_7_176));
wire output_9_176, output_9_1, output_8_176;
mixer gate_output_8_176(.a(output_9_176), .b(output_9_1), .y(output_8_176));
wire output_10_176, output_10_1, output_9_176;
mixer gate_output_9_176(.a(output_10_176), .b(output_10_1), .y(output_9_176));
wire output_11_176, output_11_1, output_10_176;
mixer gate_output_10_176(.a(output_11_176), .b(output_11_1), .y(output_10_176));
wire output_12_176, output_12_1, output_11_176;
mixer gate_output_11_176(.a(output_12_176), .b(output_12_1), .y(output_11_176));
wire output_13_176, output_13_1, output_12_176;
mixer gate_output_12_176(.a(output_13_176), .b(output_13_1), .y(output_12_176));
wire output_14_176, output_14_1, output_13_176;
mixer gate_output_13_176(.a(output_14_176), .b(output_14_1), .y(output_13_176));
wire output_15_176, output_15_1, output_14_176;
mixer gate_output_14_176(.a(output_15_176), .b(output_15_1), .y(output_14_176));
wire output_16_176, output_16_1, output_15_176;
mixer gate_output_15_176(.a(output_16_176), .b(output_16_1), .y(output_15_176));
wire output_1_177, output_1_2, output_0_177;
mixer gate_output_0_177(.a(output_1_177), .b(output_1_2), .y(output_0_177));
wire output_2_177, output_2_2, output_1_177;
mixer gate_output_1_177(.a(output_2_177), .b(output_2_2), .y(output_1_177));
wire output_3_177, output_3_2, output_2_177;
mixer gate_output_2_177(.a(output_3_177), .b(output_3_2), .y(output_2_177));
wire output_4_177, output_4_2, output_3_177;
mixer gate_output_3_177(.a(output_4_177), .b(output_4_2), .y(output_3_177));
wire output_5_177, output_5_2, output_4_177;
mixer gate_output_4_177(.a(output_5_177), .b(output_5_2), .y(output_4_177));
wire output_6_177, output_6_2, output_5_177;
mixer gate_output_5_177(.a(output_6_177), .b(output_6_2), .y(output_5_177));
wire output_7_177, output_7_2, output_6_177;
mixer gate_output_6_177(.a(output_7_177), .b(output_7_2), .y(output_6_177));
wire output_8_177, output_8_2, output_7_177;
mixer gate_output_7_177(.a(output_8_177), .b(output_8_2), .y(output_7_177));
wire output_9_177, output_9_2, output_8_177;
mixer gate_output_8_177(.a(output_9_177), .b(output_9_2), .y(output_8_177));
wire output_10_177, output_10_2, output_9_177;
mixer gate_output_9_177(.a(output_10_177), .b(output_10_2), .y(output_9_177));
wire output_11_177, output_11_2, output_10_177;
mixer gate_output_10_177(.a(output_11_177), .b(output_11_2), .y(output_10_177));
wire output_12_177, output_12_2, output_11_177;
mixer gate_output_11_177(.a(output_12_177), .b(output_12_2), .y(output_11_177));
wire output_13_177, output_13_2, output_12_177;
mixer gate_output_12_177(.a(output_13_177), .b(output_13_2), .y(output_12_177));
wire output_14_177, output_14_2, output_13_177;
mixer gate_output_13_177(.a(output_14_177), .b(output_14_2), .y(output_13_177));
wire output_15_177, output_15_2, output_14_177;
mixer gate_output_14_177(.a(output_15_177), .b(output_15_2), .y(output_14_177));
wire output_16_177, output_16_2, output_15_177;
mixer gate_output_15_177(.a(output_16_177), .b(output_16_2), .y(output_15_177));
wire output_1_178, output_1_3, output_0_178;
mixer gate_output_0_178(.a(output_1_178), .b(output_1_3), .y(output_0_178));
wire output_2_178, output_2_3, output_1_178;
mixer gate_output_1_178(.a(output_2_178), .b(output_2_3), .y(output_1_178));
wire output_3_178, output_3_3, output_2_178;
mixer gate_output_2_178(.a(output_3_178), .b(output_3_3), .y(output_2_178));
wire output_4_178, output_4_3, output_3_178;
mixer gate_output_3_178(.a(output_4_178), .b(output_4_3), .y(output_3_178));
wire output_5_178, output_5_3, output_4_178;
mixer gate_output_4_178(.a(output_5_178), .b(output_5_3), .y(output_4_178));
wire output_6_178, output_6_3, output_5_178;
mixer gate_output_5_178(.a(output_6_178), .b(output_6_3), .y(output_5_178));
wire output_7_178, output_7_3, output_6_178;
mixer gate_output_6_178(.a(output_7_178), .b(output_7_3), .y(output_6_178));
wire output_8_178, output_8_3, output_7_178;
mixer gate_output_7_178(.a(output_8_178), .b(output_8_3), .y(output_7_178));
wire output_9_178, output_9_3, output_8_178;
mixer gate_output_8_178(.a(output_9_178), .b(output_9_3), .y(output_8_178));
wire output_10_178, output_10_3, output_9_178;
mixer gate_output_9_178(.a(output_10_178), .b(output_10_3), .y(output_9_178));
wire output_11_178, output_11_3, output_10_178;
mixer gate_output_10_178(.a(output_11_178), .b(output_11_3), .y(output_10_178));
wire output_12_178, output_12_3, output_11_178;
mixer gate_output_11_178(.a(output_12_178), .b(output_12_3), .y(output_11_178));
wire output_13_178, output_13_3, output_12_178;
mixer gate_output_12_178(.a(output_13_178), .b(output_13_3), .y(output_12_178));
wire output_14_178, output_14_3, output_13_178;
mixer gate_output_13_178(.a(output_14_178), .b(output_14_3), .y(output_13_178));
wire output_15_178, output_15_3, output_14_178;
mixer gate_output_14_178(.a(output_15_178), .b(output_15_3), .y(output_14_178));
wire output_16_178, output_16_3, output_15_178;
mixer gate_output_15_178(.a(output_16_178), .b(output_16_3), .y(output_15_178));
wire output_1_179, output_1_4, output_0_179;
mixer gate_output_0_179(.a(output_1_179), .b(output_1_4), .y(output_0_179));
wire output_2_179, output_2_4, output_1_179;
mixer gate_output_1_179(.a(output_2_179), .b(output_2_4), .y(output_1_179));
wire output_3_179, output_3_4, output_2_179;
mixer gate_output_2_179(.a(output_3_179), .b(output_3_4), .y(output_2_179));
wire output_4_179, output_4_4, output_3_179;
mixer gate_output_3_179(.a(output_4_179), .b(output_4_4), .y(output_3_179));
wire output_5_179, output_5_4, output_4_179;
mixer gate_output_4_179(.a(output_5_179), .b(output_5_4), .y(output_4_179));
wire output_6_179, output_6_4, output_5_179;
mixer gate_output_5_179(.a(output_6_179), .b(output_6_4), .y(output_5_179));
wire output_7_179, output_7_4, output_6_179;
mixer gate_output_6_179(.a(output_7_179), .b(output_7_4), .y(output_6_179));
wire output_8_179, output_8_4, output_7_179;
mixer gate_output_7_179(.a(output_8_179), .b(output_8_4), .y(output_7_179));
wire output_9_179, output_9_4, output_8_179;
mixer gate_output_8_179(.a(output_9_179), .b(output_9_4), .y(output_8_179));
wire output_10_179, output_10_4, output_9_179;
mixer gate_output_9_179(.a(output_10_179), .b(output_10_4), .y(output_9_179));
wire output_11_179, output_11_4, output_10_179;
mixer gate_output_10_179(.a(output_11_179), .b(output_11_4), .y(output_10_179));
wire output_12_179, output_12_4, output_11_179;
mixer gate_output_11_179(.a(output_12_179), .b(output_12_4), .y(output_11_179));
wire output_13_179, output_13_4, output_12_179;
mixer gate_output_12_179(.a(output_13_179), .b(output_13_4), .y(output_12_179));
wire output_14_179, output_14_4, output_13_179;
mixer gate_output_13_179(.a(output_14_179), .b(output_14_4), .y(output_13_179));
wire output_15_179, output_15_4, output_14_179;
mixer gate_output_14_179(.a(output_15_179), .b(output_15_4), .y(output_14_179));
wire output_16_179, output_16_4, output_15_179;
mixer gate_output_15_179(.a(output_16_179), .b(output_16_4), .y(output_15_179));
wire output_1_180, output_1_5, output_0_180;
mixer gate_output_0_180(.a(output_1_180), .b(output_1_5), .y(output_0_180));
wire output_2_180, output_2_5, output_1_180;
mixer gate_output_1_180(.a(output_2_180), .b(output_2_5), .y(output_1_180));
wire output_3_180, output_3_5, output_2_180;
mixer gate_output_2_180(.a(output_3_180), .b(output_3_5), .y(output_2_180));
wire output_4_180, output_4_5, output_3_180;
mixer gate_output_3_180(.a(output_4_180), .b(output_4_5), .y(output_3_180));
wire output_5_180, output_5_5, output_4_180;
mixer gate_output_4_180(.a(output_5_180), .b(output_5_5), .y(output_4_180));
wire output_6_180, output_6_5, output_5_180;
mixer gate_output_5_180(.a(output_6_180), .b(output_6_5), .y(output_5_180));
wire output_7_180, output_7_5, output_6_180;
mixer gate_output_6_180(.a(output_7_180), .b(output_7_5), .y(output_6_180));
wire output_8_180, output_8_5, output_7_180;
mixer gate_output_7_180(.a(output_8_180), .b(output_8_5), .y(output_7_180));
wire output_9_180, output_9_5, output_8_180;
mixer gate_output_8_180(.a(output_9_180), .b(output_9_5), .y(output_8_180));
wire output_10_180, output_10_5, output_9_180;
mixer gate_output_9_180(.a(output_10_180), .b(output_10_5), .y(output_9_180));
wire output_11_180, output_11_5, output_10_180;
mixer gate_output_10_180(.a(output_11_180), .b(output_11_5), .y(output_10_180));
wire output_12_180, output_12_5, output_11_180;
mixer gate_output_11_180(.a(output_12_180), .b(output_12_5), .y(output_11_180));
wire output_13_180, output_13_5, output_12_180;
mixer gate_output_12_180(.a(output_13_180), .b(output_13_5), .y(output_12_180));
wire output_14_180, output_14_5, output_13_180;
mixer gate_output_13_180(.a(output_14_180), .b(output_14_5), .y(output_13_180));
wire output_15_180, output_15_5, output_14_180;
mixer gate_output_14_180(.a(output_15_180), .b(output_15_5), .y(output_14_180));
wire output_16_180, output_16_5, output_15_180;
mixer gate_output_15_180(.a(output_16_180), .b(output_16_5), .y(output_15_180));
wire output_1_181, output_1_6, output_0_181;
mixer gate_output_0_181(.a(output_1_181), .b(output_1_6), .y(output_0_181));
wire output_2_181, output_2_6, output_1_181;
mixer gate_output_1_181(.a(output_2_181), .b(output_2_6), .y(output_1_181));
wire output_3_181, output_3_6, output_2_181;
mixer gate_output_2_181(.a(output_3_181), .b(output_3_6), .y(output_2_181));
wire output_4_181, output_4_6, output_3_181;
mixer gate_output_3_181(.a(output_4_181), .b(output_4_6), .y(output_3_181));
wire output_5_181, output_5_6, output_4_181;
mixer gate_output_4_181(.a(output_5_181), .b(output_5_6), .y(output_4_181));
wire output_6_181, output_6_6, output_5_181;
mixer gate_output_5_181(.a(output_6_181), .b(output_6_6), .y(output_5_181));
wire output_7_181, output_7_6, output_6_181;
mixer gate_output_6_181(.a(output_7_181), .b(output_7_6), .y(output_6_181));
wire output_8_181, output_8_6, output_7_181;
mixer gate_output_7_181(.a(output_8_181), .b(output_8_6), .y(output_7_181));
wire output_9_181, output_9_6, output_8_181;
mixer gate_output_8_181(.a(output_9_181), .b(output_9_6), .y(output_8_181));
wire output_10_181, output_10_6, output_9_181;
mixer gate_output_9_181(.a(output_10_181), .b(output_10_6), .y(output_9_181));
wire output_11_181, output_11_6, output_10_181;
mixer gate_output_10_181(.a(output_11_181), .b(output_11_6), .y(output_10_181));
wire output_12_181, output_12_6, output_11_181;
mixer gate_output_11_181(.a(output_12_181), .b(output_12_6), .y(output_11_181));
wire output_13_181, output_13_6, output_12_181;
mixer gate_output_12_181(.a(output_13_181), .b(output_13_6), .y(output_12_181));
wire output_14_181, output_14_6, output_13_181;
mixer gate_output_13_181(.a(output_14_181), .b(output_14_6), .y(output_13_181));
wire output_15_181, output_15_6, output_14_181;
mixer gate_output_14_181(.a(output_15_181), .b(output_15_6), .y(output_14_181));
wire output_16_181, output_16_6, output_15_181;
mixer gate_output_15_181(.a(output_16_181), .b(output_16_6), .y(output_15_181));
wire output_1_182, output_1_7, output_0_182;
mixer gate_output_0_182(.a(output_1_182), .b(output_1_7), .y(output_0_182));
wire output_2_182, output_2_7, output_1_182;
mixer gate_output_1_182(.a(output_2_182), .b(output_2_7), .y(output_1_182));
wire output_3_182, output_3_7, output_2_182;
mixer gate_output_2_182(.a(output_3_182), .b(output_3_7), .y(output_2_182));
wire output_4_182, output_4_7, output_3_182;
mixer gate_output_3_182(.a(output_4_182), .b(output_4_7), .y(output_3_182));
wire output_5_182, output_5_7, output_4_182;
mixer gate_output_4_182(.a(output_5_182), .b(output_5_7), .y(output_4_182));
wire output_6_182, output_6_7, output_5_182;
mixer gate_output_5_182(.a(output_6_182), .b(output_6_7), .y(output_5_182));
wire output_7_182, output_7_7, output_6_182;
mixer gate_output_6_182(.a(output_7_182), .b(output_7_7), .y(output_6_182));
wire output_8_182, output_8_7, output_7_182;
mixer gate_output_7_182(.a(output_8_182), .b(output_8_7), .y(output_7_182));
wire output_9_182, output_9_7, output_8_182;
mixer gate_output_8_182(.a(output_9_182), .b(output_9_7), .y(output_8_182));
wire output_10_182, output_10_7, output_9_182;
mixer gate_output_9_182(.a(output_10_182), .b(output_10_7), .y(output_9_182));
wire output_11_182, output_11_7, output_10_182;
mixer gate_output_10_182(.a(output_11_182), .b(output_11_7), .y(output_10_182));
wire output_12_182, output_12_7, output_11_182;
mixer gate_output_11_182(.a(output_12_182), .b(output_12_7), .y(output_11_182));
wire output_13_182, output_13_7, output_12_182;
mixer gate_output_12_182(.a(output_13_182), .b(output_13_7), .y(output_12_182));
wire output_14_182, output_14_7, output_13_182;
mixer gate_output_13_182(.a(output_14_182), .b(output_14_7), .y(output_13_182));
wire output_15_182, output_15_7, output_14_182;
mixer gate_output_14_182(.a(output_15_182), .b(output_15_7), .y(output_14_182));
wire output_16_182, output_16_7, output_15_182;
mixer gate_output_15_182(.a(output_16_182), .b(output_16_7), .y(output_15_182));
wire output_1_183, output_1_8, output_0_183;
mixer gate_output_0_183(.a(output_1_183), .b(output_1_8), .y(output_0_183));
wire output_2_183, output_2_8, output_1_183;
mixer gate_output_1_183(.a(output_2_183), .b(output_2_8), .y(output_1_183));
wire output_3_183, output_3_8, output_2_183;
mixer gate_output_2_183(.a(output_3_183), .b(output_3_8), .y(output_2_183));
wire output_4_183, output_4_8, output_3_183;
mixer gate_output_3_183(.a(output_4_183), .b(output_4_8), .y(output_3_183));
wire output_5_183, output_5_8, output_4_183;
mixer gate_output_4_183(.a(output_5_183), .b(output_5_8), .y(output_4_183));
wire output_6_183, output_6_8, output_5_183;
mixer gate_output_5_183(.a(output_6_183), .b(output_6_8), .y(output_5_183));
wire output_7_183, output_7_8, output_6_183;
mixer gate_output_6_183(.a(output_7_183), .b(output_7_8), .y(output_6_183));
wire output_8_183, output_8_8, output_7_183;
mixer gate_output_7_183(.a(output_8_183), .b(output_8_8), .y(output_7_183));
wire output_9_183, output_9_8, output_8_183;
mixer gate_output_8_183(.a(output_9_183), .b(output_9_8), .y(output_8_183));
wire output_10_183, output_10_8, output_9_183;
mixer gate_output_9_183(.a(output_10_183), .b(output_10_8), .y(output_9_183));
wire output_11_183, output_11_8, output_10_183;
mixer gate_output_10_183(.a(output_11_183), .b(output_11_8), .y(output_10_183));
wire output_12_183, output_12_8, output_11_183;
mixer gate_output_11_183(.a(output_12_183), .b(output_12_8), .y(output_11_183));
wire output_13_183, output_13_8, output_12_183;
mixer gate_output_12_183(.a(output_13_183), .b(output_13_8), .y(output_12_183));
wire output_14_183, output_14_8, output_13_183;
mixer gate_output_13_183(.a(output_14_183), .b(output_14_8), .y(output_13_183));
wire output_15_183, output_15_8, output_14_183;
mixer gate_output_14_183(.a(output_15_183), .b(output_15_8), .y(output_14_183));
wire output_16_183, output_16_8, output_15_183;
mixer gate_output_15_183(.a(output_16_183), .b(output_16_8), .y(output_15_183));
wire output_1_184, output_1_9, output_0_184;
mixer gate_output_0_184(.a(output_1_184), .b(output_1_9), .y(output_0_184));
wire output_2_184, output_2_9, output_1_184;
mixer gate_output_1_184(.a(output_2_184), .b(output_2_9), .y(output_1_184));
wire output_3_184, output_3_9, output_2_184;
mixer gate_output_2_184(.a(output_3_184), .b(output_3_9), .y(output_2_184));
wire output_4_184, output_4_9, output_3_184;
mixer gate_output_3_184(.a(output_4_184), .b(output_4_9), .y(output_3_184));
wire output_5_184, output_5_9, output_4_184;
mixer gate_output_4_184(.a(output_5_184), .b(output_5_9), .y(output_4_184));
wire output_6_184, output_6_9, output_5_184;
mixer gate_output_5_184(.a(output_6_184), .b(output_6_9), .y(output_5_184));
wire output_7_184, output_7_9, output_6_184;
mixer gate_output_6_184(.a(output_7_184), .b(output_7_9), .y(output_6_184));
wire output_8_184, output_8_9, output_7_184;
mixer gate_output_7_184(.a(output_8_184), .b(output_8_9), .y(output_7_184));
wire output_9_184, output_9_9, output_8_184;
mixer gate_output_8_184(.a(output_9_184), .b(output_9_9), .y(output_8_184));
wire output_10_184, output_10_9, output_9_184;
mixer gate_output_9_184(.a(output_10_184), .b(output_10_9), .y(output_9_184));
wire output_11_184, output_11_9, output_10_184;
mixer gate_output_10_184(.a(output_11_184), .b(output_11_9), .y(output_10_184));
wire output_12_184, output_12_9, output_11_184;
mixer gate_output_11_184(.a(output_12_184), .b(output_12_9), .y(output_11_184));
wire output_13_184, output_13_9, output_12_184;
mixer gate_output_12_184(.a(output_13_184), .b(output_13_9), .y(output_12_184));
wire output_14_184, output_14_9, output_13_184;
mixer gate_output_13_184(.a(output_14_184), .b(output_14_9), .y(output_13_184));
wire output_15_184, output_15_9, output_14_184;
mixer gate_output_14_184(.a(output_15_184), .b(output_15_9), .y(output_14_184));
wire output_16_184, output_16_9, output_15_184;
mixer gate_output_15_184(.a(output_16_184), .b(output_16_9), .y(output_15_184));
wire output_1_185, output_1_10, output_0_185;
mixer gate_output_0_185(.a(output_1_185), .b(output_1_10), .y(output_0_185));
wire output_2_185, output_2_10, output_1_185;
mixer gate_output_1_185(.a(output_2_185), .b(output_2_10), .y(output_1_185));
wire output_3_185, output_3_10, output_2_185;
mixer gate_output_2_185(.a(output_3_185), .b(output_3_10), .y(output_2_185));
wire output_4_185, output_4_10, output_3_185;
mixer gate_output_3_185(.a(output_4_185), .b(output_4_10), .y(output_3_185));
wire output_5_185, output_5_10, output_4_185;
mixer gate_output_4_185(.a(output_5_185), .b(output_5_10), .y(output_4_185));
wire output_6_185, output_6_10, output_5_185;
mixer gate_output_5_185(.a(output_6_185), .b(output_6_10), .y(output_5_185));
wire output_7_185, output_7_10, output_6_185;
mixer gate_output_6_185(.a(output_7_185), .b(output_7_10), .y(output_6_185));
wire output_8_185, output_8_10, output_7_185;
mixer gate_output_7_185(.a(output_8_185), .b(output_8_10), .y(output_7_185));
wire output_9_185, output_9_10, output_8_185;
mixer gate_output_8_185(.a(output_9_185), .b(output_9_10), .y(output_8_185));
wire output_10_185, output_10_10, output_9_185;
mixer gate_output_9_185(.a(output_10_185), .b(output_10_10), .y(output_9_185));
wire output_11_185, output_11_10, output_10_185;
mixer gate_output_10_185(.a(output_11_185), .b(output_11_10), .y(output_10_185));
wire output_12_185, output_12_10, output_11_185;
mixer gate_output_11_185(.a(output_12_185), .b(output_12_10), .y(output_11_185));
wire output_13_185, output_13_10, output_12_185;
mixer gate_output_12_185(.a(output_13_185), .b(output_13_10), .y(output_12_185));
wire output_14_185, output_14_10, output_13_185;
mixer gate_output_13_185(.a(output_14_185), .b(output_14_10), .y(output_13_185));
wire output_15_185, output_15_10, output_14_185;
mixer gate_output_14_185(.a(output_15_185), .b(output_15_10), .y(output_14_185));
wire output_16_185, output_16_10, output_15_185;
mixer gate_output_15_185(.a(output_16_185), .b(output_16_10), .y(output_15_185));
wire output_1_186, output_1_11, output_0_186;
mixer gate_output_0_186(.a(output_1_186), .b(output_1_11), .y(output_0_186));
wire output_2_186, output_2_11, output_1_186;
mixer gate_output_1_186(.a(output_2_186), .b(output_2_11), .y(output_1_186));
wire output_3_186, output_3_11, output_2_186;
mixer gate_output_2_186(.a(output_3_186), .b(output_3_11), .y(output_2_186));
wire output_4_186, output_4_11, output_3_186;
mixer gate_output_3_186(.a(output_4_186), .b(output_4_11), .y(output_3_186));
wire output_5_186, output_5_11, output_4_186;
mixer gate_output_4_186(.a(output_5_186), .b(output_5_11), .y(output_4_186));
wire output_6_186, output_6_11, output_5_186;
mixer gate_output_5_186(.a(output_6_186), .b(output_6_11), .y(output_5_186));
wire output_7_186, output_7_11, output_6_186;
mixer gate_output_6_186(.a(output_7_186), .b(output_7_11), .y(output_6_186));
wire output_8_186, output_8_11, output_7_186;
mixer gate_output_7_186(.a(output_8_186), .b(output_8_11), .y(output_7_186));
wire output_9_186, output_9_11, output_8_186;
mixer gate_output_8_186(.a(output_9_186), .b(output_9_11), .y(output_8_186));
wire output_10_186, output_10_11, output_9_186;
mixer gate_output_9_186(.a(output_10_186), .b(output_10_11), .y(output_9_186));
wire output_11_186, output_11_11, output_10_186;
mixer gate_output_10_186(.a(output_11_186), .b(output_11_11), .y(output_10_186));
wire output_12_186, output_12_11, output_11_186;
mixer gate_output_11_186(.a(output_12_186), .b(output_12_11), .y(output_11_186));
wire output_13_186, output_13_11, output_12_186;
mixer gate_output_12_186(.a(output_13_186), .b(output_13_11), .y(output_12_186));
wire output_14_186, output_14_11, output_13_186;
mixer gate_output_13_186(.a(output_14_186), .b(output_14_11), .y(output_13_186));
wire output_15_186, output_15_11, output_14_186;
mixer gate_output_14_186(.a(output_15_186), .b(output_15_11), .y(output_14_186));
wire output_16_186, output_16_11, output_15_186;
mixer gate_output_15_186(.a(output_16_186), .b(output_16_11), .y(output_15_186));
wire output_1_187, output_1_12, output_0_187;
mixer gate_output_0_187(.a(output_1_187), .b(output_1_12), .y(output_0_187));
wire output_2_187, output_2_12, output_1_187;
mixer gate_output_1_187(.a(output_2_187), .b(output_2_12), .y(output_1_187));
wire output_3_187, output_3_12, output_2_187;
mixer gate_output_2_187(.a(output_3_187), .b(output_3_12), .y(output_2_187));
wire output_4_187, output_4_12, output_3_187;
mixer gate_output_3_187(.a(output_4_187), .b(output_4_12), .y(output_3_187));
wire output_5_187, output_5_12, output_4_187;
mixer gate_output_4_187(.a(output_5_187), .b(output_5_12), .y(output_4_187));
wire output_6_187, output_6_12, output_5_187;
mixer gate_output_5_187(.a(output_6_187), .b(output_6_12), .y(output_5_187));
wire output_7_187, output_7_12, output_6_187;
mixer gate_output_6_187(.a(output_7_187), .b(output_7_12), .y(output_6_187));
wire output_8_187, output_8_12, output_7_187;
mixer gate_output_7_187(.a(output_8_187), .b(output_8_12), .y(output_7_187));
wire output_9_187, output_9_12, output_8_187;
mixer gate_output_8_187(.a(output_9_187), .b(output_9_12), .y(output_8_187));
wire output_10_187, output_10_12, output_9_187;
mixer gate_output_9_187(.a(output_10_187), .b(output_10_12), .y(output_9_187));
wire output_11_187, output_11_12, output_10_187;
mixer gate_output_10_187(.a(output_11_187), .b(output_11_12), .y(output_10_187));
wire output_12_187, output_12_12, output_11_187;
mixer gate_output_11_187(.a(output_12_187), .b(output_12_12), .y(output_11_187));
wire output_13_187, output_13_12, output_12_187;
mixer gate_output_12_187(.a(output_13_187), .b(output_13_12), .y(output_12_187));
wire output_14_187, output_14_12, output_13_187;
mixer gate_output_13_187(.a(output_14_187), .b(output_14_12), .y(output_13_187));
wire output_15_187, output_15_12, output_14_187;
mixer gate_output_14_187(.a(output_15_187), .b(output_15_12), .y(output_14_187));
wire output_16_187, output_16_12, output_15_187;
mixer gate_output_15_187(.a(output_16_187), .b(output_16_12), .y(output_15_187));
wire output_1_188, output_1_13, output_0_188;
mixer gate_output_0_188(.a(output_1_188), .b(output_1_13), .y(output_0_188));
wire output_2_188, output_2_13, output_1_188;
mixer gate_output_1_188(.a(output_2_188), .b(output_2_13), .y(output_1_188));
wire output_3_188, output_3_13, output_2_188;
mixer gate_output_2_188(.a(output_3_188), .b(output_3_13), .y(output_2_188));
wire output_4_188, output_4_13, output_3_188;
mixer gate_output_3_188(.a(output_4_188), .b(output_4_13), .y(output_3_188));
wire output_5_188, output_5_13, output_4_188;
mixer gate_output_4_188(.a(output_5_188), .b(output_5_13), .y(output_4_188));
wire output_6_188, output_6_13, output_5_188;
mixer gate_output_5_188(.a(output_6_188), .b(output_6_13), .y(output_5_188));
wire output_7_188, output_7_13, output_6_188;
mixer gate_output_6_188(.a(output_7_188), .b(output_7_13), .y(output_6_188));
wire output_8_188, output_8_13, output_7_188;
mixer gate_output_7_188(.a(output_8_188), .b(output_8_13), .y(output_7_188));
wire output_9_188, output_9_13, output_8_188;
mixer gate_output_8_188(.a(output_9_188), .b(output_9_13), .y(output_8_188));
wire output_10_188, output_10_13, output_9_188;
mixer gate_output_9_188(.a(output_10_188), .b(output_10_13), .y(output_9_188));
wire output_11_188, output_11_13, output_10_188;
mixer gate_output_10_188(.a(output_11_188), .b(output_11_13), .y(output_10_188));
wire output_12_188, output_12_13, output_11_188;
mixer gate_output_11_188(.a(output_12_188), .b(output_12_13), .y(output_11_188));
wire output_13_188, output_13_13, output_12_188;
mixer gate_output_12_188(.a(output_13_188), .b(output_13_13), .y(output_12_188));
wire output_14_188, output_14_13, output_13_188;
mixer gate_output_13_188(.a(output_14_188), .b(output_14_13), .y(output_13_188));
wire output_15_188, output_15_13, output_14_188;
mixer gate_output_14_188(.a(output_15_188), .b(output_15_13), .y(output_14_188));
wire output_16_188, output_16_13, output_15_188;
mixer gate_output_15_188(.a(output_16_188), .b(output_16_13), .y(output_15_188));
wire output_1_189, output_1_14, output_0_189;
mixer gate_output_0_189(.a(output_1_189), .b(output_1_14), .y(output_0_189));
wire output_2_189, output_2_14, output_1_189;
mixer gate_output_1_189(.a(output_2_189), .b(output_2_14), .y(output_1_189));
wire output_3_189, output_3_14, output_2_189;
mixer gate_output_2_189(.a(output_3_189), .b(output_3_14), .y(output_2_189));
wire output_4_189, output_4_14, output_3_189;
mixer gate_output_3_189(.a(output_4_189), .b(output_4_14), .y(output_3_189));
wire output_5_189, output_5_14, output_4_189;
mixer gate_output_4_189(.a(output_5_189), .b(output_5_14), .y(output_4_189));
wire output_6_189, output_6_14, output_5_189;
mixer gate_output_5_189(.a(output_6_189), .b(output_6_14), .y(output_5_189));
wire output_7_189, output_7_14, output_6_189;
mixer gate_output_6_189(.a(output_7_189), .b(output_7_14), .y(output_6_189));
wire output_8_189, output_8_14, output_7_189;
mixer gate_output_7_189(.a(output_8_189), .b(output_8_14), .y(output_7_189));
wire output_9_189, output_9_14, output_8_189;
mixer gate_output_8_189(.a(output_9_189), .b(output_9_14), .y(output_8_189));
wire output_10_189, output_10_14, output_9_189;
mixer gate_output_9_189(.a(output_10_189), .b(output_10_14), .y(output_9_189));
wire output_11_189, output_11_14, output_10_189;
mixer gate_output_10_189(.a(output_11_189), .b(output_11_14), .y(output_10_189));
wire output_12_189, output_12_14, output_11_189;
mixer gate_output_11_189(.a(output_12_189), .b(output_12_14), .y(output_11_189));
wire output_13_189, output_13_14, output_12_189;
mixer gate_output_12_189(.a(output_13_189), .b(output_13_14), .y(output_12_189));
wire output_14_189, output_14_14, output_13_189;
mixer gate_output_13_189(.a(output_14_189), .b(output_14_14), .y(output_13_189));
wire output_15_189, output_15_14, output_14_189;
mixer gate_output_14_189(.a(output_15_189), .b(output_15_14), .y(output_14_189));
wire output_16_189, output_16_14, output_15_189;
mixer gate_output_15_189(.a(output_16_189), .b(output_16_14), .y(output_15_189));
wire output_1_190, output_1_15, output_0_190;
mixer gate_output_0_190(.a(output_1_190), .b(output_1_15), .y(output_0_190));
wire output_2_190, output_2_15, output_1_190;
mixer gate_output_1_190(.a(output_2_190), .b(output_2_15), .y(output_1_190));
wire output_3_190, output_3_15, output_2_190;
mixer gate_output_2_190(.a(output_3_190), .b(output_3_15), .y(output_2_190));
wire output_4_190, output_4_15, output_3_190;
mixer gate_output_3_190(.a(output_4_190), .b(output_4_15), .y(output_3_190));
wire output_5_190, output_5_15, output_4_190;
mixer gate_output_4_190(.a(output_5_190), .b(output_5_15), .y(output_4_190));
wire output_6_190, output_6_15, output_5_190;
mixer gate_output_5_190(.a(output_6_190), .b(output_6_15), .y(output_5_190));
wire output_7_190, output_7_15, output_6_190;
mixer gate_output_6_190(.a(output_7_190), .b(output_7_15), .y(output_6_190));
wire output_8_190, output_8_15, output_7_190;
mixer gate_output_7_190(.a(output_8_190), .b(output_8_15), .y(output_7_190));
wire output_9_190, output_9_15, output_8_190;
mixer gate_output_8_190(.a(output_9_190), .b(output_9_15), .y(output_8_190));
wire output_10_190, output_10_15, output_9_190;
mixer gate_output_9_190(.a(output_10_190), .b(output_10_15), .y(output_9_190));
wire output_11_190, output_11_15, output_10_190;
mixer gate_output_10_190(.a(output_11_190), .b(output_11_15), .y(output_10_190));
wire output_12_190, output_12_15, output_11_190;
mixer gate_output_11_190(.a(output_12_190), .b(output_12_15), .y(output_11_190));
wire output_13_190, output_13_15, output_12_190;
mixer gate_output_12_190(.a(output_13_190), .b(output_13_15), .y(output_12_190));
wire output_14_190, output_14_15, output_13_190;
mixer gate_output_13_190(.a(output_14_190), .b(output_14_15), .y(output_13_190));
wire output_15_190, output_15_15, output_14_190;
mixer gate_output_14_190(.a(output_15_190), .b(output_15_15), .y(output_14_190));
wire output_16_190, output_16_15, output_15_190;
mixer gate_output_15_190(.a(output_16_190), .b(output_16_15), .y(output_15_190));
wire output_1_191, output_1_0, output_0_191;
mixer gate_output_0_191(.a(output_1_191), .b(output_1_0), .y(output_0_191));
wire output_2_191, output_2_0, output_1_191;
mixer gate_output_1_191(.a(output_2_191), .b(output_2_0), .y(output_1_191));
wire output_3_191, output_3_0, output_2_191;
mixer gate_output_2_191(.a(output_3_191), .b(output_3_0), .y(output_2_191));
wire output_4_191, output_4_0, output_3_191;
mixer gate_output_3_191(.a(output_4_191), .b(output_4_0), .y(output_3_191));
wire output_5_191, output_5_0, output_4_191;
mixer gate_output_4_191(.a(output_5_191), .b(output_5_0), .y(output_4_191));
wire output_6_191, output_6_0, output_5_191;
mixer gate_output_5_191(.a(output_6_191), .b(output_6_0), .y(output_5_191));
wire output_7_191, output_7_0, output_6_191;
mixer gate_output_6_191(.a(output_7_191), .b(output_7_0), .y(output_6_191));
wire output_8_191, output_8_0, output_7_191;
mixer gate_output_7_191(.a(output_8_191), .b(output_8_0), .y(output_7_191));
wire output_9_191, output_9_0, output_8_191;
mixer gate_output_8_191(.a(output_9_191), .b(output_9_0), .y(output_8_191));
wire output_10_191, output_10_0, output_9_191;
mixer gate_output_9_191(.a(output_10_191), .b(output_10_0), .y(output_9_191));
wire output_11_191, output_11_0, output_10_191;
mixer gate_output_10_191(.a(output_11_191), .b(output_11_0), .y(output_10_191));
wire output_12_191, output_12_0, output_11_191;
mixer gate_output_11_191(.a(output_12_191), .b(output_12_0), .y(output_11_191));
wire output_13_191, output_13_0, output_12_191;
mixer gate_output_12_191(.a(output_13_191), .b(output_13_0), .y(output_12_191));
wire output_14_191, output_14_0, output_13_191;
mixer gate_output_13_191(.a(output_14_191), .b(output_14_0), .y(output_13_191));
wire output_15_191, output_15_0, output_14_191;
mixer gate_output_14_191(.a(output_15_191), .b(output_15_0), .y(output_14_191));
wire output_16_191, output_16_0, output_15_191;
mixer gate_output_15_191(.a(output_16_191), .b(output_16_0), .y(output_15_191));
wire output_1_192, output_1_1, output_0_192;
mixer gate_output_0_192(.a(output_1_192), .b(output_1_1), .y(output_0_192));
wire output_2_192, output_2_1, output_1_192;
mixer gate_output_1_192(.a(output_2_192), .b(output_2_1), .y(output_1_192));
wire output_3_192, output_3_1, output_2_192;
mixer gate_output_2_192(.a(output_3_192), .b(output_3_1), .y(output_2_192));
wire output_4_192, output_4_1, output_3_192;
mixer gate_output_3_192(.a(output_4_192), .b(output_4_1), .y(output_3_192));
wire output_5_192, output_5_1, output_4_192;
mixer gate_output_4_192(.a(output_5_192), .b(output_5_1), .y(output_4_192));
wire output_6_192, output_6_1, output_5_192;
mixer gate_output_5_192(.a(output_6_192), .b(output_6_1), .y(output_5_192));
wire output_7_192, output_7_1, output_6_192;
mixer gate_output_6_192(.a(output_7_192), .b(output_7_1), .y(output_6_192));
wire output_8_192, output_8_1, output_7_192;
mixer gate_output_7_192(.a(output_8_192), .b(output_8_1), .y(output_7_192));
wire output_9_192, output_9_1, output_8_192;
mixer gate_output_8_192(.a(output_9_192), .b(output_9_1), .y(output_8_192));
wire output_10_192, output_10_1, output_9_192;
mixer gate_output_9_192(.a(output_10_192), .b(output_10_1), .y(output_9_192));
wire output_11_192, output_11_1, output_10_192;
mixer gate_output_10_192(.a(output_11_192), .b(output_11_1), .y(output_10_192));
wire output_12_192, output_12_1, output_11_192;
mixer gate_output_11_192(.a(output_12_192), .b(output_12_1), .y(output_11_192));
wire output_13_192, output_13_1, output_12_192;
mixer gate_output_12_192(.a(output_13_192), .b(output_13_1), .y(output_12_192));
wire output_14_192, output_14_1, output_13_192;
mixer gate_output_13_192(.a(output_14_192), .b(output_14_1), .y(output_13_192));
wire output_15_192, output_15_1, output_14_192;
mixer gate_output_14_192(.a(output_15_192), .b(output_15_1), .y(output_14_192));
wire output_16_192, output_16_1, output_15_192;
mixer gate_output_15_192(.a(output_16_192), .b(output_16_1), .y(output_15_192));
wire output_1_193, output_1_2, output_0_193;
mixer gate_output_0_193(.a(output_1_193), .b(output_1_2), .y(output_0_193));
wire output_2_193, output_2_2, output_1_193;
mixer gate_output_1_193(.a(output_2_193), .b(output_2_2), .y(output_1_193));
wire output_3_193, output_3_2, output_2_193;
mixer gate_output_2_193(.a(output_3_193), .b(output_3_2), .y(output_2_193));
wire output_4_193, output_4_2, output_3_193;
mixer gate_output_3_193(.a(output_4_193), .b(output_4_2), .y(output_3_193));
wire output_5_193, output_5_2, output_4_193;
mixer gate_output_4_193(.a(output_5_193), .b(output_5_2), .y(output_4_193));
wire output_6_193, output_6_2, output_5_193;
mixer gate_output_5_193(.a(output_6_193), .b(output_6_2), .y(output_5_193));
wire output_7_193, output_7_2, output_6_193;
mixer gate_output_6_193(.a(output_7_193), .b(output_7_2), .y(output_6_193));
wire output_8_193, output_8_2, output_7_193;
mixer gate_output_7_193(.a(output_8_193), .b(output_8_2), .y(output_7_193));
wire output_9_193, output_9_2, output_8_193;
mixer gate_output_8_193(.a(output_9_193), .b(output_9_2), .y(output_8_193));
wire output_10_193, output_10_2, output_9_193;
mixer gate_output_9_193(.a(output_10_193), .b(output_10_2), .y(output_9_193));
wire output_11_193, output_11_2, output_10_193;
mixer gate_output_10_193(.a(output_11_193), .b(output_11_2), .y(output_10_193));
wire output_12_193, output_12_2, output_11_193;
mixer gate_output_11_193(.a(output_12_193), .b(output_12_2), .y(output_11_193));
wire output_13_193, output_13_2, output_12_193;
mixer gate_output_12_193(.a(output_13_193), .b(output_13_2), .y(output_12_193));
wire output_14_193, output_14_2, output_13_193;
mixer gate_output_13_193(.a(output_14_193), .b(output_14_2), .y(output_13_193));
wire output_15_193, output_15_2, output_14_193;
mixer gate_output_14_193(.a(output_15_193), .b(output_15_2), .y(output_14_193));
wire output_16_193, output_16_2, output_15_193;
mixer gate_output_15_193(.a(output_16_193), .b(output_16_2), .y(output_15_193));
wire output_1_194, output_1_3, output_0_194;
mixer gate_output_0_194(.a(output_1_194), .b(output_1_3), .y(output_0_194));
wire output_2_194, output_2_3, output_1_194;
mixer gate_output_1_194(.a(output_2_194), .b(output_2_3), .y(output_1_194));
wire output_3_194, output_3_3, output_2_194;
mixer gate_output_2_194(.a(output_3_194), .b(output_3_3), .y(output_2_194));
wire output_4_194, output_4_3, output_3_194;
mixer gate_output_3_194(.a(output_4_194), .b(output_4_3), .y(output_3_194));
wire output_5_194, output_5_3, output_4_194;
mixer gate_output_4_194(.a(output_5_194), .b(output_5_3), .y(output_4_194));
wire output_6_194, output_6_3, output_5_194;
mixer gate_output_5_194(.a(output_6_194), .b(output_6_3), .y(output_5_194));
wire output_7_194, output_7_3, output_6_194;
mixer gate_output_6_194(.a(output_7_194), .b(output_7_3), .y(output_6_194));
wire output_8_194, output_8_3, output_7_194;
mixer gate_output_7_194(.a(output_8_194), .b(output_8_3), .y(output_7_194));
wire output_9_194, output_9_3, output_8_194;
mixer gate_output_8_194(.a(output_9_194), .b(output_9_3), .y(output_8_194));
wire output_10_194, output_10_3, output_9_194;
mixer gate_output_9_194(.a(output_10_194), .b(output_10_3), .y(output_9_194));
wire output_11_194, output_11_3, output_10_194;
mixer gate_output_10_194(.a(output_11_194), .b(output_11_3), .y(output_10_194));
wire output_12_194, output_12_3, output_11_194;
mixer gate_output_11_194(.a(output_12_194), .b(output_12_3), .y(output_11_194));
wire output_13_194, output_13_3, output_12_194;
mixer gate_output_12_194(.a(output_13_194), .b(output_13_3), .y(output_12_194));
wire output_14_194, output_14_3, output_13_194;
mixer gate_output_13_194(.a(output_14_194), .b(output_14_3), .y(output_13_194));
wire output_15_194, output_15_3, output_14_194;
mixer gate_output_14_194(.a(output_15_194), .b(output_15_3), .y(output_14_194));
wire output_16_194, output_16_3, output_15_194;
mixer gate_output_15_194(.a(output_16_194), .b(output_16_3), .y(output_15_194));
wire output_1_195, output_1_4, output_0_195;
mixer gate_output_0_195(.a(output_1_195), .b(output_1_4), .y(output_0_195));
wire output_2_195, output_2_4, output_1_195;
mixer gate_output_1_195(.a(output_2_195), .b(output_2_4), .y(output_1_195));
wire output_3_195, output_3_4, output_2_195;
mixer gate_output_2_195(.a(output_3_195), .b(output_3_4), .y(output_2_195));
wire output_4_195, output_4_4, output_3_195;
mixer gate_output_3_195(.a(output_4_195), .b(output_4_4), .y(output_3_195));
wire output_5_195, output_5_4, output_4_195;
mixer gate_output_4_195(.a(output_5_195), .b(output_5_4), .y(output_4_195));
wire output_6_195, output_6_4, output_5_195;
mixer gate_output_5_195(.a(output_6_195), .b(output_6_4), .y(output_5_195));
wire output_7_195, output_7_4, output_6_195;
mixer gate_output_6_195(.a(output_7_195), .b(output_7_4), .y(output_6_195));
wire output_8_195, output_8_4, output_7_195;
mixer gate_output_7_195(.a(output_8_195), .b(output_8_4), .y(output_7_195));
wire output_9_195, output_9_4, output_8_195;
mixer gate_output_8_195(.a(output_9_195), .b(output_9_4), .y(output_8_195));
wire output_10_195, output_10_4, output_9_195;
mixer gate_output_9_195(.a(output_10_195), .b(output_10_4), .y(output_9_195));
wire output_11_195, output_11_4, output_10_195;
mixer gate_output_10_195(.a(output_11_195), .b(output_11_4), .y(output_10_195));
wire output_12_195, output_12_4, output_11_195;
mixer gate_output_11_195(.a(output_12_195), .b(output_12_4), .y(output_11_195));
wire output_13_195, output_13_4, output_12_195;
mixer gate_output_12_195(.a(output_13_195), .b(output_13_4), .y(output_12_195));
wire output_14_195, output_14_4, output_13_195;
mixer gate_output_13_195(.a(output_14_195), .b(output_14_4), .y(output_13_195));
wire output_15_195, output_15_4, output_14_195;
mixer gate_output_14_195(.a(output_15_195), .b(output_15_4), .y(output_14_195));
wire output_16_195, output_16_4, output_15_195;
mixer gate_output_15_195(.a(output_16_195), .b(output_16_4), .y(output_15_195));
wire output_1_196, output_1_5, output_0_196;
mixer gate_output_0_196(.a(output_1_196), .b(output_1_5), .y(output_0_196));
wire output_2_196, output_2_5, output_1_196;
mixer gate_output_1_196(.a(output_2_196), .b(output_2_5), .y(output_1_196));
wire output_3_196, output_3_5, output_2_196;
mixer gate_output_2_196(.a(output_3_196), .b(output_3_5), .y(output_2_196));
wire output_4_196, output_4_5, output_3_196;
mixer gate_output_3_196(.a(output_4_196), .b(output_4_5), .y(output_3_196));
wire output_5_196, output_5_5, output_4_196;
mixer gate_output_4_196(.a(output_5_196), .b(output_5_5), .y(output_4_196));
wire output_6_196, output_6_5, output_5_196;
mixer gate_output_5_196(.a(output_6_196), .b(output_6_5), .y(output_5_196));
wire output_7_196, output_7_5, output_6_196;
mixer gate_output_6_196(.a(output_7_196), .b(output_7_5), .y(output_6_196));
wire output_8_196, output_8_5, output_7_196;
mixer gate_output_7_196(.a(output_8_196), .b(output_8_5), .y(output_7_196));
wire output_9_196, output_9_5, output_8_196;
mixer gate_output_8_196(.a(output_9_196), .b(output_9_5), .y(output_8_196));
wire output_10_196, output_10_5, output_9_196;
mixer gate_output_9_196(.a(output_10_196), .b(output_10_5), .y(output_9_196));
wire output_11_196, output_11_5, output_10_196;
mixer gate_output_10_196(.a(output_11_196), .b(output_11_5), .y(output_10_196));
wire output_12_196, output_12_5, output_11_196;
mixer gate_output_11_196(.a(output_12_196), .b(output_12_5), .y(output_11_196));
wire output_13_196, output_13_5, output_12_196;
mixer gate_output_12_196(.a(output_13_196), .b(output_13_5), .y(output_12_196));
wire output_14_196, output_14_5, output_13_196;
mixer gate_output_13_196(.a(output_14_196), .b(output_14_5), .y(output_13_196));
wire output_15_196, output_15_5, output_14_196;
mixer gate_output_14_196(.a(output_15_196), .b(output_15_5), .y(output_14_196));
wire output_16_196, output_16_5, output_15_196;
mixer gate_output_15_196(.a(output_16_196), .b(output_16_5), .y(output_15_196));
wire output_1_197, output_1_6, output_0_197;
mixer gate_output_0_197(.a(output_1_197), .b(output_1_6), .y(output_0_197));
wire output_2_197, output_2_6, output_1_197;
mixer gate_output_1_197(.a(output_2_197), .b(output_2_6), .y(output_1_197));
wire output_3_197, output_3_6, output_2_197;
mixer gate_output_2_197(.a(output_3_197), .b(output_3_6), .y(output_2_197));
wire output_4_197, output_4_6, output_3_197;
mixer gate_output_3_197(.a(output_4_197), .b(output_4_6), .y(output_3_197));
wire output_5_197, output_5_6, output_4_197;
mixer gate_output_4_197(.a(output_5_197), .b(output_5_6), .y(output_4_197));
wire output_6_197, output_6_6, output_5_197;
mixer gate_output_5_197(.a(output_6_197), .b(output_6_6), .y(output_5_197));
wire output_7_197, output_7_6, output_6_197;
mixer gate_output_6_197(.a(output_7_197), .b(output_7_6), .y(output_6_197));
wire output_8_197, output_8_6, output_7_197;
mixer gate_output_7_197(.a(output_8_197), .b(output_8_6), .y(output_7_197));
wire output_9_197, output_9_6, output_8_197;
mixer gate_output_8_197(.a(output_9_197), .b(output_9_6), .y(output_8_197));
wire output_10_197, output_10_6, output_9_197;
mixer gate_output_9_197(.a(output_10_197), .b(output_10_6), .y(output_9_197));
wire output_11_197, output_11_6, output_10_197;
mixer gate_output_10_197(.a(output_11_197), .b(output_11_6), .y(output_10_197));
wire output_12_197, output_12_6, output_11_197;
mixer gate_output_11_197(.a(output_12_197), .b(output_12_6), .y(output_11_197));
wire output_13_197, output_13_6, output_12_197;
mixer gate_output_12_197(.a(output_13_197), .b(output_13_6), .y(output_12_197));
wire output_14_197, output_14_6, output_13_197;
mixer gate_output_13_197(.a(output_14_197), .b(output_14_6), .y(output_13_197));
wire output_15_197, output_15_6, output_14_197;
mixer gate_output_14_197(.a(output_15_197), .b(output_15_6), .y(output_14_197));
wire output_16_197, output_16_6, output_15_197;
mixer gate_output_15_197(.a(output_16_197), .b(output_16_6), .y(output_15_197));
wire output_1_198, output_1_7, output_0_198;
mixer gate_output_0_198(.a(output_1_198), .b(output_1_7), .y(output_0_198));
wire output_2_198, output_2_7, output_1_198;
mixer gate_output_1_198(.a(output_2_198), .b(output_2_7), .y(output_1_198));
wire output_3_198, output_3_7, output_2_198;
mixer gate_output_2_198(.a(output_3_198), .b(output_3_7), .y(output_2_198));
wire output_4_198, output_4_7, output_3_198;
mixer gate_output_3_198(.a(output_4_198), .b(output_4_7), .y(output_3_198));
wire output_5_198, output_5_7, output_4_198;
mixer gate_output_4_198(.a(output_5_198), .b(output_5_7), .y(output_4_198));
wire output_6_198, output_6_7, output_5_198;
mixer gate_output_5_198(.a(output_6_198), .b(output_6_7), .y(output_5_198));
wire output_7_198, output_7_7, output_6_198;
mixer gate_output_6_198(.a(output_7_198), .b(output_7_7), .y(output_6_198));
wire output_8_198, output_8_7, output_7_198;
mixer gate_output_7_198(.a(output_8_198), .b(output_8_7), .y(output_7_198));
wire output_9_198, output_9_7, output_8_198;
mixer gate_output_8_198(.a(output_9_198), .b(output_9_7), .y(output_8_198));
wire output_10_198, output_10_7, output_9_198;
mixer gate_output_9_198(.a(output_10_198), .b(output_10_7), .y(output_9_198));
wire output_11_198, output_11_7, output_10_198;
mixer gate_output_10_198(.a(output_11_198), .b(output_11_7), .y(output_10_198));
wire output_12_198, output_12_7, output_11_198;
mixer gate_output_11_198(.a(output_12_198), .b(output_12_7), .y(output_11_198));
wire output_13_198, output_13_7, output_12_198;
mixer gate_output_12_198(.a(output_13_198), .b(output_13_7), .y(output_12_198));
wire output_14_198, output_14_7, output_13_198;
mixer gate_output_13_198(.a(output_14_198), .b(output_14_7), .y(output_13_198));
wire output_15_198, output_15_7, output_14_198;
mixer gate_output_14_198(.a(output_15_198), .b(output_15_7), .y(output_14_198));
wire output_16_198, output_16_7, output_15_198;
mixer gate_output_15_198(.a(output_16_198), .b(output_16_7), .y(output_15_198));
wire output_1_199, output_1_8, output_0_199;
mixer gate_output_0_199(.a(output_1_199), .b(output_1_8), .y(output_0_199));
wire output_2_199, output_2_8, output_1_199;
mixer gate_output_1_199(.a(output_2_199), .b(output_2_8), .y(output_1_199));
wire output_3_199, output_3_8, output_2_199;
mixer gate_output_2_199(.a(output_3_199), .b(output_3_8), .y(output_2_199));
wire output_4_199, output_4_8, output_3_199;
mixer gate_output_3_199(.a(output_4_199), .b(output_4_8), .y(output_3_199));
wire output_5_199, output_5_8, output_4_199;
mixer gate_output_4_199(.a(output_5_199), .b(output_5_8), .y(output_4_199));
wire output_6_199, output_6_8, output_5_199;
mixer gate_output_5_199(.a(output_6_199), .b(output_6_8), .y(output_5_199));
wire output_7_199, output_7_8, output_6_199;
mixer gate_output_6_199(.a(output_7_199), .b(output_7_8), .y(output_6_199));
wire output_8_199, output_8_8, output_7_199;
mixer gate_output_7_199(.a(output_8_199), .b(output_8_8), .y(output_7_199));
wire output_9_199, output_9_8, output_8_199;
mixer gate_output_8_199(.a(output_9_199), .b(output_9_8), .y(output_8_199));
wire output_10_199, output_10_8, output_9_199;
mixer gate_output_9_199(.a(output_10_199), .b(output_10_8), .y(output_9_199));
wire output_11_199, output_11_8, output_10_199;
mixer gate_output_10_199(.a(output_11_199), .b(output_11_8), .y(output_10_199));
wire output_12_199, output_12_8, output_11_199;
mixer gate_output_11_199(.a(output_12_199), .b(output_12_8), .y(output_11_199));
wire output_13_199, output_13_8, output_12_199;
mixer gate_output_12_199(.a(output_13_199), .b(output_13_8), .y(output_12_199));
wire output_14_199, output_14_8, output_13_199;
mixer gate_output_13_199(.a(output_14_199), .b(output_14_8), .y(output_13_199));
wire output_15_199, output_15_8, output_14_199;
mixer gate_output_14_199(.a(output_15_199), .b(output_15_8), .y(output_14_199));
wire output_16_199, output_16_8, output_15_199;
mixer gate_output_15_199(.a(output_16_199), .b(output_16_8), .y(output_15_199));
wire output_1_200, output_1_9, output_0_200;
mixer gate_output_0_200(.a(output_1_200), .b(output_1_9), .y(output_0_200));
wire output_2_200, output_2_9, output_1_200;
mixer gate_output_1_200(.a(output_2_200), .b(output_2_9), .y(output_1_200));
wire output_3_200, output_3_9, output_2_200;
mixer gate_output_2_200(.a(output_3_200), .b(output_3_9), .y(output_2_200));
wire output_4_200, output_4_9, output_3_200;
mixer gate_output_3_200(.a(output_4_200), .b(output_4_9), .y(output_3_200));
wire output_5_200, output_5_9, output_4_200;
mixer gate_output_4_200(.a(output_5_200), .b(output_5_9), .y(output_4_200));
wire output_6_200, output_6_9, output_5_200;
mixer gate_output_5_200(.a(output_6_200), .b(output_6_9), .y(output_5_200));
wire output_7_200, output_7_9, output_6_200;
mixer gate_output_6_200(.a(output_7_200), .b(output_7_9), .y(output_6_200));
wire output_8_200, output_8_9, output_7_200;
mixer gate_output_7_200(.a(output_8_200), .b(output_8_9), .y(output_7_200));
wire output_9_200, output_9_9, output_8_200;
mixer gate_output_8_200(.a(output_9_200), .b(output_9_9), .y(output_8_200));
wire output_10_200, output_10_9, output_9_200;
mixer gate_output_9_200(.a(output_10_200), .b(output_10_9), .y(output_9_200));
wire output_11_200, output_11_9, output_10_200;
mixer gate_output_10_200(.a(output_11_200), .b(output_11_9), .y(output_10_200));
wire output_12_200, output_12_9, output_11_200;
mixer gate_output_11_200(.a(output_12_200), .b(output_12_9), .y(output_11_200));
wire output_13_200, output_13_9, output_12_200;
mixer gate_output_12_200(.a(output_13_200), .b(output_13_9), .y(output_12_200));
wire output_14_200, output_14_9, output_13_200;
mixer gate_output_13_200(.a(output_14_200), .b(output_14_9), .y(output_13_200));
wire output_15_200, output_15_9, output_14_200;
mixer gate_output_14_200(.a(output_15_200), .b(output_15_9), .y(output_14_200));
wire output_16_200, output_16_9, output_15_200;
mixer gate_output_15_200(.a(output_16_200), .b(output_16_9), .y(output_15_200));
wire output_1_201, output_1_10, output_0_201;
mixer gate_output_0_201(.a(output_1_201), .b(output_1_10), .y(output_0_201));
wire output_2_201, output_2_10, output_1_201;
mixer gate_output_1_201(.a(output_2_201), .b(output_2_10), .y(output_1_201));
wire output_3_201, output_3_10, output_2_201;
mixer gate_output_2_201(.a(output_3_201), .b(output_3_10), .y(output_2_201));
wire output_4_201, output_4_10, output_3_201;
mixer gate_output_3_201(.a(output_4_201), .b(output_4_10), .y(output_3_201));
wire output_5_201, output_5_10, output_4_201;
mixer gate_output_4_201(.a(output_5_201), .b(output_5_10), .y(output_4_201));
wire output_6_201, output_6_10, output_5_201;
mixer gate_output_5_201(.a(output_6_201), .b(output_6_10), .y(output_5_201));
wire output_7_201, output_7_10, output_6_201;
mixer gate_output_6_201(.a(output_7_201), .b(output_7_10), .y(output_6_201));
wire output_8_201, output_8_10, output_7_201;
mixer gate_output_7_201(.a(output_8_201), .b(output_8_10), .y(output_7_201));
wire output_9_201, output_9_10, output_8_201;
mixer gate_output_8_201(.a(output_9_201), .b(output_9_10), .y(output_8_201));
wire output_10_201, output_10_10, output_9_201;
mixer gate_output_9_201(.a(output_10_201), .b(output_10_10), .y(output_9_201));
wire output_11_201, output_11_10, output_10_201;
mixer gate_output_10_201(.a(output_11_201), .b(output_11_10), .y(output_10_201));
wire output_12_201, output_12_10, output_11_201;
mixer gate_output_11_201(.a(output_12_201), .b(output_12_10), .y(output_11_201));
wire output_13_201, output_13_10, output_12_201;
mixer gate_output_12_201(.a(output_13_201), .b(output_13_10), .y(output_12_201));
wire output_14_201, output_14_10, output_13_201;
mixer gate_output_13_201(.a(output_14_201), .b(output_14_10), .y(output_13_201));
wire output_15_201, output_15_10, output_14_201;
mixer gate_output_14_201(.a(output_15_201), .b(output_15_10), .y(output_14_201));
wire output_16_201, output_16_10, output_15_201;
mixer gate_output_15_201(.a(output_16_201), .b(output_16_10), .y(output_15_201));
wire output_1_202, output_1_11, output_0_202;
mixer gate_output_0_202(.a(output_1_202), .b(output_1_11), .y(output_0_202));
wire output_2_202, output_2_11, output_1_202;
mixer gate_output_1_202(.a(output_2_202), .b(output_2_11), .y(output_1_202));
wire output_3_202, output_3_11, output_2_202;
mixer gate_output_2_202(.a(output_3_202), .b(output_3_11), .y(output_2_202));
wire output_4_202, output_4_11, output_3_202;
mixer gate_output_3_202(.a(output_4_202), .b(output_4_11), .y(output_3_202));
wire output_5_202, output_5_11, output_4_202;
mixer gate_output_4_202(.a(output_5_202), .b(output_5_11), .y(output_4_202));
wire output_6_202, output_6_11, output_5_202;
mixer gate_output_5_202(.a(output_6_202), .b(output_6_11), .y(output_5_202));
wire output_7_202, output_7_11, output_6_202;
mixer gate_output_6_202(.a(output_7_202), .b(output_7_11), .y(output_6_202));
wire output_8_202, output_8_11, output_7_202;
mixer gate_output_7_202(.a(output_8_202), .b(output_8_11), .y(output_7_202));
wire output_9_202, output_9_11, output_8_202;
mixer gate_output_8_202(.a(output_9_202), .b(output_9_11), .y(output_8_202));
wire output_10_202, output_10_11, output_9_202;
mixer gate_output_9_202(.a(output_10_202), .b(output_10_11), .y(output_9_202));
wire output_11_202, output_11_11, output_10_202;
mixer gate_output_10_202(.a(output_11_202), .b(output_11_11), .y(output_10_202));
wire output_12_202, output_12_11, output_11_202;
mixer gate_output_11_202(.a(output_12_202), .b(output_12_11), .y(output_11_202));
wire output_13_202, output_13_11, output_12_202;
mixer gate_output_12_202(.a(output_13_202), .b(output_13_11), .y(output_12_202));
wire output_14_202, output_14_11, output_13_202;
mixer gate_output_13_202(.a(output_14_202), .b(output_14_11), .y(output_13_202));
wire output_15_202, output_15_11, output_14_202;
mixer gate_output_14_202(.a(output_15_202), .b(output_15_11), .y(output_14_202));
wire output_16_202, output_16_11, output_15_202;
mixer gate_output_15_202(.a(output_16_202), .b(output_16_11), .y(output_15_202));
wire output_1_203, output_1_12, output_0_203;
mixer gate_output_0_203(.a(output_1_203), .b(output_1_12), .y(output_0_203));
wire output_2_203, output_2_12, output_1_203;
mixer gate_output_1_203(.a(output_2_203), .b(output_2_12), .y(output_1_203));
wire output_3_203, output_3_12, output_2_203;
mixer gate_output_2_203(.a(output_3_203), .b(output_3_12), .y(output_2_203));
wire output_4_203, output_4_12, output_3_203;
mixer gate_output_3_203(.a(output_4_203), .b(output_4_12), .y(output_3_203));
wire output_5_203, output_5_12, output_4_203;
mixer gate_output_4_203(.a(output_5_203), .b(output_5_12), .y(output_4_203));
wire output_6_203, output_6_12, output_5_203;
mixer gate_output_5_203(.a(output_6_203), .b(output_6_12), .y(output_5_203));
wire output_7_203, output_7_12, output_6_203;
mixer gate_output_6_203(.a(output_7_203), .b(output_7_12), .y(output_6_203));
wire output_8_203, output_8_12, output_7_203;
mixer gate_output_7_203(.a(output_8_203), .b(output_8_12), .y(output_7_203));
wire output_9_203, output_9_12, output_8_203;
mixer gate_output_8_203(.a(output_9_203), .b(output_9_12), .y(output_8_203));
wire output_10_203, output_10_12, output_9_203;
mixer gate_output_9_203(.a(output_10_203), .b(output_10_12), .y(output_9_203));
wire output_11_203, output_11_12, output_10_203;
mixer gate_output_10_203(.a(output_11_203), .b(output_11_12), .y(output_10_203));
wire output_12_203, output_12_12, output_11_203;
mixer gate_output_11_203(.a(output_12_203), .b(output_12_12), .y(output_11_203));
wire output_13_203, output_13_12, output_12_203;
mixer gate_output_12_203(.a(output_13_203), .b(output_13_12), .y(output_12_203));
wire output_14_203, output_14_12, output_13_203;
mixer gate_output_13_203(.a(output_14_203), .b(output_14_12), .y(output_13_203));
wire output_15_203, output_15_12, output_14_203;
mixer gate_output_14_203(.a(output_15_203), .b(output_15_12), .y(output_14_203));
wire output_16_203, output_16_12, output_15_203;
mixer gate_output_15_203(.a(output_16_203), .b(output_16_12), .y(output_15_203));
wire output_1_204, output_1_13, output_0_204;
mixer gate_output_0_204(.a(output_1_204), .b(output_1_13), .y(output_0_204));
wire output_2_204, output_2_13, output_1_204;
mixer gate_output_1_204(.a(output_2_204), .b(output_2_13), .y(output_1_204));
wire output_3_204, output_3_13, output_2_204;
mixer gate_output_2_204(.a(output_3_204), .b(output_3_13), .y(output_2_204));
wire output_4_204, output_4_13, output_3_204;
mixer gate_output_3_204(.a(output_4_204), .b(output_4_13), .y(output_3_204));
wire output_5_204, output_5_13, output_4_204;
mixer gate_output_4_204(.a(output_5_204), .b(output_5_13), .y(output_4_204));
wire output_6_204, output_6_13, output_5_204;
mixer gate_output_5_204(.a(output_6_204), .b(output_6_13), .y(output_5_204));
wire output_7_204, output_7_13, output_6_204;
mixer gate_output_6_204(.a(output_7_204), .b(output_7_13), .y(output_6_204));
wire output_8_204, output_8_13, output_7_204;
mixer gate_output_7_204(.a(output_8_204), .b(output_8_13), .y(output_7_204));
wire output_9_204, output_9_13, output_8_204;
mixer gate_output_8_204(.a(output_9_204), .b(output_9_13), .y(output_8_204));
wire output_10_204, output_10_13, output_9_204;
mixer gate_output_9_204(.a(output_10_204), .b(output_10_13), .y(output_9_204));
wire output_11_204, output_11_13, output_10_204;
mixer gate_output_10_204(.a(output_11_204), .b(output_11_13), .y(output_10_204));
wire output_12_204, output_12_13, output_11_204;
mixer gate_output_11_204(.a(output_12_204), .b(output_12_13), .y(output_11_204));
wire output_13_204, output_13_13, output_12_204;
mixer gate_output_12_204(.a(output_13_204), .b(output_13_13), .y(output_12_204));
wire output_14_204, output_14_13, output_13_204;
mixer gate_output_13_204(.a(output_14_204), .b(output_14_13), .y(output_13_204));
wire output_15_204, output_15_13, output_14_204;
mixer gate_output_14_204(.a(output_15_204), .b(output_15_13), .y(output_14_204));
wire output_16_204, output_16_13, output_15_204;
mixer gate_output_15_204(.a(output_16_204), .b(output_16_13), .y(output_15_204));
wire output_1_205, output_1_14, output_0_205;
mixer gate_output_0_205(.a(output_1_205), .b(output_1_14), .y(output_0_205));
wire output_2_205, output_2_14, output_1_205;
mixer gate_output_1_205(.a(output_2_205), .b(output_2_14), .y(output_1_205));
wire output_3_205, output_3_14, output_2_205;
mixer gate_output_2_205(.a(output_3_205), .b(output_3_14), .y(output_2_205));
wire output_4_205, output_4_14, output_3_205;
mixer gate_output_3_205(.a(output_4_205), .b(output_4_14), .y(output_3_205));
wire output_5_205, output_5_14, output_4_205;
mixer gate_output_4_205(.a(output_5_205), .b(output_5_14), .y(output_4_205));
wire output_6_205, output_6_14, output_5_205;
mixer gate_output_5_205(.a(output_6_205), .b(output_6_14), .y(output_5_205));
wire output_7_205, output_7_14, output_6_205;
mixer gate_output_6_205(.a(output_7_205), .b(output_7_14), .y(output_6_205));
wire output_8_205, output_8_14, output_7_205;
mixer gate_output_7_205(.a(output_8_205), .b(output_8_14), .y(output_7_205));
wire output_9_205, output_9_14, output_8_205;
mixer gate_output_8_205(.a(output_9_205), .b(output_9_14), .y(output_8_205));
wire output_10_205, output_10_14, output_9_205;
mixer gate_output_9_205(.a(output_10_205), .b(output_10_14), .y(output_9_205));
wire output_11_205, output_11_14, output_10_205;
mixer gate_output_10_205(.a(output_11_205), .b(output_11_14), .y(output_10_205));
wire output_12_205, output_12_14, output_11_205;
mixer gate_output_11_205(.a(output_12_205), .b(output_12_14), .y(output_11_205));
wire output_13_205, output_13_14, output_12_205;
mixer gate_output_12_205(.a(output_13_205), .b(output_13_14), .y(output_12_205));
wire output_14_205, output_14_14, output_13_205;
mixer gate_output_13_205(.a(output_14_205), .b(output_14_14), .y(output_13_205));
wire output_15_205, output_15_14, output_14_205;
mixer gate_output_14_205(.a(output_15_205), .b(output_15_14), .y(output_14_205));
wire output_16_205, output_16_14, output_15_205;
mixer gate_output_15_205(.a(output_16_205), .b(output_16_14), .y(output_15_205));
wire output_1_206, output_1_15, output_0_206;
mixer gate_output_0_206(.a(output_1_206), .b(output_1_15), .y(output_0_206));
wire output_2_206, output_2_15, output_1_206;
mixer gate_output_1_206(.a(output_2_206), .b(output_2_15), .y(output_1_206));
wire output_3_206, output_3_15, output_2_206;
mixer gate_output_2_206(.a(output_3_206), .b(output_3_15), .y(output_2_206));
wire output_4_206, output_4_15, output_3_206;
mixer gate_output_3_206(.a(output_4_206), .b(output_4_15), .y(output_3_206));
wire output_5_206, output_5_15, output_4_206;
mixer gate_output_4_206(.a(output_5_206), .b(output_5_15), .y(output_4_206));
wire output_6_206, output_6_15, output_5_206;
mixer gate_output_5_206(.a(output_6_206), .b(output_6_15), .y(output_5_206));
wire output_7_206, output_7_15, output_6_206;
mixer gate_output_6_206(.a(output_7_206), .b(output_7_15), .y(output_6_206));
wire output_8_206, output_8_15, output_7_206;
mixer gate_output_7_206(.a(output_8_206), .b(output_8_15), .y(output_7_206));
wire output_9_206, output_9_15, output_8_206;
mixer gate_output_8_206(.a(output_9_206), .b(output_9_15), .y(output_8_206));
wire output_10_206, output_10_15, output_9_206;
mixer gate_output_9_206(.a(output_10_206), .b(output_10_15), .y(output_9_206));
wire output_11_206, output_11_15, output_10_206;
mixer gate_output_10_206(.a(output_11_206), .b(output_11_15), .y(output_10_206));
wire output_12_206, output_12_15, output_11_206;
mixer gate_output_11_206(.a(output_12_206), .b(output_12_15), .y(output_11_206));
wire output_13_206, output_13_15, output_12_206;
mixer gate_output_12_206(.a(output_13_206), .b(output_13_15), .y(output_12_206));
wire output_14_206, output_14_15, output_13_206;
mixer gate_output_13_206(.a(output_14_206), .b(output_14_15), .y(output_13_206));
wire output_15_206, output_15_15, output_14_206;
mixer gate_output_14_206(.a(output_15_206), .b(output_15_15), .y(output_14_206));
wire output_16_206, output_16_15, output_15_206;
mixer gate_output_15_206(.a(output_16_206), .b(output_16_15), .y(output_15_206));
wire output_1_207, output_1_0, output_0_207;
mixer gate_output_0_207(.a(output_1_207), .b(output_1_0), .y(output_0_207));
wire output_2_207, output_2_0, output_1_207;
mixer gate_output_1_207(.a(output_2_207), .b(output_2_0), .y(output_1_207));
wire output_3_207, output_3_0, output_2_207;
mixer gate_output_2_207(.a(output_3_207), .b(output_3_0), .y(output_2_207));
wire output_4_207, output_4_0, output_3_207;
mixer gate_output_3_207(.a(output_4_207), .b(output_4_0), .y(output_3_207));
wire output_5_207, output_5_0, output_4_207;
mixer gate_output_4_207(.a(output_5_207), .b(output_5_0), .y(output_4_207));
wire output_6_207, output_6_0, output_5_207;
mixer gate_output_5_207(.a(output_6_207), .b(output_6_0), .y(output_5_207));
wire output_7_207, output_7_0, output_6_207;
mixer gate_output_6_207(.a(output_7_207), .b(output_7_0), .y(output_6_207));
wire output_8_207, output_8_0, output_7_207;
mixer gate_output_7_207(.a(output_8_207), .b(output_8_0), .y(output_7_207));
wire output_9_207, output_9_0, output_8_207;
mixer gate_output_8_207(.a(output_9_207), .b(output_9_0), .y(output_8_207));
wire output_10_207, output_10_0, output_9_207;
mixer gate_output_9_207(.a(output_10_207), .b(output_10_0), .y(output_9_207));
wire output_11_207, output_11_0, output_10_207;
mixer gate_output_10_207(.a(output_11_207), .b(output_11_0), .y(output_10_207));
wire output_12_207, output_12_0, output_11_207;
mixer gate_output_11_207(.a(output_12_207), .b(output_12_0), .y(output_11_207));
wire output_13_207, output_13_0, output_12_207;
mixer gate_output_12_207(.a(output_13_207), .b(output_13_0), .y(output_12_207));
wire output_14_207, output_14_0, output_13_207;
mixer gate_output_13_207(.a(output_14_207), .b(output_14_0), .y(output_13_207));
wire output_15_207, output_15_0, output_14_207;
mixer gate_output_14_207(.a(output_15_207), .b(output_15_0), .y(output_14_207));
wire output_16_207, output_16_0, output_15_207;
mixer gate_output_15_207(.a(output_16_207), .b(output_16_0), .y(output_15_207));
wire output_1_208, output_1_1, output_0_208;
mixer gate_output_0_208(.a(output_1_208), .b(output_1_1), .y(output_0_208));
wire output_2_208, output_2_1, output_1_208;
mixer gate_output_1_208(.a(output_2_208), .b(output_2_1), .y(output_1_208));
wire output_3_208, output_3_1, output_2_208;
mixer gate_output_2_208(.a(output_3_208), .b(output_3_1), .y(output_2_208));
wire output_4_208, output_4_1, output_3_208;
mixer gate_output_3_208(.a(output_4_208), .b(output_4_1), .y(output_3_208));
wire output_5_208, output_5_1, output_4_208;
mixer gate_output_4_208(.a(output_5_208), .b(output_5_1), .y(output_4_208));
wire output_6_208, output_6_1, output_5_208;
mixer gate_output_5_208(.a(output_6_208), .b(output_6_1), .y(output_5_208));
wire output_7_208, output_7_1, output_6_208;
mixer gate_output_6_208(.a(output_7_208), .b(output_7_1), .y(output_6_208));
wire output_8_208, output_8_1, output_7_208;
mixer gate_output_7_208(.a(output_8_208), .b(output_8_1), .y(output_7_208));
wire output_9_208, output_9_1, output_8_208;
mixer gate_output_8_208(.a(output_9_208), .b(output_9_1), .y(output_8_208));
wire output_10_208, output_10_1, output_9_208;
mixer gate_output_9_208(.a(output_10_208), .b(output_10_1), .y(output_9_208));
wire output_11_208, output_11_1, output_10_208;
mixer gate_output_10_208(.a(output_11_208), .b(output_11_1), .y(output_10_208));
wire output_12_208, output_12_1, output_11_208;
mixer gate_output_11_208(.a(output_12_208), .b(output_12_1), .y(output_11_208));
wire output_13_208, output_13_1, output_12_208;
mixer gate_output_12_208(.a(output_13_208), .b(output_13_1), .y(output_12_208));
wire output_14_208, output_14_1, output_13_208;
mixer gate_output_13_208(.a(output_14_208), .b(output_14_1), .y(output_13_208));
wire output_15_208, output_15_1, output_14_208;
mixer gate_output_14_208(.a(output_15_208), .b(output_15_1), .y(output_14_208));
wire output_16_208, output_16_1, output_15_208;
mixer gate_output_15_208(.a(output_16_208), .b(output_16_1), .y(output_15_208));
wire output_1_209, output_1_2, output_0_209;
mixer gate_output_0_209(.a(output_1_209), .b(output_1_2), .y(output_0_209));
wire output_2_209, output_2_2, output_1_209;
mixer gate_output_1_209(.a(output_2_209), .b(output_2_2), .y(output_1_209));
wire output_3_209, output_3_2, output_2_209;
mixer gate_output_2_209(.a(output_3_209), .b(output_3_2), .y(output_2_209));
wire output_4_209, output_4_2, output_3_209;
mixer gate_output_3_209(.a(output_4_209), .b(output_4_2), .y(output_3_209));
wire output_5_209, output_5_2, output_4_209;
mixer gate_output_4_209(.a(output_5_209), .b(output_5_2), .y(output_4_209));
wire output_6_209, output_6_2, output_5_209;
mixer gate_output_5_209(.a(output_6_209), .b(output_6_2), .y(output_5_209));
wire output_7_209, output_7_2, output_6_209;
mixer gate_output_6_209(.a(output_7_209), .b(output_7_2), .y(output_6_209));
wire output_8_209, output_8_2, output_7_209;
mixer gate_output_7_209(.a(output_8_209), .b(output_8_2), .y(output_7_209));
wire output_9_209, output_9_2, output_8_209;
mixer gate_output_8_209(.a(output_9_209), .b(output_9_2), .y(output_8_209));
wire output_10_209, output_10_2, output_9_209;
mixer gate_output_9_209(.a(output_10_209), .b(output_10_2), .y(output_9_209));
wire output_11_209, output_11_2, output_10_209;
mixer gate_output_10_209(.a(output_11_209), .b(output_11_2), .y(output_10_209));
wire output_12_209, output_12_2, output_11_209;
mixer gate_output_11_209(.a(output_12_209), .b(output_12_2), .y(output_11_209));
wire output_13_209, output_13_2, output_12_209;
mixer gate_output_12_209(.a(output_13_209), .b(output_13_2), .y(output_12_209));
wire output_14_209, output_14_2, output_13_209;
mixer gate_output_13_209(.a(output_14_209), .b(output_14_2), .y(output_13_209));
wire output_15_209, output_15_2, output_14_209;
mixer gate_output_14_209(.a(output_15_209), .b(output_15_2), .y(output_14_209));
wire output_16_209, output_16_2, output_15_209;
mixer gate_output_15_209(.a(output_16_209), .b(output_16_2), .y(output_15_209));
wire output_1_210, output_1_3, output_0_210;
mixer gate_output_0_210(.a(output_1_210), .b(output_1_3), .y(output_0_210));
wire output_2_210, output_2_3, output_1_210;
mixer gate_output_1_210(.a(output_2_210), .b(output_2_3), .y(output_1_210));
wire output_3_210, output_3_3, output_2_210;
mixer gate_output_2_210(.a(output_3_210), .b(output_3_3), .y(output_2_210));
wire output_4_210, output_4_3, output_3_210;
mixer gate_output_3_210(.a(output_4_210), .b(output_4_3), .y(output_3_210));
wire output_5_210, output_5_3, output_4_210;
mixer gate_output_4_210(.a(output_5_210), .b(output_5_3), .y(output_4_210));
wire output_6_210, output_6_3, output_5_210;
mixer gate_output_5_210(.a(output_6_210), .b(output_6_3), .y(output_5_210));
wire output_7_210, output_7_3, output_6_210;
mixer gate_output_6_210(.a(output_7_210), .b(output_7_3), .y(output_6_210));
wire output_8_210, output_8_3, output_7_210;
mixer gate_output_7_210(.a(output_8_210), .b(output_8_3), .y(output_7_210));
wire output_9_210, output_9_3, output_8_210;
mixer gate_output_8_210(.a(output_9_210), .b(output_9_3), .y(output_8_210));
wire output_10_210, output_10_3, output_9_210;
mixer gate_output_9_210(.a(output_10_210), .b(output_10_3), .y(output_9_210));
wire output_11_210, output_11_3, output_10_210;
mixer gate_output_10_210(.a(output_11_210), .b(output_11_3), .y(output_10_210));
wire output_12_210, output_12_3, output_11_210;
mixer gate_output_11_210(.a(output_12_210), .b(output_12_3), .y(output_11_210));
wire output_13_210, output_13_3, output_12_210;
mixer gate_output_12_210(.a(output_13_210), .b(output_13_3), .y(output_12_210));
wire output_14_210, output_14_3, output_13_210;
mixer gate_output_13_210(.a(output_14_210), .b(output_14_3), .y(output_13_210));
wire output_15_210, output_15_3, output_14_210;
mixer gate_output_14_210(.a(output_15_210), .b(output_15_3), .y(output_14_210));
wire output_16_210, output_16_3, output_15_210;
mixer gate_output_15_210(.a(output_16_210), .b(output_16_3), .y(output_15_210));
wire output_1_211, output_1_4, output_0_211;
mixer gate_output_0_211(.a(output_1_211), .b(output_1_4), .y(output_0_211));
wire output_2_211, output_2_4, output_1_211;
mixer gate_output_1_211(.a(output_2_211), .b(output_2_4), .y(output_1_211));
wire output_3_211, output_3_4, output_2_211;
mixer gate_output_2_211(.a(output_3_211), .b(output_3_4), .y(output_2_211));
wire output_4_211, output_4_4, output_3_211;
mixer gate_output_3_211(.a(output_4_211), .b(output_4_4), .y(output_3_211));
wire output_5_211, output_5_4, output_4_211;
mixer gate_output_4_211(.a(output_5_211), .b(output_5_4), .y(output_4_211));
wire output_6_211, output_6_4, output_5_211;
mixer gate_output_5_211(.a(output_6_211), .b(output_6_4), .y(output_5_211));
wire output_7_211, output_7_4, output_6_211;
mixer gate_output_6_211(.a(output_7_211), .b(output_7_4), .y(output_6_211));
wire output_8_211, output_8_4, output_7_211;
mixer gate_output_7_211(.a(output_8_211), .b(output_8_4), .y(output_7_211));
wire output_9_211, output_9_4, output_8_211;
mixer gate_output_8_211(.a(output_9_211), .b(output_9_4), .y(output_8_211));
wire output_10_211, output_10_4, output_9_211;
mixer gate_output_9_211(.a(output_10_211), .b(output_10_4), .y(output_9_211));
wire output_11_211, output_11_4, output_10_211;
mixer gate_output_10_211(.a(output_11_211), .b(output_11_4), .y(output_10_211));
wire output_12_211, output_12_4, output_11_211;
mixer gate_output_11_211(.a(output_12_211), .b(output_12_4), .y(output_11_211));
wire output_13_211, output_13_4, output_12_211;
mixer gate_output_12_211(.a(output_13_211), .b(output_13_4), .y(output_12_211));
wire output_14_211, output_14_4, output_13_211;
mixer gate_output_13_211(.a(output_14_211), .b(output_14_4), .y(output_13_211));
wire output_15_211, output_15_4, output_14_211;
mixer gate_output_14_211(.a(output_15_211), .b(output_15_4), .y(output_14_211));
wire output_16_211, output_16_4, output_15_211;
mixer gate_output_15_211(.a(output_16_211), .b(output_16_4), .y(output_15_211));
wire output_1_212, output_1_5, output_0_212;
mixer gate_output_0_212(.a(output_1_212), .b(output_1_5), .y(output_0_212));
wire output_2_212, output_2_5, output_1_212;
mixer gate_output_1_212(.a(output_2_212), .b(output_2_5), .y(output_1_212));
wire output_3_212, output_3_5, output_2_212;
mixer gate_output_2_212(.a(output_3_212), .b(output_3_5), .y(output_2_212));
wire output_4_212, output_4_5, output_3_212;
mixer gate_output_3_212(.a(output_4_212), .b(output_4_5), .y(output_3_212));
wire output_5_212, output_5_5, output_4_212;
mixer gate_output_4_212(.a(output_5_212), .b(output_5_5), .y(output_4_212));
wire output_6_212, output_6_5, output_5_212;
mixer gate_output_5_212(.a(output_6_212), .b(output_6_5), .y(output_5_212));
wire output_7_212, output_7_5, output_6_212;
mixer gate_output_6_212(.a(output_7_212), .b(output_7_5), .y(output_6_212));
wire output_8_212, output_8_5, output_7_212;
mixer gate_output_7_212(.a(output_8_212), .b(output_8_5), .y(output_7_212));
wire output_9_212, output_9_5, output_8_212;
mixer gate_output_8_212(.a(output_9_212), .b(output_9_5), .y(output_8_212));
wire output_10_212, output_10_5, output_9_212;
mixer gate_output_9_212(.a(output_10_212), .b(output_10_5), .y(output_9_212));
wire output_11_212, output_11_5, output_10_212;
mixer gate_output_10_212(.a(output_11_212), .b(output_11_5), .y(output_10_212));
wire output_12_212, output_12_5, output_11_212;
mixer gate_output_11_212(.a(output_12_212), .b(output_12_5), .y(output_11_212));
wire output_13_212, output_13_5, output_12_212;
mixer gate_output_12_212(.a(output_13_212), .b(output_13_5), .y(output_12_212));
wire output_14_212, output_14_5, output_13_212;
mixer gate_output_13_212(.a(output_14_212), .b(output_14_5), .y(output_13_212));
wire output_15_212, output_15_5, output_14_212;
mixer gate_output_14_212(.a(output_15_212), .b(output_15_5), .y(output_14_212));
wire output_16_212, output_16_5, output_15_212;
mixer gate_output_15_212(.a(output_16_212), .b(output_16_5), .y(output_15_212));
wire output_1_213, output_1_6, output_0_213;
mixer gate_output_0_213(.a(output_1_213), .b(output_1_6), .y(output_0_213));
wire output_2_213, output_2_6, output_1_213;
mixer gate_output_1_213(.a(output_2_213), .b(output_2_6), .y(output_1_213));
wire output_3_213, output_3_6, output_2_213;
mixer gate_output_2_213(.a(output_3_213), .b(output_3_6), .y(output_2_213));
wire output_4_213, output_4_6, output_3_213;
mixer gate_output_3_213(.a(output_4_213), .b(output_4_6), .y(output_3_213));
wire output_5_213, output_5_6, output_4_213;
mixer gate_output_4_213(.a(output_5_213), .b(output_5_6), .y(output_4_213));
wire output_6_213, output_6_6, output_5_213;
mixer gate_output_5_213(.a(output_6_213), .b(output_6_6), .y(output_5_213));
wire output_7_213, output_7_6, output_6_213;
mixer gate_output_6_213(.a(output_7_213), .b(output_7_6), .y(output_6_213));
wire output_8_213, output_8_6, output_7_213;
mixer gate_output_7_213(.a(output_8_213), .b(output_8_6), .y(output_7_213));
wire output_9_213, output_9_6, output_8_213;
mixer gate_output_8_213(.a(output_9_213), .b(output_9_6), .y(output_8_213));
wire output_10_213, output_10_6, output_9_213;
mixer gate_output_9_213(.a(output_10_213), .b(output_10_6), .y(output_9_213));
wire output_11_213, output_11_6, output_10_213;
mixer gate_output_10_213(.a(output_11_213), .b(output_11_6), .y(output_10_213));
wire output_12_213, output_12_6, output_11_213;
mixer gate_output_11_213(.a(output_12_213), .b(output_12_6), .y(output_11_213));
wire output_13_213, output_13_6, output_12_213;
mixer gate_output_12_213(.a(output_13_213), .b(output_13_6), .y(output_12_213));
wire output_14_213, output_14_6, output_13_213;
mixer gate_output_13_213(.a(output_14_213), .b(output_14_6), .y(output_13_213));
wire output_15_213, output_15_6, output_14_213;
mixer gate_output_14_213(.a(output_15_213), .b(output_15_6), .y(output_14_213));
wire output_16_213, output_16_6, output_15_213;
mixer gate_output_15_213(.a(output_16_213), .b(output_16_6), .y(output_15_213));
wire output_1_214, output_1_7, output_0_214;
mixer gate_output_0_214(.a(output_1_214), .b(output_1_7), .y(output_0_214));
wire output_2_214, output_2_7, output_1_214;
mixer gate_output_1_214(.a(output_2_214), .b(output_2_7), .y(output_1_214));
wire output_3_214, output_3_7, output_2_214;
mixer gate_output_2_214(.a(output_3_214), .b(output_3_7), .y(output_2_214));
wire output_4_214, output_4_7, output_3_214;
mixer gate_output_3_214(.a(output_4_214), .b(output_4_7), .y(output_3_214));
wire output_5_214, output_5_7, output_4_214;
mixer gate_output_4_214(.a(output_5_214), .b(output_5_7), .y(output_4_214));
wire output_6_214, output_6_7, output_5_214;
mixer gate_output_5_214(.a(output_6_214), .b(output_6_7), .y(output_5_214));
wire output_7_214, output_7_7, output_6_214;
mixer gate_output_6_214(.a(output_7_214), .b(output_7_7), .y(output_6_214));
wire output_8_214, output_8_7, output_7_214;
mixer gate_output_7_214(.a(output_8_214), .b(output_8_7), .y(output_7_214));
wire output_9_214, output_9_7, output_8_214;
mixer gate_output_8_214(.a(output_9_214), .b(output_9_7), .y(output_8_214));
wire output_10_214, output_10_7, output_9_214;
mixer gate_output_9_214(.a(output_10_214), .b(output_10_7), .y(output_9_214));
wire output_11_214, output_11_7, output_10_214;
mixer gate_output_10_214(.a(output_11_214), .b(output_11_7), .y(output_10_214));
wire output_12_214, output_12_7, output_11_214;
mixer gate_output_11_214(.a(output_12_214), .b(output_12_7), .y(output_11_214));
wire output_13_214, output_13_7, output_12_214;
mixer gate_output_12_214(.a(output_13_214), .b(output_13_7), .y(output_12_214));
wire output_14_214, output_14_7, output_13_214;
mixer gate_output_13_214(.a(output_14_214), .b(output_14_7), .y(output_13_214));
wire output_15_214, output_15_7, output_14_214;
mixer gate_output_14_214(.a(output_15_214), .b(output_15_7), .y(output_14_214));
wire output_16_214, output_16_7, output_15_214;
mixer gate_output_15_214(.a(output_16_214), .b(output_16_7), .y(output_15_214));
wire output_1_215, output_1_8, output_0_215;
mixer gate_output_0_215(.a(output_1_215), .b(output_1_8), .y(output_0_215));
wire output_2_215, output_2_8, output_1_215;
mixer gate_output_1_215(.a(output_2_215), .b(output_2_8), .y(output_1_215));
wire output_3_215, output_3_8, output_2_215;
mixer gate_output_2_215(.a(output_3_215), .b(output_3_8), .y(output_2_215));
wire output_4_215, output_4_8, output_3_215;
mixer gate_output_3_215(.a(output_4_215), .b(output_4_8), .y(output_3_215));
wire output_5_215, output_5_8, output_4_215;
mixer gate_output_4_215(.a(output_5_215), .b(output_5_8), .y(output_4_215));
wire output_6_215, output_6_8, output_5_215;
mixer gate_output_5_215(.a(output_6_215), .b(output_6_8), .y(output_5_215));
wire output_7_215, output_7_8, output_6_215;
mixer gate_output_6_215(.a(output_7_215), .b(output_7_8), .y(output_6_215));
wire output_8_215, output_8_8, output_7_215;
mixer gate_output_7_215(.a(output_8_215), .b(output_8_8), .y(output_7_215));
wire output_9_215, output_9_8, output_8_215;
mixer gate_output_8_215(.a(output_9_215), .b(output_9_8), .y(output_8_215));
wire output_10_215, output_10_8, output_9_215;
mixer gate_output_9_215(.a(output_10_215), .b(output_10_8), .y(output_9_215));
wire output_11_215, output_11_8, output_10_215;
mixer gate_output_10_215(.a(output_11_215), .b(output_11_8), .y(output_10_215));
wire output_12_215, output_12_8, output_11_215;
mixer gate_output_11_215(.a(output_12_215), .b(output_12_8), .y(output_11_215));
wire output_13_215, output_13_8, output_12_215;
mixer gate_output_12_215(.a(output_13_215), .b(output_13_8), .y(output_12_215));
wire output_14_215, output_14_8, output_13_215;
mixer gate_output_13_215(.a(output_14_215), .b(output_14_8), .y(output_13_215));
wire output_15_215, output_15_8, output_14_215;
mixer gate_output_14_215(.a(output_15_215), .b(output_15_8), .y(output_14_215));
wire output_16_215, output_16_8, output_15_215;
mixer gate_output_15_215(.a(output_16_215), .b(output_16_8), .y(output_15_215));
wire output_1_216, output_1_9, output_0_216;
mixer gate_output_0_216(.a(output_1_216), .b(output_1_9), .y(output_0_216));
wire output_2_216, output_2_9, output_1_216;
mixer gate_output_1_216(.a(output_2_216), .b(output_2_9), .y(output_1_216));
wire output_3_216, output_3_9, output_2_216;
mixer gate_output_2_216(.a(output_3_216), .b(output_3_9), .y(output_2_216));
wire output_4_216, output_4_9, output_3_216;
mixer gate_output_3_216(.a(output_4_216), .b(output_4_9), .y(output_3_216));
wire output_5_216, output_5_9, output_4_216;
mixer gate_output_4_216(.a(output_5_216), .b(output_5_9), .y(output_4_216));
wire output_6_216, output_6_9, output_5_216;
mixer gate_output_5_216(.a(output_6_216), .b(output_6_9), .y(output_5_216));
wire output_7_216, output_7_9, output_6_216;
mixer gate_output_6_216(.a(output_7_216), .b(output_7_9), .y(output_6_216));
wire output_8_216, output_8_9, output_7_216;
mixer gate_output_7_216(.a(output_8_216), .b(output_8_9), .y(output_7_216));
wire output_9_216, output_9_9, output_8_216;
mixer gate_output_8_216(.a(output_9_216), .b(output_9_9), .y(output_8_216));
wire output_10_216, output_10_9, output_9_216;
mixer gate_output_9_216(.a(output_10_216), .b(output_10_9), .y(output_9_216));
wire output_11_216, output_11_9, output_10_216;
mixer gate_output_10_216(.a(output_11_216), .b(output_11_9), .y(output_10_216));
wire output_12_216, output_12_9, output_11_216;
mixer gate_output_11_216(.a(output_12_216), .b(output_12_9), .y(output_11_216));
wire output_13_216, output_13_9, output_12_216;
mixer gate_output_12_216(.a(output_13_216), .b(output_13_9), .y(output_12_216));
wire output_14_216, output_14_9, output_13_216;
mixer gate_output_13_216(.a(output_14_216), .b(output_14_9), .y(output_13_216));
wire output_15_216, output_15_9, output_14_216;
mixer gate_output_14_216(.a(output_15_216), .b(output_15_9), .y(output_14_216));
wire output_16_216, output_16_9, output_15_216;
mixer gate_output_15_216(.a(output_16_216), .b(output_16_9), .y(output_15_216));
wire output_1_217, output_1_10, output_0_217;
mixer gate_output_0_217(.a(output_1_217), .b(output_1_10), .y(output_0_217));
wire output_2_217, output_2_10, output_1_217;
mixer gate_output_1_217(.a(output_2_217), .b(output_2_10), .y(output_1_217));
wire output_3_217, output_3_10, output_2_217;
mixer gate_output_2_217(.a(output_3_217), .b(output_3_10), .y(output_2_217));
wire output_4_217, output_4_10, output_3_217;
mixer gate_output_3_217(.a(output_4_217), .b(output_4_10), .y(output_3_217));
wire output_5_217, output_5_10, output_4_217;
mixer gate_output_4_217(.a(output_5_217), .b(output_5_10), .y(output_4_217));
wire output_6_217, output_6_10, output_5_217;
mixer gate_output_5_217(.a(output_6_217), .b(output_6_10), .y(output_5_217));
wire output_7_217, output_7_10, output_6_217;
mixer gate_output_6_217(.a(output_7_217), .b(output_7_10), .y(output_6_217));
wire output_8_217, output_8_10, output_7_217;
mixer gate_output_7_217(.a(output_8_217), .b(output_8_10), .y(output_7_217));
wire output_9_217, output_9_10, output_8_217;
mixer gate_output_8_217(.a(output_9_217), .b(output_9_10), .y(output_8_217));
wire output_10_217, output_10_10, output_9_217;
mixer gate_output_9_217(.a(output_10_217), .b(output_10_10), .y(output_9_217));
wire output_11_217, output_11_10, output_10_217;
mixer gate_output_10_217(.a(output_11_217), .b(output_11_10), .y(output_10_217));
wire output_12_217, output_12_10, output_11_217;
mixer gate_output_11_217(.a(output_12_217), .b(output_12_10), .y(output_11_217));
wire output_13_217, output_13_10, output_12_217;
mixer gate_output_12_217(.a(output_13_217), .b(output_13_10), .y(output_12_217));
wire output_14_217, output_14_10, output_13_217;
mixer gate_output_13_217(.a(output_14_217), .b(output_14_10), .y(output_13_217));
wire output_15_217, output_15_10, output_14_217;
mixer gate_output_14_217(.a(output_15_217), .b(output_15_10), .y(output_14_217));
wire output_16_217, output_16_10, output_15_217;
mixer gate_output_15_217(.a(output_16_217), .b(output_16_10), .y(output_15_217));
wire output_1_218, output_1_11, output_0_218;
mixer gate_output_0_218(.a(output_1_218), .b(output_1_11), .y(output_0_218));
wire output_2_218, output_2_11, output_1_218;
mixer gate_output_1_218(.a(output_2_218), .b(output_2_11), .y(output_1_218));
wire output_3_218, output_3_11, output_2_218;
mixer gate_output_2_218(.a(output_3_218), .b(output_3_11), .y(output_2_218));
wire output_4_218, output_4_11, output_3_218;
mixer gate_output_3_218(.a(output_4_218), .b(output_4_11), .y(output_3_218));
wire output_5_218, output_5_11, output_4_218;
mixer gate_output_4_218(.a(output_5_218), .b(output_5_11), .y(output_4_218));
wire output_6_218, output_6_11, output_5_218;
mixer gate_output_5_218(.a(output_6_218), .b(output_6_11), .y(output_5_218));
wire output_7_218, output_7_11, output_6_218;
mixer gate_output_6_218(.a(output_7_218), .b(output_7_11), .y(output_6_218));
wire output_8_218, output_8_11, output_7_218;
mixer gate_output_7_218(.a(output_8_218), .b(output_8_11), .y(output_7_218));
wire output_9_218, output_9_11, output_8_218;
mixer gate_output_8_218(.a(output_9_218), .b(output_9_11), .y(output_8_218));
wire output_10_218, output_10_11, output_9_218;
mixer gate_output_9_218(.a(output_10_218), .b(output_10_11), .y(output_9_218));
wire output_11_218, output_11_11, output_10_218;
mixer gate_output_10_218(.a(output_11_218), .b(output_11_11), .y(output_10_218));
wire output_12_218, output_12_11, output_11_218;
mixer gate_output_11_218(.a(output_12_218), .b(output_12_11), .y(output_11_218));
wire output_13_218, output_13_11, output_12_218;
mixer gate_output_12_218(.a(output_13_218), .b(output_13_11), .y(output_12_218));
wire output_14_218, output_14_11, output_13_218;
mixer gate_output_13_218(.a(output_14_218), .b(output_14_11), .y(output_13_218));
wire output_15_218, output_15_11, output_14_218;
mixer gate_output_14_218(.a(output_15_218), .b(output_15_11), .y(output_14_218));
wire output_16_218, output_16_11, output_15_218;
mixer gate_output_15_218(.a(output_16_218), .b(output_16_11), .y(output_15_218));
wire output_1_219, output_1_12, output_0_219;
mixer gate_output_0_219(.a(output_1_219), .b(output_1_12), .y(output_0_219));
wire output_2_219, output_2_12, output_1_219;
mixer gate_output_1_219(.a(output_2_219), .b(output_2_12), .y(output_1_219));
wire output_3_219, output_3_12, output_2_219;
mixer gate_output_2_219(.a(output_3_219), .b(output_3_12), .y(output_2_219));
wire output_4_219, output_4_12, output_3_219;
mixer gate_output_3_219(.a(output_4_219), .b(output_4_12), .y(output_3_219));
wire output_5_219, output_5_12, output_4_219;
mixer gate_output_4_219(.a(output_5_219), .b(output_5_12), .y(output_4_219));
wire output_6_219, output_6_12, output_5_219;
mixer gate_output_5_219(.a(output_6_219), .b(output_6_12), .y(output_5_219));
wire output_7_219, output_7_12, output_6_219;
mixer gate_output_6_219(.a(output_7_219), .b(output_7_12), .y(output_6_219));
wire output_8_219, output_8_12, output_7_219;
mixer gate_output_7_219(.a(output_8_219), .b(output_8_12), .y(output_7_219));
wire output_9_219, output_9_12, output_8_219;
mixer gate_output_8_219(.a(output_9_219), .b(output_9_12), .y(output_8_219));
wire output_10_219, output_10_12, output_9_219;
mixer gate_output_9_219(.a(output_10_219), .b(output_10_12), .y(output_9_219));
wire output_11_219, output_11_12, output_10_219;
mixer gate_output_10_219(.a(output_11_219), .b(output_11_12), .y(output_10_219));
wire output_12_219, output_12_12, output_11_219;
mixer gate_output_11_219(.a(output_12_219), .b(output_12_12), .y(output_11_219));
wire output_13_219, output_13_12, output_12_219;
mixer gate_output_12_219(.a(output_13_219), .b(output_13_12), .y(output_12_219));
wire output_14_219, output_14_12, output_13_219;
mixer gate_output_13_219(.a(output_14_219), .b(output_14_12), .y(output_13_219));
wire output_15_219, output_15_12, output_14_219;
mixer gate_output_14_219(.a(output_15_219), .b(output_15_12), .y(output_14_219));
wire output_16_219, output_16_12, output_15_219;
mixer gate_output_15_219(.a(output_16_219), .b(output_16_12), .y(output_15_219));
wire output_1_220, output_1_13, output_0_220;
mixer gate_output_0_220(.a(output_1_220), .b(output_1_13), .y(output_0_220));
wire output_2_220, output_2_13, output_1_220;
mixer gate_output_1_220(.a(output_2_220), .b(output_2_13), .y(output_1_220));
wire output_3_220, output_3_13, output_2_220;
mixer gate_output_2_220(.a(output_3_220), .b(output_3_13), .y(output_2_220));
wire output_4_220, output_4_13, output_3_220;
mixer gate_output_3_220(.a(output_4_220), .b(output_4_13), .y(output_3_220));
wire output_5_220, output_5_13, output_4_220;
mixer gate_output_4_220(.a(output_5_220), .b(output_5_13), .y(output_4_220));
wire output_6_220, output_6_13, output_5_220;
mixer gate_output_5_220(.a(output_6_220), .b(output_6_13), .y(output_5_220));
wire output_7_220, output_7_13, output_6_220;
mixer gate_output_6_220(.a(output_7_220), .b(output_7_13), .y(output_6_220));
wire output_8_220, output_8_13, output_7_220;
mixer gate_output_7_220(.a(output_8_220), .b(output_8_13), .y(output_7_220));
wire output_9_220, output_9_13, output_8_220;
mixer gate_output_8_220(.a(output_9_220), .b(output_9_13), .y(output_8_220));
wire output_10_220, output_10_13, output_9_220;
mixer gate_output_9_220(.a(output_10_220), .b(output_10_13), .y(output_9_220));
wire output_11_220, output_11_13, output_10_220;
mixer gate_output_10_220(.a(output_11_220), .b(output_11_13), .y(output_10_220));
wire output_12_220, output_12_13, output_11_220;
mixer gate_output_11_220(.a(output_12_220), .b(output_12_13), .y(output_11_220));
wire output_13_220, output_13_13, output_12_220;
mixer gate_output_12_220(.a(output_13_220), .b(output_13_13), .y(output_12_220));
wire output_14_220, output_14_13, output_13_220;
mixer gate_output_13_220(.a(output_14_220), .b(output_14_13), .y(output_13_220));
wire output_15_220, output_15_13, output_14_220;
mixer gate_output_14_220(.a(output_15_220), .b(output_15_13), .y(output_14_220));
wire output_16_220, output_16_13, output_15_220;
mixer gate_output_15_220(.a(output_16_220), .b(output_16_13), .y(output_15_220));
wire output_1_221, output_1_14, output_0_221;
mixer gate_output_0_221(.a(output_1_221), .b(output_1_14), .y(output_0_221));
wire output_2_221, output_2_14, output_1_221;
mixer gate_output_1_221(.a(output_2_221), .b(output_2_14), .y(output_1_221));
wire output_3_221, output_3_14, output_2_221;
mixer gate_output_2_221(.a(output_3_221), .b(output_3_14), .y(output_2_221));
wire output_4_221, output_4_14, output_3_221;
mixer gate_output_3_221(.a(output_4_221), .b(output_4_14), .y(output_3_221));
wire output_5_221, output_5_14, output_4_221;
mixer gate_output_4_221(.a(output_5_221), .b(output_5_14), .y(output_4_221));
wire output_6_221, output_6_14, output_5_221;
mixer gate_output_5_221(.a(output_6_221), .b(output_6_14), .y(output_5_221));
wire output_7_221, output_7_14, output_6_221;
mixer gate_output_6_221(.a(output_7_221), .b(output_7_14), .y(output_6_221));
wire output_8_221, output_8_14, output_7_221;
mixer gate_output_7_221(.a(output_8_221), .b(output_8_14), .y(output_7_221));
wire output_9_221, output_9_14, output_8_221;
mixer gate_output_8_221(.a(output_9_221), .b(output_9_14), .y(output_8_221));
wire output_10_221, output_10_14, output_9_221;
mixer gate_output_9_221(.a(output_10_221), .b(output_10_14), .y(output_9_221));
wire output_11_221, output_11_14, output_10_221;
mixer gate_output_10_221(.a(output_11_221), .b(output_11_14), .y(output_10_221));
wire output_12_221, output_12_14, output_11_221;
mixer gate_output_11_221(.a(output_12_221), .b(output_12_14), .y(output_11_221));
wire output_13_221, output_13_14, output_12_221;
mixer gate_output_12_221(.a(output_13_221), .b(output_13_14), .y(output_12_221));
wire output_14_221, output_14_14, output_13_221;
mixer gate_output_13_221(.a(output_14_221), .b(output_14_14), .y(output_13_221));
wire output_15_221, output_15_14, output_14_221;
mixer gate_output_14_221(.a(output_15_221), .b(output_15_14), .y(output_14_221));
wire output_16_221, output_16_14, output_15_221;
mixer gate_output_15_221(.a(output_16_221), .b(output_16_14), .y(output_15_221));
wire output_1_222, output_1_15, output_0_222;
mixer gate_output_0_222(.a(output_1_222), .b(output_1_15), .y(output_0_222));
wire output_2_222, output_2_15, output_1_222;
mixer gate_output_1_222(.a(output_2_222), .b(output_2_15), .y(output_1_222));
wire output_3_222, output_3_15, output_2_222;
mixer gate_output_2_222(.a(output_3_222), .b(output_3_15), .y(output_2_222));
wire output_4_222, output_4_15, output_3_222;
mixer gate_output_3_222(.a(output_4_222), .b(output_4_15), .y(output_3_222));
wire output_5_222, output_5_15, output_4_222;
mixer gate_output_4_222(.a(output_5_222), .b(output_5_15), .y(output_4_222));
wire output_6_222, output_6_15, output_5_222;
mixer gate_output_5_222(.a(output_6_222), .b(output_6_15), .y(output_5_222));
wire output_7_222, output_7_15, output_6_222;
mixer gate_output_6_222(.a(output_7_222), .b(output_7_15), .y(output_6_222));
wire output_8_222, output_8_15, output_7_222;
mixer gate_output_7_222(.a(output_8_222), .b(output_8_15), .y(output_7_222));
wire output_9_222, output_9_15, output_8_222;
mixer gate_output_8_222(.a(output_9_222), .b(output_9_15), .y(output_8_222));
wire output_10_222, output_10_15, output_9_222;
mixer gate_output_9_222(.a(output_10_222), .b(output_10_15), .y(output_9_222));
wire output_11_222, output_11_15, output_10_222;
mixer gate_output_10_222(.a(output_11_222), .b(output_11_15), .y(output_10_222));
wire output_12_222, output_12_15, output_11_222;
mixer gate_output_11_222(.a(output_12_222), .b(output_12_15), .y(output_11_222));
wire output_13_222, output_13_15, output_12_222;
mixer gate_output_12_222(.a(output_13_222), .b(output_13_15), .y(output_12_222));
wire output_14_222, output_14_15, output_13_222;
mixer gate_output_13_222(.a(output_14_222), .b(output_14_15), .y(output_13_222));
wire output_15_222, output_15_15, output_14_222;
mixer gate_output_14_222(.a(output_15_222), .b(output_15_15), .y(output_14_222));
wire output_16_222, output_16_15, output_15_222;
mixer gate_output_15_222(.a(output_16_222), .b(output_16_15), .y(output_15_222));
wire output_1_223, output_1_0, output_0_223;
mixer gate_output_0_223(.a(output_1_223), .b(output_1_0), .y(output_0_223));
wire output_2_223, output_2_0, output_1_223;
mixer gate_output_1_223(.a(output_2_223), .b(output_2_0), .y(output_1_223));
wire output_3_223, output_3_0, output_2_223;
mixer gate_output_2_223(.a(output_3_223), .b(output_3_0), .y(output_2_223));
wire output_4_223, output_4_0, output_3_223;
mixer gate_output_3_223(.a(output_4_223), .b(output_4_0), .y(output_3_223));
wire output_5_223, output_5_0, output_4_223;
mixer gate_output_4_223(.a(output_5_223), .b(output_5_0), .y(output_4_223));
wire output_6_223, output_6_0, output_5_223;
mixer gate_output_5_223(.a(output_6_223), .b(output_6_0), .y(output_5_223));
wire output_7_223, output_7_0, output_6_223;
mixer gate_output_6_223(.a(output_7_223), .b(output_7_0), .y(output_6_223));
wire output_8_223, output_8_0, output_7_223;
mixer gate_output_7_223(.a(output_8_223), .b(output_8_0), .y(output_7_223));
wire output_9_223, output_9_0, output_8_223;
mixer gate_output_8_223(.a(output_9_223), .b(output_9_0), .y(output_8_223));
wire output_10_223, output_10_0, output_9_223;
mixer gate_output_9_223(.a(output_10_223), .b(output_10_0), .y(output_9_223));
wire output_11_223, output_11_0, output_10_223;
mixer gate_output_10_223(.a(output_11_223), .b(output_11_0), .y(output_10_223));
wire output_12_223, output_12_0, output_11_223;
mixer gate_output_11_223(.a(output_12_223), .b(output_12_0), .y(output_11_223));
wire output_13_223, output_13_0, output_12_223;
mixer gate_output_12_223(.a(output_13_223), .b(output_13_0), .y(output_12_223));
wire output_14_223, output_14_0, output_13_223;
mixer gate_output_13_223(.a(output_14_223), .b(output_14_0), .y(output_13_223));
wire output_15_223, output_15_0, output_14_223;
mixer gate_output_14_223(.a(output_15_223), .b(output_15_0), .y(output_14_223));
wire output_16_223, output_16_0, output_15_223;
mixer gate_output_15_223(.a(output_16_223), .b(output_16_0), .y(output_15_223));
wire output_1_224, output_1_1, output_0_224;
mixer gate_output_0_224(.a(output_1_224), .b(output_1_1), .y(output_0_224));
wire output_2_224, output_2_1, output_1_224;
mixer gate_output_1_224(.a(output_2_224), .b(output_2_1), .y(output_1_224));
wire output_3_224, output_3_1, output_2_224;
mixer gate_output_2_224(.a(output_3_224), .b(output_3_1), .y(output_2_224));
wire output_4_224, output_4_1, output_3_224;
mixer gate_output_3_224(.a(output_4_224), .b(output_4_1), .y(output_3_224));
wire output_5_224, output_5_1, output_4_224;
mixer gate_output_4_224(.a(output_5_224), .b(output_5_1), .y(output_4_224));
wire output_6_224, output_6_1, output_5_224;
mixer gate_output_5_224(.a(output_6_224), .b(output_6_1), .y(output_5_224));
wire output_7_224, output_7_1, output_6_224;
mixer gate_output_6_224(.a(output_7_224), .b(output_7_1), .y(output_6_224));
wire output_8_224, output_8_1, output_7_224;
mixer gate_output_7_224(.a(output_8_224), .b(output_8_1), .y(output_7_224));
wire output_9_224, output_9_1, output_8_224;
mixer gate_output_8_224(.a(output_9_224), .b(output_9_1), .y(output_8_224));
wire output_10_224, output_10_1, output_9_224;
mixer gate_output_9_224(.a(output_10_224), .b(output_10_1), .y(output_9_224));
wire output_11_224, output_11_1, output_10_224;
mixer gate_output_10_224(.a(output_11_224), .b(output_11_1), .y(output_10_224));
wire output_12_224, output_12_1, output_11_224;
mixer gate_output_11_224(.a(output_12_224), .b(output_12_1), .y(output_11_224));
wire output_13_224, output_13_1, output_12_224;
mixer gate_output_12_224(.a(output_13_224), .b(output_13_1), .y(output_12_224));
wire output_14_224, output_14_1, output_13_224;
mixer gate_output_13_224(.a(output_14_224), .b(output_14_1), .y(output_13_224));
wire output_15_224, output_15_1, output_14_224;
mixer gate_output_14_224(.a(output_15_224), .b(output_15_1), .y(output_14_224));
wire output_16_224, output_16_1, output_15_224;
mixer gate_output_15_224(.a(output_16_224), .b(output_16_1), .y(output_15_224));
wire output_1_225, output_1_2, output_0_225;
mixer gate_output_0_225(.a(output_1_225), .b(output_1_2), .y(output_0_225));
wire output_2_225, output_2_2, output_1_225;
mixer gate_output_1_225(.a(output_2_225), .b(output_2_2), .y(output_1_225));
wire output_3_225, output_3_2, output_2_225;
mixer gate_output_2_225(.a(output_3_225), .b(output_3_2), .y(output_2_225));
wire output_4_225, output_4_2, output_3_225;
mixer gate_output_3_225(.a(output_4_225), .b(output_4_2), .y(output_3_225));
wire output_5_225, output_5_2, output_4_225;
mixer gate_output_4_225(.a(output_5_225), .b(output_5_2), .y(output_4_225));
wire output_6_225, output_6_2, output_5_225;
mixer gate_output_5_225(.a(output_6_225), .b(output_6_2), .y(output_5_225));
wire output_7_225, output_7_2, output_6_225;
mixer gate_output_6_225(.a(output_7_225), .b(output_7_2), .y(output_6_225));
wire output_8_225, output_8_2, output_7_225;
mixer gate_output_7_225(.a(output_8_225), .b(output_8_2), .y(output_7_225));
wire output_9_225, output_9_2, output_8_225;
mixer gate_output_8_225(.a(output_9_225), .b(output_9_2), .y(output_8_225));
wire output_10_225, output_10_2, output_9_225;
mixer gate_output_9_225(.a(output_10_225), .b(output_10_2), .y(output_9_225));
wire output_11_225, output_11_2, output_10_225;
mixer gate_output_10_225(.a(output_11_225), .b(output_11_2), .y(output_10_225));
wire output_12_225, output_12_2, output_11_225;
mixer gate_output_11_225(.a(output_12_225), .b(output_12_2), .y(output_11_225));
wire output_13_225, output_13_2, output_12_225;
mixer gate_output_12_225(.a(output_13_225), .b(output_13_2), .y(output_12_225));
wire output_14_225, output_14_2, output_13_225;
mixer gate_output_13_225(.a(output_14_225), .b(output_14_2), .y(output_13_225));
wire output_15_225, output_15_2, output_14_225;
mixer gate_output_14_225(.a(output_15_225), .b(output_15_2), .y(output_14_225));
wire output_16_225, output_16_2, output_15_225;
mixer gate_output_15_225(.a(output_16_225), .b(output_16_2), .y(output_15_225));
wire output_1_226, output_1_3, output_0_226;
mixer gate_output_0_226(.a(output_1_226), .b(output_1_3), .y(output_0_226));
wire output_2_226, output_2_3, output_1_226;
mixer gate_output_1_226(.a(output_2_226), .b(output_2_3), .y(output_1_226));
wire output_3_226, output_3_3, output_2_226;
mixer gate_output_2_226(.a(output_3_226), .b(output_3_3), .y(output_2_226));
wire output_4_226, output_4_3, output_3_226;
mixer gate_output_3_226(.a(output_4_226), .b(output_4_3), .y(output_3_226));
wire output_5_226, output_5_3, output_4_226;
mixer gate_output_4_226(.a(output_5_226), .b(output_5_3), .y(output_4_226));
wire output_6_226, output_6_3, output_5_226;
mixer gate_output_5_226(.a(output_6_226), .b(output_6_3), .y(output_5_226));
wire output_7_226, output_7_3, output_6_226;
mixer gate_output_6_226(.a(output_7_226), .b(output_7_3), .y(output_6_226));
wire output_8_226, output_8_3, output_7_226;
mixer gate_output_7_226(.a(output_8_226), .b(output_8_3), .y(output_7_226));
wire output_9_226, output_9_3, output_8_226;
mixer gate_output_8_226(.a(output_9_226), .b(output_9_3), .y(output_8_226));
wire output_10_226, output_10_3, output_9_226;
mixer gate_output_9_226(.a(output_10_226), .b(output_10_3), .y(output_9_226));
wire output_11_226, output_11_3, output_10_226;
mixer gate_output_10_226(.a(output_11_226), .b(output_11_3), .y(output_10_226));
wire output_12_226, output_12_3, output_11_226;
mixer gate_output_11_226(.a(output_12_226), .b(output_12_3), .y(output_11_226));
wire output_13_226, output_13_3, output_12_226;
mixer gate_output_12_226(.a(output_13_226), .b(output_13_3), .y(output_12_226));
wire output_14_226, output_14_3, output_13_226;
mixer gate_output_13_226(.a(output_14_226), .b(output_14_3), .y(output_13_226));
wire output_15_226, output_15_3, output_14_226;
mixer gate_output_14_226(.a(output_15_226), .b(output_15_3), .y(output_14_226));
wire output_16_226, output_16_3, output_15_226;
mixer gate_output_15_226(.a(output_16_226), .b(output_16_3), .y(output_15_226));
wire output_1_227, output_1_4, output_0_227;
mixer gate_output_0_227(.a(output_1_227), .b(output_1_4), .y(output_0_227));
wire output_2_227, output_2_4, output_1_227;
mixer gate_output_1_227(.a(output_2_227), .b(output_2_4), .y(output_1_227));
wire output_3_227, output_3_4, output_2_227;
mixer gate_output_2_227(.a(output_3_227), .b(output_3_4), .y(output_2_227));
wire output_4_227, output_4_4, output_3_227;
mixer gate_output_3_227(.a(output_4_227), .b(output_4_4), .y(output_3_227));
wire output_5_227, output_5_4, output_4_227;
mixer gate_output_4_227(.a(output_5_227), .b(output_5_4), .y(output_4_227));
wire output_6_227, output_6_4, output_5_227;
mixer gate_output_5_227(.a(output_6_227), .b(output_6_4), .y(output_5_227));
wire output_7_227, output_7_4, output_6_227;
mixer gate_output_6_227(.a(output_7_227), .b(output_7_4), .y(output_6_227));
wire output_8_227, output_8_4, output_7_227;
mixer gate_output_7_227(.a(output_8_227), .b(output_8_4), .y(output_7_227));
wire output_9_227, output_9_4, output_8_227;
mixer gate_output_8_227(.a(output_9_227), .b(output_9_4), .y(output_8_227));
wire output_10_227, output_10_4, output_9_227;
mixer gate_output_9_227(.a(output_10_227), .b(output_10_4), .y(output_9_227));
wire output_11_227, output_11_4, output_10_227;
mixer gate_output_10_227(.a(output_11_227), .b(output_11_4), .y(output_10_227));
wire output_12_227, output_12_4, output_11_227;
mixer gate_output_11_227(.a(output_12_227), .b(output_12_4), .y(output_11_227));
wire output_13_227, output_13_4, output_12_227;
mixer gate_output_12_227(.a(output_13_227), .b(output_13_4), .y(output_12_227));
wire output_14_227, output_14_4, output_13_227;
mixer gate_output_13_227(.a(output_14_227), .b(output_14_4), .y(output_13_227));
wire output_15_227, output_15_4, output_14_227;
mixer gate_output_14_227(.a(output_15_227), .b(output_15_4), .y(output_14_227));
wire output_16_227, output_16_4, output_15_227;
mixer gate_output_15_227(.a(output_16_227), .b(output_16_4), .y(output_15_227));
wire output_1_228, output_1_5, output_0_228;
mixer gate_output_0_228(.a(output_1_228), .b(output_1_5), .y(output_0_228));
wire output_2_228, output_2_5, output_1_228;
mixer gate_output_1_228(.a(output_2_228), .b(output_2_5), .y(output_1_228));
wire output_3_228, output_3_5, output_2_228;
mixer gate_output_2_228(.a(output_3_228), .b(output_3_5), .y(output_2_228));
wire output_4_228, output_4_5, output_3_228;
mixer gate_output_3_228(.a(output_4_228), .b(output_4_5), .y(output_3_228));
wire output_5_228, output_5_5, output_4_228;
mixer gate_output_4_228(.a(output_5_228), .b(output_5_5), .y(output_4_228));
wire output_6_228, output_6_5, output_5_228;
mixer gate_output_5_228(.a(output_6_228), .b(output_6_5), .y(output_5_228));
wire output_7_228, output_7_5, output_6_228;
mixer gate_output_6_228(.a(output_7_228), .b(output_7_5), .y(output_6_228));
wire output_8_228, output_8_5, output_7_228;
mixer gate_output_7_228(.a(output_8_228), .b(output_8_5), .y(output_7_228));
wire output_9_228, output_9_5, output_8_228;
mixer gate_output_8_228(.a(output_9_228), .b(output_9_5), .y(output_8_228));
wire output_10_228, output_10_5, output_9_228;
mixer gate_output_9_228(.a(output_10_228), .b(output_10_5), .y(output_9_228));
wire output_11_228, output_11_5, output_10_228;
mixer gate_output_10_228(.a(output_11_228), .b(output_11_5), .y(output_10_228));
wire output_12_228, output_12_5, output_11_228;
mixer gate_output_11_228(.a(output_12_228), .b(output_12_5), .y(output_11_228));
wire output_13_228, output_13_5, output_12_228;
mixer gate_output_12_228(.a(output_13_228), .b(output_13_5), .y(output_12_228));
wire output_14_228, output_14_5, output_13_228;
mixer gate_output_13_228(.a(output_14_228), .b(output_14_5), .y(output_13_228));
wire output_15_228, output_15_5, output_14_228;
mixer gate_output_14_228(.a(output_15_228), .b(output_15_5), .y(output_14_228));
wire output_16_228, output_16_5, output_15_228;
mixer gate_output_15_228(.a(output_16_228), .b(output_16_5), .y(output_15_228));
wire output_1_229, output_1_6, output_0_229;
mixer gate_output_0_229(.a(output_1_229), .b(output_1_6), .y(output_0_229));
wire output_2_229, output_2_6, output_1_229;
mixer gate_output_1_229(.a(output_2_229), .b(output_2_6), .y(output_1_229));
wire output_3_229, output_3_6, output_2_229;
mixer gate_output_2_229(.a(output_3_229), .b(output_3_6), .y(output_2_229));
wire output_4_229, output_4_6, output_3_229;
mixer gate_output_3_229(.a(output_4_229), .b(output_4_6), .y(output_3_229));
wire output_5_229, output_5_6, output_4_229;
mixer gate_output_4_229(.a(output_5_229), .b(output_5_6), .y(output_4_229));
wire output_6_229, output_6_6, output_5_229;
mixer gate_output_5_229(.a(output_6_229), .b(output_6_6), .y(output_5_229));
wire output_7_229, output_7_6, output_6_229;
mixer gate_output_6_229(.a(output_7_229), .b(output_7_6), .y(output_6_229));
wire output_8_229, output_8_6, output_7_229;
mixer gate_output_7_229(.a(output_8_229), .b(output_8_6), .y(output_7_229));
wire output_9_229, output_9_6, output_8_229;
mixer gate_output_8_229(.a(output_9_229), .b(output_9_6), .y(output_8_229));
wire output_10_229, output_10_6, output_9_229;
mixer gate_output_9_229(.a(output_10_229), .b(output_10_6), .y(output_9_229));
wire output_11_229, output_11_6, output_10_229;
mixer gate_output_10_229(.a(output_11_229), .b(output_11_6), .y(output_10_229));
wire output_12_229, output_12_6, output_11_229;
mixer gate_output_11_229(.a(output_12_229), .b(output_12_6), .y(output_11_229));
wire output_13_229, output_13_6, output_12_229;
mixer gate_output_12_229(.a(output_13_229), .b(output_13_6), .y(output_12_229));
wire output_14_229, output_14_6, output_13_229;
mixer gate_output_13_229(.a(output_14_229), .b(output_14_6), .y(output_13_229));
wire output_15_229, output_15_6, output_14_229;
mixer gate_output_14_229(.a(output_15_229), .b(output_15_6), .y(output_14_229));
wire output_16_229, output_16_6, output_15_229;
mixer gate_output_15_229(.a(output_16_229), .b(output_16_6), .y(output_15_229));
wire output_1_230, output_1_7, output_0_230;
mixer gate_output_0_230(.a(output_1_230), .b(output_1_7), .y(output_0_230));
wire output_2_230, output_2_7, output_1_230;
mixer gate_output_1_230(.a(output_2_230), .b(output_2_7), .y(output_1_230));
wire output_3_230, output_3_7, output_2_230;
mixer gate_output_2_230(.a(output_3_230), .b(output_3_7), .y(output_2_230));
wire output_4_230, output_4_7, output_3_230;
mixer gate_output_3_230(.a(output_4_230), .b(output_4_7), .y(output_3_230));
wire output_5_230, output_5_7, output_4_230;
mixer gate_output_4_230(.a(output_5_230), .b(output_5_7), .y(output_4_230));
wire output_6_230, output_6_7, output_5_230;
mixer gate_output_5_230(.a(output_6_230), .b(output_6_7), .y(output_5_230));
wire output_7_230, output_7_7, output_6_230;
mixer gate_output_6_230(.a(output_7_230), .b(output_7_7), .y(output_6_230));
wire output_8_230, output_8_7, output_7_230;
mixer gate_output_7_230(.a(output_8_230), .b(output_8_7), .y(output_7_230));
wire output_9_230, output_9_7, output_8_230;
mixer gate_output_8_230(.a(output_9_230), .b(output_9_7), .y(output_8_230));
wire output_10_230, output_10_7, output_9_230;
mixer gate_output_9_230(.a(output_10_230), .b(output_10_7), .y(output_9_230));
wire output_11_230, output_11_7, output_10_230;
mixer gate_output_10_230(.a(output_11_230), .b(output_11_7), .y(output_10_230));
wire output_12_230, output_12_7, output_11_230;
mixer gate_output_11_230(.a(output_12_230), .b(output_12_7), .y(output_11_230));
wire output_13_230, output_13_7, output_12_230;
mixer gate_output_12_230(.a(output_13_230), .b(output_13_7), .y(output_12_230));
wire output_14_230, output_14_7, output_13_230;
mixer gate_output_13_230(.a(output_14_230), .b(output_14_7), .y(output_13_230));
wire output_15_230, output_15_7, output_14_230;
mixer gate_output_14_230(.a(output_15_230), .b(output_15_7), .y(output_14_230));
wire output_16_230, output_16_7, output_15_230;
mixer gate_output_15_230(.a(output_16_230), .b(output_16_7), .y(output_15_230));
wire output_1_231, output_1_8, output_0_231;
mixer gate_output_0_231(.a(output_1_231), .b(output_1_8), .y(output_0_231));
wire output_2_231, output_2_8, output_1_231;
mixer gate_output_1_231(.a(output_2_231), .b(output_2_8), .y(output_1_231));
wire output_3_231, output_3_8, output_2_231;
mixer gate_output_2_231(.a(output_3_231), .b(output_3_8), .y(output_2_231));
wire output_4_231, output_4_8, output_3_231;
mixer gate_output_3_231(.a(output_4_231), .b(output_4_8), .y(output_3_231));
wire output_5_231, output_5_8, output_4_231;
mixer gate_output_4_231(.a(output_5_231), .b(output_5_8), .y(output_4_231));
wire output_6_231, output_6_8, output_5_231;
mixer gate_output_5_231(.a(output_6_231), .b(output_6_8), .y(output_5_231));
wire output_7_231, output_7_8, output_6_231;
mixer gate_output_6_231(.a(output_7_231), .b(output_7_8), .y(output_6_231));
wire output_8_231, output_8_8, output_7_231;
mixer gate_output_7_231(.a(output_8_231), .b(output_8_8), .y(output_7_231));
wire output_9_231, output_9_8, output_8_231;
mixer gate_output_8_231(.a(output_9_231), .b(output_9_8), .y(output_8_231));
wire output_10_231, output_10_8, output_9_231;
mixer gate_output_9_231(.a(output_10_231), .b(output_10_8), .y(output_9_231));
wire output_11_231, output_11_8, output_10_231;
mixer gate_output_10_231(.a(output_11_231), .b(output_11_8), .y(output_10_231));
wire output_12_231, output_12_8, output_11_231;
mixer gate_output_11_231(.a(output_12_231), .b(output_12_8), .y(output_11_231));
wire output_13_231, output_13_8, output_12_231;
mixer gate_output_12_231(.a(output_13_231), .b(output_13_8), .y(output_12_231));
wire output_14_231, output_14_8, output_13_231;
mixer gate_output_13_231(.a(output_14_231), .b(output_14_8), .y(output_13_231));
wire output_15_231, output_15_8, output_14_231;
mixer gate_output_14_231(.a(output_15_231), .b(output_15_8), .y(output_14_231));
wire output_16_231, output_16_8, output_15_231;
mixer gate_output_15_231(.a(output_16_231), .b(output_16_8), .y(output_15_231));
wire output_1_232, output_1_9, output_0_232;
mixer gate_output_0_232(.a(output_1_232), .b(output_1_9), .y(output_0_232));
wire output_2_232, output_2_9, output_1_232;
mixer gate_output_1_232(.a(output_2_232), .b(output_2_9), .y(output_1_232));
wire output_3_232, output_3_9, output_2_232;
mixer gate_output_2_232(.a(output_3_232), .b(output_3_9), .y(output_2_232));
wire output_4_232, output_4_9, output_3_232;
mixer gate_output_3_232(.a(output_4_232), .b(output_4_9), .y(output_3_232));
wire output_5_232, output_5_9, output_4_232;
mixer gate_output_4_232(.a(output_5_232), .b(output_5_9), .y(output_4_232));
wire output_6_232, output_6_9, output_5_232;
mixer gate_output_5_232(.a(output_6_232), .b(output_6_9), .y(output_5_232));
wire output_7_232, output_7_9, output_6_232;
mixer gate_output_6_232(.a(output_7_232), .b(output_7_9), .y(output_6_232));
wire output_8_232, output_8_9, output_7_232;
mixer gate_output_7_232(.a(output_8_232), .b(output_8_9), .y(output_7_232));
wire output_9_232, output_9_9, output_8_232;
mixer gate_output_8_232(.a(output_9_232), .b(output_9_9), .y(output_8_232));
wire output_10_232, output_10_9, output_9_232;
mixer gate_output_9_232(.a(output_10_232), .b(output_10_9), .y(output_9_232));
wire output_11_232, output_11_9, output_10_232;
mixer gate_output_10_232(.a(output_11_232), .b(output_11_9), .y(output_10_232));
wire output_12_232, output_12_9, output_11_232;
mixer gate_output_11_232(.a(output_12_232), .b(output_12_9), .y(output_11_232));
wire output_13_232, output_13_9, output_12_232;
mixer gate_output_12_232(.a(output_13_232), .b(output_13_9), .y(output_12_232));
wire output_14_232, output_14_9, output_13_232;
mixer gate_output_13_232(.a(output_14_232), .b(output_14_9), .y(output_13_232));
wire output_15_232, output_15_9, output_14_232;
mixer gate_output_14_232(.a(output_15_232), .b(output_15_9), .y(output_14_232));
wire output_16_232, output_16_9, output_15_232;
mixer gate_output_15_232(.a(output_16_232), .b(output_16_9), .y(output_15_232));
wire output_1_233, output_1_10, output_0_233;
mixer gate_output_0_233(.a(output_1_233), .b(output_1_10), .y(output_0_233));
wire output_2_233, output_2_10, output_1_233;
mixer gate_output_1_233(.a(output_2_233), .b(output_2_10), .y(output_1_233));
wire output_3_233, output_3_10, output_2_233;
mixer gate_output_2_233(.a(output_3_233), .b(output_3_10), .y(output_2_233));
wire output_4_233, output_4_10, output_3_233;
mixer gate_output_3_233(.a(output_4_233), .b(output_4_10), .y(output_3_233));
wire output_5_233, output_5_10, output_4_233;
mixer gate_output_4_233(.a(output_5_233), .b(output_5_10), .y(output_4_233));
wire output_6_233, output_6_10, output_5_233;
mixer gate_output_5_233(.a(output_6_233), .b(output_6_10), .y(output_5_233));
wire output_7_233, output_7_10, output_6_233;
mixer gate_output_6_233(.a(output_7_233), .b(output_7_10), .y(output_6_233));
wire output_8_233, output_8_10, output_7_233;
mixer gate_output_7_233(.a(output_8_233), .b(output_8_10), .y(output_7_233));
wire output_9_233, output_9_10, output_8_233;
mixer gate_output_8_233(.a(output_9_233), .b(output_9_10), .y(output_8_233));
wire output_10_233, output_10_10, output_9_233;
mixer gate_output_9_233(.a(output_10_233), .b(output_10_10), .y(output_9_233));
wire output_11_233, output_11_10, output_10_233;
mixer gate_output_10_233(.a(output_11_233), .b(output_11_10), .y(output_10_233));
wire output_12_233, output_12_10, output_11_233;
mixer gate_output_11_233(.a(output_12_233), .b(output_12_10), .y(output_11_233));
wire output_13_233, output_13_10, output_12_233;
mixer gate_output_12_233(.a(output_13_233), .b(output_13_10), .y(output_12_233));
wire output_14_233, output_14_10, output_13_233;
mixer gate_output_13_233(.a(output_14_233), .b(output_14_10), .y(output_13_233));
wire output_15_233, output_15_10, output_14_233;
mixer gate_output_14_233(.a(output_15_233), .b(output_15_10), .y(output_14_233));
wire output_16_233, output_16_10, output_15_233;
mixer gate_output_15_233(.a(output_16_233), .b(output_16_10), .y(output_15_233));
wire output_1_234, output_1_11, output_0_234;
mixer gate_output_0_234(.a(output_1_234), .b(output_1_11), .y(output_0_234));
wire output_2_234, output_2_11, output_1_234;
mixer gate_output_1_234(.a(output_2_234), .b(output_2_11), .y(output_1_234));
wire output_3_234, output_3_11, output_2_234;
mixer gate_output_2_234(.a(output_3_234), .b(output_3_11), .y(output_2_234));
wire output_4_234, output_4_11, output_3_234;
mixer gate_output_3_234(.a(output_4_234), .b(output_4_11), .y(output_3_234));
wire output_5_234, output_5_11, output_4_234;
mixer gate_output_4_234(.a(output_5_234), .b(output_5_11), .y(output_4_234));
wire output_6_234, output_6_11, output_5_234;
mixer gate_output_5_234(.a(output_6_234), .b(output_6_11), .y(output_5_234));
wire output_7_234, output_7_11, output_6_234;
mixer gate_output_6_234(.a(output_7_234), .b(output_7_11), .y(output_6_234));
wire output_8_234, output_8_11, output_7_234;
mixer gate_output_7_234(.a(output_8_234), .b(output_8_11), .y(output_7_234));
wire output_9_234, output_9_11, output_8_234;
mixer gate_output_8_234(.a(output_9_234), .b(output_9_11), .y(output_8_234));
wire output_10_234, output_10_11, output_9_234;
mixer gate_output_9_234(.a(output_10_234), .b(output_10_11), .y(output_9_234));
wire output_11_234, output_11_11, output_10_234;
mixer gate_output_10_234(.a(output_11_234), .b(output_11_11), .y(output_10_234));
wire output_12_234, output_12_11, output_11_234;
mixer gate_output_11_234(.a(output_12_234), .b(output_12_11), .y(output_11_234));
wire output_13_234, output_13_11, output_12_234;
mixer gate_output_12_234(.a(output_13_234), .b(output_13_11), .y(output_12_234));
wire output_14_234, output_14_11, output_13_234;
mixer gate_output_13_234(.a(output_14_234), .b(output_14_11), .y(output_13_234));
wire output_15_234, output_15_11, output_14_234;
mixer gate_output_14_234(.a(output_15_234), .b(output_15_11), .y(output_14_234));
wire output_16_234, output_16_11, output_15_234;
mixer gate_output_15_234(.a(output_16_234), .b(output_16_11), .y(output_15_234));
wire output_1_235, output_1_12, output_0_235;
mixer gate_output_0_235(.a(output_1_235), .b(output_1_12), .y(output_0_235));
wire output_2_235, output_2_12, output_1_235;
mixer gate_output_1_235(.a(output_2_235), .b(output_2_12), .y(output_1_235));
wire output_3_235, output_3_12, output_2_235;
mixer gate_output_2_235(.a(output_3_235), .b(output_3_12), .y(output_2_235));
wire output_4_235, output_4_12, output_3_235;
mixer gate_output_3_235(.a(output_4_235), .b(output_4_12), .y(output_3_235));
wire output_5_235, output_5_12, output_4_235;
mixer gate_output_4_235(.a(output_5_235), .b(output_5_12), .y(output_4_235));
wire output_6_235, output_6_12, output_5_235;
mixer gate_output_5_235(.a(output_6_235), .b(output_6_12), .y(output_5_235));
wire output_7_235, output_7_12, output_6_235;
mixer gate_output_6_235(.a(output_7_235), .b(output_7_12), .y(output_6_235));
wire output_8_235, output_8_12, output_7_235;
mixer gate_output_7_235(.a(output_8_235), .b(output_8_12), .y(output_7_235));
wire output_9_235, output_9_12, output_8_235;
mixer gate_output_8_235(.a(output_9_235), .b(output_9_12), .y(output_8_235));
wire output_10_235, output_10_12, output_9_235;
mixer gate_output_9_235(.a(output_10_235), .b(output_10_12), .y(output_9_235));
wire output_11_235, output_11_12, output_10_235;
mixer gate_output_10_235(.a(output_11_235), .b(output_11_12), .y(output_10_235));
wire output_12_235, output_12_12, output_11_235;
mixer gate_output_11_235(.a(output_12_235), .b(output_12_12), .y(output_11_235));
wire output_13_235, output_13_12, output_12_235;
mixer gate_output_12_235(.a(output_13_235), .b(output_13_12), .y(output_12_235));
wire output_14_235, output_14_12, output_13_235;
mixer gate_output_13_235(.a(output_14_235), .b(output_14_12), .y(output_13_235));
wire output_15_235, output_15_12, output_14_235;
mixer gate_output_14_235(.a(output_15_235), .b(output_15_12), .y(output_14_235));
wire output_16_235, output_16_12, output_15_235;
mixer gate_output_15_235(.a(output_16_235), .b(output_16_12), .y(output_15_235));
wire output_1_236, output_1_13, output_0_236;
mixer gate_output_0_236(.a(output_1_236), .b(output_1_13), .y(output_0_236));
wire output_2_236, output_2_13, output_1_236;
mixer gate_output_1_236(.a(output_2_236), .b(output_2_13), .y(output_1_236));
wire output_3_236, output_3_13, output_2_236;
mixer gate_output_2_236(.a(output_3_236), .b(output_3_13), .y(output_2_236));
wire output_4_236, output_4_13, output_3_236;
mixer gate_output_3_236(.a(output_4_236), .b(output_4_13), .y(output_3_236));
wire output_5_236, output_5_13, output_4_236;
mixer gate_output_4_236(.a(output_5_236), .b(output_5_13), .y(output_4_236));
wire output_6_236, output_6_13, output_5_236;
mixer gate_output_5_236(.a(output_6_236), .b(output_6_13), .y(output_5_236));
wire output_7_236, output_7_13, output_6_236;
mixer gate_output_6_236(.a(output_7_236), .b(output_7_13), .y(output_6_236));
wire output_8_236, output_8_13, output_7_236;
mixer gate_output_7_236(.a(output_8_236), .b(output_8_13), .y(output_7_236));
wire output_9_236, output_9_13, output_8_236;
mixer gate_output_8_236(.a(output_9_236), .b(output_9_13), .y(output_8_236));
wire output_10_236, output_10_13, output_9_236;
mixer gate_output_9_236(.a(output_10_236), .b(output_10_13), .y(output_9_236));
wire output_11_236, output_11_13, output_10_236;
mixer gate_output_10_236(.a(output_11_236), .b(output_11_13), .y(output_10_236));
wire output_12_236, output_12_13, output_11_236;
mixer gate_output_11_236(.a(output_12_236), .b(output_12_13), .y(output_11_236));
wire output_13_236, output_13_13, output_12_236;
mixer gate_output_12_236(.a(output_13_236), .b(output_13_13), .y(output_12_236));
wire output_14_236, output_14_13, output_13_236;
mixer gate_output_13_236(.a(output_14_236), .b(output_14_13), .y(output_13_236));
wire output_15_236, output_15_13, output_14_236;
mixer gate_output_14_236(.a(output_15_236), .b(output_15_13), .y(output_14_236));
wire output_16_236, output_16_13, output_15_236;
mixer gate_output_15_236(.a(output_16_236), .b(output_16_13), .y(output_15_236));
wire output_1_237, output_1_14, output_0_237;
mixer gate_output_0_237(.a(output_1_237), .b(output_1_14), .y(output_0_237));
wire output_2_237, output_2_14, output_1_237;
mixer gate_output_1_237(.a(output_2_237), .b(output_2_14), .y(output_1_237));
wire output_3_237, output_3_14, output_2_237;
mixer gate_output_2_237(.a(output_3_237), .b(output_3_14), .y(output_2_237));
wire output_4_237, output_4_14, output_3_237;
mixer gate_output_3_237(.a(output_4_237), .b(output_4_14), .y(output_3_237));
wire output_5_237, output_5_14, output_4_237;
mixer gate_output_4_237(.a(output_5_237), .b(output_5_14), .y(output_4_237));
wire output_6_237, output_6_14, output_5_237;
mixer gate_output_5_237(.a(output_6_237), .b(output_6_14), .y(output_5_237));
wire output_7_237, output_7_14, output_6_237;
mixer gate_output_6_237(.a(output_7_237), .b(output_7_14), .y(output_6_237));
wire output_8_237, output_8_14, output_7_237;
mixer gate_output_7_237(.a(output_8_237), .b(output_8_14), .y(output_7_237));
wire output_9_237, output_9_14, output_8_237;
mixer gate_output_8_237(.a(output_9_237), .b(output_9_14), .y(output_8_237));
wire output_10_237, output_10_14, output_9_237;
mixer gate_output_9_237(.a(output_10_237), .b(output_10_14), .y(output_9_237));
wire output_11_237, output_11_14, output_10_237;
mixer gate_output_10_237(.a(output_11_237), .b(output_11_14), .y(output_10_237));
wire output_12_237, output_12_14, output_11_237;
mixer gate_output_11_237(.a(output_12_237), .b(output_12_14), .y(output_11_237));
wire output_13_237, output_13_14, output_12_237;
mixer gate_output_12_237(.a(output_13_237), .b(output_13_14), .y(output_12_237));
wire output_14_237, output_14_14, output_13_237;
mixer gate_output_13_237(.a(output_14_237), .b(output_14_14), .y(output_13_237));
wire output_15_237, output_15_14, output_14_237;
mixer gate_output_14_237(.a(output_15_237), .b(output_15_14), .y(output_14_237));
wire output_16_237, output_16_14, output_15_237;
mixer gate_output_15_237(.a(output_16_237), .b(output_16_14), .y(output_15_237));
wire output_1_238, output_1_15, output_0_238;
mixer gate_output_0_238(.a(output_1_238), .b(output_1_15), .y(output_0_238));
wire output_2_238, output_2_15, output_1_238;
mixer gate_output_1_238(.a(output_2_238), .b(output_2_15), .y(output_1_238));
wire output_3_238, output_3_15, output_2_238;
mixer gate_output_2_238(.a(output_3_238), .b(output_3_15), .y(output_2_238));
wire output_4_238, output_4_15, output_3_238;
mixer gate_output_3_238(.a(output_4_238), .b(output_4_15), .y(output_3_238));
wire output_5_238, output_5_15, output_4_238;
mixer gate_output_4_238(.a(output_5_238), .b(output_5_15), .y(output_4_238));
wire output_6_238, output_6_15, output_5_238;
mixer gate_output_5_238(.a(output_6_238), .b(output_6_15), .y(output_5_238));
wire output_7_238, output_7_15, output_6_238;
mixer gate_output_6_238(.a(output_7_238), .b(output_7_15), .y(output_6_238));
wire output_8_238, output_8_15, output_7_238;
mixer gate_output_7_238(.a(output_8_238), .b(output_8_15), .y(output_7_238));
wire output_9_238, output_9_15, output_8_238;
mixer gate_output_8_238(.a(output_9_238), .b(output_9_15), .y(output_8_238));
wire output_10_238, output_10_15, output_9_238;
mixer gate_output_9_238(.a(output_10_238), .b(output_10_15), .y(output_9_238));
wire output_11_238, output_11_15, output_10_238;
mixer gate_output_10_238(.a(output_11_238), .b(output_11_15), .y(output_10_238));
wire output_12_238, output_12_15, output_11_238;
mixer gate_output_11_238(.a(output_12_238), .b(output_12_15), .y(output_11_238));
wire output_13_238, output_13_15, output_12_238;
mixer gate_output_12_238(.a(output_13_238), .b(output_13_15), .y(output_12_238));
wire output_14_238, output_14_15, output_13_238;
mixer gate_output_13_238(.a(output_14_238), .b(output_14_15), .y(output_13_238));
wire output_15_238, output_15_15, output_14_238;
mixer gate_output_14_238(.a(output_15_238), .b(output_15_15), .y(output_14_238));
wire output_16_238, output_16_15, output_15_238;
mixer gate_output_15_238(.a(output_16_238), .b(output_16_15), .y(output_15_238));
wire output_1_239, output_1_0, output_0_239;
mixer gate_output_0_239(.a(output_1_239), .b(output_1_0), .y(output_0_239));
wire output_2_239, output_2_0, output_1_239;
mixer gate_output_1_239(.a(output_2_239), .b(output_2_0), .y(output_1_239));
wire output_3_239, output_3_0, output_2_239;
mixer gate_output_2_239(.a(output_3_239), .b(output_3_0), .y(output_2_239));
wire output_4_239, output_4_0, output_3_239;
mixer gate_output_3_239(.a(output_4_239), .b(output_4_0), .y(output_3_239));
wire output_5_239, output_5_0, output_4_239;
mixer gate_output_4_239(.a(output_5_239), .b(output_5_0), .y(output_4_239));
wire output_6_239, output_6_0, output_5_239;
mixer gate_output_5_239(.a(output_6_239), .b(output_6_0), .y(output_5_239));
wire output_7_239, output_7_0, output_6_239;
mixer gate_output_6_239(.a(output_7_239), .b(output_7_0), .y(output_6_239));
wire output_8_239, output_8_0, output_7_239;
mixer gate_output_7_239(.a(output_8_239), .b(output_8_0), .y(output_7_239));
wire output_9_239, output_9_0, output_8_239;
mixer gate_output_8_239(.a(output_9_239), .b(output_9_0), .y(output_8_239));
wire output_10_239, output_10_0, output_9_239;
mixer gate_output_9_239(.a(output_10_239), .b(output_10_0), .y(output_9_239));
wire output_11_239, output_11_0, output_10_239;
mixer gate_output_10_239(.a(output_11_239), .b(output_11_0), .y(output_10_239));
wire output_12_239, output_12_0, output_11_239;
mixer gate_output_11_239(.a(output_12_239), .b(output_12_0), .y(output_11_239));
wire output_13_239, output_13_0, output_12_239;
mixer gate_output_12_239(.a(output_13_239), .b(output_13_0), .y(output_12_239));
wire output_14_239, output_14_0, output_13_239;
mixer gate_output_13_239(.a(output_14_239), .b(output_14_0), .y(output_13_239));
wire output_15_239, output_15_0, output_14_239;
mixer gate_output_14_239(.a(output_15_239), .b(output_15_0), .y(output_14_239));
wire output_16_239, output_16_0, output_15_239;
mixer gate_output_15_239(.a(output_16_239), .b(output_16_0), .y(output_15_239));
wire output_1_240, output_1_1, output_0_240;
mixer gate_output_0_240(.a(output_1_240), .b(output_1_1), .y(output_0_240));
wire output_2_240, output_2_1, output_1_240;
mixer gate_output_1_240(.a(output_2_240), .b(output_2_1), .y(output_1_240));
wire output_3_240, output_3_1, output_2_240;
mixer gate_output_2_240(.a(output_3_240), .b(output_3_1), .y(output_2_240));
wire output_4_240, output_4_1, output_3_240;
mixer gate_output_3_240(.a(output_4_240), .b(output_4_1), .y(output_3_240));
wire output_5_240, output_5_1, output_4_240;
mixer gate_output_4_240(.a(output_5_240), .b(output_5_1), .y(output_4_240));
wire output_6_240, output_6_1, output_5_240;
mixer gate_output_5_240(.a(output_6_240), .b(output_6_1), .y(output_5_240));
wire output_7_240, output_7_1, output_6_240;
mixer gate_output_6_240(.a(output_7_240), .b(output_7_1), .y(output_6_240));
wire output_8_240, output_8_1, output_7_240;
mixer gate_output_7_240(.a(output_8_240), .b(output_8_1), .y(output_7_240));
wire output_9_240, output_9_1, output_8_240;
mixer gate_output_8_240(.a(output_9_240), .b(output_9_1), .y(output_8_240));
wire output_10_240, output_10_1, output_9_240;
mixer gate_output_9_240(.a(output_10_240), .b(output_10_1), .y(output_9_240));
wire output_11_240, output_11_1, output_10_240;
mixer gate_output_10_240(.a(output_11_240), .b(output_11_1), .y(output_10_240));
wire output_12_240, output_12_1, output_11_240;
mixer gate_output_11_240(.a(output_12_240), .b(output_12_1), .y(output_11_240));
wire output_13_240, output_13_1, output_12_240;
mixer gate_output_12_240(.a(output_13_240), .b(output_13_1), .y(output_12_240));
wire output_14_240, output_14_1, output_13_240;
mixer gate_output_13_240(.a(output_14_240), .b(output_14_1), .y(output_13_240));
wire output_15_240, output_15_1, output_14_240;
mixer gate_output_14_240(.a(output_15_240), .b(output_15_1), .y(output_14_240));
wire output_16_240, output_16_1, output_15_240;
mixer gate_output_15_240(.a(output_16_240), .b(output_16_1), .y(output_15_240));
wire output_1_241, output_1_2, output_0_241;
mixer gate_output_0_241(.a(output_1_241), .b(output_1_2), .y(output_0_241));
wire output_2_241, output_2_2, output_1_241;
mixer gate_output_1_241(.a(output_2_241), .b(output_2_2), .y(output_1_241));
wire output_3_241, output_3_2, output_2_241;
mixer gate_output_2_241(.a(output_3_241), .b(output_3_2), .y(output_2_241));
wire output_4_241, output_4_2, output_3_241;
mixer gate_output_3_241(.a(output_4_241), .b(output_4_2), .y(output_3_241));
wire output_5_241, output_5_2, output_4_241;
mixer gate_output_4_241(.a(output_5_241), .b(output_5_2), .y(output_4_241));
wire output_6_241, output_6_2, output_5_241;
mixer gate_output_5_241(.a(output_6_241), .b(output_6_2), .y(output_5_241));
wire output_7_241, output_7_2, output_6_241;
mixer gate_output_6_241(.a(output_7_241), .b(output_7_2), .y(output_6_241));
wire output_8_241, output_8_2, output_7_241;
mixer gate_output_7_241(.a(output_8_241), .b(output_8_2), .y(output_7_241));
wire output_9_241, output_9_2, output_8_241;
mixer gate_output_8_241(.a(output_9_241), .b(output_9_2), .y(output_8_241));
wire output_10_241, output_10_2, output_9_241;
mixer gate_output_9_241(.a(output_10_241), .b(output_10_2), .y(output_9_241));
wire output_11_241, output_11_2, output_10_241;
mixer gate_output_10_241(.a(output_11_241), .b(output_11_2), .y(output_10_241));
wire output_12_241, output_12_2, output_11_241;
mixer gate_output_11_241(.a(output_12_241), .b(output_12_2), .y(output_11_241));
wire output_13_241, output_13_2, output_12_241;
mixer gate_output_12_241(.a(output_13_241), .b(output_13_2), .y(output_12_241));
wire output_14_241, output_14_2, output_13_241;
mixer gate_output_13_241(.a(output_14_241), .b(output_14_2), .y(output_13_241));
wire output_15_241, output_15_2, output_14_241;
mixer gate_output_14_241(.a(output_15_241), .b(output_15_2), .y(output_14_241));
wire output_16_241, output_16_2, output_15_241;
mixer gate_output_15_241(.a(output_16_241), .b(output_16_2), .y(output_15_241));
wire output_1_242, output_1_3, output_0_242;
mixer gate_output_0_242(.a(output_1_242), .b(output_1_3), .y(output_0_242));
wire output_2_242, output_2_3, output_1_242;
mixer gate_output_1_242(.a(output_2_242), .b(output_2_3), .y(output_1_242));
wire output_3_242, output_3_3, output_2_242;
mixer gate_output_2_242(.a(output_3_242), .b(output_3_3), .y(output_2_242));
wire output_4_242, output_4_3, output_3_242;
mixer gate_output_3_242(.a(output_4_242), .b(output_4_3), .y(output_3_242));
wire output_5_242, output_5_3, output_4_242;
mixer gate_output_4_242(.a(output_5_242), .b(output_5_3), .y(output_4_242));
wire output_6_242, output_6_3, output_5_242;
mixer gate_output_5_242(.a(output_6_242), .b(output_6_3), .y(output_5_242));
wire output_7_242, output_7_3, output_6_242;
mixer gate_output_6_242(.a(output_7_242), .b(output_7_3), .y(output_6_242));
wire output_8_242, output_8_3, output_7_242;
mixer gate_output_7_242(.a(output_8_242), .b(output_8_3), .y(output_7_242));
wire output_9_242, output_9_3, output_8_242;
mixer gate_output_8_242(.a(output_9_242), .b(output_9_3), .y(output_8_242));
wire output_10_242, output_10_3, output_9_242;
mixer gate_output_9_242(.a(output_10_242), .b(output_10_3), .y(output_9_242));
wire output_11_242, output_11_3, output_10_242;
mixer gate_output_10_242(.a(output_11_242), .b(output_11_3), .y(output_10_242));
wire output_12_242, output_12_3, output_11_242;
mixer gate_output_11_242(.a(output_12_242), .b(output_12_3), .y(output_11_242));
wire output_13_242, output_13_3, output_12_242;
mixer gate_output_12_242(.a(output_13_242), .b(output_13_3), .y(output_12_242));
wire output_14_242, output_14_3, output_13_242;
mixer gate_output_13_242(.a(output_14_242), .b(output_14_3), .y(output_13_242));
wire output_15_242, output_15_3, output_14_242;
mixer gate_output_14_242(.a(output_15_242), .b(output_15_3), .y(output_14_242));
wire output_16_242, output_16_3, output_15_242;
mixer gate_output_15_242(.a(output_16_242), .b(output_16_3), .y(output_15_242));
wire output_1_243, output_1_4, output_0_243;
mixer gate_output_0_243(.a(output_1_243), .b(output_1_4), .y(output_0_243));
wire output_2_243, output_2_4, output_1_243;
mixer gate_output_1_243(.a(output_2_243), .b(output_2_4), .y(output_1_243));
wire output_3_243, output_3_4, output_2_243;
mixer gate_output_2_243(.a(output_3_243), .b(output_3_4), .y(output_2_243));
wire output_4_243, output_4_4, output_3_243;
mixer gate_output_3_243(.a(output_4_243), .b(output_4_4), .y(output_3_243));
wire output_5_243, output_5_4, output_4_243;
mixer gate_output_4_243(.a(output_5_243), .b(output_5_4), .y(output_4_243));
wire output_6_243, output_6_4, output_5_243;
mixer gate_output_5_243(.a(output_6_243), .b(output_6_4), .y(output_5_243));
wire output_7_243, output_7_4, output_6_243;
mixer gate_output_6_243(.a(output_7_243), .b(output_7_4), .y(output_6_243));
wire output_8_243, output_8_4, output_7_243;
mixer gate_output_7_243(.a(output_8_243), .b(output_8_4), .y(output_7_243));
wire output_9_243, output_9_4, output_8_243;
mixer gate_output_8_243(.a(output_9_243), .b(output_9_4), .y(output_8_243));
wire output_10_243, output_10_4, output_9_243;
mixer gate_output_9_243(.a(output_10_243), .b(output_10_4), .y(output_9_243));
wire output_11_243, output_11_4, output_10_243;
mixer gate_output_10_243(.a(output_11_243), .b(output_11_4), .y(output_10_243));
wire output_12_243, output_12_4, output_11_243;
mixer gate_output_11_243(.a(output_12_243), .b(output_12_4), .y(output_11_243));
wire output_13_243, output_13_4, output_12_243;
mixer gate_output_12_243(.a(output_13_243), .b(output_13_4), .y(output_12_243));
wire output_14_243, output_14_4, output_13_243;
mixer gate_output_13_243(.a(output_14_243), .b(output_14_4), .y(output_13_243));
wire output_15_243, output_15_4, output_14_243;
mixer gate_output_14_243(.a(output_15_243), .b(output_15_4), .y(output_14_243));
wire output_16_243, output_16_4, output_15_243;
mixer gate_output_15_243(.a(output_16_243), .b(output_16_4), .y(output_15_243));
wire output_1_244, output_1_5, output_0_244;
mixer gate_output_0_244(.a(output_1_244), .b(output_1_5), .y(output_0_244));
wire output_2_244, output_2_5, output_1_244;
mixer gate_output_1_244(.a(output_2_244), .b(output_2_5), .y(output_1_244));
wire output_3_244, output_3_5, output_2_244;
mixer gate_output_2_244(.a(output_3_244), .b(output_3_5), .y(output_2_244));
wire output_4_244, output_4_5, output_3_244;
mixer gate_output_3_244(.a(output_4_244), .b(output_4_5), .y(output_3_244));
wire output_5_244, output_5_5, output_4_244;
mixer gate_output_4_244(.a(output_5_244), .b(output_5_5), .y(output_4_244));
wire output_6_244, output_6_5, output_5_244;
mixer gate_output_5_244(.a(output_6_244), .b(output_6_5), .y(output_5_244));
wire output_7_244, output_7_5, output_6_244;
mixer gate_output_6_244(.a(output_7_244), .b(output_7_5), .y(output_6_244));
wire output_8_244, output_8_5, output_7_244;
mixer gate_output_7_244(.a(output_8_244), .b(output_8_5), .y(output_7_244));
wire output_9_244, output_9_5, output_8_244;
mixer gate_output_8_244(.a(output_9_244), .b(output_9_5), .y(output_8_244));
wire output_10_244, output_10_5, output_9_244;
mixer gate_output_9_244(.a(output_10_244), .b(output_10_5), .y(output_9_244));
wire output_11_244, output_11_5, output_10_244;
mixer gate_output_10_244(.a(output_11_244), .b(output_11_5), .y(output_10_244));
wire output_12_244, output_12_5, output_11_244;
mixer gate_output_11_244(.a(output_12_244), .b(output_12_5), .y(output_11_244));
wire output_13_244, output_13_5, output_12_244;
mixer gate_output_12_244(.a(output_13_244), .b(output_13_5), .y(output_12_244));
wire output_14_244, output_14_5, output_13_244;
mixer gate_output_13_244(.a(output_14_244), .b(output_14_5), .y(output_13_244));
wire output_15_244, output_15_5, output_14_244;
mixer gate_output_14_244(.a(output_15_244), .b(output_15_5), .y(output_14_244));
wire output_16_244, output_16_5, output_15_244;
mixer gate_output_15_244(.a(output_16_244), .b(output_16_5), .y(output_15_244));
wire output_1_245, output_1_6, output_0_245;
mixer gate_output_0_245(.a(output_1_245), .b(output_1_6), .y(output_0_245));
wire output_2_245, output_2_6, output_1_245;
mixer gate_output_1_245(.a(output_2_245), .b(output_2_6), .y(output_1_245));
wire output_3_245, output_3_6, output_2_245;
mixer gate_output_2_245(.a(output_3_245), .b(output_3_6), .y(output_2_245));
wire output_4_245, output_4_6, output_3_245;
mixer gate_output_3_245(.a(output_4_245), .b(output_4_6), .y(output_3_245));
wire output_5_245, output_5_6, output_4_245;
mixer gate_output_4_245(.a(output_5_245), .b(output_5_6), .y(output_4_245));
wire output_6_245, output_6_6, output_5_245;
mixer gate_output_5_245(.a(output_6_245), .b(output_6_6), .y(output_5_245));
wire output_7_245, output_7_6, output_6_245;
mixer gate_output_6_245(.a(output_7_245), .b(output_7_6), .y(output_6_245));
wire output_8_245, output_8_6, output_7_245;
mixer gate_output_7_245(.a(output_8_245), .b(output_8_6), .y(output_7_245));
wire output_9_245, output_9_6, output_8_245;
mixer gate_output_8_245(.a(output_9_245), .b(output_9_6), .y(output_8_245));
wire output_10_245, output_10_6, output_9_245;
mixer gate_output_9_245(.a(output_10_245), .b(output_10_6), .y(output_9_245));
wire output_11_245, output_11_6, output_10_245;
mixer gate_output_10_245(.a(output_11_245), .b(output_11_6), .y(output_10_245));
wire output_12_245, output_12_6, output_11_245;
mixer gate_output_11_245(.a(output_12_245), .b(output_12_6), .y(output_11_245));
wire output_13_245, output_13_6, output_12_245;
mixer gate_output_12_245(.a(output_13_245), .b(output_13_6), .y(output_12_245));
wire output_14_245, output_14_6, output_13_245;
mixer gate_output_13_245(.a(output_14_245), .b(output_14_6), .y(output_13_245));
wire output_15_245, output_15_6, output_14_245;
mixer gate_output_14_245(.a(output_15_245), .b(output_15_6), .y(output_14_245));
wire output_16_245, output_16_6, output_15_245;
mixer gate_output_15_245(.a(output_16_245), .b(output_16_6), .y(output_15_245));
wire output_1_246, output_1_7, output_0_246;
mixer gate_output_0_246(.a(output_1_246), .b(output_1_7), .y(output_0_246));
wire output_2_246, output_2_7, output_1_246;
mixer gate_output_1_246(.a(output_2_246), .b(output_2_7), .y(output_1_246));
wire output_3_246, output_3_7, output_2_246;
mixer gate_output_2_246(.a(output_3_246), .b(output_3_7), .y(output_2_246));
wire output_4_246, output_4_7, output_3_246;
mixer gate_output_3_246(.a(output_4_246), .b(output_4_7), .y(output_3_246));
wire output_5_246, output_5_7, output_4_246;
mixer gate_output_4_246(.a(output_5_246), .b(output_5_7), .y(output_4_246));
wire output_6_246, output_6_7, output_5_246;
mixer gate_output_5_246(.a(output_6_246), .b(output_6_7), .y(output_5_246));
wire output_7_246, output_7_7, output_6_246;
mixer gate_output_6_246(.a(output_7_246), .b(output_7_7), .y(output_6_246));
wire output_8_246, output_8_7, output_7_246;
mixer gate_output_7_246(.a(output_8_246), .b(output_8_7), .y(output_7_246));
wire output_9_246, output_9_7, output_8_246;
mixer gate_output_8_246(.a(output_9_246), .b(output_9_7), .y(output_8_246));
wire output_10_246, output_10_7, output_9_246;
mixer gate_output_9_246(.a(output_10_246), .b(output_10_7), .y(output_9_246));
wire output_11_246, output_11_7, output_10_246;
mixer gate_output_10_246(.a(output_11_246), .b(output_11_7), .y(output_10_246));
wire output_12_246, output_12_7, output_11_246;
mixer gate_output_11_246(.a(output_12_246), .b(output_12_7), .y(output_11_246));
wire output_13_246, output_13_7, output_12_246;
mixer gate_output_12_246(.a(output_13_246), .b(output_13_7), .y(output_12_246));
wire output_14_246, output_14_7, output_13_246;
mixer gate_output_13_246(.a(output_14_246), .b(output_14_7), .y(output_13_246));
wire output_15_246, output_15_7, output_14_246;
mixer gate_output_14_246(.a(output_15_246), .b(output_15_7), .y(output_14_246));
wire output_16_246, output_16_7, output_15_246;
mixer gate_output_15_246(.a(output_16_246), .b(output_16_7), .y(output_15_246));
wire output_1_247, output_1_8, output_0_247;
mixer gate_output_0_247(.a(output_1_247), .b(output_1_8), .y(output_0_247));
wire output_2_247, output_2_8, output_1_247;
mixer gate_output_1_247(.a(output_2_247), .b(output_2_8), .y(output_1_247));
wire output_3_247, output_3_8, output_2_247;
mixer gate_output_2_247(.a(output_3_247), .b(output_3_8), .y(output_2_247));
wire output_4_247, output_4_8, output_3_247;
mixer gate_output_3_247(.a(output_4_247), .b(output_4_8), .y(output_3_247));
wire output_5_247, output_5_8, output_4_247;
mixer gate_output_4_247(.a(output_5_247), .b(output_5_8), .y(output_4_247));
wire output_6_247, output_6_8, output_5_247;
mixer gate_output_5_247(.a(output_6_247), .b(output_6_8), .y(output_5_247));
wire output_7_247, output_7_8, output_6_247;
mixer gate_output_6_247(.a(output_7_247), .b(output_7_8), .y(output_6_247));
wire output_8_247, output_8_8, output_7_247;
mixer gate_output_7_247(.a(output_8_247), .b(output_8_8), .y(output_7_247));
wire output_9_247, output_9_8, output_8_247;
mixer gate_output_8_247(.a(output_9_247), .b(output_9_8), .y(output_8_247));
wire output_10_247, output_10_8, output_9_247;
mixer gate_output_9_247(.a(output_10_247), .b(output_10_8), .y(output_9_247));
wire output_11_247, output_11_8, output_10_247;
mixer gate_output_10_247(.a(output_11_247), .b(output_11_8), .y(output_10_247));
wire output_12_247, output_12_8, output_11_247;
mixer gate_output_11_247(.a(output_12_247), .b(output_12_8), .y(output_11_247));
wire output_13_247, output_13_8, output_12_247;
mixer gate_output_12_247(.a(output_13_247), .b(output_13_8), .y(output_12_247));
wire output_14_247, output_14_8, output_13_247;
mixer gate_output_13_247(.a(output_14_247), .b(output_14_8), .y(output_13_247));
wire output_15_247, output_15_8, output_14_247;
mixer gate_output_14_247(.a(output_15_247), .b(output_15_8), .y(output_14_247));
wire output_16_247, output_16_8, output_15_247;
mixer gate_output_15_247(.a(output_16_247), .b(output_16_8), .y(output_15_247));
wire output_1_248, output_1_9, output_0_248;
mixer gate_output_0_248(.a(output_1_248), .b(output_1_9), .y(output_0_248));
wire output_2_248, output_2_9, output_1_248;
mixer gate_output_1_248(.a(output_2_248), .b(output_2_9), .y(output_1_248));
wire output_3_248, output_3_9, output_2_248;
mixer gate_output_2_248(.a(output_3_248), .b(output_3_9), .y(output_2_248));
wire output_4_248, output_4_9, output_3_248;
mixer gate_output_3_248(.a(output_4_248), .b(output_4_9), .y(output_3_248));
wire output_5_248, output_5_9, output_4_248;
mixer gate_output_4_248(.a(output_5_248), .b(output_5_9), .y(output_4_248));
wire output_6_248, output_6_9, output_5_248;
mixer gate_output_5_248(.a(output_6_248), .b(output_6_9), .y(output_5_248));
wire output_7_248, output_7_9, output_6_248;
mixer gate_output_6_248(.a(output_7_248), .b(output_7_9), .y(output_6_248));
wire output_8_248, output_8_9, output_7_248;
mixer gate_output_7_248(.a(output_8_248), .b(output_8_9), .y(output_7_248));
wire output_9_248, output_9_9, output_8_248;
mixer gate_output_8_248(.a(output_9_248), .b(output_9_9), .y(output_8_248));
wire output_10_248, output_10_9, output_9_248;
mixer gate_output_9_248(.a(output_10_248), .b(output_10_9), .y(output_9_248));
wire output_11_248, output_11_9, output_10_248;
mixer gate_output_10_248(.a(output_11_248), .b(output_11_9), .y(output_10_248));
wire output_12_248, output_12_9, output_11_248;
mixer gate_output_11_248(.a(output_12_248), .b(output_12_9), .y(output_11_248));
wire output_13_248, output_13_9, output_12_248;
mixer gate_output_12_248(.a(output_13_248), .b(output_13_9), .y(output_12_248));
wire output_14_248, output_14_9, output_13_248;
mixer gate_output_13_248(.a(output_14_248), .b(output_14_9), .y(output_13_248));
wire output_15_248, output_15_9, output_14_248;
mixer gate_output_14_248(.a(output_15_248), .b(output_15_9), .y(output_14_248));
wire output_16_248, output_16_9, output_15_248;
mixer gate_output_15_248(.a(output_16_248), .b(output_16_9), .y(output_15_248));
wire output_1_249, output_1_10, output_0_249;
mixer gate_output_0_249(.a(output_1_249), .b(output_1_10), .y(output_0_249));
wire output_2_249, output_2_10, output_1_249;
mixer gate_output_1_249(.a(output_2_249), .b(output_2_10), .y(output_1_249));
wire output_3_249, output_3_10, output_2_249;
mixer gate_output_2_249(.a(output_3_249), .b(output_3_10), .y(output_2_249));
wire output_4_249, output_4_10, output_3_249;
mixer gate_output_3_249(.a(output_4_249), .b(output_4_10), .y(output_3_249));
wire output_5_249, output_5_10, output_4_249;
mixer gate_output_4_249(.a(output_5_249), .b(output_5_10), .y(output_4_249));
wire output_6_249, output_6_10, output_5_249;
mixer gate_output_5_249(.a(output_6_249), .b(output_6_10), .y(output_5_249));
wire output_7_249, output_7_10, output_6_249;
mixer gate_output_6_249(.a(output_7_249), .b(output_7_10), .y(output_6_249));
wire output_8_249, output_8_10, output_7_249;
mixer gate_output_7_249(.a(output_8_249), .b(output_8_10), .y(output_7_249));
wire output_9_249, output_9_10, output_8_249;
mixer gate_output_8_249(.a(output_9_249), .b(output_9_10), .y(output_8_249));
wire output_10_249, output_10_10, output_9_249;
mixer gate_output_9_249(.a(output_10_249), .b(output_10_10), .y(output_9_249));
wire output_11_249, output_11_10, output_10_249;
mixer gate_output_10_249(.a(output_11_249), .b(output_11_10), .y(output_10_249));
wire output_12_249, output_12_10, output_11_249;
mixer gate_output_11_249(.a(output_12_249), .b(output_12_10), .y(output_11_249));
wire output_13_249, output_13_10, output_12_249;
mixer gate_output_12_249(.a(output_13_249), .b(output_13_10), .y(output_12_249));
wire output_14_249, output_14_10, output_13_249;
mixer gate_output_13_249(.a(output_14_249), .b(output_14_10), .y(output_13_249));
wire output_15_249, output_15_10, output_14_249;
mixer gate_output_14_249(.a(output_15_249), .b(output_15_10), .y(output_14_249));
wire output_16_249, output_16_10, output_15_249;
mixer gate_output_15_249(.a(output_16_249), .b(output_16_10), .y(output_15_249));
wire output_1_250, output_1_11, output_0_250;
mixer gate_output_0_250(.a(output_1_250), .b(output_1_11), .y(output_0_250));
wire output_2_250, output_2_11, output_1_250;
mixer gate_output_1_250(.a(output_2_250), .b(output_2_11), .y(output_1_250));
wire output_3_250, output_3_11, output_2_250;
mixer gate_output_2_250(.a(output_3_250), .b(output_3_11), .y(output_2_250));
wire output_4_250, output_4_11, output_3_250;
mixer gate_output_3_250(.a(output_4_250), .b(output_4_11), .y(output_3_250));
wire output_5_250, output_5_11, output_4_250;
mixer gate_output_4_250(.a(output_5_250), .b(output_5_11), .y(output_4_250));
wire output_6_250, output_6_11, output_5_250;
mixer gate_output_5_250(.a(output_6_250), .b(output_6_11), .y(output_5_250));
wire output_7_250, output_7_11, output_6_250;
mixer gate_output_6_250(.a(output_7_250), .b(output_7_11), .y(output_6_250));
wire output_8_250, output_8_11, output_7_250;
mixer gate_output_7_250(.a(output_8_250), .b(output_8_11), .y(output_7_250));
wire output_9_250, output_9_11, output_8_250;
mixer gate_output_8_250(.a(output_9_250), .b(output_9_11), .y(output_8_250));
wire output_10_250, output_10_11, output_9_250;
mixer gate_output_9_250(.a(output_10_250), .b(output_10_11), .y(output_9_250));
wire output_11_250, output_11_11, output_10_250;
mixer gate_output_10_250(.a(output_11_250), .b(output_11_11), .y(output_10_250));
wire output_12_250, output_12_11, output_11_250;
mixer gate_output_11_250(.a(output_12_250), .b(output_12_11), .y(output_11_250));
wire output_13_250, output_13_11, output_12_250;
mixer gate_output_12_250(.a(output_13_250), .b(output_13_11), .y(output_12_250));
wire output_14_250, output_14_11, output_13_250;
mixer gate_output_13_250(.a(output_14_250), .b(output_14_11), .y(output_13_250));
wire output_15_250, output_15_11, output_14_250;
mixer gate_output_14_250(.a(output_15_250), .b(output_15_11), .y(output_14_250));
wire output_16_250, output_16_11, output_15_250;
mixer gate_output_15_250(.a(output_16_250), .b(output_16_11), .y(output_15_250));
wire output_1_251, output_1_12, output_0_251;
mixer gate_output_0_251(.a(output_1_251), .b(output_1_12), .y(output_0_251));
wire output_2_251, output_2_12, output_1_251;
mixer gate_output_1_251(.a(output_2_251), .b(output_2_12), .y(output_1_251));
wire output_3_251, output_3_12, output_2_251;
mixer gate_output_2_251(.a(output_3_251), .b(output_3_12), .y(output_2_251));
wire output_4_251, output_4_12, output_3_251;
mixer gate_output_3_251(.a(output_4_251), .b(output_4_12), .y(output_3_251));
wire output_5_251, output_5_12, output_4_251;
mixer gate_output_4_251(.a(output_5_251), .b(output_5_12), .y(output_4_251));
wire output_6_251, output_6_12, output_5_251;
mixer gate_output_5_251(.a(output_6_251), .b(output_6_12), .y(output_5_251));
wire output_7_251, output_7_12, output_6_251;
mixer gate_output_6_251(.a(output_7_251), .b(output_7_12), .y(output_6_251));
wire output_8_251, output_8_12, output_7_251;
mixer gate_output_7_251(.a(output_8_251), .b(output_8_12), .y(output_7_251));
wire output_9_251, output_9_12, output_8_251;
mixer gate_output_8_251(.a(output_9_251), .b(output_9_12), .y(output_8_251));
wire output_10_251, output_10_12, output_9_251;
mixer gate_output_9_251(.a(output_10_251), .b(output_10_12), .y(output_9_251));
wire output_11_251, output_11_12, output_10_251;
mixer gate_output_10_251(.a(output_11_251), .b(output_11_12), .y(output_10_251));
wire output_12_251, output_12_12, output_11_251;
mixer gate_output_11_251(.a(output_12_251), .b(output_12_12), .y(output_11_251));
wire output_13_251, output_13_12, output_12_251;
mixer gate_output_12_251(.a(output_13_251), .b(output_13_12), .y(output_12_251));
wire output_14_251, output_14_12, output_13_251;
mixer gate_output_13_251(.a(output_14_251), .b(output_14_12), .y(output_13_251));
wire output_15_251, output_15_12, output_14_251;
mixer gate_output_14_251(.a(output_15_251), .b(output_15_12), .y(output_14_251));
wire output_16_251, output_16_12, output_15_251;
mixer gate_output_15_251(.a(output_16_251), .b(output_16_12), .y(output_15_251));
wire output_1_252, output_1_13, output_0_252;
mixer gate_output_0_252(.a(output_1_252), .b(output_1_13), .y(output_0_252));
wire output_2_252, output_2_13, output_1_252;
mixer gate_output_1_252(.a(output_2_252), .b(output_2_13), .y(output_1_252));
wire output_3_252, output_3_13, output_2_252;
mixer gate_output_2_252(.a(output_3_252), .b(output_3_13), .y(output_2_252));
wire output_4_252, output_4_13, output_3_252;
mixer gate_output_3_252(.a(output_4_252), .b(output_4_13), .y(output_3_252));
wire output_5_252, output_5_13, output_4_252;
mixer gate_output_4_252(.a(output_5_252), .b(output_5_13), .y(output_4_252));
wire output_6_252, output_6_13, output_5_252;
mixer gate_output_5_252(.a(output_6_252), .b(output_6_13), .y(output_5_252));
wire output_7_252, output_7_13, output_6_252;
mixer gate_output_6_252(.a(output_7_252), .b(output_7_13), .y(output_6_252));
wire output_8_252, output_8_13, output_7_252;
mixer gate_output_7_252(.a(output_8_252), .b(output_8_13), .y(output_7_252));
wire output_9_252, output_9_13, output_8_252;
mixer gate_output_8_252(.a(output_9_252), .b(output_9_13), .y(output_8_252));
wire output_10_252, output_10_13, output_9_252;
mixer gate_output_9_252(.a(output_10_252), .b(output_10_13), .y(output_9_252));
wire output_11_252, output_11_13, output_10_252;
mixer gate_output_10_252(.a(output_11_252), .b(output_11_13), .y(output_10_252));
wire output_12_252, output_12_13, output_11_252;
mixer gate_output_11_252(.a(output_12_252), .b(output_12_13), .y(output_11_252));
wire output_13_252, output_13_13, output_12_252;
mixer gate_output_12_252(.a(output_13_252), .b(output_13_13), .y(output_12_252));
wire output_14_252, output_14_13, output_13_252;
mixer gate_output_13_252(.a(output_14_252), .b(output_14_13), .y(output_13_252));
wire output_15_252, output_15_13, output_14_252;
mixer gate_output_14_252(.a(output_15_252), .b(output_15_13), .y(output_14_252));
wire output_16_252, output_16_13, output_15_252;
mixer gate_output_15_252(.a(output_16_252), .b(output_16_13), .y(output_15_252));
wire output_1_253, output_1_14, output_0_253;
mixer gate_output_0_253(.a(output_1_253), .b(output_1_14), .y(output_0_253));
wire output_2_253, output_2_14, output_1_253;
mixer gate_output_1_253(.a(output_2_253), .b(output_2_14), .y(output_1_253));
wire output_3_253, output_3_14, output_2_253;
mixer gate_output_2_253(.a(output_3_253), .b(output_3_14), .y(output_2_253));
wire output_4_253, output_4_14, output_3_253;
mixer gate_output_3_253(.a(output_4_253), .b(output_4_14), .y(output_3_253));
wire output_5_253, output_5_14, output_4_253;
mixer gate_output_4_253(.a(output_5_253), .b(output_5_14), .y(output_4_253));
wire output_6_253, output_6_14, output_5_253;
mixer gate_output_5_253(.a(output_6_253), .b(output_6_14), .y(output_5_253));
wire output_7_253, output_7_14, output_6_253;
mixer gate_output_6_253(.a(output_7_253), .b(output_7_14), .y(output_6_253));
wire output_8_253, output_8_14, output_7_253;
mixer gate_output_7_253(.a(output_8_253), .b(output_8_14), .y(output_7_253));
wire output_9_253, output_9_14, output_8_253;
mixer gate_output_8_253(.a(output_9_253), .b(output_9_14), .y(output_8_253));
wire output_10_253, output_10_14, output_9_253;
mixer gate_output_9_253(.a(output_10_253), .b(output_10_14), .y(output_9_253));
wire output_11_253, output_11_14, output_10_253;
mixer gate_output_10_253(.a(output_11_253), .b(output_11_14), .y(output_10_253));
wire output_12_253, output_12_14, output_11_253;
mixer gate_output_11_253(.a(output_12_253), .b(output_12_14), .y(output_11_253));
wire output_13_253, output_13_14, output_12_253;
mixer gate_output_12_253(.a(output_13_253), .b(output_13_14), .y(output_12_253));
wire output_14_253, output_14_14, output_13_253;
mixer gate_output_13_253(.a(output_14_253), .b(output_14_14), .y(output_13_253));
wire output_15_253, output_15_14, output_14_253;
mixer gate_output_14_253(.a(output_15_253), .b(output_15_14), .y(output_14_253));
wire output_16_253, output_16_14, output_15_253;
mixer gate_output_15_253(.a(output_16_253), .b(output_16_14), .y(output_15_253));
wire output_1_254, output_1_15, output_0_254;
mixer gate_output_0_254(.a(output_1_254), .b(output_1_15), .y(output_0_254));
wire output_2_254, output_2_15, output_1_254;
mixer gate_output_1_254(.a(output_2_254), .b(output_2_15), .y(output_1_254));
wire output_3_254, output_3_15, output_2_254;
mixer gate_output_2_254(.a(output_3_254), .b(output_3_15), .y(output_2_254));
wire output_4_254, output_4_15, output_3_254;
mixer gate_output_3_254(.a(output_4_254), .b(output_4_15), .y(output_3_254));
wire output_5_254, output_5_15, output_4_254;
mixer gate_output_4_254(.a(output_5_254), .b(output_5_15), .y(output_4_254));
wire output_6_254, output_6_15, output_5_254;
mixer gate_output_5_254(.a(output_6_254), .b(output_6_15), .y(output_5_254));
wire output_7_254, output_7_15, output_6_254;
mixer gate_output_6_254(.a(output_7_254), .b(output_7_15), .y(output_6_254));
wire output_8_254, output_8_15, output_7_254;
mixer gate_output_7_254(.a(output_8_254), .b(output_8_15), .y(output_7_254));
wire output_9_254, output_9_15, output_8_254;
mixer gate_output_8_254(.a(output_9_254), .b(output_9_15), .y(output_8_254));
wire output_10_254, output_10_15, output_9_254;
mixer gate_output_9_254(.a(output_10_254), .b(output_10_15), .y(output_9_254));
wire output_11_254, output_11_15, output_10_254;
mixer gate_output_10_254(.a(output_11_254), .b(output_11_15), .y(output_10_254));
wire output_12_254, output_12_15, output_11_254;
mixer gate_output_11_254(.a(output_12_254), .b(output_12_15), .y(output_11_254));
wire output_13_254, output_13_15, output_12_254;
mixer gate_output_12_254(.a(output_13_254), .b(output_13_15), .y(output_12_254));
wire output_14_254, output_14_15, output_13_254;
mixer gate_output_13_254(.a(output_14_254), .b(output_14_15), .y(output_13_254));
wire output_15_254, output_15_15, output_14_254;
mixer gate_output_14_254(.a(output_15_254), .b(output_15_15), .y(output_14_254));
wire output_16_254, output_16_15, output_15_254;
mixer gate_output_15_254(.a(output_16_254), .b(output_16_15), .y(output_15_254));
wire output_1_255, output_1_0, output_0_255;
mixer gate_output_0_255(.a(output_1_255), .b(output_1_0), .y(output_0_255));
wire output_2_255, output_2_0, output_1_255;
mixer gate_output_1_255(.a(output_2_255), .b(output_2_0), .y(output_1_255));
wire output_3_255, output_3_0, output_2_255;
mixer gate_output_2_255(.a(output_3_255), .b(output_3_0), .y(output_2_255));
wire output_4_255, output_4_0, output_3_255;
mixer gate_output_3_255(.a(output_4_255), .b(output_4_0), .y(output_3_255));
wire output_5_255, output_5_0, output_4_255;
mixer gate_output_4_255(.a(output_5_255), .b(output_5_0), .y(output_4_255));
wire output_6_255, output_6_0, output_5_255;
mixer gate_output_5_255(.a(output_6_255), .b(output_6_0), .y(output_5_255));
wire output_7_255, output_7_0, output_6_255;
mixer gate_output_6_255(.a(output_7_255), .b(output_7_0), .y(output_6_255));
wire output_8_255, output_8_0, output_7_255;
mixer gate_output_7_255(.a(output_8_255), .b(output_8_0), .y(output_7_255));
wire output_9_255, output_9_0, output_8_255;
mixer gate_output_8_255(.a(output_9_255), .b(output_9_0), .y(output_8_255));
wire output_10_255, output_10_0, output_9_255;
mixer gate_output_9_255(.a(output_10_255), .b(output_10_0), .y(output_9_255));
wire output_11_255, output_11_0, output_10_255;
mixer gate_output_10_255(.a(output_11_255), .b(output_11_0), .y(output_10_255));
wire output_12_255, output_12_0, output_11_255;
mixer gate_output_11_255(.a(output_12_255), .b(output_12_0), .y(output_11_255));
wire output_13_255, output_13_0, output_12_255;
mixer gate_output_12_255(.a(output_13_255), .b(output_13_0), .y(output_12_255));
wire output_14_255, output_14_0, output_13_255;
mixer gate_output_13_255(.a(output_14_255), .b(output_14_0), .y(output_13_255));
wire output_15_255, output_15_0, output_14_255;
mixer gate_output_14_255(.a(output_15_255), .b(output_15_0), .y(output_14_255));
wire output_16_255, output_16_0, output_15_255;
mixer gate_output_15_255(.a(output_16_255), .b(output_16_0), .y(output_15_255));
wire output_1_256, output_1_1, output_0_256;
mixer gate_output_0_256(.a(output_1_256), .b(output_1_1), .y(output_0_256));
wire output_2_256, output_2_1, output_1_256;
mixer gate_output_1_256(.a(output_2_256), .b(output_2_1), .y(output_1_256));
wire output_3_256, output_3_1, output_2_256;
mixer gate_output_2_256(.a(output_3_256), .b(output_3_1), .y(output_2_256));
wire output_4_256, output_4_1, output_3_256;
mixer gate_output_3_256(.a(output_4_256), .b(output_4_1), .y(output_3_256));
wire output_5_256, output_5_1, output_4_256;
mixer gate_output_4_256(.a(output_5_256), .b(output_5_1), .y(output_4_256));
wire output_6_256, output_6_1, output_5_256;
mixer gate_output_5_256(.a(output_6_256), .b(output_6_1), .y(output_5_256));
wire output_7_256, output_7_1, output_6_256;
mixer gate_output_6_256(.a(output_7_256), .b(output_7_1), .y(output_6_256));
wire output_8_256, output_8_1, output_7_256;
mixer gate_output_7_256(.a(output_8_256), .b(output_8_1), .y(output_7_256));
wire output_9_256, output_9_1, output_8_256;
mixer gate_output_8_256(.a(output_9_256), .b(output_9_1), .y(output_8_256));
wire output_10_256, output_10_1, output_9_256;
mixer gate_output_9_256(.a(output_10_256), .b(output_10_1), .y(output_9_256));
wire output_11_256, output_11_1, output_10_256;
mixer gate_output_10_256(.a(output_11_256), .b(output_11_1), .y(output_10_256));
wire output_12_256, output_12_1, output_11_256;
mixer gate_output_11_256(.a(output_12_256), .b(output_12_1), .y(output_11_256));
wire output_13_256, output_13_1, output_12_256;
mixer gate_output_12_256(.a(output_13_256), .b(output_13_1), .y(output_12_256));
wire output_14_256, output_14_1, output_13_256;
mixer gate_output_13_256(.a(output_14_256), .b(output_14_1), .y(output_13_256));
wire output_15_256, output_15_1, output_14_256;
mixer gate_output_14_256(.a(output_15_256), .b(output_15_1), .y(output_14_256));
wire output_16_256, output_16_1, output_15_256;
mixer gate_output_15_256(.a(output_16_256), .b(output_16_1), .y(output_15_256));
wire output_1_257, output_1_2, output_0_257;
mixer gate_output_0_257(.a(output_1_257), .b(output_1_2), .y(output_0_257));
wire output_2_257, output_2_2, output_1_257;
mixer gate_output_1_257(.a(output_2_257), .b(output_2_2), .y(output_1_257));
wire output_3_257, output_3_2, output_2_257;
mixer gate_output_2_257(.a(output_3_257), .b(output_3_2), .y(output_2_257));
wire output_4_257, output_4_2, output_3_257;
mixer gate_output_3_257(.a(output_4_257), .b(output_4_2), .y(output_3_257));
wire output_5_257, output_5_2, output_4_257;
mixer gate_output_4_257(.a(output_5_257), .b(output_5_2), .y(output_4_257));
wire output_6_257, output_6_2, output_5_257;
mixer gate_output_5_257(.a(output_6_257), .b(output_6_2), .y(output_5_257));
wire output_7_257, output_7_2, output_6_257;
mixer gate_output_6_257(.a(output_7_257), .b(output_7_2), .y(output_6_257));
wire output_8_257, output_8_2, output_7_257;
mixer gate_output_7_257(.a(output_8_257), .b(output_8_2), .y(output_7_257));
wire output_9_257, output_9_2, output_8_257;
mixer gate_output_8_257(.a(output_9_257), .b(output_9_2), .y(output_8_257));
wire output_10_257, output_10_2, output_9_257;
mixer gate_output_9_257(.a(output_10_257), .b(output_10_2), .y(output_9_257));
wire output_11_257, output_11_2, output_10_257;
mixer gate_output_10_257(.a(output_11_257), .b(output_11_2), .y(output_10_257));
wire output_12_257, output_12_2, output_11_257;
mixer gate_output_11_257(.a(output_12_257), .b(output_12_2), .y(output_11_257));
wire output_13_257, output_13_2, output_12_257;
mixer gate_output_12_257(.a(output_13_257), .b(output_13_2), .y(output_12_257));
wire output_14_257, output_14_2, output_13_257;
mixer gate_output_13_257(.a(output_14_257), .b(output_14_2), .y(output_13_257));
wire output_15_257, output_15_2, output_14_257;
mixer gate_output_14_257(.a(output_15_257), .b(output_15_2), .y(output_14_257));
wire output_16_257, output_16_2, output_15_257;
mixer gate_output_15_257(.a(output_16_257), .b(output_16_2), .y(output_15_257));
wire output_1_258, output_1_3, output_0_258;
mixer gate_output_0_258(.a(output_1_258), .b(output_1_3), .y(output_0_258));
wire output_2_258, output_2_3, output_1_258;
mixer gate_output_1_258(.a(output_2_258), .b(output_2_3), .y(output_1_258));
wire output_3_258, output_3_3, output_2_258;
mixer gate_output_2_258(.a(output_3_258), .b(output_3_3), .y(output_2_258));
wire output_4_258, output_4_3, output_3_258;
mixer gate_output_3_258(.a(output_4_258), .b(output_4_3), .y(output_3_258));
wire output_5_258, output_5_3, output_4_258;
mixer gate_output_4_258(.a(output_5_258), .b(output_5_3), .y(output_4_258));
wire output_6_258, output_6_3, output_5_258;
mixer gate_output_5_258(.a(output_6_258), .b(output_6_3), .y(output_5_258));
wire output_7_258, output_7_3, output_6_258;
mixer gate_output_6_258(.a(output_7_258), .b(output_7_3), .y(output_6_258));
wire output_8_258, output_8_3, output_7_258;
mixer gate_output_7_258(.a(output_8_258), .b(output_8_3), .y(output_7_258));
wire output_9_258, output_9_3, output_8_258;
mixer gate_output_8_258(.a(output_9_258), .b(output_9_3), .y(output_8_258));
wire output_10_258, output_10_3, output_9_258;
mixer gate_output_9_258(.a(output_10_258), .b(output_10_3), .y(output_9_258));
wire output_11_258, output_11_3, output_10_258;
mixer gate_output_10_258(.a(output_11_258), .b(output_11_3), .y(output_10_258));
wire output_12_258, output_12_3, output_11_258;
mixer gate_output_11_258(.a(output_12_258), .b(output_12_3), .y(output_11_258));
wire output_13_258, output_13_3, output_12_258;
mixer gate_output_12_258(.a(output_13_258), .b(output_13_3), .y(output_12_258));
wire output_14_258, output_14_3, output_13_258;
mixer gate_output_13_258(.a(output_14_258), .b(output_14_3), .y(output_13_258));
wire output_15_258, output_15_3, output_14_258;
mixer gate_output_14_258(.a(output_15_258), .b(output_15_3), .y(output_14_258));
wire output_16_258, output_16_3, output_15_258;
mixer gate_output_15_258(.a(output_16_258), .b(output_16_3), .y(output_15_258));
wire output_1_259, output_1_4, output_0_259;
mixer gate_output_0_259(.a(output_1_259), .b(output_1_4), .y(output_0_259));
wire output_2_259, output_2_4, output_1_259;
mixer gate_output_1_259(.a(output_2_259), .b(output_2_4), .y(output_1_259));
wire output_3_259, output_3_4, output_2_259;
mixer gate_output_2_259(.a(output_3_259), .b(output_3_4), .y(output_2_259));
wire output_4_259, output_4_4, output_3_259;
mixer gate_output_3_259(.a(output_4_259), .b(output_4_4), .y(output_3_259));
wire output_5_259, output_5_4, output_4_259;
mixer gate_output_4_259(.a(output_5_259), .b(output_5_4), .y(output_4_259));
wire output_6_259, output_6_4, output_5_259;
mixer gate_output_5_259(.a(output_6_259), .b(output_6_4), .y(output_5_259));
wire output_7_259, output_7_4, output_6_259;
mixer gate_output_6_259(.a(output_7_259), .b(output_7_4), .y(output_6_259));
wire output_8_259, output_8_4, output_7_259;
mixer gate_output_7_259(.a(output_8_259), .b(output_8_4), .y(output_7_259));
wire output_9_259, output_9_4, output_8_259;
mixer gate_output_8_259(.a(output_9_259), .b(output_9_4), .y(output_8_259));
wire output_10_259, output_10_4, output_9_259;
mixer gate_output_9_259(.a(output_10_259), .b(output_10_4), .y(output_9_259));
wire output_11_259, output_11_4, output_10_259;
mixer gate_output_10_259(.a(output_11_259), .b(output_11_4), .y(output_10_259));
wire output_12_259, output_12_4, output_11_259;
mixer gate_output_11_259(.a(output_12_259), .b(output_12_4), .y(output_11_259));
wire output_13_259, output_13_4, output_12_259;
mixer gate_output_12_259(.a(output_13_259), .b(output_13_4), .y(output_12_259));
wire output_14_259, output_14_4, output_13_259;
mixer gate_output_13_259(.a(output_14_259), .b(output_14_4), .y(output_13_259));
wire output_15_259, output_15_4, output_14_259;
mixer gate_output_14_259(.a(output_15_259), .b(output_15_4), .y(output_14_259));
wire output_16_259, output_16_4, output_15_259;
mixer gate_output_15_259(.a(output_16_259), .b(output_16_4), .y(output_15_259));
wire output_1_260, output_1_5, output_0_260;
mixer gate_output_0_260(.a(output_1_260), .b(output_1_5), .y(output_0_260));
wire output_2_260, output_2_5, output_1_260;
mixer gate_output_1_260(.a(output_2_260), .b(output_2_5), .y(output_1_260));
wire output_3_260, output_3_5, output_2_260;
mixer gate_output_2_260(.a(output_3_260), .b(output_3_5), .y(output_2_260));
wire output_4_260, output_4_5, output_3_260;
mixer gate_output_3_260(.a(output_4_260), .b(output_4_5), .y(output_3_260));
wire output_5_260, output_5_5, output_4_260;
mixer gate_output_4_260(.a(output_5_260), .b(output_5_5), .y(output_4_260));
wire output_6_260, output_6_5, output_5_260;
mixer gate_output_5_260(.a(output_6_260), .b(output_6_5), .y(output_5_260));
wire output_7_260, output_7_5, output_6_260;
mixer gate_output_6_260(.a(output_7_260), .b(output_7_5), .y(output_6_260));
wire output_8_260, output_8_5, output_7_260;
mixer gate_output_7_260(.a(output_8_260), .b(output_8_5), .y(output_7_260));
wire output_9_260, output_9_5, output_8_260;
mixer gate_output_8_260(.a(output_9_260), .b(output_9_5), .y(output_8_260));
wire output_10_260, output_10_5, output_9_260;
mixer gate_output_9_260(.a(output_10_260), .b(output_10_5), .y(output_9_260));
wire output_11_260, output_11_5, output_10_260;
mixer gate_output_10_260(.a(output_11_260), .b(output_11_5), .y(output_10_260));
wire output_12_260, output_12_5, output_11_260;
mixer gate_output_11_260(.a(output_12_260), .b(output_12_5), .y(output_11_260));
wire output_13_260, output_13_5, output_12_260;
mixer gate_output_12_260(.a(output_13_260), .b(output_13_5), .y(output_12_260));
wire output_14_260, output_14_5, output_13_260;
mixer gate_output_13_260(.a(output_14_260), .b(output_14_5), .y(output_13_260));
wire output_15_260, output_15_5, output_14_260;
mixer gate_output_14_260(.a(output_15_260), .b(output_15_5), .y(output_14_260));
wire output_16_260, output_16_5, output_15_260;
mixer gate_output_15_260(.a(output_16_260), .b(output_16_5), .y(output_15_260));
wire output_1_261, output_1_6, output_0_261;
mixer gate_output_0_261(.a(output_1_261), .b(output_1_6), .y(output_0_261));
wire output_2_261, output_2_6, output_1_261;
mixer gate_output_1_261(.a(output_2_261), .b(output_2_6), .y(output_1_261));
wire output_3_261, output_3_6, output_2_261;
mixer gate_output_2_261(.a(output_3_261), .b(output_3_6), .y(output_2_261));
wire output_4_261, output_4_6, output_3_261;
mixer gate_output_3_261(.a(output_4_261), .b(output_4_6), .y(output_3_261));
wire output_5_261, output_5_6, output_4_261;
mixer gate_output_4_261(.a(output_5_261), .b(output_5_6), .y(output_4_261));
wire output_6_261, output_6_6, output_5_261;
mixer gate_output_5_261(.a(output_6_261), .b(output_6_6), .y(output_5_261));
wire output_7_261, output_7_6, output_6_261;
mixer gate_output_6_261(.a(output_7_261), .b(output_7_6), .y(output_6_261));
wire output_8_261, output_8_6, output_7_261;
mixer gate_output_7_261(.a(output_8_261), .b(output_8_6), .y(output_7_261));
wire output_9_261, output_9_6, output_8_261;
mixer gate_output_8_261(.a(output_9_261), .b(output_9_6), .y(output_8_261));
wire output_10_261, output_10_6, output_9_261;
mixer gate_output_9_261(.a(output_10_261), .b(output_10_6), .y(output_9_261));
wire output_11_261, output_11_6, output_10_261;
mixer gate_output_10_261(.a(output_11_261), .b(output_11_6), .y(output_10_261));
wire output_12_261, output_12_6, output_11_261;
mixer gate_output_11_261(.a(output_12_261), .b(output_12_6), .y(output_11_261));
wire output_13_261, output_13_6, output_12_261;
mixer gate_output_12_261(.a(output_13_261), .b(output_13_6), .y(output_12_261));
wire output_14_261, output_14_6, output_13_261;
mixer gate_output_13_261(.a(output_14_261), .b(output_14_6), .y(output_13_261));
wire output_15_261, output_15_6, output_14_261;
mixer gate_output_14_261(.a(output_15_261), .b(output_15_6), .y(output_14_261));
wire output_16_261, output_16_6, output_15_261;
mixer gate_output_15_261(.a(output_16_261), .b(output_16_6), .y(output_15_261));
wire output_1_262, output_1_7, output_0_262;
mixer gate_output_0_262(.a(output_1_262), .b(output_1_7), .y(output_0_262));
wire output_2_262, output_2_7, output_1_262;
mixer gate_output_1_262(.a(output_2_262), .b(output_2_7), .y(output_1_262));
wire output_3_262, output_3_7, output_2_262;
mixer gate_output_2_262(.a(output_3_262), .b(output_3_7), .y(output_2_262));
wire output_4_262, output_4_7, output_3_262;
mixer gate_output_3_262(.a(output_4_262), .b(output_4_7), .y(output_3_262));
wire output_5_262, output_5_7, output_4_262;
mixer gate_output_4_262(.a(output_5_262), .b(output_5_7), .y(output_4_262));
wire output_6_262, output_6_7, output_5_262;
mixer gate_output_5_262(.a(output_6_262), .b(output_6_7), .y(output_5_262));
wire output_7_262, output_7_7, output_6_262;
mixer gate_output_6_262(.a(output_7_262), .b(output_7_7), .y(output_6_262));
wire output_8_262, output_8_7, output_7_262;
mixer gate_output_7_262(.a(output_8_262), .b(output_8_7), .y(output_7_262));
wire output_9_262, output_9_7, output_8_262;
mixer gate_output_8_262(.a(output_9_262), .b(output_9_7), .y(output_8_262));
wire output_10_262, output_10_7, output_9_262;
mixer gate_output_9_262(.a(output_10_262), .b(output_10_7), .y(output_9_262));
wire output_11_262, output_11_7, output_10_262;
mixer gate_output_10_262(.a(output_11_262), .b(output_11_7), .y(output_10_262));
wire output_12_262, output_12_7, output_11_262;
mixer gate_output_11_262(.a(output_12_262), .b(output_12_7), .y(output_11_262));
wire output_13_262, output_13_7, output_12_262;
mixer gate_output_12_262(.a(output_13_262), .b(output_13_7), .y(output_12_262));
wire output_14_262, output_14_7, output_13_262;
mixer gate_output_13_262(.a(output_14_262), .b(output_14_7), .y(output_13_262));
wire output_15_262, output_15_7, output_14_262;
mixer gate_output_14_262(.a(output_15_262), .b(output_15_7), .y(output_14_262));
wire output_16_262, output_16_7, output_15_262;
mixer gate_output_15_262(.a(output_16_262), .b(output_16_7), .y(output_15_262));
wire output_1_263, output_1_8, output_0_263;
mixer gate_output_0_263(.a(output_1_263), .b(output_1_8), .y(output_0_263));
wire output_2_263, output_2_8, output_1_263;
mixer gate_output_1_263(.a(output_2_263), .b(output_2_8), .y(output_1_263));
wire output_3_263, output_3_8, output_2_263;
mixer gate_output_2_263(.a(output_3_263), .b(output_3_8), .y(output_2_263));
wire output_4_263, output_4_8, output_3_263;
mixer gate_output_3_263(.a(output_4_263), .b(output_4_8), .y(output_3_263));
wire output_5_263, output_5_8, output_4_263;
mixer gate_output_4_263(.a(output_5_263), .b(output_5_8), .y(output_4_263));
wire output_6_263, output_6_8, output_5_263;
mixer gate_output_5_263(.a(output_6_263), .b(output_6_8), .y(output_5_263));
wire output_7_263, output_7_8, output_6_263;
mixer gate_output_6_263(.a(output_7_263), .b(output_7_8), .y(output_6_263));
wire output_8_263, output_8_8, output_7_263;
mixer gate_output_7_263(.a(output_8_263), .b(output_8_8), .y(output_7_263));
wire output_9_263, output_9_8, output_8_263;
mixer gate_output_8_263(.a(output_9_263), .b(output_9_8), .y(output_8_263));
wire output_10_263, output_10_8, output_9_263;
mixer gate_output_9_263(.a(output_10_263), .b(output_10_8), .y(output_9_263));
wire output_11_263, output_11_8, output_10_263;
mixer gate_output_10_263(.a(output_11_263), .b(output_11_8), .y(output_10_263));
wire output_12_263, output_12_8, output_11_263;
mixer gate_output_11_263(.a(output_12_263), .b(output_12_8), .y(output_11_263));
wire output_13_263, output_13_8, output_12_263;
mixer gate_output_12_263(.a(output_13_263), .b(output_13_8), .y(output_12_263));
wire output_14_263, output_14_8, output_13_263;
mixer gate_output_13_263(.a(output_14_263), .b(output_14_8), .y(output_13_263));
wire output_15_263, output_15_8, output_14_263;
mixer gate_output_14_263(.a(output_15_263), .b(output_15_8), .y(output_14_263));
wire output_16_263, output_16_8, output_15_263;
mixer gate_output_15_263(.a(output_16_263), .b(output_16_8), .y(output_15_263));
wire output_1_264, output_1_9, output_0_264;
mixer gate_output_0_264(.a(output_1_264), .b(output_1_9), .y(output_0_264));
wire output_2_264, output_2_9, output_1_264;
mixer gate_output_1_264(.a(output_2_264), .b(output_2_9), .y(output_1_264));
wire output_3_264, output_3_9, output_2_264;
mixer gate_output_2_264(.a(output_3_264), .b(output_3_9), .y(output_2_264));
wire output_4_264, output_4_9, output_3_264;
mixer gate_output_3_264(.a(output_4_264), .b(output_4_9), .y(output_3_264));
wire output_5_264, output_5_9, output_4_264;
mixer gate_output_4_264(.a(output_5_264), .b(output_5_9), .y(output_4_264));
wire output_6_264, output_6_9, output_5_264;
mixer gate_output_5_264(.a(output_6_264), .b(output_6_9), .y(output_5_264));
wire output_7_264, output_7_9, output_6_264;
mixer gate_output_6_264(.a(output_7_264), .b(output_7_9), .y(output_6_264));
wire output_8_264, output_8_9, output_7_264;
mixer gate_output_7_264(.a(output_8_264), .b(output_8_9), .y(output_7_264));
wire output_9_264, output_9_9, output_8_264;
mixer gate_output_8_264(.a(output_9_264), .b(output_9_9), .y(output_8_264));
wire output_10_264, output_10_9, output_9_264;
mixer gate_output_9_264(.a(output_10_264), .b(output_10_9), .y(output_9_264));
wire output_11_264, output_11_9, output_10_264;
mixer gate_output_10_264(.a(output_11_264), .b(output_11_9), .y(output_10_264));
wire output_12_264, output_12_9, output_11_264;
mixer gate_output_11_264(.a(output_12_264), .b(output_12_9), .y(output_11_264));
wire output_13_264, output_13_9, output_12_264;
mixer gate_output_12_264(.a(output_13_264), .b(output_13_9), .y(output_12_264));
wire output_14_264, output_14_9, output_13_264;
mixer gate_output_13_264(.a(output_14_264), .b(output_14_9), .y(output_13_264));
wire output_15_264, output_15_9, output_14_264;
mixer gate_output_14_264(.a(output_15_264), .b(output_15_9), .y(output_14_264));
wire output_16_264, output_16_9, output_15_264;
mixer gate_output_15_264(.a(output_16_264), .b(output_16_9), .y(output_15_264));
wire output_1_265, output_1_10, output_0_265;
mixer gate_output_0_265(.a(output_1_265), .b(output_1_10), .y(output_0_265));
wire output_2_265, output_2_10, output_1_265;
mixer gate_output_1_265(.a(output_2_265), .b(output_2_10), .y(output_1_265));
wire output_3_265, output_3_10, output_2_265;
mixer gate_output_2_265(.a(output_3_265), .b(output_3_10), .y(output_2_265));
wire output_4_265, output_4_10, output_3_265;
mixer gate_output_3_265(.a(output_4_265), .b(output_4_10), .y(output_3_265));
wire output_5_265, output_5_10, output_4_265;
mixer gate_output_4_265(.a(output_5_265), .b(output_5_10), .y(output_4_265));
wire output_6_265, output_6_10, output_5_265;
mixer gate_output_5_265(.a(output_6_265), .b(output_6_10), .y(output_5_265));
wire output_7_265, output_7_10, output_6_265;
mixer gate_output_6_265(.a(output_7_265), .b(output_7_10), .y(output_6_265));
wire output_8_265, output_8_10, output_7_265;
mixer gate_output_7_265(.a(output_8_265), .b(output_8_10), .y(output_7_265));
wire output_9_265, output_9_10, output_8_265;
mixer gate_output_8_265(.a(output_9_265), .b(output_9_10), .y(output_8_265));
wire output_10_265, output_10_10, output_9_265;
mixer gate_output_9_265(.a(output_10_265), .b(output_10_10), .y(output_9_265));
wire output_11_265, output_11_10, output_10_265;
mixer gate_output_10_265(.a(output_11_265), .b(output_11_10), .y(output_10_265));
wire output_12_265, output_12_10, output_11_265;
mixer gate_output_11_265(.a(output_12_265), .b(output_12_10), .y(output_11_265));
wire output_13_265, output_13_10, output_12_265;
mixer gate_output_12_265(.a(output_13_265), .b(output_13_10), .y(output_12_265));
wire output_14_265, output_14_10, output_13_265;
mixer gate_output_13_265(.a(output_14_265), .b(output_14_10), .y(output_13_265));
wire output_15_265, output_15_10, output_14_265;
mixer gate_output_14_265(.a(output_15_265), .b(output_15_10), .y(output_14_265));
wire output_16_265, output_16_10, output_15_265;
mixer gate_output_15_265(.a(output_16_265), .b(output_16_10), .y(output_15_265));
wire output_1_266, output_1_11, output_0_266;
mixer gate_output_0_266(.a(output_1_266), .b(output_1_11), .y(output_0_266));
wire output_2_266, output_2_11, output_1_266;
mixer gate_output_1_266(.a(output_2_266), .b(output_2_11), .y(output_1_266));
wire output_3_266, output_3_11, output_2_266;
mixer gate_output_2_266(.a(output_3_266), .b(output_3_11), .y(output_2_266));
wire output_4_266, output_4_11, output_3_266;
mixer gate_output_3_266(.a(output_4_266), .b(output_4_11), .y(output_3_266));
wire output_5_266, output_5_11, output_4_266;
mixer gate_output_4_266(.a(output_5_266), .b(output_5_11), .y(output_4_266));
wire output_6_266, output_6_11, output_5_266;
mixer gate_output_5_266(.a(output_6_266), .b(output_6_11), .y(output_5_266));
wire output_7_266, output_7_11, output_6_266;
mixer gate_output_6_266(.a(output_7_266), .b(output_7_11), .y(output_6_266));
wire output_8_266, output_8_11, output_7_266;
mixer gate_output_7_266(.a(output_8_266), .b(output_8_11), .y(output_7_266));
wire output_9_266, output_9_11, output_8_266;
mixer gate_output_8_266(.a(output_9_266), .b(output_9_11), .y(output_8_266));
wire output_10_266, output_10_11, output_9_266;
mixer gate_output_9_266(.a(output_10_266), .b(output_10_11), .y(output_9_266));
wire output_11_266, output_11_11, output_10_266;
mixer gate_output_10_266(.a(output_11_266), .b(output_11_11), .y(output_10_266));
wire output_12_266, output_12_11, output_11_266;
mixer gate_output_11_266(.a(output_12_266), .b(output_12_11), .y(output_11_266));
wire output_13_266, output_13_11, output_12_266;
mixer gate_output_12_266(.a(output_13_266), .b(output_13_11), .y(output_12_266));
wire output_14_266, output_14_11, output_13_266;
mixer gate_output_13_266(.a(output_14_266), .b(output_14_11), .y(output_13_266));
wire output_15_266, output_15_11, output_14_266;
mixer gate_output_14_266(.a(output_15_266), .b(output_15_11), .y(output_14_266));
wire output_16_266, output_16_11, output_15_266;
mixer gate_output_15_266(.a(output_16_266), .b(output_16_11), .y(output_15_266));
wire output_1_267, output_1_12, output_0_267;
mixer gate_output_0_267(.a(output_1_267), .b(output_1_12), .y(output_0_267));
wire output_2_267, output_2_12, output_1_267;
mixer gate_output_1_267(.a(output_2_267), .b(output_2_12), .y(output_1_267));
wire output_3_267, output_3_12, output_2_267;
mixer gate_output_2_267(.a(output_3_267), .b(output_3_12), .y(output_2_267));
wire output_4_267, output_4_12, output_3_267;
mixer gate_output_3_267(.a(output_4_267), .b(output_4_12), .y(output_3_267));
wire output_5_267, output_5_12, output_4_267;
mixer gate_output_4_267(.a(output_5_267), .b(output_5_12), .y(output_4_267));
wire output_6_267, output_6_12, output_5_267;
mixer gate_output_5_267(.a(output_6_267), .b(output_6_12), .y(output_5_267));
wire output_7_267, output_7_12, output_6_267;
mixer gate_output_6_267(.a(output_7_267), .b(output_7_12), .y(output_6_267));
wire output_8_267, output_8_12, output_7_267;
mixer gate_output_7_267(.a(output_8_267), .b(output_8_12), .y(output_7_267));
wire output_9_267, output_9_12, output_8_267;
mixer gate_output_8_267(.a(output_9_267), .b(output_9_12), .y(output_8_267));
wire output_10_267, output_10_12, output_9_267;
mixer gate_output_9_267(.a(output_10_267), .b(output_10_12), .y(output_9_267));
wire output_11_267, output_11_12, output_10_267;
mixer gate_output_10_267(.a(output_11_267), .b(output_11_12), .y(output_10_267));
wire output_12_267, output_12_12, output_11_267;
mixer gate_output_11_267(.a(output_12_267), .b(output_12_12), .y(output_11_267));
wire output_13_267, output_13_12, output_12_267;
mixer gate_output_12_267(.a(output_13_267), .b(output_13_12), .y(output_12_267));
wire output_14_267, output_14_12, output_13_267;
mixer gate_output_13_267(.a(output_14_267), .b(output_14_12), .y(output_13_267));
wire output_15_267, output_15_12, output_14_267;
mixer gate_output_14_267(.a(output_15_267), .b(output_15_12), .y(output_14_267));
wire output_16_267, output_16_12, output_15_267;
mixer gate_output_15_267(.a(output_16_267), .b(output_16_12), .y(output_15_267));
wire output_1_268, output_1_13, output_0_268;
mixer gate_output_0_268(.a(output_1_268), .b(output_1_13), .y(output_0_268));
wire output_2_268, output_2_13, output_1_268;
mixer gate_output_1_268(.a(output_2_268), .b(output_2_13), .y(output_1_268));
wire output_3_268, output_3_13, output_2_268;
mixer gate_output_2_268(.a(output_3_268), .b(output_3_13), .y(output_2_268));
wire output_4_268, output_4_13, output_3_268;
mixer gate_output_3_268(.a(output_4_268), .b(output_4_13), .y(output_3_268));
wire output_5_268, output_5_13, output_4_268;
mixer gate_output_4_268(.a(output_5_268), .b(output_5_13), .y(output_4_268));
wire output_6_268, output_6_13, output_5_268;
mixer gate_output_5_268(.a(output_6_268), .b(output_6_13), .y(output_5_268));
wire output_7_268, output_7_13, output_6_268;
mixer gate_output_6_268(.a(output_7_268), .b(output_7_13), .y(output_6_268));
wire output_8_268, output_8_13, output_7_268;
mixer gate_output_7_268(.a(output_8_268), .b(output_8_13), .y(output_7_268));
wire output_9_268, output_9_13, output_8_268;
mixer gate_output_8_268(.a(output_9_268), .b(output_9_13), .y(output_8_268));
wire output_10_268, output_10_13, output_9_268;
mixer gate_output_9_268(.a(output_10_268), .b(output_10_13), .y(output_9_268));
wire output_11_268, output_11_13, output_10_268;
mixer gate_output_10_268(.a(output_11_268), .b(output_11_13), .y(output_10_268));
wire output_12_268, output_12_13, output_11_268;
mixer gate_output_11_268(.a(output_12_268), .b(output_12_13), .y(output_11_268));
wire output_13_268, output_13_13, output_12_268;
mixer gate_output_12_268(.a(output_13_268), .b(output_13_13), .y(output_12_268));
wire output_14_268, output_14_13, output_13_268;
mixer gate_output_13_268(.a(output_14_268), .b(output_14_13), .y(output_13_268));
wire output_15_268, output_15_13, output_14_268;
mixer gate_output_14_268(.a(output_15_268), .b(output_15_13), .y(output_14_268));
wire output_16_268, output_16_13, output_15_268;
mixer gate_output_15_268(.a(output_16_268), .b(output_16_13), .y(output_15_268));
wire output_1_269, output_1_14, output_0_269;
mixer gate_output_0_269(.a(output_1_269), .b(output_1_14), .y(output_0_269));
wire output_2_269, output_2_14, output_1_269;
mixer gate_output_1_269(.a(output_2_269), .b(output_2_14), .y(output_1_269));
wire output_3_269, output_3_14, output_2_269;
mixer gate_output_2_269(.a(output_3_269), .b(output_3_14), .y(output_2_269));
wire output_4_269, output_4_14, output_3_269;
mixer gate_output_3_269(.a(output_4_269), .b(output_4_14), .y(output_3_269));
wire output_5_269, output_5_14, output_4_269;
mixer gate_output_4_269(.a(output_5_269), .b(output_5_14), .y(output_4_269));
wire output_6_269, output_6_14, output_5_269;
mixer gate_output_5_269(.a(output_6_269), .b(output_6_14), .y(output_5_269));
wire output_7_269, output_7_14, output_6_269;
mixer gate_output_6_269(.a(output_7_269), .b(output_7_14), .y(output_6_269));
wire output_8_269, output_8_14, output_7_269;
mixer gate_output_7_269(.a(output_8_269), .b(output_8_14), .y(output_7_269));
wire output_9_269, output_9_14, output_8_269;
mixer gate_output_8_269(.a(output_9_269), .b(output_9_14), .y(output_8_269));
wire output_10_269, output_10_14, output_9_269;
mixer gate_output_9_269(.a(output_10_269), .b(output_10_14), .y(output_9_269));
wire output_11_269, output_11_14, output_10_269;
mixer gate_output_10_269(.a(output_11_269), .b(output_11_14), .y(output_10_269));
wire output_12_269, output_12_14, output_11_269;
mixer gate_output_11_269(.a(output_12_269), .b(output_12_14), .y(output_11_269));
wire output_13_269, output_13_14, output_12_269;
mixer gate_output_12_269(.a(output_13_269), .b(output_13_14), .y(output_12_269));
wire output_14_269, output_14_14, output_13_269;
mixer gate_output_13_269(.a(output_14_269), .b(output_14_14), .y(output_13_269));
wire output_15_269, output_15_14, output_14_269;
mixer gate_output_14_269(.a(output_15_269), .b(output_15_14), .y(output_14_269));
wire output_16_269, output_16_14, output_15_269;
mixer gate_output_15_269(.a(output_16_269), .b(output_16_14), .y(output_15_269));
wire output_1_270, output_1_15, output_0_270;
mixer gate_output_0_270(.a(output_1_270), .b(output_1_15), .y(output_0_270));
wire output_2_270, output_2_15, output_1_270;
mixer gate_output_1_270(.a(output_2_270), .b(output_2_15), .y(output_1_270));
wire output_3_270, output_3_15, output_2_270;
mixer gate_output_2_270(.a(output_3_270), .b(output_3_15), .y(output_2_270));
wire output_4_270, output_4_15, output_3_270;
mixer gate_output_3_270(.a(output_4_270), .b(output_4_15), .y(output_3_270));
wire output_5_270, output_5_15, output_4_270;
mixer gate_output_4_270(.a(output_5_270), .b(output_5_15), .y(output_4_270));
wire output_6_270, output_6_15, output_5_270;
mixer gate_output_5_270(.a(output_6_270), .b(output_6_15), .y(output_5_270));
wire output_7_270, output_7_15, output_6_270;
mixer gate_output_6_270(.a(output_7_270), .b(output_7_15), .y(output_6_270));
wire output_8_270, output_8_15, output_7_270;
mixer gate_output_7_270(.a(output_8_270), .b(output_8_15), .y(output_7_270));
wire output_9_270, output_9_15, output_8_270;
mixer gate_output_8_270(.a(output_9_270), .b(output_9_15), .y(output_8_270));
wire output_10_270, output_10_15, output_9_270;
mixer gate_output_9_270(.a(output_10_270), .b(output_10_15), .y(output_9_270));
wire output_11_270, output_11_15, output_10_270;
mixer gate_output_10_270(.a(output_11_270), .b(output_11_15), .y(output_10_270));
wire output_12_270, output_12_15, output_11_270;
mixer gate_output_11_270(.a(output_12_270), .b(output_12_15), .y(output_11_270));
wire output_13_270, output_13_15, output_12_270;
mixer gate_output_12_270(.a(output_13_270), .b(output_13_15), .y(output_12_270));
wire output_14_270, output_14_15, output_13_270;
mixer gate_output_13_270(.a(output_14_270), .b(output_14_15), .y(output_13_270));
wire output_15_270, output_15_15, output_14_270;
mixer gate_output_14_270(.a(output_15_270), .b(output_15_15), .y(output_14_270));
wire output_16_270, output_16_15, output_15_270;
mixer gate_output_15_270(.a(output_16_270), .b(output_16_15), .y(output_15_270));
wire output_1_271, output_1_0, output_0_271;
mixer gate_output_0_271(.a(output_1_271), .b(output_1_0), .y(output_0_271));
wire output_2_271, output_2_0, output_1_271;
mixer gate_output_1_271(.a(output_2_271), .b(output_2_0), .y(output_1_271));
wire output_3_271, output_3_0, output_2_271;
mixer gate_output_2_271(.a(output_3_271), .b(output_3_0), .y(output_2_271));
wire output_4_271, output_4_0, output_3_271;
mixer gate_output_3_271(.a(output_4_271), .b(output_4_0), .y(output_3_271));
wire output_5_271, output_5_0, output_4_271;
mixer gate_output_4_271(.a(output_5_271), .b(output_5_0), .y(output_4_271));
wire output_6_271, output_6_0, output_5_271;
mixer gate_output_5_271(.a(output_6_271), .b(output_6_0), .y(output_5_271));
wire output_7_271, output_7_0, output_6_271;
mixer gate_output_6_271(.a(output_7_271), .b(output_7_0), .y(output_6_271));
wire output_8_271, output_8_0, output_7_271;
mixer gate_output_7_271(.a(output_8_271), .b(output_8_0), .y(output_7_271));
wire output_9_271, output_9_0, output_8_271;
mixer gate_output_8_271(.a(output_9_271), .b(output_9_0), .y(output_8_271));
wire output_10_271, output_10_0, output_9_271;
mixer gate_output_9_271(.a(output_10_271), .b(output_10_0), .y(output_9_271));
wire output_11_271, output_11_0, output_10_271;
mixer gate_output_10_271(.a(output_11_271), .b(output_11_0), .y(output_10_271));
wire output_12_271, output_12_0, output_11_271;
mixer gate_output_11_271(.a(output_12_271), .b(output_12_0), .y(output_11_271));
wire output_13_271, output_13_0, output_12_271;
mixer gate_output_12_271(.a(output_13_271), .b(output_13_0), .y(output_12_271));
wire output_14_271, output_14_0, output_13_271;
mixer gate_output_13_271(.a(output_14_271), .b(output_14_0), .y(output_13_271));
wire output_15_271, output_15_0, output_14_271;
mixer gate_output_14_271(.a(output_15_271), .b(output_15_0), .y(output_14_271));
wire output_16_271, output_16_0, output_15_271;
mixer gate_output_15_271(.a(output_16_271), .b(output_16_0), .y(output_15_271));
wire output_1_272, output_1_1, output_0_272;
mixer gate_output_0_272(.a(output_1_272), .b(output_1_1), .y(output_0_272));
wire output_2_272, output_2_1, output_1_272;
mixer gate_output_1_272(.a(output_2_272), .b(output_2_1), .y(output_1_272));
wire output_3_272, output_3_1, output_2_272;
mixer gate_output_2_272(.a(output_3_272), .b(output_3_1), .y(output_2_272));
wire output_4_272, output_4_1, output_3_272;
mixer gate_output_3_272(.a(output_4_272), .b(output_4_1), .y(output_3_272));
wire output_5_272, output_5_1, output_4_272;
mixer gate_output_4_272(.a(output_5_272), .b(output_5_1), .y(output_4_272));
wire output_6_272, output_6_1, output_5_272;
mixer gate_output_5_272(.a(output_6_272), .b(output_6_1), .y(output_5_272));
wire output_7_272, output_7_1, output_6_272;
mixer gate_output_6_272(.a(output_7_272), .b(output_7_1), .y(output_6_272));
wire output_8_272, output_8_1, output_7_272;
mixer gate_output_7_272(.a(output_8_272), .b(output_8_1), .y(output_7_272));
wire output_9_272, output_9_1, output_8_272;
mixer gate_output_8_272(.a(output_9_272), .b(output_9_1), .y(output_8_272));
wire output_10_272, output_10_1, output_9_272;
mixer gate_output_9_272(.a(output_10_272), .b(output_10_1), .y(output_9_272));
wire output_11_272, output_11_1, output_10_272;
mixer gate_output_10_272(.a(output_11_272), .b(output_11_1), .y(output_10_272));
wire output_12_272, output_12_1, output_11_272;
mixer gate_output_11_272(.a(output_12_272), .b(output_12_1), .y(output_11_272));
wire output_13_272, output_13_1, output_12_272;
mixer gate_output_12_272(.a(output_13_272), .b(output_13_1), .y(output_12_272));
wire output_14_272, output_14_1, output_13_272;
mixer gate_output_13_272(.a(output_14_272), .b(output_14_1), .y(output_13_272));
wire output_15_272, output_15_1, output_14_272;
mixer gate_output_14_272(.a(output_15_272), .b(output_15_1), .y(output_14_272));
wire output_16_272, output_16_1, output_15_272;
mixer gate_output_15_272(.a(output_16_272), .b(output_16_1), .y(output_15_272));
wire output_1_273, output_1_2, output_0_273;
mixer gate_output_0_273(.a(output_1_273), .b(output_1_2), .y(output_0_273));
wire output_2_273, output_2_2, output_1_273;
mixer gate_output_1_273(.a(output_2_273), .b(output_2_2), .y(output_1_273));
wire output_3_273, output_3_2, output_2_273;
mixer gate_output_2_273(.a(output_3_273), .b(output_3_2), .y(output_2_273));
wire output_4_273, output_4_2, output_3_273;
mixer gate_output_3_273(.a(output_4_273), .b(output_4_2), .y(output_3_273));
wire output_5_273, output_5_2, output_4_273;
mixer gate_output_4_273(.a(output_5_273), .b(output_5_2), .y(output_4_273));
wire output_6_273, output_6_2, output_5_273;
mixer gate_output_5_273(.a(output_6_273), .b(output_6_2), .y(output_5_273));
wire output_7_273, output_7_2, output_6_273;
mixer gate_output_6_273(.a(output_7_273), .b(output_7_2), .y(output_6_273));
wire output_8_273, output_8_2, output_7_273;
mixer gate_output_7_273(.a(output_8_273), .b(output_8_2), .y(output_7_273));
wire output_9_273, output_9_2, output_8_273;
mixer gate_output_8_273(.a(output_9_273), .b(output_9_2), .y(output_8_273));
wire output_10_273, output_10_2, output_9_273;
mixer gate_output_9_273(.a(output_10_273), .b(output_10_2), .y(output_9_273));
wire output_11_273, output_11_2, output_10_273;
mixer gate_output_10_273(.a(output_11_273), .b(output_11_2), .y(output_10_273));
wire output_12_273, output_12_2, output_11_273;
mixer gate_output_11_273(.a(output_12_273), .b(output_12_2), .y(output_11_273));
wire output_13_273, output_13_2, output_12_273;
mixer gate_output_12_273(.a(output_13_273), .b(output_13_2), .y(output_12_273));
wire output_14_273, output_14_2, output_13_273;
mixer gate_output_13_273(.a(output_14_273), .b(output_14_2), .y(output_13_273));
wire output_15_273, output_15_2, output_14_273;
mixer gate_output_14_273(.a(output_15_273), .b(output_15_2), .y(output_14_273));
wire output_16_273, output_16_2, output_15_273;
mixer gate_output_15_273(.a(output_16_273), .b(output_16_2), .y(output_15_273));
wire output_1_274, output_1_3, output_0_274;
mixer gate_output_0_274(.a(output_1_274), .b(output_1_3), .y(output_0_274));
wire output_2_274, output_2_3, output_1_274;
mixer gate_output_1_274(.a(output_2_274), .b(output_2_3), .y(output_1_274));
wire output_3_274, output_3_3, output_2_274;
mixer gate_output_2_274(.a(output_3_274), .b(output_3_3), .y(output_2_274));
wire output_4_274, output_4_3, output_3_274;
mixer gate_output_3_274(.a(output_4_274), .b(output_4_3), .y(output_3_274));
wire output_5_274, output_5_3, output_4_274;
mixer gate_output_4_274(.a(output_5_274), .b(output_5_3), .y(output_4_274));
wire output_6_274, output_6_3, output_5_274;
mixer gate_output_5_274(.a(output_6_274), .b(output_6_3), .y(output_5_274));
wire output_7_274, output_7_3, output_6_274;
mixer gate_output_6_274(.a(output_7_274), .b(output_7_3), .y(output_6_274));
wire output_8_274, output_8_3, output_7_274;
mixer gate_output_7_274(.a(output_8_274), .b(output_8_3), .y(output_7_274));
wire output_9_274, output_9_3, output_8_274;
mixer gate_output_8_274(.a(output_9_274), .b(output_9_3), .y(output_8_274));
wire output_10_274, output_10_3, output_9_274;
mixer gate_output_9_274(.a(output_10_274), .b(output_10_3), .y(output_9_274));
wire output_11_274, output_11_3, output_10_274;
mixer gate_output_10_274(.a(output_11_274), .b(output_11_3), .y(output_10_274));
wire output_12_274, output_12_3, output_11_274;
mixer gate_output_11_274(.a(output_12_274), .b(output_12_3), .y(output_11_274));
wire output_13_274, output_13_3, output_12_274;
mixer gate_output_12_274(.a(output_13_274), .b(output_13_3), .y(output_12_274));
wire output_14_274, output_14_3, output_13_274;
mixer gate_output_13_274(.a(output_14_274), .b(output_14_3), .y(output_13_274));
wire output_15_274, output_15_3, output_14_274;
mixer gate_output_14_274(.a(output_15_274), .b(output_15_3), .y(output_14_274));
wire output_16_274, output_16_3, output_15_274;
mixer gate_output_15_274(.a(output_16_274), .b(output_16_3), .y(output_15_274));
wire output_1_275, output_1_4, output_0_275;
mixer gate_output_0_275(.a(output_1_275), .b(output_1_4), .y(output_0_275));
wire output_2_275, output_2_4, output_1_275;
mixer gate_output_1_275(.a(output_2_275), .b(output_2_4), .y(output_1_275));
wire output_3_275, output_3_4, output_2_275;
mixer gate_output_2_275(.a(output_3_275), .b(output_3_4), .y(output_2_275));
wire output_4_275, output_4_4, output_3_275;
mixer gate_output_3_275(.a(output_4_275), .b(output_4_4), .y(output_3_275));
wire output_5_275, output_5_4, output_4_275;
mixer gate_output_4_275(.a(output_5_275), .b(output_5_4), .y(output_4_275));
wire output_6_275, output_6_4, output_5_275;
mixer gate_output_5_275(.a(output_6_275), .b(output_6_4), .y(output_5_275));
wire output_7_275, output_7_4, output_6_275;
mixer gate_output_6_275(.a(output_7_275), .b(output_7_4), .y(output_6_275));
wire output_8_275, output_8_4, output_7_275;
mixer gate_output_7_275(.a(output_8_275), .b(output_8_4), .y(output_7_275));
wire output_9_275, output_9_4, output_8_275;
mixer gate_output_8_275(.a(output_9_275), .b(output_9_4), .y(output_8_275));
wire output_10_275, output_10_4, output_9_275;
mixer gate_output_9_275(.a(output_10_275), .b(output_10_4), .y(output_9_275));
wire output_11_275, output_11_4, output_10_275;
mixer gate_output_10_275(.a(output_11_275), .b(output_11_4), .y(output_10_275));
wire output_12_275, output_12_4, output_11_275;
mixer gate_output_11_275(.a(output_12_275), .b(output_12_4), .y(output_11_275));
wire output_13_275, output_13_4, output_12_275;
mixer gate_output_12_275(.a(output_13_275), .b(output_13_4), .y(output_12_275));
wire output_14_275, output_14_4, output_13_275;
mixer gate_output_13_275(.a(output_14_275), .b(output_14_4), .y(output_13_275));
wire output_15_275, output_15_4, output_14_275;
mixer gate_output_14_275(.a(output_15_275), .b(output_15_4), .y(output_14_275));
wire output_16_275, output_16_4, output_15_275;
mixer gate_output_15_275(.a(output_16_275), .b(output_16_4), .y(output_15_275));
wire output_1_276, output_1_5, output_0_276;
mixer gate_output_0_276(.a(output_1_276), .b(output_1_5), .y(output_0_276));
wire output_2_276, output_2_5, output_1_276;
mixer gate_output_1_276(.a(output_2_276), .b(output_2_5), .y(output_1_276));
wire output_3_276, output_3_5, output_2_276;
mixer gate_output_2_276(.a(output_3_276), .b(output_3_5), .y(output_2_276));
wire output_4_276, output_4_5, output_3_276;
mixer gate_output_3_276(.a(output_4_276), .b(output_4_5), .y(output_3_276));
wire output_5_276, output_5_5, output_4_276;
mixer gate_output_4_276(.a(output_5_276), .b(output_5_5), .y(output_4_276));
wire output_6_276, output_6_5, output_5_276;
mixer gate_output_5_276(.a(output_6_276), .b(output_6_5), .y(output_5_276));
wire output_7_276, output_7_5, output_6_276;
mixer gate_output_6_276(.a(output_7_276), .b(output_7_5), .y(output_6_276));
wire output_8_276, output_8_5, output_7_276;
mixer gate_output_7_276(.a(output_8_276), .b(output_8_5), .y(output_7_276));
wire output_9_276, output_9_5, output_8_276;
mixer gate_output_8_276(.a(output_9_276), .b(output_9_5), .y(output_8_276));
wire output_10_276, output_10_5, output_9_276;
mixer gate_output_9_276(.a(output_10_276), .b(output_10_5), .y(output_9_276));
wire output_11_276, output_11_5, output_10_276;
mixer gate_output_10_276(.a(output_11_276), .b(output_11_5), .y(output_10_276));
wire output_12_276, output_12_5, output_11_276;
mixer gate_output_11_276(.a(output_12_276), .b(output_12_5), .y(output_11_276));
wire output_13_276, output_13_5, output_12_276;
mixer gate_output_12_276(.a(output_13_276), .b(output_13_5), .y(output_12_276));
wire output_14_276, output_14_5, output_13_276;
mixer gate_output_13_276(.a(output_14_276), .b(output_14_5), .y(output_13_276));
wire output_15_276, output_15_5, output_14_276;
mixer gate_output_14_276(.a(output_15_276), .b(output_15_5), .y(output_14_276));
wire output_16_276, output_16_5, output_15_276;
mixer gate_output_15_276(.a(output_16_276), .b(output_16_5), .y(output_15_276));
wire output_1_277, output_1_6, output_0_277;
mixer gate_output_0_277(.a(output_1_277), .b(output_1_6), .y(output_0_277));
wire output_2_277, output_2_6, output_1_277;
mixer gate_output_1_277(.a(output_2_277), .b(output_2_6), .y(output_1_277));
wire output_3_277, output_3_6, output_2_277;
mixer gate_output_2_277(.a(output_3_277), .b(output_3_6), .y(output_2_277));
wire output_4_277, output_4_6, output_3_277;
mixer gate_output_3_277(.a(output_4_277), .b(output_4_6), .y(output_3_277));
wire output_5_277, output_5_6, output_4_277;
mixer gate_output_4_277(.a(output_5_277), .b(output_5_6), .y(output_4_277));
wire output_6_277, output_6_6, output_5_277;
mixer gate_output_5_277(.a(output_6_277), .b(output_6_6), .y(output_5_277));
wire output_7_277, output_7_6, output_6_277;
mixer gate_output_6_277(.a(output_7_277), .b(output_7_6), .y(output_6_277));
wire output_8_277, output_8_6, output_7_277;
mixer gate_output_7_277(.a(output_8_277), .b(output_8_6), .y(output_7_277));
wire output_9_277, output_9_6, output_8_277;
mixer gate_output_8_277(.a(output_9_277), .b(output_9_6), .y(output_8_277));
wire output_10_277, output_10_6, output_9_277;
mixer gate_output_9_277(.a(output_10_277), .b(output_10_6), .y(output_9_277));
wire output_11_277, output_11_6, output_10_277;
mixer gate_output_10_277(.a(output_11_277), .b(output_11_6), .y(output_10_277));
wire output_12_277, output_12_6, output_11_277;
mixer gate_output_11_277(.a(output_12_277), .b(output_12_6), .y(output_11_277));
wire output_13_277, output_13_6, output_12_277;
mixer gate_output_12_277(.a(output_13_277), .b(output_13_6), .y(output_12_277));
wire output_14_277, output_14_6, output_13_277;
mixer gate_output_13_277(.a(output_14_277), .b(output_14_6), .y(output_13_277));
wire output_15_277, output_15_6, output_14_277;
mixer gate_output_14_277(.a(output_15_277), .b(output_15_6), .y(output_14_277));
wire output_16_277, output_16_6, output_15_277;
mixer gate_output_15_277(.a(output_16_277), .b(output_16_6), .y(output_15_277));
wire output_1_278, output_1_7, output_0_278;
mixer gate_output_0_278(.a(output_1_278), .b(output_1_7), .y(output_0_278));
wire output_2_278, output_2_7, output_1_278;
mixer gate_output_1_278(.a(output_2_278), .b(output_2_7), .y(output_1_278));
wire output_3_278, output_3_7, output_2_278;
mixer gate_output_2_278(.a(output_3_278), .b(output_3_7), .y(output_2_278));
wire output_4_278, output_4_7, output_3_278;
mixer gate_output_3_278(.a(output_4_278), .b(output_4_7), .y(output_3_278));
wire output_5_278, output_5_7, output_4_278;
mixer gate_output_4_278(.a(output_5_278), .b(output_5_7), .y(output_4_278));
wire output_6_278, output_6_7, output_5_278;
mixer gate_output_5_278(.a(output_6_278), .b(output_6_7), .y(output_5_278));
wire output_7_278, output_7_7, output_6_278;
mixer gate_output_6_278(.a(output_7_278), .b(output_7_7), .y(output_6_278));
wire output_8_278, output_8_7, output_7_278;
mixer gate_output_7_278(.a(output_8_278), .b(output_8_7), .y(output_7_278));
wire output_9_278, output_9_7, output_8_278;
mixer gate_output_8_278(.a(output_9_278), .b(output_9_7), .y(output_8_278));
wire output_10_278, output_10_7, output_9_278;
mixer gate_output_9_278(.a(output_10_278), .b(output_10_7), .y(output_9_278));
wire output_11_278, output_11_7, output_10_278;
mixer gate_output_10_278(.a(output_11_278), .b(output_11_7), .y(output_10_278));
wire output_12_278, output_12_7, output_11_278;
mixer gate_output_11_278(.a(output_12_278), .b(output_12_7), .y(output_11_278));
wire output_13_278, output_13_7, output_12_278;
mixer gate_output_12_278(.a(output_13_278), .b(output_13_7), .y(output_12_278));
wire output_14_278, output_14_7, output_13_278;
mixer gate_output_13_278(.a(output_14_278), .b(output_14_7), .y(output_13_278));
wire output_15_278, output_15_7, output_14_278;
mixer gate_output_14_278(.a(output_15_278), .b(output_15_7), .y(output_14_278));
wire output_16_278, output_16_7, output_15_278;
mixer gate_output_15_278(.a(output_16_278), .b(output_16_7), .y(output_15_278));
wire output_1_279, output_1_8, output_0_279;
mixer gate_output_0_279(.a(output_1_279), .b(output_1_8), .y(output_0_279));
wire output_2_279, output_2_8, output_1_279;
mixer gate_output_1_279(.a(output_2_279), .b(output_2_8), .y(output_1_279));
wire output_3_279, output_3_8, output_2_279;
mixer gate_output_2_279(.a(output_3_279), .b(output_3_8), .y(output_2_279));
wire output_4_279, output_4_8, output_3_279;
mixer gate_output_3_279(.a(output_4_279), .b(output_4_8), .y(output_3_279));
wire output_5_279, output_5_8, output_4_279;
mixer gate_output_4_279(.a(output_5_279), .b(output_5_8), .y(output_4_279));
wire output_6_279, output_6_8, output_5_279;
mixer gate_output_5_279(.a(output_6_279), .b(output_6_8), .y(output_5_279));
wire output_7_279, output_7_8, output_6_279;
mixer gate_output_6_279(.a(output_7_279), .b(output_7_8), .y(output_6_279));
wire output_8_279, output_8_8, output_7_279;
mixer gate_output_7_279(.a(output_8_279), .b(output_8_8), .y(output_7_279));
wire output_9_279, output_9_8, output_8_279;
mixer gate_output_8_279(.a(output_9_279), .b(output_9_8), .y(output_8_279));
wire output_10_279, output_10_8, output_9_279;
mixer gate_output_9_279(.a(output_10_279), .b(output_10_8), .y(output_9_279));
wire output_11_279, output_11_8, output_10_279;
mixer gate_output_10_279(.a(output_11_279), .b(output_11_8), .y(output_10_279));
wire output_12_279, output_12_8, output_11_279;
mixer gate_output_11_279(.a(output_12_279), .b(output_12_8), .y(output_11_279));
wire output_13_279, output_13_8, output_12_279;
mixer gate_output_12_279(.a(output_13_279), .b(output_13_8), .y(output_12_279));
wire output_14_279, output_14_8, output_13_279;
mixer gate_output_13_279(.a(output_14_279), .b(output_14_8), .y(output_13_279));
wire output_15_279, output_15_8, output_14_279;
mixer gate_output_14_279(.a(output_15_279), .b(output_15_8), .y(output_14_279));
wire output_16_279, output_16_8, output_15_279;
mixer gate_output_15_279(.a(output_16_279), .b(output_16_8), .y(output_15_279));
wire output_1_280, output_1_9, output_0_280;
mixer gate_output_0_280(.a(output_1_280), .b(output_1_9), .y(output_0_280));
wire output_2_280, output_2_9, output_1_280;
mixer gate_output_1_280(.a(output_2_280), .b(output_2_9), .y(output_1_280));
wire output_3_280, output_3_9, output_2_280;
mixer gate_output_2_280(.a(output_3_280), .b(output_3_9), .y(output_2_280));
wire output_4_280, output_4_9, output_3_280;
mixer gate_output_3_280(.a(output_4_280), .b(output_4_9), .y(output_3_280));
wire output_5_280, output_5_9, output_4_280;
mixer gate_output_4_280(.a(output_5_280), .b(output_5_9), .y(output_4_280));
wire output_6_280, output_6_9, output_5_280;
mixer gate_output_5_280(.a(output_6_280), .b(output_6_9), .y(output_5_280));
wire output_7_280, output_7_9, output_6_280;
mixer gate_output_6_280(.a(output_7_280), .b(output_7_9), .y(output_6_280));
wire output_8_280, output_8_9, output_7_280;
mixer gate_output_7_280(.a(output_8_280), .b(output_8_9), .y(output_7_280));
wire output_9_280, output_9_9, output_8_280;
mixer gate_output_8_280(.a(output_9_280), .b(output_9_9), .y(output_8_280));
wire output_10_280, output_10_9, output_9_280;
mixer gate_output_9_280(.a(output_10_280), .b(output_10_9), .y(output_9_280));
wire output_11_280, output_11_9, output_10_280;
mixer gate_output_10_280(.a(output_11_280), .b(output_11_9), .y(output_10_280));
wire output_12_280, output_12_9, output_11_280;
mixer gate_output_11_280(.a(output_12_280), .b(output_12_9), .y(output_11_280));
wire output_13_280, output_13_9, output_12_280;
mixer gate_output_12_280(.a(output_13_280), .b(output_13_9), .y(output_12_280));
wire output_14_280, output_14_9, output_13_280;
mixer gate_output_13_280(.a(output_14_280), .b(output_14_9), .y(output_13_280));
wire output_15_280, output_15_9, output_14_280;
mixer gate_output_14_280(.a(output_15_280), .b(output_15_9), .y(output_14_280));
wire output_16_280, output_16_9, output_15_280;
mixer gate_output_15_280(.a(output_16_280), .b(output_16_9), .y(output_15_280));
wire output_1_281, output_1_10, output_0_281;
mixer gate_output_0_281(.a(output_1_281), .b(output_1_10), .y(output_0_281));
wire output_2_281, output_2_10, output_1_281;
mixer gate_output_1_281(.a(output_2_281), .b(output_2_10), .y(output_1_281));
wire output_3_281, output_3_10, output_2_281;
mixer gate_output_2_281(.a(output_3_281), .b(output_3_10), .y(output_2_281));
wire output_4_281, output_4_10, output_3_281;
mixer gate_output_3_281(.a(output_4_281), .b(output_4_10), .y(output_3_281));
wire output_5_281, output_5_10, output_4_281;
mixer gate_output_4_281(.a(output_5_281), .b(output_5_10), .y(output_4_281));
wire output_6_281, output_6_10, output_5_281;
mixer gate_output_5_281(.a(output_6_281), .b(output_6_10), .y(output_5_281));
wire output_7_281, output_7_10, output_6_281;
mixer gate_output_6_281(.a(output_7_281), .b(output_7_10), .y(output_6_281));
wire output_8_281, output_8_10, output_7_281;
mixer gate_output_7_281(.a(output_8_281), .b(output_8_10), .y(output_7_281));
wire output_9_281, output_9_10, output_8_281;
mixer gate_output_8_281(.a(output_9_281), .b(output_9_10), .y(output_8_281));
wire output_10_281, output_10_10, output_9_281;
mixer gate_output_9_281(.a(output_10_281), .b(output_10_10), .y(output_9_281));
wire output_11_281, output_11_10, output_10_281;
mixer gate_output_10_281(.a(output_11_281), .b(output_11_10), .y(output_10_281));
wire output_12_281, output_12_10, output_11_281;
mixer gate_output_11_281(.a(output_12_281), .b(output_12_10), .y(output_11_281));
wire output_13_281, output_13_10, output_12_281;
mixer gate_output_12_281(.a(output_13_281), .b(output_13_10), .y(output_12_281));
wire output_14_281, output_14_10, output_13_281;
mixer gate_output_13_281(.a(output_14_281), .b(output_14_10), .y(output_13_281));
wire output_15_281, output_15_10, output_14_281;
mixer gate_output_14_281(.a(output_15_281), .b(output_15_10), .y(output_14_281));
wire output_16_281, output_16_10, output_15_281;
mixer gate_output_15_281(.a(output_16_281), .b(output_16_10), .y(output_15_281));
wire output_1_282, output_1_11, output_0_282;
mixer gate_output_0_282(.a(output_1_282), .b(output_1_11), .y(output_0_282));
wire output_2_282, output_2_11, output_1_282;
mixer gate_output_1_282(.a(output_2_282), .b(output_2_11), .y(output_1_282));
wire output_3_282, output_3_11, output_2_282;
mixer gate_output_2_282(.a(output_3_282), .b(output_3_11), .y(output_2_282));
wire output_4_282, output_4_11, output_3_282;
mixer gate_output_3_282(.a(output_4_282), .b(output_4_11), .y(output_3_282));
wire output_5_282, output_5_11, output_4_282;
mixer gate_output_4_282(.a(output_5_282), .b(output_5_11), .y(output_4_282));
wire output_6_282, output_6_11, output_5_282;
mixer gate_output_5_282(.a(output_6_282), .b(output_6_11), .y(output_5_282));
wire output_7_282, output_7_11, output_6_282;
mixer gate_output_6_282(.a(output_7_282), .b(output_7_11), .y(output_6_282));
wire output_8_282, output_8_11, output_7_282;
mixer gate_output_7_282(.a(output_8_282), .b(output_8_11), .y(output_7_282));
wire output_9_282, output_9_11, output_8_282;
mixer gate_output_8_282(.a(output_9_282), .b(output_9_11), .y(output_8_282));
wire output_10_282, output_10_11, output_9_282;
mixer gate_output_9_282(.a(output_10_282), .b(output_10_11), .y(output_9_282));
wire output_11_282, output_11_11, output_10_282;
mixer gate_output_10_282(.a(output_11_282), .b(output_11_11), .y(output_10_282));
wire output_12_282, output_12_11, output_11_282;
mixer gate_output_11_282(.a(output_12_282), .b(output_12_11), .y(output_11_282));
wire output_13_282, output_13_11, output_12_282;
mixer gate_output_12_282(.a(output_13_282), .b(output_13_11), .y(output_12_282));
wire output_14_282, output_14_11, output_13_282;
mixer gate_output_13_282(.a(output_14_282), .b(output_14_11), .y(output_13_282));
wire output_15_282, output_15_11, output_14_282;
mixer gate_output_14_282(.a(output_15_282), .b(output_15_11), .y(output_14_282));
wire output_16_282, output_16_11, output_15_282;
mixer gate_output_15_282(.a(output_16_282), .b(output_16_11), .y(output_15_282));
wire output_1_283, output_1_12, output_0_283;
mixer gate_output_0_283(.a(output_1_283), .b(output_1_12), .y(output_0_283));
wire output_2_283, output_2_12, output_1_283;
mixer gate_output_1_283(.a(output_2_283), .b(output_2_12), .y(output_1_283));
wire output_3_283, output_3_12, output_2_283;
mixer gate_output_2_283(.a(output_3_283), .b(output_3_12), .y(output_2_283));
wire output_4_283, output_4_12, output_3_283;
mixer gate_output_3_283(.a(output_4_283), .b(output_4_12), .y(output_3_283));
wire output_5_283, output_5_12, output_4_283;
mixer gate_output_4_283(.a(output_5_283), .b(output_5_12), .y(output_4_283));
wire output_6_283, output_6_12, output_5_283;
mixer gate_output_5_283(.a(output_6_283), .b(output_6_12), .y(output_5_283));
wire output_7_283, output_7_12, output_6_283;
mixer gate_output_6_283(.a(output_7_283), .b(output_7_12), .y(output_6_283));
wire output_8_283, output_8_12, output_7_283;
mixer gate_output_7_283(.a(output_8_283), .b(output_8_12), .y(output_7_283));
wire output_9_283, output_9_12, output_8_283;
mixer gate_output_8_283(.a(output_9_283), .b(output_9_12), .y(output_8_283));
wire output_10_283, output_10_12, output_9_283;
mixer gate_output_9_283(.a(output_10_283), .b(output_10_12), .y(output_9_283));
wire output_11_283, output_11_12, output_10_283;
mixer gate_output_10_283(.a(output_11_283), .b(output_11_12), .y(output_10_283));
wire output_12_283, output_12_12, output_11_283;
mixer gate_output_11_283(.a(output_12_283), .b(output_12_12), .y(output_11_283));
wire output_13_283, output_13_12, output_12_283;
mixer gate_output_12_283(.a(output_13_283), .b(output_13_12), .y(output_12_283));
wire output_14_283, output_14_12, output_13_283;
mixer gate_output_13_283(.a(output_14_283), .b(output_14_12), .y(output_13_283));
wire output_15_283, output_15_12, output_14_283;
mixer gate_output_14_283(.a(output_15_283), .b(output_15_12), .y(output_14_283));
wire output_16_283, output_16_12, output_15_283;
mixer gate_output_15_283(.a(output_16_283), .b(output_16_12), .y(output_15_283));
wire output_1_284, output_1_13, output_0_284;
mixer gate_output_0_284(.a(output_1_284), .b(output_1_13), .y(output_0_284));
wire output_2_284, output_2_13, output_1_284;
mixer gate_output_1_284(.a(output_2_284), .b(output_2_13), .y(output_1_284));
wire output_3_284, output_3_13, output_2_284;
mixer gate_output_2_284(.a(output_3_284), .b(output_3_13), .y(output_2_284));
wire output_4_284, output_4_13, output_3_284;
mixer gate_output_3_284(.a(output_4_284), .b(output_4_13), .y(output_3_284));
wire output_5_284, output_5_13, output_4_284;
mixer gate_output_4_284(.a(output_5_284), .b(output_5_13), .y(output_4_284));
wire output_6_284, output_6_13, output_5_284;
mixer gate_output_5_284(.a(output_6_284), .b(output_6_13), .y(output_5_284));
wire output_7_284, output_7_13, output_6_284;
mixer gate_output_6_284(.a(output_7_284), .b(output_7_13), .y(output_6_284));
wire output_8_284, output_8_13, output_7_284;
mixer gate_output_7_284(.a(output_8_284), .b(output_8_13), .y(output_7_284));
wire output_9_284, output_9_13, output_8_284;
mixer gate_output_8_284(.a(output_9_284), .b(output_9_13), .y(output_8_284));
wire output_10_284, output_10_13, output_9_284;
mixer gate_output_9_284(.a(output_10_284), .b(output_10_13), .y(output_9_284));
wire output_11_284, output_11_13, output_10_284;
mixer gate_output_10_284(.a(output_11_284), .b(output_11_13), .y(output_10_284));
wire output_12_284, output_12_13, output_11_284;
mixer gate_output_11_284(.a(output_12_284), .b(output_12_13), .y(output_11_284));
wire output_13_284, output_13_13, output_12_284;
mixer gate_output_12_284(.a(output_13_284), .b(output_13_13), .y(output_12_284));
wire output_14_284, output_14_13, output_13_284;
mixer gate_output_13_284(.a(output_14_284), .b(output_14_13), .y(output_13_284));
wire output_15_284, output_15_13, output_14_284;
mixer gate_output_14_284(.a(output_15_284), .b(output_15_13), .y(output_14_284));
wire output_16_284, output_16_13, output_15_284;
mixer gate_output_15_284(.a(output_16_284), .b(output_16_13), .y(output_15_284));
wire output_1_285, output_1_14, output_0_285;
mixer gate_output_0_285(.a(output_1_285), .b(output_1_14), .y(output_0_285));
wire output_2_285, output_2_14, output_1_285;
mixer gate_output_1_285(.a(output_2_285), .b(output_2_14), .y(output_1_285));
wire output_3_285, output_3_14, output_2_285;
mixer gate_output_2_285(.a(output_3_285), .b(output_3_14), .y(output_2_285));
wire output_4_285, output_4_14, output_3_285;
mixer gate_output_3_285(.a(output_4_285), .b(output_4_14), .y(output_3_285));
wire output_5_285, output_5_14, output_4_285;
mixer gate_output_4_285(.a(output_5_285), .b(output_5_14), .y(output_4_285));
wire output_6_285, output_6_14, output_5_285;
mixer gate_output_5_285(.a(output_6_285), .b(output_6_14), .y(output_5_285));
wire output_7_285, output_7_14, output_6_285;
mixer gate_output_6_285(.a(output_7_285), .b(output_7_14), .y(output_6_285));
wire output_8_285, output_8_14, output_7_285;
mixer gate_output_7_285(.a(output_8_285), .b(output_8_14), .y(output_7_285));
wire output_9_285, output_9_14, output_8_285;
mixer gate_output_8_285(.a(output_9_285), .b(output_9_14), .y(output_8_285));
wire output_10_285, output_10_14, output_9_285;
mixer gate_output_9_285(.a(output_10_285), .b(output_10_14), .y(output_9_285));
wire output_11_285, output_11_14, output_10_285;
mixer gate_output_10_285(.a(output_11_285), .b(output_11_14), .y(output_10_285));
wire output_12_285, output_12_14, output_11_285;
mixer gate_output_11_285(.a(output_12_285), .b(output_12_14), .y(output_11_285));
wire output_13_285, output_13_14, output_12_285;
mixer gate_output_12_285(.a(output_13_285), .b(output_13_14), .y(output_12_285));
wire output_14_285, output_14_14, output_13_285;
mixer gate_output_13_285(.a(output_14_285), .b(output_14_14), .y(output_13_285));
wire output_15_285, output_15_14, output_14_285;
mixer gate_output_14_285(.a(output_15_285), .b(output_15_14), .y(output_14_285));
wire output_16_285, output_16_14, output_15_285;
mixer gate_output_15_285(.a(output_16_285), .b(output_16_14), .y(output_15_285));
wire output_1_286, output_1_15, output_0_286;
mixer gate_output_0_286(.a(output_1_286), .b(output_1_15), .y(output_0_286));
wire output_2_286, output_2_15, output_1_286;
mixer gate_output_1_286(.a(output_2_286), .b(output_2_15), .y(output_1_286));
wire output_3_286, output_3_15, output_2_286;
mixer gate_output_2_286(.a(output_3_286), .b(output_3_15), .y(output_2_286));
wire output_4_286, output_4_15, output_3_286;
mixer gate_output_3_286(.a(output_4_286), .b(output_4_15), .y(output_3_286));
wire output_5_286, output_5_15, output_4_286;
mixer gate_output_4_286(.a(output_5_286), .b(output_5_15), .y(output_4_286));
wire output_6_286, output_6_15, output_5_286;
mixer gate_output_5_286(.a(output_6_286), .b(output_6_15), .y(output_5_286));
wire output_7_286, output_7_15, output_6_286;
mixer gate_output_6_286(.a(output_7_286), .b(output_7_15), .y(output_6_286));
wire output_8_286, output_8_15, output_7_286;
mixer gate_output_7_286(.a(output_8_286), .b(output_8_15), .y(output_7_286));
wire output_9_286, output_9_15, output_8_286;
mixer gate_output_8_286(.a(output_9_286), .b(output_9_15), .y(output_8_286));
wire output_10_286, output_10_15, output_9_286;
mixer gate_output_9_286(.a(output_10_286), .b(output_10_15), .y(output_9_286));
wire output_11_286, output_11_15, output_10_286;
mixer gate_output_10_286(.a(output_11_286), .b(output_11_15), .y(output_10_286));
wire output_12_286, output_12_15, output_11_286;
mixer gate_output_11_286(.a(output_12_286), .b(output_12_15), .y(output_11_286));
wire output_13_286, output_13_15, output_12_286;
mixer gate_output_12_286(.a(output_13_286), .b(output_13_15), .y(output_12_286));
wire output_14_286, output_14_15, output_13_286;
mixer gate_output_13_286(.a(output_14_286), .b(output_14_15), .y(output_13_286));
wire output_15_286, output_15_15, output_14_286;
mixer gate_output_14_286(.a(output_15_286), .b(output_15_15), .y(output_14_286));
wire output_16_286, output_16_15, output_15_286;
mixer gate_output_15_286(.a(output_16_286), .b(output_16_15), .y(output_15_286));
wire output_1_287, output_1_0, output_0_287;
mixer gate_output_0_287(.a(output_1_287), .b(output_1_0), .y(output_0_287));
wire output_2_287, output_2_0, output_1_287;
mixer gate_output_1_287(.a(output_2_287), .b(output_2_0), .y(output_1_287));
wire output_3_287, output_3_0, output_2_287;
mixer gate_output_2_287(.a(output_3_287), .b(output_3_0), .y(output_2_287));
wire output_4_287, output_4_0, output_3_287;
mixer gate_output_3_287(.a(output_4_287), .b(output_4_0), .y(output_3_287));
wire output_5_287, output_5_0, output_4_287;
mixer gate_output_4_287(.a(output_5_287), .b(output_5_0), .y(output_4_287));
wire output_6_287, output_6_0, output_5_287;
mixer gate_output_5_287(.a(output_6_287), .b(output_6_0), .y(output_5_287));
wire output_7_287, output_7_0, output_6_287;
mixer gate_output_6_287(.a(output_7_287), .b(output_7_0), .y(output_6_287));
wire output_8_287, output_8_0, output_7_287;
mixer gate_output_7_287(.a(output_8_287), .b(output_8_0), .y(output_7_287));
wire output_9_287, output_9_0, output_8_287;
mixer gate_output_8_287(.a(output_9_287), .b(output_9_0), .y(output_8_287));
wire output_10_287, output_10_0, output_9_287;
mixer gate_output_9_287(.a(output_10_287), .b(output_10_0), .y(output_9_287));
wire output_11_287, output_11_0, output_10_287;
mixer gate_output_10_287(.a(output_11_287), .b(output_11_0), .y(output_10_287));
wire output_12_287, output_12_0, output_11_287;
mixer gate_output_11_287(.a(output_12_287), .b(output_12_0), .y(output_11_287));
wire output_13_287, output_13_0, output_12_287;
mixer gate_output_12_287(.a(output_13_287), .b(output_13_0), .y(output_12_287));
wire output_14_287, output_14_0, output_13_287;
mixer gate_output_13_287(.a(output_14_287), .b(output_14_0), .y(output_13_287));
wire output_15_287, output_15_0, output_14_287;
mixer gate_output_14_287(.a(output_15_287), .b(output_15_0), .y(output_14_287));
wire output_16_287, output_16_0, output_15_287;
mixer gate_output_15_287(.a(output_16_287), .b(output_16_0), .y(output_15_287));
wire output_1_288, output_1_1, output_0_288;
mixer gate_output_0_288(.a(output_1_288), .b(output_1_1), .y(output_0_288));
wire output_2_288, output_2_1, output_1_288;
mixer gate_output_1_288(.a(output_2_288), .b(output_2_1), .y(output_1_288));
wire output_3_288, output_3_1, output_2_288;
mixer gate_output_2_288(.a(output_3_288), .b(output_3_1), .y(output_2_288));
wire output_4_288, output_4_1, output_3_288;
mixer gate_output_3_288(.a(output_4_288), .b(output_4_1), .y(output_3_288));
wire output_5_288, output_5_1, output_4_288;
mixer gate_output_4_288(.a(output_5_288), .b(output_5_1), .y(output_4_288));
wire output_6_288, output_6_1, output_5_288;
mixer gate_output_5_288(.a(output_6_288), .b(output_6_1), .y(output_5_288));
wire output_7_288, output_7_1, output_6_288;
mixer gate_output_6_288(.a(output_7_288), .b(output_7_1), .y(output_6_288));
wire output_8_288, output_8_1, output_7_288;
mixer gate_output_7_288(.a(output_8_288), .b(output_8_1), .y(output_7_288));
wire output_9_288, output_9_1, output_8_288;
mixer gate_output_8_288(.a(output_9_288), .b(output_9_1), .y(output_8_288));
wire output_10_288, output_10_1, output_9_288;
mixer gate_output_9_288(.a(output_10_288), .b(output_10_1), .y(output_9_288));
wire output_11_288, output_11_1, output_10_288;
mixer gate_output_10_288(.a(output_11_288), .b(output_11_1), .y(output_10_288));
wire output_12_288, output_12_1, output_11_288;
mixer gate_output_11_288(.a(output_12_288), .b(output_12_1), .y(output_11_288));
wire output_13_288, output_13_1, output_12_288;
mixer gate_output_12_288(.a(output_13_288), .b(output_13_1), .y(output_12_288));
wire output_14_288, output_14_1, output_13_288;
mixer gate_output_13_288(.a(output_14_288), .b(output_14_1), .y(output_13_288));
wire output_15_288, output_15_1, output_14_288;
mixer gate_output_14_288(.a(output_15_288), .b(output_15_1), .y(output_14_288));
wire output_16_288, output_16_1, output_15_288;
mixer gate_output_15_288(.a(output_16_288), .b(output_16_1), .y(output_15_288));
wire output_1_289, output_1_2, output_0_289;
mixer gate_output_0_289(.a(output_1_289), .b(output_1_2), .y(output_0_289));
wire output_2_289, output_2_2, output_1_289;
mixer gate_output_1_289(.a(output_2_289), .b(output_2_2), .y(output_1_289));
wire output_3_289, output_3_2, output_2_289;
mixer gate_output_2_289(.a(output_3_289), .b(output_3_2), .y(output_2_289));
wire output_4_289, output_4_2, output_3_289;
mixer gate_output_3_289(.a(output_4_289), .b(output_4_2), .y(output_3_289));
wire output_5_289, output_5_2, output_4_289;
mixer gate_output_4_289(.a(output_5_289), .b(output_5_2), .y(output_4_289));
wire output_6_289, output_6_2, output_5_289;
mixer gate_output_5_289(.a(output_6_289), .b(output_6_2), .y(output_5_289));
wire output_7_289, output_7_2, output_6_289;
mixer gate_output_6_289(.a(output_7_289), .b(output_7_2), .y(output_6_289));
wire output_8_289, output_8_2, output_7_289;
mixer gate_output_7_289(.a(output_8_289), .b(output_8_2), .y(output_7_289));
wire output_9_289, output_9_2, output_8_289;
mixer gate_output_8_289(.a(output_9_289), .b(output_9_2), .y(output_8_289));
wire output_10_289, output_10_2, output_9_289;
mixer gate_output_9_289(.a(output_10_289), .b(output_10_2), .y(output_9_289));
wire output_11_289, output_11_2, output_10_289;
mixer gate_output_10_289(.a(output_11_289), .b(output_11_2), .y(output_10_289));
wire output_12_289, output_12_2, output_11_289;
mixer gate_output_11_289(.a(output_12_289), .b(output_12_2), .y(output_11_289));
wire output_13_289, output_13_2, output_12_289;
mixer gate_output_12_289(.a(output_13_289), .b(output_13_2), .y(output_12_289));
wire output_14_289, output_14_2, output_13_289;
mixer gate_output_13_289(.a(output_14_289), .b(output_14_2), .y(output_13_289));
wire output_15_289, output_15_2, output_14_289;
mixer gate_output_14_289(.a(output_15_289), .b(output_15_2), .y(output_14_289));
wire output_16_289, output_16_2, output_15_289;
mixer gate_output_15_289(.a(output_16_289), .b(output_16_2), .y(output_15_289));
wire output_1_290, output_1_3, output_0_290;
mixer gate_output_0_290(.a(output_1_290), .b(output_1_3), .y(output_0_290));
wire output_2_290, output_2_3, output_1_290;
mixer gate_output_1_290(.a(output_2_290), .b(output_2_3), .y(output_1_290));
wire output_3_290, output_3_3, output_2_290;
mixer gate_output_2_290(.a(output_3_290), .b(output_3_3), .y(output_2_290));
wire output_4_290, output_4_3, output_3_290;
mixer gate_output_3_290(.a(output_4_290), .b(output_4_3), .y(output_3_290));
wire output_5_290, output_5_3, output_4_290;
mixer gate_output_4_290(.a(output_5_290), .b(output_5_3), .y(output_4_290));
wire output_6_290, output_6_3, output_5_290;
mixer gate_output_5_290(.a(output_6_290), .b(output_6_3), .y(output_5_290));
wire output_7_290, output_7_3, output_6_290;
mixer gate_output_6_290(.a(output_7_290), .b(output_7_3), .y(output_6_290));
wire output_8_290, output_8_3, output_7_290;
mixer gate_output_7_290(.a(output_8_290), .b(output_8_3), .y(output_7_290));
wire output_9_290, output_9_3, output_8_290;
mixer gate_output_8_290(.a(output_9_290), .b(output_9_3), .y(output_8_290));
wire output_10_290, output_10_3, output_9_290;
mixer gate_output_9_290(.a(output_10_290), .b(output_10_3), .y(output_9_290));
wire output_11_290, output_11_3, output_10_290;
mixer gate_output_10_290(.a(output_11_290), .b(output_11_3), .y(output_10_290));
wire output_12_290, output_12_3, output_11_290;
mixer gate_output_11_290(.a(output_12_290), .b(output_12_3), .y(output_11_290));
wire output_13_290, output_13_3, output_12_290;
mixer gate_output_12_290(.a(output_13_290), .b(output_13_3), .y(output_12_290));
wire output_14_290, output_14_3, output_13_290;
mixer gate_output_13_290(.a(output_14_290), .b(output_14_3), .y(output_13_290));
wire output_15_290, output_15_3, output_14_290;
mixer gate_output_14_290(.a(output_15_290), .b(output_15_3), .y(output_14_290));
wire output_16_290, output_16_3, output_15_290;
mixer gate_output_15_290(.a(output_16_290), .b(output_16_3), .y(output_15_290));
wire output_1_291, output_1_4, output_0_291;
mixer gate_output_0_291(.a(output_1_291), .b(output_1_4), .y(output_0_291));
wire output_2_291, output_2_4, output_1_291;
mixer gate_output_1_291(.a(output_2_291), .b(output_2_4), .y(output_1_291));
wire output_3_291, output_3_4, output_2_291;
mixer gate_output_2_291(.a(output_3_291), .b(output_3_4), .y(output_2_291));
wire output_4_291, output_4_4, output_3_291;
mixer gate_output_3_291(.a(output_4_291), .b(output_4_4), .y(output_3_291));
wire output_5_291, output_5_4, output_4_291;
mixer gate_output_4_291(.a(output_5_291), .b(output_5_4), .y(output_4_291));
wire output_6_291, output_6_4, output_5_291;
mixer gate_output_5_291(.a(output_6_291), .b(output_6_4), .y(output_5_291));
wire output_7_291, output_7_4, output_6_291;
mixer gate_output_6_291(.a(output_7_291), .b(output_7_4), .y(output_6_291));
wire output_8_291, output_8_4, output_7_291;
mixer gate_output_7_291(.a(output_8_291), .b(output_8_4), .y(output_7_291));
wire output_9_291, output_9_4, output_8_291;
mixer gate_output_8_291(.a(output_9_291), .b(output_9_4), .y(output_8_291));
wire output_10_291, output_10_4, output_9_291;
mixer gate_output_9_291(.a(output_10_291), .b(output_10_4), .y(output_9_291));
wire output_11_291, output_11_4, output_10_291;
mixer gate_output_10_291(.a(output_11_291), .b(output_11_4), .y(output_10_291));
wire output_12_291, output_12_4, output_11_291;
mixer gate_output_11_291(.a(output_12_291), .b(output_12_4), .y(output_11_291));
wire output_13_291, output_13_4, output_12_291;
mixer gate_output_12_291(.a(output_13_291), .b(output_13_4), .y(output_12_291));
wire output_14_291, output_14_4, output_13_291;
mixer gate_output_13_291(.a(output_14_291), .b(output_14_4), .y(output_13_291));
wire output_15_291, output_15_4, output_14_291;
mixer gate_output_14_291(.a(output_15_291), .b(output_15_4), .y(output_14_291));
wire output_16_291, output_16_4, output_15_291;
mixer gate_output_15_291(.a(output_16_291), .b(output_16_4), .y(output_15_291));
wire output_1_292, output_1_5, output_0_292;
mixer gate_output_0_292(.a(output_1_292), .b(output_1_5), .y(output_0_292));
wire output_2_292, output_2_5, output_1_292;
mixer gate_output_1_292(.a(output_2_292), .b(output_2_5), .y(output_1_292));
wire output_3_292, output_3_5, output_2_292;
mixer gate_output_2_292(.a(output_3_292), .b(output_3_5), .y(output_2_292));
wire output_4_292, output_4_5, output_3_292;
mixer gate_output_3_292(.a(output_4_292), .b(output_4_5), .y(output_3_292));
wire output_5_292, output_5_5, output_4_292;
mixer gate_output_4_292(.a(output_5_292), .b(output_5_5), .y(output_4_292));
wire output_6_292, output_6_5, output_5_292;
mixer gate_output_5_292(.a(output_6_292), .b(output_6_5), .y(output_5_292));
wire output_7_292, output_7_5, output_6_292;
mixer gate_output_6_292(.a(output_7_292), .b(output_7_5), .y(output_6_292));
wire output_8_292, output_8_5, output_7_292;
mixer gate_output_7_292(.a(output_8_292), .b(output_8_5), .y(output_7_292));
wire output_9_292, output_9_5, output_8_292;
mixer gate_output_8_292(.a(output_9_292), .b(output_9_5), .y(output_8_292));
wire output_10_292, output_10_5, output_9_292;
mixer gate_output_9_292(.a(output_10_292), .b(output_10_5), .y(output_9_292));
wire output_11_292, output_11_5, output_10_292;
mixer gate_output_10_292(.a(output_11_292), .b(output_11_5), .y(output_10_292));
wire output_12_292, output_12_5, output_11_292;
mixer gate_output_11_292(.a(output_12_292), .b(output_12_5), .y(output_11_292));
wire output_13_292, output_13_5, output_12_292;
mixer gate_output_12_292(.a(output_13_292), .b(output_13_5), .y(output_12_292));
wire output_14_292, output_14_5, output_13_292;
mixer gate_output_13_292(.a(output_14_292), .b(output_14_5), .y(output_13_292));
wire output_15_292, output_15_5, output_14_292;
mixer gate_output_14_292(.a(output_15_292), .b(output_15_5), .y(output_14_292));
wire output_16_292, output_16_5, output_15_292;
mixer gate_output_15_292(.a(output_16_292), .b(output_16_5), .y(output_15_292));
wire output_1_293, output_1_6, output_0_293;
mixer gate_output_0_293(.a(output_1_293), .b(output_1_6), .y(output_0_293));
wire output_2_293, output_2_6, output_1_293;
mixer gate_output_1_293(.a(output_2_293), .b(output_2_6), .y(output_1_293));
wire output_3_293, output_3_6, output_2_293;
mixer gate_output_2_293(.a(output_3_293), .b(output_3_6), .y(output_2_293));
wire output_4_293, output_4_6, output_3_293;
mixer gate_output_3_293(.a(output_4_293), .b(output_4_6), .y(output_3_293));
wire output_5_293, output_5_6, output_4_293;
mixer gate_output_4_293(.a(output_5_293), .b(output_5_6), .y(output_4_293));
wire output_6_293, output_6_6, output_5_293;
mixer gate_output_5_293(.a(output_6_293), .b(output_6_6), .y(output_5_293));
wire output_7_293, output_7_6, output_6_293;
mixer gate_output_6_293(.a(output_7_293), .b(output_7_6), .y(output_6_293));
wire output_8_293, output_8_6, output_7_293;
mixer gate_output_7_293(.a(output_8_293), .b(output_8_6), .y(output_7_293));
wire output_9_293, output_9_6, output_8_293;
mixer gate_output_8_293(.a(output_9_293), .b(output_9_6), .y(output_8_293));
wire output_10_293, output_10_6, output_9_293;
mixer gate_output_9_293(.a(output_10_293), .b(output_10_6), .y(output_9_293));
wire output_11_293, output_11_6, output_10_293;
mixer gate_output_10_293(.a(output_11_293), .b(output_11_6), .y(output_10_293));
wire output_12_293, output_12_6, output_11_293;
mixer gate_output_11_293(.a(output_12_293), .b(output_12_6), .y(output_11_293));
wire output_13_293, output_13_6, output_12_293;
mixer gate_output_12_293(.a(output_13_293), .b(output_13_6), .y(output_12_293));
wire output_14_293, output_14_6, output_13_293;
mixer gate_output_13_293(.a(output_14_293), .b(output_14_6), .y(output_13_293));
wire output_15_293, output_15_6, output_14_293;
mixer gate_output_14_293(.a(output_15_293), .b(output_15_6), .y(output_14_293));
wire output_16_293, output_16_6, output_15_293;
mixer gate_output_15_293(.a(output_16_293), .b(output_16_6), .y(output_15_293));
wire output_1_294, output_1_7, output_0_294;
mixer gate_output_0_294(.a(output_1_294), .b(output_1_7), .y(output_0_294));
wire output_2_294, output_2_7, output_1_294;
mixer gate_output_1_294(.a(output_2_294), .b(output_2_7), .y(output_1_294));
wire output_3_294, output_3_7, output_2_294;
mixer gate_output_2_294(.a(output_3_294), .b(output_3_7), .y(output_2_294));
wire output_4_294, output_4_7, output_3_294;
mixer gate_output_3_294(.a(output_4_294), .b(output_4_7), .y(output_3_294));
wire output_5_294, output_5_7, output_4_294;
mixer gate_output_4_294(.a(output_5_294), .b(output_5_7), .y(output_4_294));
wire output_6_294, output_6_7, output_5_294;
mixer gate_output_5_294(.a(output_6_294), .b(output_6_7), .y(output_5_294));
wire output_7_294, output_7_7, output_6_294;
mixer gate_output_6_294(.a(output_7_294), .b(output_7_7), .y(output_6_294));
wire output_8_294, output_8_7, output_7_294;
mixer gate_output_7_294(.a(output_8_294), .b(output_8_7), .y(output_7_294));
wire output_9_294, output_9_7, output_8_294;
mixer gate_output_8_294(.a(output_9_294), .b(output_9_7), .y(output_8_294));
wire output_10_294, output_10_7, output_9_294;
mixer gate_output_9_294(.a(output_10_294), .b(output_10_7), .y(output_9_294));
wire output_11_294, output_11_7, output_10_294;
mixer gate_output_10_294(.a(output_11_294), .b(output_11_7), .y(output_10_294));
wire output_12_294, output_12_7, output_11_294;
mixer gate_output_11_294(.a(output_12_294), .b(output_12_7), .y(output_11_294));
wire output_13_294, output_13_7, output_12_294;
mixer gate_output_12_294(.a(output_13_294), .b(output_13_7), .y(output_12_294));
wire output_14_294, output_14_7, output_13_294;
mixer gate_output_13_294(.a(output_14_294), .b(output_14_7), .y(output_13_294));
wire output_15_294, output_15_7, output_14_294;
mixer gate_output_14_294(.a(output_15_294), .b(output_15_7), .y(output_14_294));
wire output_16_294, output_16_7, output_15_294;
mixer gate_output_15_294(.a(output_16_294), .b(output_16_7), .y(output_15_294));
wire output_1_295, output_1_8, output_0_295;
mixer gate_output_0_295(.a(output_1_295), .b(output_1_8), .y(output_0_295));
wire output_2_295, output_2_8, output_1_295;
mixer gate_output_1_295(.a(output_2_295), .b(output_2_8), .y(output_1_295));
wire output_3_295, output_3_8, output_2_295;
mixer gate_output_2_295(.a(output_3_295), .b(output_3_8), .y(output_2_295));
wire output_4_295, output_4_8, output_3_295;
mixer gate_output_3_295(.a(output_4_295), .b(output_4_8), .y(output_3_295));
wire output_5_295, output_5_8, output_4_295;
mixer gate_output_4_295(.a(output_5_295), .b(output_5_8), .y(output_4_295));
wire output_6_295, output_6_8, output_5_295;
mixer gate_output_5_295(.a(output_6_295), .b(output_6_8), .y(output_5_295));
wire output_7_295, output_7_8, output_6_295;
mixer gate_output_6_295(.a(output_7_295), .b(output_7_8), .y(output_6_295));
wire output_8_295, output_8_8, output_7_295;
mixer gate_output_7_295(.a(output_8_295), .b(output_8_8), .y(output_7_295));
wire output_9_295, output_9_8, output_8_295;
mixer gate_output_8_295(.a(output_9_295), .b(output_9_8), .y(output_8_295));
wire output_10_295, output_10_8, output_9_295;
mixer gate_output_9_295(.a(output_10_295), .b(output_10_8), .y(output_9_295));
wire output_11_295, output_11_8, output_10_295;
mixer gate_output_10_295(.a(output_11_295), .b(output_11_8), .y(output_10_295));
wire output_12_295, output_12_8, output_11_295;
mixer gate_output_11_295(.a(output_12_295), .b(output_12_8), .y(output_11_295));
wire output_13_295, output_13_8, output_12_295;
mixer gate_output_12_295(.a(output_13_295), .b(output_13_8), .y(output_12_295));
wire output_14_295, output_14_8, output_13_295;
mixer gate_output_13_295(.a(output_14_295), .b(output_14_8), .y(output_13_295));
wire output_15_295, output_15_8, output_14_295;
mixer gate_output_14_295(.a(output_15_295), .b(output_15_8), .y(output_14_295));
wire output_16_295, output_16_8, output_15_295;
mixer gate_output_15_295(.a(output_16_295), .b(output_16_8), .y(output_15_295));
wire output_1_296, output_1_9, output_0_296;
mixer gate_output_0_296(.a(output_1_296), .b(output_1_9), .y(output_0_296));
wire output_2_296, output_2_9, output_1_296;
mixer gate_output_1_296(.a(output_2_296), .b(output_2_9), .y(output_1_296));
wire output_3_296, output_3_9, output_2_296;
mixer gate_output_2_296(.a(output_3_296), .b(output_3_9), .y(output_2_296));
wire output_4_296, output_4_9, output_3_296;
mixer gate_output_3_296(.a(output_4_296), .b(output_4_9), .y(output_3_296));
wire output_5_296, output_5_9, output_4_296;
mixer gate_output_4_296(.a(output_5_296), .b(output_5_9), .y(output_4_296));
wire output_6_296, output_6_9, output_5_296;
mixer gate_output_5_296(.a(output_6_296), .b(output_6_9), .y(output_5_296));
wire output_7_296, output_7_9, output_6_296;
mixer gate_output_6_296(.a(output_7_296), .b(output_7_9), .y(output_6_296));
wire output_8_296, output_8_9, output_7_296;
mixer gate_output_7_296(.a(output_8_296), .b(output_8_9), .y(output_7_296));
wire output_9_296, output_9_9, output_8_296;
mixer gate_output_8_296(.a(output_9_296), .b(output_9_9), .y(output_8_296));
wire output_10_296, output_10_9, output_9_296;
mixer gate_output_9_296(.a(output_10_296), .b(output_10_9), .y(output_9_296));
wire output_11_296, output_11_9, output_10_296;
mixer gate_output_10_296(.a(output_11_296), .b(output_11_9), .y(output_10_296));
wire output_12_296, output_12_9, output_11_296;
mixer gate_output_11_296(.a(output_12_296), .b(output_12_9), .y(output_11_296));
wire output_13_296, output_13_9, output_12_296;
mixer gate_output_12_296(.a(output_13_296), .b(output_13_9), .y(output_12_296));
wire output_14_296, output_14_9, output_13_296;
mixer gate_output_13_296(.a(output_14_296), .b(output_14_9), .y(output_13_296));
wire output_15_296, output_15_9, output_14_296;
mixer gate_output_14_296(.a(output_15_296), .b(output_15_9), .y(output_14_296));
wire output_16_296, output_16_9, output_15_296;
mixer gate_output_15_296(.a(output_16_296), .b(output_16_9), .y(output_15_296));
wire output_1_297, output_1_10, output_0_297;
mixer gate_output_0_297(.a(output_1_297), .b(output_1_10), .y(output_0_297));
wire output_2_297, output_2_10, output_1_297;
mixer gate_output_1_297(.a(output_2_297), .b(output_2_10), .y(output_1_297));
wire output_3_297, output_3_10, output_2_297;
mixer gate_output_2_297(.a(output_3_297), .b(output_3_10), .y(output_2_297));
wire output_4_297, output_4_10, output_3_297;
mixer gate_output_3_297(.a(output_4_297), .b(output_4_10), .y(output_3_297));
wire output_5_297, output_5_10, output_4_297;
mixer gate_output_4_297(.a(output_5_297), .b(output_5_10), .y(output_4_297));
wire output_6_297, output_6_10, output_5_297;
mixer gate_output_5_297(.a(output_6_297), .b(output_6_10), .y(output_5_297));
wire output_7_297, output_7_10, output_6_297;
mixer gate_output_6_297(.a(output_7_297), .b(output_7_10), .y(output_6_297));
wire output_8_297, output_8_10, output_7_297;
mixer gate_output_7_297(.a(output_8_297), .b(output_8_10), .y(output_7_297));
wire output_9_297, output_9_10, output_8_297;
mixer gate_output_8_297(.a(output_9_297), .b(output_9_10), .y(output_8_297));
wire output_10_297, output_10_10, output_9_297;
mixer gate_output_9_297(.a(output_10_297), .b(output_10_10), .y(output_9_297));
wire output_11_297, output_11_10, output_10_297;
mixer gate_output_10_297(.a(output_11_297), .b(output_11_10), .y(output_10_297));
wire output_12_297, output_12_10, output_11_297;
mixer gate_output_11_297(.a(output_12_297), .b(output_12_10), .y(output_11_297));
wire output_13_297, output_13_10, output_12_297;
mixer gate_output_12_297(.a(output_13_297), .b(output_13_10), .y(output_12_297));
wire output_14_297, output_14_10, output_13_297;
mixer gate_output_13_297(.a(output_14_297), .b(output_14_10), .y(output_13_297));
wire output_15_297, output_15_10, output_14_297;
mixer gate_output_14_297(.a(output_15_297), .b(output_15_10), .y(output_14_297));
wire output_16_297, output_16_10, output_15_297;
mixer gate_output_15_297(.a(output_16_297), .b(output_16_10), .y(output_15_297));
wire output_1_298, output_1_11, output_0_298;
mixer gate_output_0_298(.a(output_1_298), .b(output_1_11), .y(output_0_298));
wire output_2_298, output_2_11, output_1_298;
mixer gate_output_1_298(.a(output_2_298), .b(output_2_11), .y(output_1_298));
wire output_3_298, output_3_11, output_2_298;
mixer gate_output_2_298(.a(output_3_298), .b(output_3_11), .y(output_2_298));
wire output_4_298, output_4_11, output_3_298;
mixer gate_output_3_298(.a(output_4_298), .b(output_4_11), .y(output_3_298));
wire output_5_298, output_5_11, output_4_298;
mixer gate_output_4_298(.a(output_5_298), .b(output_5_11), .y(output_4_298));
wire output_6_298, output_6_11, output_5_298;
mixer gate_output_5_298(.a(output_6_298), .b(output_6_11), .y(output_5_298));
wire output_7_298, output_7_11, output_6_298;
mixer gate_output_6_298(.a(output_7_298), .b(output_7_11), .y(output_6_298));
wire output_8_298, output_8_11, output_7_298;
mixer gate_output_7_298(.a(output_8_298), .b(output_8_11), .y(output_7_298));
wire output_9_298, output_9_11, output_8_298;
mixer gate_output_8_298(.a(output_9_298), .b(output_9_11), .y(output_8_298));
wire output_10_298, output_10_11, output_9_298;
mixer gate_output_9_298(.a(output_10_298), .b(output_10_11), .y(output_9_298));
wire output_11_298, output_11_11, output_10_298;
mixer gate_output_10_298(.a(output_11_298), .b(output_11_11), .y(output_10_298));
wire output_12_298, output_12_11, output_11_298;
mixer gate_output_11_298(.a(output_12_298), .b(output_12_11), .y(output_11_298));
wire output_13_298, output_13_11, output_12_298;
mixer gate_output_12_298(.a(output_13_298), .b(output_13_11), .y(output_12_298));
wire output_14_298, output_14_11, output_13_298;
mixer gate_output_13_298(.a(output_14_298), .b(output_14_11), .y(output_13_298));
wire output_15_298, output_15_11, output_14_298;
mixer gate_output_14_298(.a(output_15_298), .b(output_15_11), .y(output_14_298));
wire output_16_298, output_16_11, output_15_298;
mixer gate_output_15_298(.a(output_16_298), .b(output_16_11), .y(output_15_298));
wire output_1_299, output_1_12, output_0_299;
mixer gate_output_0_299(.a(output_1_299), .b(output_1_12), .y(output_0_299));
wire output_2_299, output_2_12, output_1_299;
mixer gate_output_1_299(.a(output_2_299), .b(output_2_12), .y(output_1_299));
wire output_3_299, output_3_12, output_2_299;
mixer gate_output_2_299(.a(output_3_299), .b(output_3_12), .y(output_2_299));
wire output_4_299, output_4_12, output_3_299;
mixer gate_output_3_299(.a(output_4_299), .b(output_4_12), .y(output_3_299));
wire output_5_299, output_5_12, output_4_299;
mixer gate_output_4_299(.a(output_5_299), .b(output_5_12), .y(output_4_299));
wire output_6_299, output_6_12, output_5_299;
mixer gate_output_5_299(.a(output_6_299), .b(output_6_12), .y(output_5_299));
wire output_7_299, output_7_12, output_6_299;
mixer gate_output_6_299(.a(output_7_299), .b(output_7_12), .y(output_6_299));
wire output_8_299, output_8_12, output_7_299;
mixer gate_output_7_299(.a(output_8_299), .b(output_8_12), .y(output_7_299));
wire output_9_299, output_9_12, output_8_299;
mixer gate_output_8_299(.a(output_9_299), .b(output_9_12), .y(output_8_299));
wire output_10_299, output_10_12, output_9_299;
mixer gate_output_9_299(.a(output_10_299), .b(output_10_12), .y(output_9_299));
wire output_11_299, output_11_12, output_10_299;
mixer gate_output_10_299(.a(output_11_299), .b(output_11_12), .y(output_10_299));
wire output_12_299, output_12_12, output_11_299;
mixer gate_output_11_299(.a(output_12_299), .b(output_12_12), .y(output_11_299));
wire output_13_299, output_13_12, output_12_299;
mixer gate_output_12_299(.a(output_13_299), .b(output_13_12), .y(output_12_299));
wire output_14_299, output_14_12, output_13_299;
mixer gate_output_13_299(.a(output_14_299), .b(output_14_12), .y(output_13_299));
wire output_15_299, output_15_12, output_14_299;
mixer gate_output_14_299(.a(output_15_299), .b(output_15_12), .y(output_14_299));
wire output_16_299, output_16_12, output_15_299;
mixer gate_output_15_299(.a(output_16_299), .b(output_16_12), .y(output_15_299));
wire output_1_300, output_1_13, output_0_300;
mixer gate_output_0_300(.a(output_1_300), .b(output_1_13), .y(output_0_300));
wire output_2_300, output_2_13, output_1_300;
mixer gate_output_1_300(.a(output_2_300), .b(output_2_13), .y(output_1_300));
wire output_3_300, output_3_13, output_2_300;
mixer gate_output_2_300(.a(output_3_300), .b(output_3_13), .y(output_2_300));
wire output_4_300, output_4_13, output_3_300;
mixer gate_output_3_300(.a(output_4_300), .b(output_4_13), .y(output_3_300));
wire output_5_300, output_5_13, output_4_300;
mixer gate_output_4_300(.a(output_5_300), .b(output_5_13), .y(output_4_300));
wire output_6_300, output_6_13, output_5_300;
mixer gate_output_5_300(.a(output_6_300), .b(output_6_13), .y(output_5_300));
wire output_7_300, output_7_13, output_6_300;
mixer gate_output_6_300(.a(output_7_300), .b(output_7_13), .y(output_6_300));
wire output_8_300, output_8_13, output_7_300;
mixer gate_output_7_300(.a(output_8_300), .b(output_8_13), .y(output_7_300));
wire output_9_300, output_9_13, output_8_300;
mixer gate_output_8_300(.a(output_9_300), .b(output_9_13), .y(output_8_300));
wire output_10_300, output_10_13, output_9_300;
mixer gate_output_9_300(.a(output_10_300), .b(output_10_13), .y(output_9_300));
wire output_11_300, output_11_13, output_10_300;
mixer gate_output_10_300(.a(output_11_300), .b(output_11_13), .y(output_10_300));
wire output_12_300, output_12_13, output_11_300;
mixer gate_output_11_300(.a(output_12_300), .b(output_12_13), .y(output_11_300));
wire output_13_300, output_13_13, output_12_300;
mixer gate_output_12_300(.a(output_13_300), .b(output_13_13), .y(output_12_300));
wire output_14_300, output_14_13, output_13_300;
mixer gate_output_13_300(.a(output_14_300), .b(output_14_13), .y(output_13_300));
wire output_15_300, output_15_13, output_14_300;
mixer gate_output_14_300(.a(output_15_300), .b(output_15_13), .y(output_14_300));
wire output_16_300, output_16_13, output_15_300;
mixer gate_output_15_300(.a(output_16_300), .b(output_16_13), .y(output_15_300));
wire output_1_301, output_1_14, output_0_301;
mixer gate_output_0_301(.a(output_1_301), .b(output_1_14), .y(output_0_301));
wire output_2_301, output_2_14, output_1_301;
mixer gate_output_1_301(.a(output_2_301), .b(output_2_14), .y(output_1_301));
wire output_3_301, output_3_14, output_2_301;
mixer gate_output_2_301(.a(output_3_301), .b(output_3_14), .y(output_2_301));
wire output_4_301, output_4_14, output_3_301;
mixer gate_output_3_301(.a(output_4_301), .b(output_4_14), .y(output_3_301));
wire output_5_301, output_5_14, output_4_301;
mixer gate_output_4_301(.a(output_5_301), .b(output_5_14), .y(output_4_301));
wire output_6_301, output_6_14, output_5_301;
mixer gate_output_5_301(.a(output_6_301), .b(output_6_14), .y(output_5_301));
wire output_7_301, output_7_14, output_6_301;
mixer gate_output_6_301(.a(output_7_301), .b(output_7_14), .y(output_6_301));
wire output_8_301, output_8_14, output_7_301;
mixer gate_output_7_301(.a(output_8_301), .b(output_8_14), .y(output_7_301));
wire output_9_301, output_9_14, output_8_301;
mixer gate_output_8_301(.a(output_9_301), .b(output_9_14), .y(output_8_301));
wire output_10_301, output_10_14, output_9_301;
mixer gate_output_9_301(.a(output_10_301), .b(output_10_14), .y(output_9_301));
wire output_11_301, output_11_14, output_10_301;
mixer gate_output_10_301(.a(output_11_301), .b(output_11_14), .y(output_10_301));
wire output_12_301, output_12_14, output_11_301;
mixer gate_output_11_301(.a(output_12_301), .b(output_12_14), .y(output_11_301));
wire output_13_301, output_13_14, output_12_301;
mixer gate_output_12_301(.a(output_13_301), .b(output_13_14), .y(output_12_301));
wire output_14_301, output_14_14, output_13_301;
mixer gate_output_13_301(.a(output_14_301), .b(output_14_14), .y(output_13_301));
wire output_15_301, output_15_14, output_14_301;
mixer gate_output_14_301(.a(output_15_301), .b(output_15_14), .y(output_14_301));
wire output_16_301, output_16_14, output_15_301;
mixer gate_output_15_301(.a(output_16_301), .b(output_16_14), .y(output_15_301));
wire output_1_302, output_1_15, output_0_302;
mixer gate_output_0_302(.a(output_1_302), .b(output_1_15), .y(output_0_302));
wire output_2_302, output_2_15, output_1_302;
mixer gate_output_1_302(.a(output_2_302), .b(output_2_15), .y(output_1_302));
wire output_3_302, output_3_15, output_2_302;
mixer gate_output_2_302(.a(output_3_302), .b(output_3_15), .y(output_2_302));
wire output_4_302, output_4_15, output_3_302;
mixer gate_output_3_302(.a(output_4_302), .b(output_4_15), .y(output_3_302));
wire output_5_302, output_5_15, output_4_302;
mixer gate_output_4_302(.a(output_5_302), .b(output_5_15), .y(output_4_302));
wire output_6_302, output_6_15, output_5_302;
mixer gate_output_5_302(.a(output_6_302), .b(output_6_15), .y(output_5_302));
wire output_7_302, output_7_15, output_6_302;
mixer gate_output_6_302(.a(output_7_302), .b(output_7_15), .y(output_6_302));
wire output_8_302, output_8_15, output_7_302;
mixer gate_output_7_302(.a(output_8_302), .b(output_8_15), .y(output_7_302));
wire output_9_302, output_9_15, output_8_302;
mixer gate_output_8_302(.a(output_9_302), .b(output_9_15), .y(output_8_302));
wire output_10_302, output_10_15, output_9_302;
mixer gate_output_9_302(.a(output_10_302), .b(output_10_15), .y(output_9_302));
wire output_11_302, output_11_15, output_10_302;
mixer gate_output_10_302(.a(output_11_302), .b(output_11_15), .y(output_10_302));
wire output_12_302, output_12_15, output_11_302;
mixer gate_output_11_302(.a(output_12_302), .b(output_12_15), .y(output_11_302));
wire output_13_302, output_13_15, output_12_302;
mixer gate_output_12_302(.a(output_13_302), .b(output_13_15), .y(output_12_302));
wire output_14_302, output_14_15, output_13_302;
mixer gate_output_13_302(.a(output_14_302), .b(output_14_15), .y(output_13_302));
wire output_15_302, output_15_15, output_14_302;
mixer gate_output_14_302(.a(output_15_302), .b(output_15_15), .y(output_14_302));
wire output_16_302, output_16_15, output_15_302;
mixer gate_output_15_302(.a(output_16_302), .b(output_16_15), .y(output_15_302));
wire output_1_303, output_1_0, output_0_303;
mixer gate_output_0_303(.a(output_1_303), .b(output_1_0), .y(output_0_303));
wire output_2_303, output_2_0, output_1_303;
mixer gate_output_1_303(.a(output_2_303), .b(output_2_0), .y(output_1_303));
wire output_3_303, output_3_0, output_2_303;
mixer gate_output_2_303(.a(output_3_303), .b(output_3_0), .y(output_2_303));
wire output_4_303, output_4_0, output_3_303;
mixer gate_output_3_303(.a(output_4_303), .b(output_4_0), .y(output_3_303));
wire output_5_303, output_5_0, output_4_303;
mixer gate_output_4_303(.a(output_5_303), .b(output_5_0), .y(output_4_303));
wire output_6_303, output_6_0, output_5_303;
mixer gate_output_5_303(.a(output_6_303), .b(output_6_0), .y(output_5_303));
wire output_7_303, output_7_0, output_6_303;
mixer gate_output_6_303(.a(output_7_303), .b(output_7_0), .y(output_6_303));
wire output_8_303, output_8_0, output_7_303;
mixer gate_output_7_303(.a(output_8_303), .b(output_8_0), .y(output_7_303));
wire output_9_303, output_9_0, output_8_303;
mixer gate_output_8_303(.a(output_9_303), .b(output_9_0), .y(output_8_303));
wire output_10_303, output_10_0, output_9_303;
mixer gate_output_9_303(.a(output_10_303), .b(output_10_0), .y(output_9_303));
wire output_11_303, output_11_0, output_10_303;
mixer gate_output_10_303(.a(output_11_303), .b(output_11_0), .y(output_10_303));
wire output_12_303, output_12_0, output_11_303;
mixer gate_output_11_303(.a(output_12_303), .b(output_12_0), .y(output_11_303));
wire output_13_303, output_13_0, output_12_303;
mixer gate_output_12_303(.a(output_13_303), .b(output_13_0), .y(output_12_303));
wire output_14_303, output_14_0, output_13_303;
mixer gate_output_13_303(.a(output_14_303), .b(output_14_0), .y(output_13_303));
wire output_15_303, output_15_0, output_14_303;
mixer gate_output_14_303(.a(output_15_303), .b(output_15_0), .y(output_14_303));
wire output_16_303, output_16_0, output_15_303;
mixer gate_output_15_303(.a(output_16_303), .b(output_16_0), .y(output_15_303));
wire output_1_304, output_1_1, output_0_304;
mixer gate_output_0_304(.a(output_1_304), .b(output_1_1), .y(output_0_304));
wire output_2_304, output_2_1, output_1_304;
mixer gate_output_1_304(.a(output_2_304), .b(output_2_1), .y(output_1_304));
wire output_3_304, output_3_1, output_2_304;
mixer gate_output_2_304(.a(output_3_304), .b(output_3_1), .y(output_2_304));
wire output_4_304, output_4_1, output_3_304;
mixer gate_output_3_304(.a(output_4_304), .b(output_4_1), .y(output_3_304));
wire output_5_304, output_5_1, output_4_304;
mixer gate_output_4_304(.a(output_5_304), .b(output_5_1), .y(output_4_304));
wire output_6_304, output_6_1, output_5_304;
mixer gate_output_5_304(.a(output_6_304), .b(output_6_1), .y(output_5_304));
wire output_7_304, output_7_1, output_6_304;
mixer gate_output_6_304(.a(output_7_304), .b(output_7_1), .y(output_6_304));
wire output_8_304, output_8_1, output_7_304;
mixer gate_output_7_304(.a(output_8_304), .b(output_8_1), .y(output_7_304));
wire output_9_304, output_9_1, output_8_304;
mixer gate_output_8_304(.a(output_9_304), .b(output_9_1), .y(output_8_304));
wire output_10_304, output_10_1, output_9_304;
mixer gate_output_9_304(.a(output_10_304), .b(output_10_1), .y(output_9_304));
wire output_11_304, output_11_1, output_10_304;
mixer gate_output_10_304(.a(output_11_304), .b(output_11_1), .y(output_10_304));
wire output_12_304, output_12_1, output_11_304;
mixer gate_output_11_304(.a(output_12_304), .b(output_12_1), .y(output_11_304));
wire output_13_304, output_13_1, output_12_304;
mixer gate_output_12_304(.a(output_13_304), .b(output_13_1), .y(output_12_304));
wire output_14_304, output_14_1, output_13_304;
mixer gate_output_13_304(.a(output_14_304), .b(output_14_1), .y(output_13_304));
wire output_15_304, output_15_1, output_14_304;
mixer gate_output_14_304(.a(output_15_304), .b(output_15_1), .y(output_14_304));
wire output_16_304, output_16_1, output_15_304;
mixer gate_output_15_304(.a(output_16_304), .b(output_16_1), .y(output_15_304));
wire output_1_305, output_1_2, output_0_305;
mixer gate_output_0_305(.a(output_1_305), .b(output_1_2), .y(output_0_305));
wire output_2_305, output_2_2, output_1_305;
mixer gate_output_1_305(.a(output_2_305), .b(output_2_2), .y(output_1_305));
wire output_3_305, output_3_2, output_2_305;
mixer gate_output_2_305(.a(output_3_305), .b(output_3_2), .y(output_2_305));
wire output_4_305, output_4_2, output_3_305;
mixer gate_output_3_305(.a(output_4_305), .b(output_4_2), .y(output_3_305));
wire output_5_305, output_5_2, output_4_305;
mixer gate_output_4_305(.a(output_5_305), .b(output_5_2), .y(output_4_305));
wire output_6_305, output_6_2, output_5_305;
mixer gate_output_5_305(.a(output_6_305), .b(output_6_2), .y(output_5_305));
wire output_7_305, output_7_2, output_6_305;
mixer gate_output_6_305(.a(output_7_305), .b(output_7_2), .y(output_6_305));
wire output_8_305, output_8_2, output_7_305;
mixer gate_output_7_305(.a(output_8_305), .b(output_8_2), .y(output_7_305));
wire output_9_305, output_9_2, output_8_305;
mixer gate_output_8_305(.a(output_9_305), .b(output_9_2), .y(output_8_305));
wire output_10_305, output_10_2, output_9_305;
mixer gate_output_9_305(.a(output_10_305), .b(output_10_2), .y(output_9_305));
wire output_11_305, output_11_2, output_10_305;
mixer gate_output_10_305(.a(output_11_305), .b(output_11_2), .y(output_10_305));
wire output_12_305, output_12_2, output_11_305;
mixer gate_output_11_305(.a(output_12_305), .b(output_12_2), .y(output_11_305));
wire output_13_305, output_13_2, output_12_305;
mixer gate_output_12_305(.a(output_13_305), .b(output_13_2), .y(output_12_305));
wire output_14_305, output_14_2, output_13_305;
mixer gate_output_13_305(.a(output_14_305), .b(output_14_2), .y(output_13_305));
wire output_15_305, output_15_2, output_14_305;
mixer gate_output_14_305(.a(output_15_305), .b(output_15_2), .y(output_14_305));
wire output_16_305, output_16_2, output_15_305;
mixer gate_output_15_305(.a(output_16_305), .b(output_16_2), .y(output_15_305));
wire output_1_306, output_1_3, output_0_306;
mixer gate_output_0_306(.a(output_1_306), .b(output_1_3), .y(output_0_306));
wire output_2_306, output_2_3, output_1_306;
mixer gate_output_1_306(.a(output_2_306), .b(output_2_3), .y(output_1_306));
wire output_3_306, output_3_3, output_2_306;
mixer gate_output_2_306(.a(output_3_306), .b(output_3_3), .y(output_2_306));
wire output_4_306, output_4_3, output_3_306;
mixer gate_output_3_306(.a(output_4_306), .b(output_4_3), .y(output_3_306));
wire output_5_306, output_5_3, output_4_306;
mixer gate_output_4_306(.a(output_5_306), .b(output_5_3), .y(output_4_306));
wire output_6_306, output_6_3, output_5_306;
mixer gate_output_5_306(.a(output_6_306), .b(output_6_3), .y(output_5_306));
wire output_7_306, output_7_3, output_6_306;
mixer gate_output_6_306(.a(output_7_306), .b(output_7_3), .y(output_6_306));
wire output_8_306, output_8_3, output_7_306;
mixer gate_output_7_306(.a(output_8_306), .b(output_8_3), .y(output_7_306));
wire output_9_306, output_9_3, output_8_306;
mixer gate_output_8_306(.a(output_9_306), .b(output_9_3), .y(output_8_306));
wire output_10_306, output_10_3, output_9_306;
mixer gate_output_9_306(.a(output_10_306), .b(output_10_3), .y(output_9_306));
wire output_11_306, output_11_3, output_10_306;
mixer gate_output_10_306(.a(output_11_306), .b(output_11_3), .y(output_10_306));
wire output_12_306, output_12_3, output_11_306;
mixer gate_output_11_306(.a(output_12_306), .b(output_12_3), .y(output_11_306));
wire output_13_306, output_13_3, output_12_306;
mixer gate_output_12_306(.a(output_13_306), .b(output_13_3), .y(output_12_306));
wire output_14_306, output_14_3, output_13_306;
mixer gate_output_13_306(.a(output_14_306), .b(output_14_3), .y(output_13_306));
wire output_15_306, output_15_3, output_14_306;
mixer gate_output_14_306(.a(output_15_306), .b(output_15_3), .y(output_14_306));
wire output_16_306, output_16_3, output_15_306;
mixer gate_output_15_306(.a(output_16_306), .b(output_16_3), .y(output_15_306));
wire output_1_307, output_1_4, output_0_307;
mixer gate_output_0_307(.a(output_1_307), .b(output_1_4), .y(output_0_307));
wire output_2_307, output_2_4, output_1_307;
mixer gate_output_1_307(.a(output_2_307), .b(output_2_4), .y(output_1_307));
wire output_3_307, output_3_4, output_2_307;
mixer gate_output_2_307(.a(output_3_307), .b(output_3_4), .y(output_2_307));
wire output_4_307, output_4_4, output_3_307;
mixer gate_output_3_307(.a(output_4_307), .b(output_4_4), .y(output_3_307));
wire output_5_307, output_5_4, output_4_307;
mixer gate_output_4_307(.a(output_5_307), .b(output_5_4), .y(output_4_307));
wire output_6_307, output_6_4, output_5_307;
mixer gate_output_5_307(.a(output_6_307), .b(output_6_4), .y(output_5_307));
wire output_7_307, output_7_4, output_6_307;
mixer gate_output_6_307(.a(output_7_307), .b(output_7_4), .y(output_6_307));
wire output_8_307, output_8_4, output_7_307;
mixer gate_output_7_307(.a(output_8_307), .b(output_8_4), .y(output_7_307));
wire output_9_307, output_9_4, output_8_307;
mixer gate_output_8_307(.a(output_9_307), .b(output_9_4), .y(output_8_307));
wire output_10_307, output_10_4, output_9_307;
mixer gate_output_9_307(.a(output_10_307), .b(output_10_4), .y(output_9_307));
wire output_11_307, output_11_4, output_10_307;
mixer gate_output_10_307(.a(output_11_307), .b(output_11_4), .y(output_10_307));
wire output_12_307, output_12_4, output_11_307;
mixer gate_output_11_307(.a(output_12_307), .b(output_12_4), .y(output_11_307));
wire output_13_307, output_13_4, output_12_307;
mixer gate_output_12_307(.a(output_13_307), .b(output_13_4), .y(output_12_307));
wire output_14_307, output_14_4, output_13_307;
mixer gate_output_13_307(.a(output_14_307), .b(output_14_4), .y(output_13_307));
wire output_15_307, output_15_4, output_14_307;
mixer gate_output_14_307(.a(output_15_307), .b(output_15_4), .y(output_14_307));
wire output_16_307, output_16_4, output_15_307;
mixer gate_output_15_307(.a(output_16_307), .b(output_16_4), .y(output_15_307));
wire output_1_308, output_1_5, output_0_308;
mixer gate_output_0_308(.a(output_1_308), .b(output_1_5), .y(output_0_308));
wire output_2_308, output_2_5, output_1_308;
mixer gate_output_1_308(.a(output_2_308), .b(output_2_5), .y(output_1_308));
wire output_3_308, output_3_5, output_2_308;
mixer gate_output_2_308(.a(output_3_308), .b(output_3_5), .y(output_2_308));
wire output_4_308, output_4_5, output_3_308;
mixer gate_output_3_308(.a(output_4_308), .b(output_4_5), .y(output_3_308));
wire output_5_308, output_5_5, output_4_308;
mixer gate_output_4_308(.a(output_5_308), .b(output_5_5), .y(output_4_308));
wire output_6_308, output_6_5, output_5_308;
mixer gate_output_5_308(.a(output_6_308), .b(output_6_5), .y(output_5_308));
wire output_7_308, output_7_5, output_6_308;
mixer gate_output_6_308(.a(output_7_308), .b(output_7_5), .y(output_6_308));
wire output_8_308, output_8_5, output_7_308;
mixer gate_output_7_308(.a(output_8_308), .b(output_8_5), .y(output_7_308));
wire output_9_308, output_9_5, output_8_308;
mixer gate_output_8_308(.a(output_9_308), .b(output_9_5), .y(output_8_308));
wire output_10_308, output_10_5, output_9_308;
mixer gate_output_9_308(.a(output_10_308), .b(output_10_5), .y(output_9_308));
wire output_11_308, output_11_5, output_10_308;
mixer gate_output_10_308(.a(output_11_308), .b(output_11_5), .y(output_10_308));
wire output_12_308, output_12_5, output_11_308;
mixer gate_output_11_308(.a(output_12_308), .b(output_12_5), .y(output_11_308));
wire output_13_308, output_13_5, output_12_308;
mixer gate_output_12_308(.a(output_13_308), .b(output_13_5), .y(output_12_308));
wire output_14_308, output_14_5, output_13_308;
mixer gate_output_13_308(.a(output_14_308), .b(output_14_5), .y(output_13_308));
wire output_15_308, output_15_5, output_14_308;
mixer gate_output_14_308(.a(output_15_308), .b(output_15_5), .y(output_14_308));
wire output_16_308, output_16_5, output_15_308;
mixer gate_output_15_308(.a(output_16_308), .b(output_16_5), .y(output_15_308));
wire output_1_309, output_1_6, output_0_309;
mixer gate_output_0_309(.a(output_1_309), .b(output_1_6), .y(output_0_309));
wire output_2_309, output_2_6, output_1_309;
mixer gate_output_1_309(.a(output_2_309), .b(output_2_6), .y(output_1_309));
wire output_3_309, output_3_6, output_2_309;
mixer gate_output_2_309(.a(output_3_309), .b(output_3_6), .y(output_2_309));
wire output_4_309, output_4_6, output_3_309;
mixer gate_output_3_309(.a(output_4_309), .b(output_4_6), .y(output_3_309));
wire output_5_309, output_5_6, output_4_309;
mixer gate_output_4_309(.a(output_5_309), .b(output_5_6), .y(output_4_309));
wire output_6_309, output_6_6, output_5_309;
mixer gate_output_5_309(.a(output_6_309), .b(output_6_6), .y(output_5_309));
wire output_7_309, output_7_6, output_6_309;
mixer gate_output_6_309(.a(output_7_309), .b(output_7_6), .y(output_6_309));
wire output_8_309, output_8_6, output_7_309;
mixer gate_output_7_309(.a(output_8_309), .b(output_8_6), .y(output_7_309));
wire output_9_309, output_9_6, output_8_309;
mixer gate_output_8_309(.a(output_9_309), .b(output_9_6), .y(output_8_309));
wire output_10_309, output_10_6, output_9_309;
mixer gate_output_9_309(.a(output_10_309), .b(output_10_6), .y(output_9_309));
wire output_11_309, output_11_6, output_10_309;
mixer gate_output_10_309(.a(output_11_309), .b(output_11_6), .y(output_10_309));
wire output_12_309, output_12_6, output_11_309;
mixer gate_output_11_309(.a(output_12_309), .b(output_12_6), .y(output_11_309));
wire output_13_309, output_13_6, output_12_309;
mixer gate_output_12_309(.a(output_13_309), .b(output_13_6), .y(output_12_309));
wire output_14_309, output_14_6, output_13_309;
mixer gate_output_13_309(.a(output_14_309), .b(output_14_6), .y(output_13_309));
wire output_15_309, output_15_6, output_14_309;
mixer gate_output_14_309(.a(output_15_309), .b(output_15_6), .y(output_14_309));
wire output_16_309, output_16_6, output_15_309;
mixer gate_output_15_309(.a(output_16_309), .b(output_16_6), .y(output_15_309));
wire output_1_310, output_1_7, output_0_310;
mixer gate_output_0_310(.a(output_1_310), .b(output_1_7), .y(output_0_310));
wire output_2_310, output_2_7, output_1_310;
mixer gate_output_1_310(.a(output_2_310), .b(output_2_7), .y(output_1_310));
wire output_3_310, output_3_7, output_2_310;
mixer gate_output_2_310(.a(output_3_310), .b(output_3_7), .y(output_2_310));
wire output_4_310, output_4_7, output_3_310;
mixer gate_output_3_310(.a(output_4_310), .b(output_4_7), .y(output_3_310));
wire output_5_310, output_5_7, output_4_310;
mixer gate_output_4_310(.a(output_5_310), .b(output_5_7), .y(output_4_310));
wire output_6_310, output_6_7, output_5_310;
mixer gate_output_5_310(.a(output_6_310), .b(output_6_7), .y(output_5_310));
wire output_7_310, output_7_7, output_6_310;
mixer gate_output_6_310(.a(output_7_310), .b(output_7_7), .y(output_6_310));
wire output_8_310, output_8_7, output_7_310;
mixer gate_output_7_310(.a(output_8_310), .b(output_8_7), .y(output_7_310));
wire output_9_310, output_9_7, output_8_310;
mixer gate_output_8_310(.a(output_9_310), .b(output_9_7), .y(output_8_310));
wire output_10_310, output_10_7, output_9_310;
mixer gate_output_9_310(.a(output_10_310), .b(output_10_7), .y(output_9_310));
wire output_11_310, output_11_7, output_10_310;
mixer gate_output_10_310(.a(output_11_310), .b(output_11_7), .y(output_10_310));
wire output_12_310, output_12_7, output_11_310;
mixer gate_output_11_310(.a(output_12_310), .b(output_12_7), .y(output_11_310));
wire output_13_310, output_13_7, output_12_310;
mixer gate_output_12_310(.a(output_13_310), .b(output_13_7), .y(output_12_310));
wire output_14_310, output_14_7, output_13_310;
mixer gate_output_13_310(.a(output_14_310), .b(output_14_7), .y(output_13_310));
wire output_15_310, output_15_7, output_14_310;
mixer gate_output_14_310(.a(output_15_310), .b(output_15_7), .y(output_14_310));
wire output_16_310, output_16_7, output_15_310;
mixer gate_output_15_310(.a(output_16_310), .b(output_16_7), .y(output_15_310));
wire output_1_311, output_1_8, output_0_311;
mixer gate_output_0_311(.a(output_1_311), .b(output_1_8), .y(output_0_311));
wire output_2_311, output_2_8, output_1_311;
mixer gate_output_1_311(.a(output_2_311), .b(output_2_8), .y(output_1_311));
wire output_3_311, output_3_8, output_2_311;
mixer gate_output_2_311(.a(output_3_311), .b(output_3_8), .y(output_2_311));
wire output_4_311, output_4_8, output_3_311;
mixer gate_output_3_311(.a(output_4_311), .b(output_4_8), .y(output_3_311));
wire output_5_311, output_5_8, output_4_311;
mixer gate_output_4_311(.a(output_5_311), .b(output_5_8), .y(output_4_311));
wire output_6_311, output_6_8, output_5_311;
mixer gate_output_5_311(.a(output_6_311), .b(output_6_8), .y(output_5_311));
wire output_7_311, output_7_8, output_6_311;
mixer gate_output_6_311(.a(output_7_311), .b(output_7_8), .y(output_6_311));
wire output_8_311, output_8_8, output_7_311;
mixer gate_output_7_311(.a(output_8_311), .b(output_8_8), .y(output_7_311));
wire output_9_311, output_9_8, output_8_311;
mixer gate_output_8_311(.a(output_9_311), .b(output_9_8), .y(output_8_311));
wire output_10_311, output_10_8, output_9_311;
mixer gate_output_9_311(.a(output_10_311), .b(output_10_8), .y(output_9_311));
wire output_11_311, output_11_8, output_10_311;
mixer gate_output_10_311(.a(output_11_311), .b(output_11_8), .y(output_10_311));
wire output_12_311, output_12_8, output_11_311;
mixer gate_output_11_311(.a(output_12_311), .b(output_12_8), .y(output_11_311));
wire output_13_311, output_13_8, output_12_311;
mixer gate_output_12_311(.a(output_13_311), .b(output_13_8), .y(output_12_311));
wire output_14_311, output_14_8, output_13_311;
mixer gate_output_13_311(.a(output_14_311), .b(output_14_8), .y(output_13_311));
wire output_15_311, output_15_8, output_14_311;
mixer gate_output_14_311(.a(output_15_311), .b(output_15_8), .y(output_14_311));
wire output_16_311, output_16_8, output_15_311;
mixer gate_output_15_311(.a(output_16_311), .b(output_16_8), .y(output_15_311));
wire output_1_312, output_1_9, output_0_312;
mixer gate_output_0_312(.a(output_1_312), .b(output_1_9), .y(output_0_312));
wire output_2_312, output_2_9, output_1_312;
mixer gate_output_1_312(.a(output_2_312), .b(output_2_9), .y(output_1_312));
wire output_3_312, output_3_9, output_2_312;
mixer gate_output_2_312(.a(output_3_312), .b(output_3_9), .y(output_2_312));
wire output_4_312, output_4_9, output_3_312;
mixer gate_output_3_312(.a(output_4_312), .b(output_4_9), .y(output_3_312));
wire output_5_312, output_5_9, output_4_312;
mixer gate_output_4_312(.a(output_5_312), .b(output_5_9), .y(output_4_312));
wire output_6_312, output_6_9, output_5_312;
mixer gate_output_5_312(.a(output_6_312), .b(output_6_9), .y(output_5_312));
wire output_7_312, output_7_9, output_6_312;
mixer gate_output_6_312(.a(output_7_312), .b(output_7_9), .y(output_6_312));
wire output_8_312, output_8_9, output_7_312;
mixer gate_output_7_312(.a(output_8_312), .b(output_8_9), .y(output_7_312));
wire output_9_312, output_9_9, output_8_312;
mixer gate_output_8_312(.a(output_9_312), .b(output_9_9), .y(output_8_312));
wire output_10_312, output_10_9, output_9_312;
mixer gate_output_9_312(.a(output_10_312), .b(output_10_9), .y(output_9_312));
wire output_11_312, output_11_9, output_10_312;
mixer gate_output_10_312(.a(output_11_312), .b(output_11_9), .y(output_10_312));
wire output_12_312, output_12_9, output_11_312;
mixer gate_output_11_312(.a(output_12_312), .b(output_12_9), .y(output_11_312));
wire output_13_312, output_13_9, output_12_312;
mixer gate_output_12_312(.a(output_13_312), .b(output_13_9), .y(output_12_312));
wire output_14_312, output_14_9, output_13_312;
mixer gate_output_13_312(.a(output_14_312), .b(output_14_9), .y(output_13_312));
wire output_15_312, output_15_9, output_14_312;
mixer gate_output_14_312(.a(output_15_312), .b(output_15_9), .y(output_14_312));
wire output_16_312, output_16_9, output_15_312;
mixer gate_output_15_312(.a(output_16_312), .b(output_16_9), .y(output_15_312));
wire output_1_313, output_1_10, output_0_313;
mixer gate_output_0_313(.a(output_1_313), .b(output_1_10), .y(output_0_313));
wire output_2_313, output_2_10, output_1_313;
mixer gate_output_1_313(.a(output_2_313), .b(output_2_10), .y(output_1_313));
wire output_3_313, output_3_10, output_2_313;
mixer gate_output_2_313(.a(output_3_313), .b(output_3_10), .y(output_2_313));
wire output_4_313, output_4_10, output_3_313;
mixer gate_output_3_313(.a(output_4_313), .b(output_4_10), .y(output_3_313));
wire output_5_313, output_5_10, output_4_313;
mixer gate_output_4_313(.a(output_5_313), .b(output_5_10), .y(output_4_313));
wire output_6_313, output_6_10, output_5_313;
mixer gate_output_5_313(.a(output_6_313), .b(output_6_10), .y(output_5_313));
wire output_7_313, output_7_10, output_6_313;
mixer gate_output_6_313(.a(output_7_313), .b(output_7_10), .y(output_6_313));
wire output_8_313, output_8_10, output_7_313;
mixer gate_output_7_313(.a(output_8_313), .b(output_8_10), .y(output_7_313));
wire output_9_313, output_9_10, output_8_313;
mixer gate_output_8_313(.a(output_9_313), .b(output_9_10), .y(output_8_313));
wire output_10_313, output_10_10, output_9_313;
mixer gate_output_9_313(.a(output_10_313), .b(output_10_10), .y(output_9_313));
wire output_11_313, output_11_10, output_10_313;
mixer gate_output_10_313(.a(output_11_313), .b(output_11_10), .y(output_10_313));
wire output_12_313, output_12_10, output_11_313;
mixer gate_output_11_313(.a(output_12_313), .b(output_12_10), .y(output_11_313));
wire output_13_313, output_13_10, output_12_313;
mixer gate_output_12_313(.a(output_13_313), .b(output_13_10), .y(output_12_313));
wire output_14_313, output_14_10, output_13_313;
mixer gate_output_13_313(.a(output_14_313), .b(output_14_10), .y(output_13_313));
wire output_15_313, output_15_10, output_14_313;
mixer gate_output_14_313(.a(output_15_313), .b(output_15_10), .y(output_14_313));
wire output_16_313, output_16_10, output_15_313;
mixer gate_output_15_313(.a(output_16_313), .b(output_16_10), .y(output_15_313));
wire output_1_314, output_1_11, output_0_314;
mixer gate_output_0_314(.a(output_1_314), .b(output_1_11), .y(output_0_314));
wire output_2_314, output_2_11, output_1_314;
mixer gate_output_1_314(.a(output_2_314), .b(output_2_11), .y(output_1_314));
wire output_3_314, output_3_11, output_2_314;
mixer gate_output_2_314(.a(output_3_314), .b(output_3_11), .y(output_2_314));
wire output_4_314, output_4_11, output_3_314;
mixer gate_output_3_314(.a(output_4_314), .b(output_4_11), .y(output_3_314));
wire output_5_314, output_5_11, output_4_314;
mixer gate_output_4_314(.a(output_5_314), .b(output_5_11), .y(output_4_314));
wire output_6_314, output_6_11, output_5_314;
mixer gate_output_5_314(.a(output_6_314), .b(output_6_11), .y(output_5_314));
wire output_7_314, output_7_11, output_6_314;
mixer gate_output_6_314(.a(output_7_314), .b(output_7_11), .y(output_6_314));
wire output_8_314, output_8_11, output_7_314;
mixer gate_output_7_314(.a(output_8_314), .b(output_8_11), .y(output_7_314));
wire output_9_314, output_9_11, output_8_314;
mixer gate_output_8_314(.a(output_9_314), .b(output_9_11), .y(output_8_314));
wire output_10_314, output_10_11, output_9_314;
mixer gate_output_9_314(.a(output_10_314), .b(output_10_11), .y(output_9_314));
wire output_11_314, output_11_11, output_10_314;
mixer gate_output_10_314(.a(output_11_314), .b(output_11_11), .y(output_10_314));
wire output_12_314, output_12_11, output_11_314;
mixer gate_output_11_314(.a(output_12_314), .b(output_12_11), .y(output_11_314));
wire output_13_314, output_13_11, output_12_314;
mixer gate_output_12_314(.a(output_13_314), .b(output_13_11), .y(output_12_314));
wire output_14_314, output_14_11, output_13_314;
mixer gate_output_13_314(.a(output_14_314), .b(output_14_11), .y(output_13_314));
wire output_15_314, output_15_11, output_14_314;
mixer gate_output_14_314(.a(output_15_314), .b(output_15_11), .y(output_14_314));
wire output_16_314, output_16_11, output_15_314;
mixer gate_output_15_314(.a(output_16_314), .b(output_16_11), .y(output_15_314));
wire output_1_315, output_1_12, output_0_315;
mixer gate_output_0_315(.a(output_1_315), .b(output_1_12), .y(output_0_315));
wire output_2_315, output_2_12, output_1_315;
mixer gate_output_1_315(.a(output_2_315), .b(output_2_12), .y(output_1_315));
wire output_3_315, output_3_12, output_2_315;
mixer gate_output_2_315(.a(output_3_315), .b(output_3_12), .y(output_2_315));
wire output_4_315, output_4_12, output_3_315;
mixer gate_output_3_315(.a(output_4_315), .b(output_4_12), .y(output_3_315));
wire output_5_315, output_5_12, output_4_315;
mixer gate_output_4_315(.a(output_5_315), .b(output_5_12), .y(output_4_315));
wire output_6_315, output_6_12, output_5_315;
mixer gate_output_5_315(.a(output_6_315), .b(output_6_12), .y(output_5_315));
wire output_7_315, output_7_12, output_6_315;
mixer gate_output_6_315(.a(output_7_315), .b(output_7_12), .y(output_6_315));
wire output_8_315, output_8_12, output_7_315;
mixer gate_output_7_315(.a(output_8_315), .b(output_8_12), .y(output_7_315));
wire output_9_315, output_9_12, output_8_315;
mixer gate_output_8_315(.a(output_9_315), .b(output_9_12), .y(output_8_315));
wire output_10_315, output_10_12, output_9_315;
mixer gate_output_9_315(.a(output_10_315), .b(output_10_12), .y(output_9_315));
wire output_11_315, output_11_12, output_10_315;
mixer gate_output_10_315(.a(output_11_315), .b(output_11_12), .y(output_10_315));
wire output_12_315, output_12_12, output_11_315;
mixer gate_output_11_315(.a(output_12_315), .b(output_12_12), .y(output_11_315));
wire output_13_315, output_13_12, output_12_315;
mixer gate_output_12_315(.a(output_13_315), .b(output_13_12), .y(output_12_315));
wire output_14_315, output_14_12, output_13_315;
mixer gate_output_13_315(.a(output_14_315), .b(output_14_12), .y(output_13_315));
wire output_15_315, output_15_12, output_14_315;
mixer gate_output_14_315(.a(output_15_315), .b(output_15_12), .y(output_14_315));
wire output_16_315, output_16_12, output_15_315;
mixer gate_output_15_315(.a(output_16_315), .b(output_16_12), .y(output_15_315));
wire output_1_316, output_1_13, output_0_316;
mixer gate_output_0_316(.a(output_1_316), .b(output_1_13), .y(output_0_316));
wire output_2_316, output_2_13, output_1_316;
mixer gate_output_1_316(.a(output_2_316), .b(output_2_13), .y(output_1_316));
wire output_3_316, output_3_13, output_2_316;
mixer gate_output_2_316(.a(output_3_316), .b(output_3_13), .y(output_2_316));
wire output_4_316, output_4_13, output_3_316;
mixer gate_output_3_316(.a(output_4_316), .b(output_4_13), .y(output_3_316));
wire output_5_316, output_5_13, output_4_316;
mixer gate_output_4_316(.a(output_5_316), .b(output_5_13), .y(output_4_316));
wire output_6_316, output_6_13, output_5_316;
mixer gate_output_5_316(.a(output_6_316), .b(output_6_13), .y(output_5_316));
wire output_7_316, output_7_13, output_6_316;
mixer gate_output_6_316(.a(output_7_316), .b(output_7_13), .y(output_6_316));
wire output_8_316, output_8_13, output_7_316;
mixer gate_output_7_316(.a(output_8_316), .b(output_8_13), .y(output_7_316));
wire output_9_316, output_9_13, output_8_316;
mixer gate_output_8_316(.a(output_9_316), .b(output_9_13), .y(output_8_316));
wire output_10_316, output_10_13, output_9_316;
mixer gate_output_9_316(.a(output_10_316), .b(output_10_13), .y(output_9_316));
wire output_11_316, output_11_13, output_10_316;
mixer gate_output_10_316(.a(output_11_316), .b(output_11_13), .y(output_10_316));
wire output_12_316, output_12_13, output_11_316;
mixer gate_output_11_316(.a(output_12_316), .b(output_12_13), .y(output_11_316));
wire output_13_316, output_13_13, output_12_316;
mixer gate_output_12_316(.a(output_13_316), .b(output_13_13), .y(output_12_316));
wire output_14_316, output_14_13, output_13_316;
mixer gate_output_13_316(.a(output_14_316), .b(output_14_13), .y(output_13_316));
wire output_15_316, output_15_13, output_14_316;
mixer gate_output_14_316(.a(output_15_316), .b(output_15_13), .y(output_14_316));
wire output_16_316, output_16_13, output_15_316;
mixer gate_output_15_316(.a(output_16_316), .b(output_16_13), .y(output_15_316));
wire output_1_317, output_1_14, output_0_317;
mixer gate_output_0_317(.a(output_1_317), .b(output_1_14), .y(output_0_317));
wire output_2_317, output_2_14, output_1_317;
mixer gate_output_1_317(.a(output_2_317), .b(output_2_14), .y(output_1_317));
wire output_3_317, output_3_14, output_2_317;
mixer gate_output_2_317(.a(output_3_317), .b(output_3_14), .y(output_2_317));
wire output_4_317, output_4_14, output_3_317;
mixer gate_output_3_317(.a(output_4_317), .b(output_4_14), .y(output_3_317));
wire output_5_317, output_5_14, output_4_317;
mixer gate_output_4_317(.a(output_5_317), .b(output_5_14), .y(output_4_317));
wire output_6_317, output_6_14, output_5_317;
mixer gate_output_5_317(.a(output_6_317), .b(output_6_14), .y(output_5_317));
wire output_7_317, output_7_14, output_6_317;
mixer gate_output_6_317(.a(output_7_317), .b(output_7_14), .y(output_6_317));
wire output_8_317, output_8_14, output_7_317;
mixer gate_output_7_317(.a(output_8_317), .b(output_8_14), .y(output_7_317));
wire output_9_317, output_9_14, output_8_317;
mixer gate_output_8_317(.a(output_9_317), .b(output_9_14), .y(output_8_317));
wire output_10_317, output_10_14, output_9_317;
mixer gate_output_9_317(.a(output_10_317), .b(output_10_14), .y(output_9_317));
wire output_11_317, output_11_14, output_10_317;
mixer gate_output_10_317(.a(output_11_317), .b(output_11_14), .y(output_10_317));
wire output_12_317, output_12_14, output_11_317;
mixer gate_output_11_317(.a(output_12_317), .b(output_12_14), .y(output_11_317));
wire output_13_317, output_13_14, output_12_317;
mixer gate_output_12_317(.a(output_13_317), .b(output_13_14), .y(output_12_317));
wire output_14_317, output_14_14, output_13_317;
mixer gate_output_13_317(.a(output_14_317), .b(output_14_14), .y(output_13_317));
wire output_15_317, output_15_14, output_14_317;
mixer gate_output_14_317(.a(output_15_317), .b(output_15_14), .y(output_14_317));
wire output_16_317, output_16_14, output_15_317;
mixer gate_output_15_317(.a(output_16_317), .b(output_16_14), .y(output_15_317));
wire output_1_318, output_1_15, output_0_318;
mixer gate_output_0_318(.a(output_1_318), .b(output_1_15), .y(output_0_318));
wire output_2_318, output_2_15, output_1_318;
mixer gate_output_1_318(.a(output_2_318), .b(output_2_15), .y(output_1_318));
wire output_3_318, output_3_15, output_2_318;
mixer gate_output_2_318(.a(output_3_318), .b(output_3_15), .y(output_2_318));
wire output_4_318, output_4_15, output_3_318;
mixer gate_output_3_318(.a(output_4_318), .b(output_4_15), .y(output_3_318));
wire output_5_318, output_5_15, output_4_318;
mixer gate_output_4_318(.a(output_5_318), .b(output_5_15), .y(output_4_318));
wire output_6_318, output_6_15, output_5_318;
mixer gate_output_5_318(.a(output_6_318), .b(output_6_15), .y(output_5_318));
wire output_7_318, output_7_15, output_6_318;
mixer gate_output_6_318(.a(output_7_318), .b(output_7_15), .y(output_6_318));
wire output_8_318, output_8_15, output_7_318;
mixer gate_output_7_318(.a(output_8_318), .b(output_8_15), .y(output_7_318));
wire output_9_318, output_9_15, output_8_318;
mixer gate_output_8_318(.a(output_9_318), .b(output_9_15), .y(output_8_318));
wire output_10_318, output_10_15, output_9_318;
mixer gate_output_9_318(.a(output_10_318), .b(output_10_15), .y(output_9_318));
wire output_11_318, output_11_15, output_10_318;
mixer gate_output_10_318(.a(output_11_318), .b(output_11_15), .y(output_10_318));
wire output_12_318, output_12_15, output_11_318;
mixer gate_output_11_318(.a(output_12_318), .b(output_12_15), .y(output_11_318));
wire output_13_318, output_13_15, output_12_318;
mixer gate_output_12_318(.a(output_13_318), .b(output_13_15), .y(output_12_318));
wire output_14_318, output_14_15, output_13_318;
mixer gate_output_13_318(.a(output_14_318), .b(output_14_15), .y(output_13_318));
wire output_15_318, output_15_15, output_14_318;
mixer gate_output_14_318(.a(output_15_318), .b(output_15_15), .y(output_14_318));
wire output_16_318, output_16_15, output_15_318;
mixer gate_output_15_318(.a(output_16_318), .b(output_16_15), .y(output_15_318));
wire output_1_319, output_1_0, output_0_319;
mixer gate_output_0_319(.a(output_1_319), .b(output_1_0), .y(output_0_319));
wire output_2_319, output_2_0, output_1_319;
mixer gate_output_1_319(.a(output_2_319), .b(output_2_0), .y(output_1_319));
wire output_3_319, output_3_0, output_2_319;
mixer gate_output_2_319(.a(output_3_319), .b(output_3_0), .y(output_2_319));
wire output_4_319, output_4_0, output_3_319;
mixer gate_output_3_319(.a(output_4_319), .b(output_4_0), .y(output_3_319));
wire output_5_319, output_5_0, output_4_319;
mixer gate_output_4_319(.a(output_5_319), .b(output_5_0), .y(output_4_319));
wire output_6_319, output_6_0, output_5_319;
mixer gate_output_5_319(.a(output_6_319), .b(output_6_0), .y(output_5_319));
wire output_7_319, output_7_0, output_6_319;
mixer gate_output_6_319(.a(output_7_319), .b(output_7_0), .y(output_6_319));
wire output_8_319, output_8_0, output_7_319;
mixer gate_output_7_319(.a(output_8_319), .b(output_8_0), .y(output_7_319));
wire output_9_319, output_9_0, output_8_319;
mixer gate_output_8_319(.a(output_9_319), .b(output_9_0), .y(output_8_319));
wire output_10_319, output_10_0, output_9_319;
mixer gate_output_9_319(.a(output_10_319), .b(output_10_0), .y(output_9_319));
wire output_11_319, output_11_0, output_10_319;
mixer gate_output_10_319(.a(output_11_319), .b(output_11_0), .y(output_10_319));
wire output_12_319, output_12_0, output_11_319;
mixer gate_output_11_319(.a(output_12_319), .b(output_12_0), .y(output_11_319));
wire output_13_319, output_13_0, output_12_319;
mixer gate_output_12_319(.a(output_13_319), .b(output_13_0), .y(output_12_319));
wire output_14_319, output_14_0, output_13_319;
mixer gate_output_13_319(.a(output_14_319), .b(output_14_0), .y(output_13_319));
wire output_15_319, output_15_0, output_14_319;
mixer gate_output_14_319(.a(output_15_319), .b(output_15_0), .y(output_14_319));
wire output_16_319, output_16_0, output_15_319;
mixer gate_output_15_319(.a(output_16_319), .b(output_16_0), .y(output_15_319));
wire output_1_320, output_1_1, output_0_320;
mixer gate_output_0_320(.a(output_1_320), .b(output_1_1), .y(output_0_320));
wire output_2_320, output_2_1, output_1_320;
mixer gate_output_1_320(.a(output_2_320), .b(output_2_1), .y(output_1_320));
wire output_3_320, output_3_1, output_2_320;
mixer gate_output_2_320(.a(output_3_320), .b(output_3_1), .y(output_2_320));
wire output_4_320, output_4_1, output_3_320;
mixer gate_output_3_320(.a(output_4_320), .b(output_4_1), .y(output_3_320));
wire output_5_320, output_5_1, output_4_320;
mixer gate_output_4_320(.a(output_5_320), .b(output_5_1), .y(output_4_320));
wire output_6_320, output_6_1, output_5_320;
mixer gate_output_5_320(.a(output_6_320), .b(output_6_1), .y(output_5_320));
wire output_7_320, output_7_1, output_6_320;
mixer gate_output_6_320(.a(output_7_320), .b(output_7_1), .y(output_6_320));
wire output_8_320, output_8_1, output_7_320;
mixer gate_output_7_320(.a(output_8_320), .b(output_8_1), .y(output_7_320));
wire output_9_320, output_9_1, output_8_320;
mixer gate_output_8_320(.a(output_9_320), .b(output_9_1), .y(output_8_320));
wire output_10_320, output_10_1, output_9_320;
mixer gate_output_9_320(.a(output_10_320), .b(output_10_1), .y(output_9_320));
wire output_11_320, output_11_1, output_10_320;
mixer gate_output_10_320(.a(output_11_320), .b(output_11_1), .y(output_10_320));
wire output_12_320, output_12_1, output_11_320;
mixer gate_output_11_320(.a(output_12_320), .b(output_12_1), .y(output_11_320));
wire output_13_320, output_13_1, output_12_320;
mixer gate_output_12_320(.a(output_13_320), .b(output_13_1), .y(output_12_320));
wire output_14_320, output_14_1, output_13_320;
mixer gate_output_13_320(.a(output_14_320), .b(output_14_1), .y(output_13_320));
wire output_15_320, output_15_1, output_14_320;
mixer gate_output_14_320(.a(output_15_320), .b(output_15_1), .y(output_14_320));
wire output_16_320, output_16_1, output_15_320;
mixer gate_output_15_320(.a(output_16_320), .b(output_16_1), .y(output_15_320));
wire output_1_321, output_1_2, output_0_321;
mixer gate_output_0_321(.a(output_1_321), .b(output_1_2), .y(output_0_321));
wire output_2_321, output_2_2, output_1_321;
mixer gate_output_1_321(.a(output_2_321), .b(output_2_2), .y(output_1_321));
wire output_3_321, output_3_2, output_2_321;
mixer gate_output_2_321(.a(output_3_321), .b(output_3_2), .y(output_2_321));
wire output_4_321, output_4_2, output_3_321;
mixer gate_output_3_321(.a(output_4_321), .b(output_4_2), .y(output_3_321));
wire output_5_321, output_5_2, output_4_321;
mixer gate_output_4_321(.a(output_5_321), .b(output_5_2), .y(output_4_321));
wire output_6_321, output_6_2, output_5_321;
mixer gate_output_5_321(.a(output_6_321), .b(output_6_2), .y(output_5_321));
wire output_7_321, output_7_2, output_6_321;
mixer gate_output_6_321(.a(output_7_321), .b(output_7_2), .y(output_6_321));
wire output_8_321, output_8_2, output_7_321;
mixer gate_output_7_321(.a(output_8_321), .b(output_8_2), .y(output_7_321));
wire output_9_321, output_9_2, output_8_321;
mixer gate_output_8_321(.a(output_9_321), .b(output_9_2), .y(output_8_321));
wire output_10_321, output_10_2, output_9_321;
mixer gate_output_9_321(.a(output_10_321), .b(output_10_2), .y(output_9_321));
wire output_11_321, output_11_2, output_10_321;
mixer gate_output_10_321(.a(output_11_321), .b(output_11_2), .y(output_10_321));
wire output_12_321, output_12_2, output_11_321;
mixer gate_output_11_321(.a(output_12_321), .b(output_12_2), .y(output_11_321));
wire output_13_321, output_13_2, output_12_321;
mixer gate_output_12_321(.a(output_13_321), .b(output_13_2), .y(output_12_321));
wire output_14_321, output_14_2, output_13_321;
mixer gate_output_13_321(.a(output_14_321), .b(output_14_2), .y(output_13_321));
wire output_15_321, output_15_2, output_14_321;
mixer gate_output_14_321(.a(output_15_321), .b(output_15_2), .y(output_14_321));
wire output_16_321, output_16_2, output_15_321;
mixer gate_output_15_321(.a(output_16_321), .b(output_16_2), .y(output_15_321));
wire output_1_322, output_1_3, output_0_322;
mixer gate_output_0_322(.a(output_1_322), .b(output_1_3), .y(output_0_322));
wire output_2_322, output_2_3, output_1_322;
mixer gate_output_1_322(.a(output_2_322), .b(output_2_3), .y(output_1_322));
wire output_3_322, output_3_3, output_2_322;
mixer gate_output_2_322(.a(output_3_322), .b(output_3_3), .y(output_2_322));
wire output_4_322, output_4_3, output_3_322;
mixer gate_output_3_322(.a(output_4_322), .b(output_4_3), .y(output_3_322));
wire output_5_322, output_5_3, output_4_322;
mixer gate_output_4_322(.a(output_5_322), .b(output_5_3), .y(output_4_322));
wire output_6_322, output_6_3, output_5_322;
mixer gate_output_5_322(.a(output_6_322), .b(output_6_3), .y(output_5_322));
wire output_7_322, output_7_3, output_6_322;
mixer gate_output_6_322(.a(output_7_322), .b(output_7_3), .y(output_6_322));
wire output_8_322, output_8_3, output_7_322;
mixer gate_output_7_322(.a(output_8_322), .b(output_8_3), .y(output_7_322));
wire output_9_322, output_9_3, output_8_322;
mixer gate_output_8_322(.a(output_9_322), .b(output_9_3), .y(output_8_322));
wire output_10_322, output_10_3, output_9_322;
mixer gate_output_9_322(.a(output_10_322), .b(output_10_3), .y(output_9_322));
wire output_11_322, output_11_3, output_10_322;
mixer gate_output_10_322(.a(output_11_322), .b(output_11_3), .y(output_10_322));
wire output_12_322, output_12_3, output_11_322;
mixer gate_output_11_322(.a(output_12_322), .b(output_12_3), .y(output_11_322));
wire output_13_322, output_13_3, output_12_322;
mixer gate_output_12_322(.a(output_13_322), .b(output_13_3), .y(output_12_322));
wire output_14_322, output_14_3, output_13_322;
mixer gate_output_13_322(.a(output_14_322), .b(output_14_3), .y(output_13_322));
wire output_15_322, output_15_3, output_14_322;
mixer gate_output_14_322(.a(output_15_322), .b(output_15_3), .y(output_14_322));
wire output_16_322, output_16_3, output_15_322;
mixer gate_output_15_322(.a(output_16_322), .b(output_16_3), .y(output_15_322));
wire output_1_323, output_1_4, output_0_323;
mixer gate_output_0_323(.a(output_1_323), .b(output_1_4), .y(output_0_323));
wire output_2_323, output_2_4, output_1_323;
mixer gate_output_1_323(.a(output_2_323), .b(output_2_4), .y(output_1_323));
wire output_3_323, output_3_4, output_2_323;
mixer gate_output_2_323(.a(output_3_323), .b(output_3_4), .y(output_2_323));
wire output_4_323, output_4_4, output_3_323;
mixer gate_output_3_323(.a(output_4_323), .b(output_4_4), .y(output_3_323));
wire output_5_323, output_5_4, output_4_323;
mixer gate_output_4_323(.a(output_5_323), .b(output_5_4), .y(output_4_323));
wire output_6_323, output_6_4, output_5_323;
mixer gate_output_5_323(.a(output_6_323), .b(output_6_4), .y(output_5_323));
wire output_7_323, output_7_4, output_6_323;
mixer gate_output_6_323(.a(output_7_323), .b(output_7_4), .y(output_6_323));
wire output_8_323, output_8_4, output_7_323;
mixer gate_output_7_323(.a(output_8_323), .b(output_8_4), .y(output_7_323));
wire output_9_323, output_9_4, output_8_323;
mixer gate_output_8_323(.a(output_9_323), .b(output_9_4), .y(output_8_323));
wire output_10_323, output_10_4, output_9_323;
mixer gate_output_9_323(.a(output_10_323), .b(output_10_4), .y(output_9_323));
wire output_11_323, output_11_4, output_10_323;
mixer gate_output_10_323(.a(output_11_323), .b(output_11_4), .y(output_10_323));
wire output_12_323, output_12_4, output_11_323;
mixer gate_output_11_323(.a(output_12_323), .b(output_12_4), .y(output_11_323));
wire output_13_323, output_13_4, output_12_323;
mixer gate_output_12_323(.a(output_13_323), .b(output_13_4), .y(output_12_323));
wire output_14_323, output_14_4, output_13_323;
mixer gate_output_13_323(.a(output_14_323), .b(output_14_4), .y(output_13_323));
wire output_15_323, output_15_4, output_14_323;
mixer gate_output_14_323(.a(output_15_323), .b(output_15_4), .y(output_14_323));
wire output_16_323, output_16_4, output_15_323;
mixer gate_output_15_323(.a(output_16_323), .b(output_16_4), .y(output_15_323));
wire output_1_324, output_1_5, output_0_324;
mixer gate_output_0_324(.a(output_1_324), .b(output_1_5), .y(output_0_324));
wire output_2_324, output_2_5, output_1_324;
mixer gate_output_1_324(.a(output_2_324), .b(output_2_5), .y(output_1_324));
wire output_3_324, output_3_5, output_2_324;
mixer gate_output_2_324(.a(output_3_324), .b(output_3_5), .y(output_2_324));
wire output_4_324, output_4_5, output_3_324;
mixer gate_output_3_324(.a(output_4_324), .b(output_4_5), .y(output_3_324));
wire output_5_324, output_5_5, output_4_324;
mixer gate_output_4_324(.a(output_5_324), .b(output_5_5), .y(output_4_324));
wire output_6_324, output_6_5, output_5_324;
mixer gate_output_5_324(.a(output_6_324), .b(output_6_5), .y(output_5_324));
wire output_7_324, output_7_5, output_6_324;
mixer gate_output_6_324(.a(output_7_324), .b(output_7_5), .y(output_6_324));
wire output_8_324, output_8_5, output_7_324;
mixer gate_output_7_324(.a(output_8_324), .b(output_8_5), .y(output_7_324));
wire output_9_324, output_9_5, output_8_324;
mixer gate_output_8_324(.a(output_9_324), .b(output_9_5), .y(output_8_324));
wire output_10_324, output_10_5, output_9_324;
mixer gate_output_9_324(.a(output_10_324), .b(output_10_5), .y(output_9_324));
wire output_11_324, output_11_5, output_10_324;
mixer gate_output_10_324(.a(output_11_324), .b(output_11_5), .y(output_10_324));
wire output_12_324, output_12_5, output_11_324;
mixer gate_output_11_324(.a(output_12_324), .b(output_12_5), .y(output_11_324));
wire output_13_324, output_13_5, output_12_324;
mixer gate_output_12_324(.a(output_13_324), .b(output_13_5), .y(output_12_324));
wire output_14_324, output_14_5, output_13_324;
mixer gate_output_13_324(.a(output_14_324), .b(output_14_5), .y(output_13_324));
wire output_15_324, output_15_5, output_14_324;
mixer gate_output_14_324(.a(output_15_324), .b(output_15_5), .y(output_14_324));
wire output_16_324, output_16_5, output_15_324;
mixer gate_output_15_324(.a(output_16_324), .b(output_16_5), .y(output_15_324));
wire output_1_325, output_1_6, output_0_325;
mixer gate_output_0_325(.a(output_1_325), .b(output_1_6), .y(output_0_325));
wire output_2_325, output_2_6, output_1_325;
mixer gate_output_1_325(.a(output_2_325), .b(output_2_6), .y(output_1_325));
wire output_3_325, output_3_6, output_2_325;
mixer gate_output_2_325(.a(output_3_325), .b(output_3_6), .y(output_2_325));
wire output_4_325, output_4_6, output_3_325;
mixer gate_output_3_325(.a(output_4_325), .b(output_4_6), .y(output_3_325));
wire output_5_325, output_5_6, output_4_325;
mixer gate_output_4_325(.a(output_5_325), .b(output_5_6), .y(output_4_325));
wire output_6_325, output_6_6, output_5_325;
mixer gate_output_5_325(.a(output_6_325), .b(output_6_6), .y(output_5_325));
wire output_7_325, output_7_6, output_6_325;
mixer gate_output_6_325(.a(output_7_325), .b(output_7_6), .y(output_6_325));
wire output_8_325, output_8_6, output_7_325;
mixer gate_output_7_325(.a(output_8_325), .b(output_8_6), .y(output_7_325));
wire output_9_325, output_9_6, output_8_325;
mixer gate_output_8_325(.a(output_9_325), .b(output_9_6), .y(output_8_325));
wire output_10_325, output_10_6, output_9_325;
mixer gate_output_9_325(.a(output_10_325), .b(output_10_6), .y(output_9_325));
wire output_11_325, output_11_6, output_10_325;
mixer gate_output_10_325(.a(output_11_325), .b(output_11_6), .y(output_10_325));
wire output_12_325, output_12_6, output_11_325;
mixer gate_output_11_325(.a(output_12_325), .b(output_12_6), .y(output_11_325));
wire output_13_325, output_13_6, output_12_325;
mixer gate_output_12_325(.a(output_13_325), .b(output_13_6), .y(output_12_325));
wire output_14_325, output_14_6, output_13_325;
mixer gate_output_13_325(.a(output_14_325), .b(output_14_6), .y(output_13_325));
wire output_15_325, output_15_6, output_14_325;
mixer gate_output_14_325(.a(output_15_325), .b(output_15_6), .y(output_14_325));
wire output_16_325, output_16_6, output_15_325;
mixer gate_output_15_325(.a(output_16_325), .b(output_16_6), .y(output_15_325));
wire output_1_326, output_1_7, output_0_326;
mixer gate_output_0_326(.a(output_1_326), .b(output_1_7), .y(output_0_326));
wire output_2_326, output_2_7, output_1_326;
mixer gate_output_1_326(.a(output_2_326), .b(output_2_7), .y(output_1_326));
wire output_3_326, output_3_7, output_2_326;
mixer gate_output_2_326(.a(output_3_326), .b(output_3_7), .y(output_2_326));
wire output_4_326, output_4_7, output_3_326;
mixer gate_output_3_326(.a(output_4_326), .b(output_4_7), .y(output_3_326));
wire output_5_326, output_5_7, output_4_326;
mixer gate_output_4_326(.a(output_5_326), .b(output_5_7), .y(output_4_326));
wire output_6_326, output_6_7, output_5_326;
mixer gate_output_5_326(.a(output_6_326), .b(output_6_7), .y(output_5_326));
wire output_7_326, output_7_7, output_6_326;
mixer gate_output_6_326(.a(output_7_326), .b(output_7_7), .y(output_6_326));
wire output_8_326, output_8_7, output_7_326;
mixer gate_output_7_326(.a(output_8_326), .b(output_8_7), .y(output_7_326));
wire output_9_326, output_9_7, output_8_326;
mixer gate_output_8_326(.a(output_9_326), .b(output_9_7), .y(output_8_326));
wire output_10_326, output_10_7, output_9_326;
mixer gate_output_9_326(.a(output_10_326), .b(output_10_7), .y(output_9_326));
wire output_11_326, output_11_7, output_10_326;
mixer gate_output_10_326(.a(output_11_326), .b(output_11_7), .y(output_10_326));
wire output_12_326, output_12_7, output_11_326;
mixer gate_output_11_326(.a(output_12_326), .b(output_12_7), .y(output_11_326));
wire output_13_326, output_13_7, output_12_326;
mixer gate_output_12_326(.a(output_13_326), .b(output_13_7), .y(output_12_326));
wire output_14_326, output_14_7, output_13_326;
mixer gate_output_13_326(.a(output_14_326), .b(output_14_7), .y(output_13_326));
wire output_15_326, output_15_7, output_14_326;
mixer gate_output_14_326(.a(output_15_326), .b(output_15_7), .y(output_14_326));
wire output_16_326, output_16_7, output_15_326;
mixer gate_output_15_326(.a(output_16_326), .b(output_16_7), .y(output_15_326));
wire output_1_327, output_1_8, output_0_327;
mixer gate_output_0_327(.a(output_1_327), .b(output_1_8), .y(output_0_327));
wire output_2_327, output_2_8, output_1_327;
mixer gate_output_1_327(.a(output_2_327), .b(output_2_8), .y(output_1_327));
wire output_3_327, output_3_8, output_2_327;
mixer gate_output_2_327(.a(output_3_327), .b(output_3_8), .y(output_2_327));
wire output_4_327, output_4_8, output_3_327;
mixer gate_output_3_327(.a(output_4_327), .b(output_4_8), .y(output_3_327));
wire output_5_327, output_5_8, output_4_327;
mixer gate_output_4_327(.a(output_5_327), .b(output_5_8), .y(output_4_327));
wire output_6_327, output_6_8, output_5_327;
mixer gate_output_5_327(.a(output_6_327), .b(output_6_8), .y(output_5_327));
wire output_7_327, output_7_8, output_6_327;
mixer gate_output_6_327(.a(output_7_327), .b(output_7_8), .y(output_6_327));
wire output_8_327, output_8_8, output_7_327;
mixer gate_output_7_327(.a(output_8_327), .b(output_8_8), .y(output_7_327));
wire output_9_327, output_9_8, output_8_327;
mixer gate_output_8_327(.a(output_9_327), .b(output_9_8), .y(output_8_327));
wire output_10_327, output_10_8, output_9_327;
mixer gate_output_9_327(.a(output_10_327), .b(output_10_8), .y(output_9_327));
wire output_11_327, output_11_8, output_10_327;
mixer gate_output_10_327(.a(output_11_327), .b(output_11_8), .y(output_10_327));
wire output_12_327, output_12_8, output_11_327;
mixer gate_output_11_327(.a(output_12_327), .b(output_12_8), .y(output_11_327));
wire output_13_327, output_13_8, output_12_327;
mixer gate_output_12_327(.a(output_13_327), .b(output_13_8), .y(output_12_327));
wire output_14_327, output_14_8, output_13_327;
mixer gate_output_13_327(.a(output_14_327), .b(output_14_8), .y(output_13_327));
wire output_15_327, output_15_8, output_14_327;
mixer gate_output_14_327(.a(output_15_327), .b(output_15_8), .y(output_14_327));
wire output_16_327, output_16_8, output_15_327;
mixer gate_output_15_327(.a(output_16_327), .b(output_16_8), .y(output_15_327));
wire output_1_328, output_1_9, output_0_328;
mixer gate_output_0_328(.a(output_1_328), .b(output_1_9), .y(output_0_328));
wire output_2_328, output_2_9, output_1_328;
mixer gate_output_1_328(.a(output_2_328), .b(output_2_9), .y(output_1_328));
wire output_3_328, output_3_9, output_2_328;
mixer gate_output_2_328(.a(output_3_328), .b(output_3_9), .y(output_2_328));
wire output_4_328, output_4_9, output_3_328;
mixer gate_output_3_328(.a(output_4_328), .b(output_4_9), .y(output_3_328));
wire output_5_328, output_5_9, output_4_328;
mixer gate_output_4_328(.a(output_5_328), .b(output_5_9), .y(output_4_328));
wire output_6_328, output_6_9, output_5_328;
mixer gate_output_5_328(.a(output_6_328), .b(output_6_9), .y(output_5_328));
wire output_7_328, output_7_9, output_6_328;
mixer gate_output_6_328(.a(output_7_328), .b(output_7_9), .y(output_6_328));
wire output_8_328, output_8_9, output_7_328;
mixer gate_output_7_328(.a(output_8_328), .b(output_8_9), .y(output_7_328));
wire output_9_328, output_9_9, output_8_328;
mixer gate_output_8_328(.a(output_9_328), .b(output_9_9), .y(output_8_328));
wire output_10_328, output_10_9, output_9_328;
mixer gate_output_9_328(.a(output_10_328), .b(output_10_9), .y(output_9_328));
wire output_11_328, output_11_9, output_10_328;
mixer gate_output_10_328(.a(output_11_328), .b(output_11_9), .y(output_10_328));
wire output_12_328, output_12_9, output_11_328;
mixer gate_output_11_328(.a(output_12_328), .b(output_12_9), .y(output_11_328));
wire output_13_328, output_13_9, output_12_328;
mixer gate_output_12_328(.a(output_13_328), .b(output_13_9), .y(output_12_328));
wire output_14_328, output_14_9, output_13_328;
mixer gate_output_13_328(.a(output_14_328), .b(output_14_9), .y(output_13_328));
wire output_15_328, output_15_9, output_14_328;
mixer gate_output_14_328(.a(output_15_328), .b(output_15_9), .y(output_14_328));
wire output_16_328, output_16_9, output_15_328;
mixer gate_output_15_328(.a(output_16_328), .b(output_16_9), .y(output_15_328));
wire output_1_329, output_1_10, output_0_329;
mixer gate_output_0_329(.a(output_1_329), .b(output_1_10), .y(output_0_329));
wire output_2_329, output_2_10, output_1_329;
mixer gate_output_1_329(.a(output_2_329), .b(output_2_10), .y(output_1_329));
wire output_3_329, output_3_10, output_2_329;
mixer gate_output_2_329(.a(output_3_329), .b(output_3_10), .y(output_2_329));
wire output_4_329, output_4_10, output_3_329;
mixer gate_output_3_329(.a(output_4_329), .b(output_4_10), .y(output_3_329));
wire output_5_329, output_5_10, output_4_329;
mixer gate_output_4_329(.a(output_5_329), .b(output_5_10), .y(output_4_329));
wire output_6_329, output_6_10, output_5_329;
mixer gate_output_5_329(.a(output_6_329), .b(output_6_10), .y(output_5_329));
wire output_7_329, output_7_10, output_6_329;
mixer gate_output_6_329(.a(output_7_329), .b(output_7_10), .y(output_6_329));
wire output_8_329, output_8_10, output_7_329;
mixer gate_output_7_329(.a(output_8_329), .b(output_8_10), .y(output_7_329));
wire output_9_329, output_9_10, output_8_329;
mixer gate_output_8_329(.a(output_9_329), .b(output_9_10), .y(output_8_329));
wire output_10_329, output_10_10, output_9_329;
mixer gate_output_9_329(.a(output_10_329), .b(output_10_10), .y(output_9_329));
wire output_11_329, output_11_10, output_10_329;
mixer gate_output_10_329(.a(output_11_329), .b(output_11_10), .y(output_10_329));
wire output_12_329, output_12_10, output_11_329;
mixer gate_output_11_329(.a(output_12_329), .b(output_12_10), .y(output_11_329));
wire output_13_329, output_13_10, output_12_329;
mixer gate_output_12_329(.a(output_13_329), .b(output_13_10), .y(output_12_329));
wire output_14_329, output_14_10, output_13_329;
mixer gate_output_13_329(.a(output_14_329), .b(output_14_10), .y(output_13_329));
wire output_15_329, output_15_10, output_14_329;
mixer gate_output_14_329(.a(output_15_329), .b(output_15_10), .y(output_14_329));
wire output_16_329, output_16_10, output_15_329;
mixer gate_output_15_329(.a(output_16_329), .b(output_16_10), .y(output_15_329));
wire output_1_330, output_1_11, output_0_330;
mixer gate_output_0_330(.a(output_1_330), .b(output_1_11), .y(output_0_330));
wire output_2_330, output_2_11, output_1_330;
mixer gate_output_1_330(.a(output_2_330), .b(output_2_11), .y(output_1_330));
wire output_3_330, output_3_11, output_2_330;
mixer gate_output_2_330(.a(output_3_330), .b(output_3_11), .y(output_2_330));
wire output_4_330, output_4_11, output_3_330;
mixer gate_output_3_330(.a(output_4_330), .b(output_4_11), .y(output_3_330));
wire output_5_330, output_5_11, output_4_330;
mixer gate_output_4_330(.a(output_5_330), .b(output_5_11), .y(output_4_330));
wire output_6_330, output_6_11, output_5_330;
mixer gate_output_5_330(.a(output_6_330), .b(output_6_11), .y(output_5_330));
wire output_7_330, output_7_11, output_6_330;
mixer gate_output_6_330(.a(output_7_330), .b(output_7_11), .y(output_6_330));
wire output_8_330, output_8_11, output_7_330;
mixer gate_output_7_330(.a(output_8_330), .b(output_8_11), .y(output_7_330));
wire output_9_330, output_9_11, output_8_330;
mixer gate_output_8_330(.a(output_9_330), .b(output_9_11), .y(output_8_330));
wire output_10_330, output_10_11, output_9_330;
mixer gate_output_9_330(.a(output_10_330), .b(output_10_11), .y(output_9_330));
wire output_11_330, output_11_11, output_10_330;
mixer gate_output_10_330(.a(output_11_330), .b(output_11_11), .y(output_10_330));
wire output_12_330, output_12_11, output_11_330;
mixer gate_output_11_330(.a(output_12_330), .b(output_12_11), .y(output_11_330));
wire output_13_330, output_13_11, output_12_330;
mixer gate_output_12_330(.a(output_13_330), .b(output_13_11), .y(output_12_330));
wire output_14_330, output_14_11, output_13_330;
mixer gate_output_13_330(.a(output_14_330), .b(output_14_11), .y(output_13_330));
wire output_15_330, output_15_11, output_14_330;
mixer gate_output_14_330(.a(output_15_330), .b(output_15_11), .y(output_14_330));
wire output_16_330, output_16_11, output_15_330;
mixer gate_output_15_330(.a(output_16_330), .b(output_16_11), .y(output_15_330));
wire output_1_331, output_1_12, output_0_331;
mixer gate_output_0_331(.a(output_1_331), .b(output_1_12), .y(output_0_331));
wire output_2_331, output_2_12, output_1_331;
mixer gate_output_1_331(.a(output_2_331), .b(output_2_12), .y(output_1_331));
wire output_3_331, output_3_12, output_2_331;
mixer gate_output_2_331(.a(output_3_331), .b(output_3_12), .y(output_2_331));
wire output_4_331, output_4_12, output_3_331;
mixer gate_output_3_331(.a(output_4_331), .b(output_4_12), .y(output_3_331));
wire output_5_331, output_5_12, output_4_331;
mixer gate_output_4_331(.a(output_5_331), .b(output_5_12), .y(output_4_331));
wire output_6_331, output_6_12, output_5_331;
mixer gate_output_5_331(.a(output_6_331), .b(output_6_12), .y(output_5_331));
wire output_7_331, output_7_12, output_6_331;
mixer gate_output_6_331(.a(output_7_331), .b(output_7_12), .y(output_6_331));
wire output_8_331, output_8_12, output_7_331;
mixer gate_output_7_331(.a(output_8_331), .b(output_8_12), .y(output_7_331));
wire output_9_331, output_9_12, output_8_331;
mixer gate_output_8_331(.a(output_9_331), .b(output_9_12), .y(output_8_331));
wire output_10_331, output_10_12, output_9_331;
mixer gate_output_9_331(.a(output_10_331), .b(output_10_12), .y(output_9_331));
wire output_11_331, output_11_12, output_10_331;
mixer gate_output_10_331(.a(output_11_331), .b(output_11_12), .y(output_10_331));
wire output_12_331, output_12_12, output_11_331;
mixer gate_output_11_331(.a(output_12_331), .b(output_12_12), .y(output_11_331));
wire output_13_331, output_13_12, output_12_331;
mixer gate_output_12_331(.a(output_13_331), .b(output_13_12), .y(output_12_331));
wire output_14_331, output_14_12, output_13_331;
mixer gate_output_13_331(.a(output_14_331), .b(output_14_12), .y(output_13_331));
wire output_15_331, output_15_12, output_14_331;
mixer gate_output_14_331(.a(output_15_331), .b(output_15_12), .y(output_14_331));
wire output_16_331, output_16_12, output_15_331;
mixer gate_output_15_331(.a(output_16_331), .b(output_16_12), .y(output_15_331));
wire output_1_332, output_1_13, output_0_332;
mixer gate_output_0_332(.a(output_1_332), .b(output_1_13), .y(output_0_332));
wire output_2_332, output_2_13, output_1_332;
mixer gate_output_1_332(.a(output_2_332), .b(output_2_13), .y(output_1_332));
wire output_3_332, output_3_13, output_2_332;
mixer gate_output_2_332(.a(output_3_332), .b(output_3_13), .y(output_2_332));
wire output_4_332, output_4_13, output_3_332;
mixer gate_output_3_332(.a(output_4_332), .b(output_4_13), .y(output_3_332));
wire output_5_332, output_5_13, output_4_332;
mixer gate_output_4_332(.a(output_5_332), .b(output_5_13), .y(output_4_332));
wire output_6_332, output_6_13, output_5_332;
mixer gate_output_5_332(.a(output_6_332), .b(output_6_13), .y(output_5_332));
wire output_7_332, output_7_13, output_6_332;
mixer gate_output_6_332(.a(output_7_332), .b(output_7_13), .y(output_6_332));
wire output_8_332, output_8_13, output_7_332;
mixer gate_output_7_332(.a(output_8_332), .b(output_8_13), .y(output_7_332));
wire output_9_332, output_9_13, output_8_332;
mixer gate_output_8_332(.a(output_9_332), .b(output_9_13), .y(output_8_332));
wire output_10_332, output_10_13, output_9_332;
mixer gate_output_9_332(.a(output_10_332), .b(output_10_13), .y(output_9_332));
wire output_11_332, output_11_13, output_10_332;
mixer gate_output_10_332(.a(output_11_332), .b(output_11_13), .y(output_10_332));
wire output_12_332, output_12_13, output_11_332;
mixer gate_output_11_332(.a(output_12_332), .b(output_12_13), .y(output_11_332));
wire output_13_332, output_13_13, output_12_332;
mixer gate_output_12_332(.a(output_13_332), .b(output_13_13), .y(output_12_332));
wire output_14_332, output_14_13, output_13_332;
mixer gate_output_13_332(.a(output_14_332), .b(output_14_13), .y(output_13_332));
wire output_15_332, output_15_13, output_14_332;
mixer gate_output_14_332(.a(output_15_332), .b(output_15_13), .y(output_14_332));
wire output_16_332, output_16_13, output_15_332;
mixer gate_output_15_332(.a(output_16_332), .b(output_16_13), .y(output_15_332));
wire output_1_333, output_1_14, output_0_333;
mixer gate_output_0_333(.a(output_1_333), .b(output_1_14), .y(output_0_333));
wire output_2_333, output_2_14, output_1_333;
mixer gate_output_1_333(.a(output_2_333), .b(output_2_14), .y(output_1_333));
wire output_3_333, output_3_14, output_2_333;
mixer gate_output_2_333(.a(output_3_333), .b(output_3_14), .y(output_2_333));
wire output_4_333, output_4_14, output_3_333;
mixer gate_output_3_333(.a(output_4_333), .b(output_4_14), .y(output_3_333));
wire output_5_333, output_5_14, output_4_333;
mixer gate_output_4_333(.a(output_5_333), .b(output_5_14), .y(output_4_333));
wire output_6_333, output_6_14, output_5_333;
mixer gate_output_5_333(.a(output_6_333), .b(output_6_14), .y(output_5_333));
wire output_7_333, output_7_14, output_6_333;
mixer gate_output_6_333(.a(output_7_333), .b(output_7_14), .y(output_6_333));
wire output_8_333, output_8_14, output_7_333;
mixer gate_output_7_333(.a(output_8_333), .b(output_8_14), .y(output_7_333));
wire output_9_333, output_9_14, output_8_333;
mixer gate_output_8_333(.a(output_9_333), .b(output_9_14), .y(output_8_333));
wire output_10_333, output_10_14, output_9_333;
mixer gate_output_9_333(.a(output_10_333), .b(output_10_14), .y(output_9_333));
wire output_11_333, output_11_14, output_10_333;
mixer gate_output_10_333(.a(output_11_333), .b(output_11_14), .y(output_10_333));
wire output_12_333, output_12_14, output_11_333;
mixer gate_output_11_333(.a(output_12_333), .b(output_12_14), .y(output_11_333));
wire output_13_333, output_13_14, output_12_333;
mixer gate_output_12_333(.a(output_13_333), .b(output_13_14), .y(output_12_333));
wire output_14_333, output_14_14, output_13_333;
mixer gate_output_13_333(.a(output_14_333), .b(output_14_14), .y(output_13_333));
wire output_15_333, output_15_14, output_14_333;
mixer gate_output_14_333(.a(output_15_333), .b(output_15_14), .y(output_14_333));
wire output_16_333, output_16_14, output_15_333;
mixer gate_output_15_333(.a(output_16_333), .b(output_16_14), .y(output_15_333));
wire output_1_334, output_1_15, output_0_334;
mixer gate_output_0_334(.a(output_1_334), .b(output_1_15), .y(output_0_334));
wire output_2_334, output_2_15, output_1_334;
mixer gate_output_1_334(.a(output_2_334), .b(output_2_15), .y(output_1_334));
wire output_3_334, output_3_15, output_2_334;
mixer gate_output_2_334(.a(output_3_334), .b(output_3_15), .y(output_2_334));
wire output_4_334, output_4_15, output_3_334;
mixer gate_output_3_334(.a(output_4_334), .b(output_4_15), .y(output_3_334));
wire output_5_334, output_5_15, output_4_334;
mixer gate_output_4_334(.a(output_5_334), .b(output_5_15), .y(output_4_334));
wire output_6_334, output_6_15, output_5_334;
mixer gate_output_5_334(.a(output_6_334), .b(output_6_15), .y(output_5_334));
wire output_7_334, output_7_15, output_6_334;
mixer gate_output_6_334(.a(output_7_334), .b(output_7_15), .y(output_6_334));
wire output_8_334, output_8_15, output_7_334;
mixer gate_output_7_334(.a(output_8_334), .b(output_8_15), .y(output_7_334));
wire output_9_334, output_9_15, output_8_334;
mixer gate_output_8_334(.a(output_9_334), .b(output_9_15), .y(output_8_334));
wire output_10_334, output_10_15, output_9_334;
mixer gate_output_9_334(.a(output_10_334), .b(output_10_15), .y(output_9_334));
wire output_11_334, output_11_15, output_10_334;
mixer gate_output_10_334(.a(output_11_334), .b(output_11_15), .y(output_10_334));
wire output_12_334, output_12_15, output_11_334;
mixer gate_output_11_334(.a(output_12_334), .b(output_12_15), .y(output_11_334));
wire output_13_334, output_13_15, output_12_334;
mixer gate_output_12_334(.a(output_13_334), .b(output_13_15), .y(output_12_334));
wire output_14_334, output_14_15, output_13_334;
mixer gate_output_13_334(.a(output_14_334), .b(output_14_15), .y(output_13_334));
wire output_15_334, output_15_15, output_14_334;
mixer gate_output_14_334(.a(output_15_334), .b(output_15_15), .y(output_14_334));
wire output_16_334, output_16_15, output_15_334;
mixer gate_output_15_334(.a(output_16_334), .b(output_16_15), .y(output_15_334));
wire output_1_335, output_1_0, output_0_335;
mixer gate_output_0_335(.a(output_1_335), .b(output_1_0), .y(output_0_335));
wire output_2_335, output_2_0, output_1_335;
mixer gate_output_1_335(.a(output_2_335), .b(output_2_0), .y(output_1_335));
wire output_3_335, output_3_0, output_2_335;
mixer gate_output_2_335(.a(output_3_335), .b(output_3_0), .y(output_2_335));
wire output_4_335, output_4_0, output_3_335;
mixer gate_output_3_335(.a(output_4_335), .b(output_4_0), .y(output_3_335));
wire output_5_335, output_5_0, output_4_335;
mixer gate_output_4_335(.a(output_5_335), .b(output_5_0), .y(output_4_335));
wire output_6_335, output_6_0, output_5_335;
mixer gate_output_5_335(.a(output_6_335), .b(output_6_0), .y(output_5_335));
wire output_7_335, output_7_0, output_6_335;
mixer gate_output_6_335(.a(output_7_335), .b(output_7_0), .y(output_6_335));
wire output_8_335, output_8_0, output_7_335;
mixer gate_output_7_335(.a(output_8_335), .b(output_8_0), .y(output_7_335));
wire output_9_335, output_9_0, output_8_335;
mixer gate_output_8_335(.a(output_9_335), .b(output_9_0), .y(output_8_335));
wire output_10_335, output_10_0, output_9_335;
mixer gate_output_9_335(.a(output_10_335), .b(output_10_0), .y(output_9_335));
wire output_11_335, output_11_0, output_10_335;
mixer gate_output_10_335(.a(output_11_335), .b(output_11_0), .y(output_10_335));
wire output_12_335, output_12_0, output_11_335;
mixer gate_output_11_335(.a(output_12_335), .b(output_12_0), .y(output_11_335));
wire output_13_335, output_13_0, output_12_335;
mixer gate_output_12_335(.a(output_13_335), .b(output_13_0), .y(output_12_335));
wire output_14_335, output_14_0, output_13_335;
mixer gate_output_13_335(.a(output_14_335), .b(output_14_0), .y(output_13_335));
wire output_15_335, output_15_0, output_14_335;
mixer gate_output_14_335(.a(output_15_335), .b(output_15_0), .y(output_14_335));
wire output_16_335, output_16_0, output_15_335;
mixer gate_output_15_335(.a(output_16_335), .b(output_16_0), .y(output_15_335));
wire output_1_336, output_1_1, output_0_336;
mixer gate_output_0_336(.a(output_1_336), .b(output_1_1), .y(output_0_336));
wire output_2_336, output_2_1, output_1_336;
mixer gate_output_1_336(.a(output_2_336), .b(output_2_1), .y(output_1_336));
wire output_3_336, output_3_1, output_2_336;
mixer gate_output_2_336(.a(output_3_336), .b(output_3_1), .y(output_2_336));
wire output_4_336, output_4_1, output_3_336;
mixer gate_output_3_336(.a(output_4_336), .b(output_4_1), .y(output_3_336));
wire output_5_336, output_5_1, output_4_336;
mixer gate_output_4_336(.a(output_5_336), .b(output_5_1), .y(output_4_336));
wire output_6_336, output_6_1, output_5_336;
mixer gate_output_5_336(.a(output_6_336), .b(output_6_1), .y(output_5_336));
wire output_7_336, output_7_1, output_6_336;
mixer gate_output_6_336(.a(output_7_336), .b(output_7_1), .y(output_6_336));
wire output_8_336, output_8_1, output_7_336;
mixer gate_output_7_336(.a(output_8_336), .b(output_8_1), .y(output_7_336));
wire output_9_336, output_9_1, output_8_336;
mixer gate_output_8_336(.a(output_9_336), .b(output_9_1), .y(output_8_336));
wire output_10_336, output_10_1, output_9_336;
mixer gate_output_9_336(.a(output_10_336), .b(output_10_1), .y(output_9_336));
wire output_11_336, output_11_1, output_10_336;
mixer gate_output_10_336(.a(output_11_336), .b(output_11_1), .y(output_10_336));
wire output_12_336, output_12_1, output_11_336;
mixer gate_output_11_336(.a(output_12_336), .b(output_12_1), .y(output_11_336));
wire output_13_336, output_13_1, output_12_336;
mixer gate_output_12_336(.a(output_13_336), .b(output_13_1), .y(output_12_336));
wire output_14_336, output_14_1, output_13_336;
mixer gate_output_13_336(.a(output_14_336), .b(output_14_1), .y(output_13_336));
wire output_15_336, output_15_1, output_14_336;
mixer gate_output_14_336(.a(output_15_336), .b(output_15_1), .y(output_14_336));
wire output_16_336, output_16_1, output_15_336;
mixer gate_output_15_336(.a(output_16_336), .b(output_16_1), .y(output_15_336));
wire output_1_337, output_1_2, output_0_337;
mixer gate_output_0_337(.a(output_1_337), .b(output_1_2), .y(output_0_337));
wire output_2_337, output_2_2, output_1_337;
mixer gate_output_1_337(.a(output_2_337), .b(output_2_2), .y(output_1_337));
wire output_3_337, output_3_2, output_2_337;
mixer gate_output_2_337(.a(output_3_337), .b(output_3_2), .y(output_2_337));
wire output_4_337, output_4_2, output_3_337;
mixer gate_output_3_337(.a(output_4_337), .b(output_4_2), .y(output_3_337));
wire output_5_337, output_5_2, output_4_337;
mixer gate_output_4_337(.a(output_5_337), .b(output_5_2), .y(output_4_337));
wire output_6_337, output_6_2, output_5_337;
mixer gate_output_5_337(.a(output_6_337), .b(output_6_2), .y(output_5_337));
wire output_7_337, output_7_2, output_6_337;
mixer gate_output_6_337(.a(output_7_337), .b(output_7_2), .y(output_6_337));
wire output_8_337, output_8_2, output_7_337;
mixer gate_output_7_337(.a(output_8_337), .b(output_8_2), .y(output_7_337));
wire output_9_337, output_9_2, output_8_337;
mixer gate_output_8_337(.a(output_9_337), .b(output_9_2), .y(output_8_337));
wire output_10_337, output_10_2, output_9_337;
mixer gate_output_9_337(.a(output_10_337), .b(output_10_2), .y(output_9_337));
wire output_11_337, output_11_2, output_10_337;
mixer gate_output_10_337(.a(output_11_337), .b(output_11_2), .y(output_10_337));
wire output_12_337, output_12_2, output_11_337;
mixer gate_output_11_337(.a(output_12_337), .b(output_12_2), .y(output_11_337));
wire output_13_337, output_13_2, output_12_337;
mixer gate_output_12_337(.a(output_13_337), .b(output_13_2), .y(output_12_337));
wire output_14_337, output_14_2, output_13_337;
mixer gate_output_13_337(.a(output_14_337), .b(output_14_2), .y(output_13_337));
wire output_15_337, output_15_2, output_14_337;
mixer gate_output_14_337(.a(output_15_337), .b(output_15_2), .y(output_14_337));
wire output_16_337, output_16_2, output_15_337;
mixer gate_output_15_337(.a(output_16_337), .b(output_16_2), .y(output_15_337));
wire output_1_338, output_1_3, output_0_338;
mixer gate_output_0_338(.a(output_1_338), .b(output_1_3), .y(output_0_338));
wire output_2_338, output_2_3, output_1_338;
mixer gate_output_1_338(.a(output_2_338), .b(output_2_3), .y(output_1_338));
wire output_3_338, output_3_3, output_2_338;
mixer gate_output_2_338(.a(output_3_338), .b(output_3_3), .y(output_2_338));
wire output_4_338, output_4_3, output_3_338;
mixer gate_output_3_338(.a(output_4_338), .b(output_4_3), .y(output_3_338));
wire output_5_338, output_5_3, output_4_338;
mixer gate_output_4_338(.a(output_5_338), .b(output_5_3), .y(output_4_338));
wire output_6_338, output_6_3, output_5_338;
mixer gate_output_5_338(.a(output_6_338), .b(output_6_3), .y(output_5_338));
wire output_7_338, output_7_3, output_6_338;
mixer gate_output_6_338(.a(output_7_338), .b(output_7_3), .y(output_6_338));
wire output_8_338, output_8_3, output_7_338;
mixer gate_output_7_338(.a(output_8_338), .b(output_8_3), .y(output_7_338));
wire output_9_338, output_9_3, output_8_338;
mixer gate_output_8_338(.a(output_9_338), .b(output_9_3), .y(output_8_338));
wire output_10_338, output_10_3, output_9_338;
mixer gate_output_9_338(.a(output_10_338), .b(output_10_3), .y(output_9_338));
wire output_11_338, output_11_3, output_10_338;
mixer gate_output_10_338(.a(output_11_338), .b(output_11_3), .y(output_10_338));
wire output_12_338, output_12_3, output_11_338;
mixer gate_output_11_338(.a(output_12_338), .b(output_12_3), .y(output_11_338));
wire output_13_338, output_13_3, output_12_338;
mixer gate_output_12_338(.a(output_13_338), .b(output_13_3), .y(output_12_338));
wire output_14_338, output_14_3, output_13_338;
mixer gate_output_13_338(.a(output_14_338), .b(output_14_3), .y(output_13_338));
wire output_15_338, output_15_3, output_14_338;
mixer gate_output_14_338(.a(output_15_338), .b(output_15_3), .y(output_14_338));
wire output_16_338, output_16_3, output_15_338;
mixer gate_output_15_338(.a(output_16_338), .b(output_16_3), .y(output_15_338));
wire output_1_339, output_1_4, output_0_339;
mixer gate_output_0_339(.a(output_1_339), .b(output_1_4), .y(output_0_339));
wire output_2_339, output_2_4, output_1_339;
mixer gate_output_1_339(.a(output_2_339), .b(output_2_4), .y(output_1_339));
wire output_3_339, output_3_4, output_2_339;
mixer gate_output_2_339(.a(output_3_339), .b(output_3_4), .y(output_2_339));
wire output_4_339, output_4_4, output_3_339;
mixer gate_output_3_339(.a(output_4_339), .b(output_4_4), .y(output_3_339));
wire output_5_339, output_5_4, output_4_339;
mixer gate_output_4_339(.a(output_5_339), .b(output_5_4), .y(output_4_339));
wire output_6_339, output_6_4, output_5_339;
mixer gate_output_5_339(.a(output_6_339), .b(output_6_4), .y(output_5_339));
wire output_7_339, output_7_4, output_6_339;
mixer gate_output_6_339(.a(output_7_339), .b(output_7_4), .y(output_6_339));
wire output_8_339, output_8_4, output_7_339;
mixer gate_output_7_339(.a(output_8_339), .b(output_8_4), .y(output_7_339));
wire output_9_339, output_9_4, output_8_339;
mixer gate_output_8_339(.a(output_9_339), .b(output_9_4), .y(output_8_339));
wire output_10_339, output_10_4, output_9_339;
mixer gate_output_9_339(.a(output_10_339), .b(output_10_4), .y(output_9_339));
wire output_11_339, output_11_4, output_10_339;
mixer gate_output_10_339(.a(output_11_339), .b(output_11_4), .y(output_10_339));
wire output_12_339, output_12_4, output_11_339;
mixer gate_output_11_339(.a(output_12_339), .b(output_12_4), .y(output_11_339));
wire output_13_339, output_13_4, output_12_339;
mixer gate_output_12_339(.a(output_13_339), .b(output_13_4), .y(output_12_339));
wire output_14_339, output_14_4, output_13_339;
mixer gate_output_13_339(.a(output_14_339), .b(output_14_4), .y(output_13_339));
wire output_15_339, output_15_4, output_14_339;
mixer gate_output_14_339(.a(output_15_339), .b(output_15_4), .y(output_14_339));
wire output_16_339, output_16_4, output_15_339;
mixer gate_output_15_339(.a(output_16_339), .b(output_16_4), .y(output_15_339));
wire output_1_340, output_1_5, output_0_340;
mixer gate_output_0_340(.a(output_1_340), .b(output_1_5), .y(output_0_340));
wire output_2_340, output_2_5, output_1_340;
mixer gate_output_1_340(.a(output_2_340), .b(output_2_5), .y(output_1_340));
wire output_3_340, output_3_5, output_2_340;
mixer gate_output_2_340(.a(output_3_340), .b(output_3_5), .y(output_2_340));
wire output_4_340, output_4_5, output_3_340;
mixer gate_output_3_340(.a(output_4_340), .b(output_4_5), .y(output_3_340));
wire output_5_340, output_5_5, output_4_340;
mixer gate_output_4_340(.a(output_5_340), .b(output_5_5), .y(output_4_340));
wire output_6_340, output_6_5, output_5_340;
mixer gate_output_5_340(.a(output_6_340), .b(output_6_5), .y(output_5_340));
wire output_7_340, output_7_5, output_6_340;
mixer gate_output_6_340(.a(output_7_340), .b(output_7_5), .y(output_6_340));
wire output_8_340, output_8_5, output_7_340;
mixer gate_output_7_340(.a(output_8_340), .b(output_8_5), .y(output_7_340));
wire output_9_340, output_9_5, output_8_340;
mixer gate_output_8_340(.a(output_9_340), .b(output_9_5), .y(output_8_340));
wire output_10_340, output_10_5, output_9_340;
mixer gate_output_9_340(.a(output_10_340), .b(output_10_5), .y(output_9_340));
wire output_11_340, output_11_5, output_10_340;
mixer gate_output_10_340(.a(output_11_340), .b(output_11_5), .y(output_10_340));
wire output_12_340, output_12_5, output_11_340;
mixer gate_output_11_340(.a(output_12_340), .b(output_12_5), .y(output_11_340));
wire output_13_340, output_13_5, output_12_340;
mixer gate_output_12_340(.a(output_13_340), .b(output_13_5), .y(output_12_340));
wire output_14_340, output_14_5, output_13_340;
mixer gate_output_13_340(.a(output_14_340), .b(output_14_5), .y(output_13_340));
wire output_15_340, output_15_5, output_14_340;
mixer gate_output_14_340(.a(output_15_340), .b(output_15_5), .y(output_14_340));
wire output_16_340, output_16_5, output_15_340;
mixer gate_output_15_340(.a(output_16_340), .b(output_16_5), .y(output_15_340));
wire output_1_341, output_1_6, output_0_341;
mixer gate_output_0_341(.a(output_1_341), .b(output_1_6), .y(output_0_341));
wire output_2_341, output_2_6, output_1_341;
mixer gate_output_1_341(.a(output_2_341), .b(output_2_6), .y(output_1_341));
wire output_3_341, output_3_6, output_2_341;
mixer gate_output_2_341(.a(output_3_341), .b(output_3_6), .y(output_2_341));
wire output_4_341, output_4_6, output_3_341;
mixer gate_output_3_341(.a(output_4_341), .b(output_4_6), .y(output_3_341));
wire output_5_341, output_5_6, output_4_341;
mixer gate_output_4_341(.a(output_5_341), .b(output_5_6), .y(output_4_341));
wire output_6_341, output_6_6, output_5_341;
mixer gate_output_5_341(.a(output_6_341), .b(output_6_6), .y(output_5_341));
wire output_7_341, output_7_6, output_6_341;
mixer gate_output_6_341(.a(output_7_341), .b(output_7_6), .y(output_6_341));
wire output_8_341, output_8_6, output_7_341;
mixer gate_output_7_341(.a(output_8_341), .b(output_8_6), .y(output_7_341));
wire output_9_341, output_9_6, output_8_341;
mixer gate_output_8_341(.a(output_9_341), .b(output_9_6), .y(output_8_341));
wire output_10_341, output_10_6, output_9_341;
mixer gate_output_9_341(.a(output_10_341), .b(output_10_6), .y(output_9_341));
wire output_11_341, output_11_6, output_10_341;
mixer gate_output_10_341(.a(output_11_341), .b(output_11_6), .y(output_10_341));
wire output_12_341, output_12_6, output_11_341;
mixer gate_output_11_341(.a(output_12_341), .b(output_12_6), .y(output_11_341));
wire output_13_341, output_13_6, output_12_341;
mixer gate_output_12_341(.a(output_13_341), .b(output_13_6), .y(output_12_341));
wire output_14_341, output_14_6, output_13_341;
mixer gate_output_13_341(.a(output_14_341), .b(output_14_6), .y(output_13_341));
wire output_15_341, output_15_6, output_14_341;
mixer gate_output_14_341(.a(output_15_341), .b(output_15_6), .y(output_14_341));
wire output_16_341, output_16_6, output_15_341;
mixer gate_output_15_341(.a(output_16_341), .b(output_16_6), .y(output_15_341));
wire output_1_342, output_1_7, output_0_342;
mixer gate_output_0_342(.a(output_1_342), .b(output_1_7), .y(output_0_342));
wire output_2_342, output_2_7, output_1_342;
mixer gate_output_1_342(.a(output_2_342), .b(output_2_7), .y(output_1_342));
wire output_3_342, output_3_7, output_2_342;
mixer gate_output_2_342(.a(output_3_342), .b(output_3_7), .y(output_2_342));
wire output_4_342, output_4_7, output_3_342;
mixer gate_output_3_342(.a(output_4_342), .b(output_4_7), .y(output_3_342));
wire output_5_342, output_5_7, output_4_342;
mixer gate_output_4_342(.a(output_5_342), .b(output_5_7), .y(output_4_342));
wire output_6_342, output_6_7, output_5_342;
mixer gate_output_5_342(.a(output_6_342), .b(output_6_7), .y(output_5_342));
wire output_7_342, output_7_7, output_6_342;
mixer gate_output_6_342(.a(output_7_342), .b(output_7_7), .y(output_6_342));
wire output_8_342, output_8_7, output_7_342;
mixer gate_output_7_342(.a(output_8_342), .b(output_8_7), .y(output_7_342));
wire output_9_342, output_9_7, output_8_342;
mixer gate_output_8_342(.a(output_9_342), .b(output_9_7), .y(output_8_342));
wire output_10_342, output_10_7, output_9_342;
mixer gate_output_9_342(.a(output_10_342), .b(output_10_7), .y(output_9_342));
wire output_11_342, output_11_7, output_10_342;
mixer gate_output_10_342(.a(output_11_342), .b(output_11_7), .y(output_10_342));
wire output_12_342, output_12_7, output_11_342;
mixer gate_output_11_342(.a(output_12_342), .b(output_12_7), .y(output_11_342));
wire output_13_342, output_13_7, output_12_342;
mixer gate_output_12_342(.a(output_13_342), .b(output_13_7), .y(output_12_342));
wire output_14_342, output_14_7, output_13_342;
mixer gate_output_13_342(.a(output_14_342), .b(output_14_7), .y(output_13_342));
wire output_15_342, output_15_7, output_14_342;
mixer gate_output_14_342(.a(output_15_342), .b(output_15_7), .y(output_14_342));
wire output_16_342, output_16_7, output_15_342;
mixer gate_output_15_342(.a(output_16_342), .b(output_16_7), .y(output_15_342));
wire output_1_343, output_1_8, output_0_343;
mixer gate_output_0_343(.a(output_1_343), .b(output_1_8), .y(output_0_343));
wire output_2_343, output_2_8, output_1_343;
mixer gate_output_1_343(.a(output_2_343), .b(output_2_8), .y(output_1_343));
wire output_3_343, output_3_8, output_2_343;
mixer gate_output_2_343(.a(output_3_343), .b(output_3_8), .y(output_2_343));
wire output_4_343, output_4_8, output_3_343;
mixer gate_output_3_343(.a(output_4_343), .b(output_4_8), .y(output_3_343));
wire output_5_343, output_5_8, output_4_343;
mixer gate_output_4_343(.a(output_5_343), .b(output_5_8), .y(output_4_343));
wire output_6_343, output_6_8, output_5_343;
mixer gate_output_5_343(.a(output_6_343), .b(output_6_8), .y(output_5_343));
wire output_7_343, output_7_8, output_6_343;
mixer gate_output_6_343(.a(output_7_343), .b(output_7_8), .y(output_6_343));
wire output_8_343, output_8_8, output_7_343;
mixer gate_output_7_343(.a(output_8_343), .b(output_8_8), .y(output_7_343));
wire output_9_343, output_9_8, output_8_343;
mixer gate_output_8_343(.a(output_9_343), .b(output_9_8), .y(output_8_343));
wire output_10_343, output_10_8, output_9_343;
mixer gate_output_9_343(.a(output_10_343), .b(output_10_8), .y(output_9_343));
wire output_11_343, output_11_8, output_10_343;
mixer gate_output_10_343(.a(output_11_343), .b(output_11_8), .y(output_10_343));
wire output_12_343, output_12_8, output_11_343;
mixer gate_output_11_343(.a(output_12_343), .b(output_12_8), .y(output_11_343));
wire output_13_343, output_13_8, output_12_343;
mixer gate_output_12_343(.a(output_13_343), .b(output_13_8), .y(output_12_343));
wire output_14_343, output_14_8, output_13_343;
mixer gate_output_13_343(.a(output_14_343), .b(output_14_8), .y(output_13_343));
wire output_15_343, output_15_8, output_14_343;
mixer gate_output_14_343(.a(output_15_343), .b(output_15_8), .y(output_14_343));
wire output_16_343, output_16_8, output_15_343;
mixer gate_output_15_343(.a(output_16_343), .b(output_16_8), .y(output_15_343));
wire output_1_344, output_1_9, output_0_344;
mixer gate_output_0_344(.a(output_1_344), .b(output_1_9), .y(output_0_344));
wire output_2_344, output_2_9, output_1_344;
mixer gate_output_1_344(.a(output_2_344), .b(output_2_9), .y(output_1_344));
wire output_3_344, output_3_9, output_2_344;
mixer gate_output_2_344(.a(output_3_344), .b(output_3_9), .y(output_2_344));
wire output_4_344, output_4_9, output_3_344;
mixer gate_output_3_344(.a(output_4_344), .b(output_4_9), .y(output_3_344));
wire output_5_344, output_5_9, output_4_344;
mixer gate_output_4_344(.a(output_5_344), .b(output_5_9), .y(output_4_344));
wire output_6_344, output_6_9, output_5_344;
mixer gate_output_5_344(.a(output_6_344), .b(output_6_9), .y(output_5_344));
wire output_7_344, output_7_9, output_6_344;
mixer gate_output_6_344(.a(output_7_344), .b(output_7_9), .y(output_6_344));
wire output_8_344, output_8_9, output_7_344;
mixer gate_output_7_344(.a(output_8_344), .b(output_8_9), .y(output_7_344));
wire output_9_344, output_9_9, output_8_344;
mixer gate_output_8_344(.a(output_9_344), .b(output_9_9), .y(output_8_344));
wire output_10_344, output_10_9, output_9_344;
mixer gate_output_9_344(.a(output_10_344), .b(output_10_9), .y(output_9_344));
wire output_11_344, output_11_9, output_10_344;
mixer gate_output_10_344(.a(output_11_344), .b(output_11_9), .y(output_10_344));
wire output_12_344, output_12_9, output_11_344;
mixer gate_output_11_344(.a(output_12_344), .b(output_12_9), .y(output_11_344));
wire output_13_344, output_13_9, output_12_344;
mixer gate_output_12_344(.a(output_13_344), .b(output_13_9), .y(output_12_344));
wire output_14_344, output_14_9, output_13_344;
mixer gate_output_13_344(.a(output_14_344), .b(output_14_9), .y(output_13_344));
wire output_15_344, output_15_9, output_14_344;
mixer gate_output_14_344(.a(output_15_344), .b(output_15_9), .y(output_14_344));
wire output_16_344, output_16_9, output_15_344;
mixer gate_output_15_344(.a(output_16_344), .b(output_16_9), .y(output_15_344));
wire output_1_345, output_1_10, output_0_345;
mixer gate_output_0_345(.a(output_1_345), .b(output_1_10), .y(output_0_345));
wire output_2_345, output_2_10, output_1_345;
mixer gate_output_1_345(.a(output_2_345), .b(output_2_10), .y(output_1_345));
wire output_3_345, output_3_10, output_2_345;
mixer gate_output_2_345(.a(output_3_345), .b(output_3_10), .y(output_2_345));
wire output_4_345, output_4_10, output_3_345;
mixer gate_output_3_345(.a(output_4_345), .b(output_4_10), .y(output_3_345));
wire output_5_345, output_5_10, output_4_345;
mixer gate_output_4_345(.a(output_5_345), .b(output_5_10), .y(output_4_345));
wire output_6_345, output_6_10, output_5_345;
mixer gate_output_5_345(.a(output_6_345), .b(output_6_10), .y(output_5_345));
wire output_7_345, output_7_10, output_6_345;
mixer gate_output_6_345(.a(output_7_345), .b(output_7_10), .y(output_6_345));
wire output_8_345, output_8_10, output_7_345;
mixer gate_output_7_345(.a(output_8_345), .b(output_8_10), .y(output_7_345));
wire output_9_345, output_9_10, output_8_345;
mixer gate_output_8_345(.a(output_9_345), .b(output_9_10), .y(output_8_345));
wire output_10_345, output_10_10, output_9_345;
mixer gate_output_9_345(.a(output_10_345), .b(output_10_10), .y(output_9_345));
wire output_11_345, output_11_10, output_10_345;
mixer gate_output_10_345(.a(output_11_345), .b(output_11_10), .y(output_10_345));
wire output_12_345, output_12_10, output_11_345;
mixer gate_output_11_345(.a(output_12_345), .b(output_12_10), .y(output_11_345));
wire output_13_345, output_13_10, output_12_345;
mixer gate_output_12_345(.a(output_13_345), .b(output_13_10), .y(output_12_345));
wire output_14_345, output_14_10, output_13_345;
mixer gate_output_13_345(.a(output_14_345), .b(output_14_10), .y(output_13_345));
wire output_15_345, output_15_10, output_14_345;
mixer gate_output_14_345(.a(output_15_345), .b(output_15_10), .y(output_14_345));
wire output_16_345, output_16_10, output_15_345;
mixer gate_output_15_345(.a(output_16_345), .b(output_16_10), .y(output_15_345));
wire output_1_346, output_1_11, output_0_346;
mixer gate_output_0_346(.a(output_1_346), .b(output_1_11), .y(output_0_346));
wire output_2_346, output_2_11, output_1_346;
mixer gate_output_1_346(.a(output_2_346), .b(output_2_11), .y(output_1_346));
wire output_3_346, output_3_11, output_2_346;
mixer gate_output_2_346(.a(output_3_346), .b(output_3_11), .y(output_2_346));
wire output_4_346, output_4_11, output_3_346;
mixer gate_output_3_346(.a(output_4_346), .b(output_4_11), .y(output_3_346));
wire output_5_346, output_5_11, output_4_346;
mixer gate_output_4_346(.a(output_5_346), .b(output_5_11), .y(output_4_346));
wire output_6_346, output_6_11, output_5_346;
mixer gate_output_5_346(.a(output_6_346), .b(output_6_11), .y(output_5_346));
wire output_7_346, output_7_11, output_6_346;
mixer gate_output_6_346(.a(output_7_346), .b(output_7_11), .y(output_6_346));
wire output_8_346, output_8_11, output_7_346;
mixer gate_output_7_346(.a(output_8_346), .b(output_8_11), .y(output_7_346));
wire output_9_346, output_9_11, output_8_346;
mixer gate_output_8_346(.a(output_9_346), .b(output_9_11), .y(output_8_346));
wire output_10_346, output_10_11, output_9_346;
mixer gate_output_9_346(.a(output_10_346), .b(output_10_11), .y(output_9_346));
wire output_11_346, output_11_11, output_10_346;
mixer gate_output_10_346(.a(output_11_346), .b(output_11_11), .y(output_10_346));
wire output_12_346, output_12_11, output_11_346;
mixer gate_output_11_346(.a(output_12_346), .b(output_12_11), .y(output_11_346));
wire output_13_346, output_13_11, output_12_346;
mixer gate_output_12_346(.a(output_13_346), .b(output_13_11), .y(output_12_346));
wire output_14_346, output_14_11, output_13_346;
mixer gate_output_13_346(.a(output_14_346), .b(output_14_11), .y(output_13_346));
wire output_15_346, output_15_11, output_14_346;
mixer gate_output_14_346(.a(output_15_346), .b(output_15_11), .y(output_14_346));
wire output_16_346, output_16_11, output_15_346;
mixer gate_output_15_346(.a(output_16_346), .b(output_16_11), .y(output_15_346));
wire output_1_347, output_1_12, output_0_347;
mixer gate_output_0_347(.a(output_1_347), .b(output_1_12), .y(output_0_347));
wire output_2_347, output_2_12, output_1_347;
mixer gate_output_1_347(.a(output_2_347), .b(output_2_12), .y(output_1_347));
wire output_3_347, output_3_12, output_2_347;
mixer gate_output_2_347(.a(output_3_347), .b(output_3_12), .y(output_2_347));
wire output_4_347, output_4_12, output_3_347;
mixer gate_output_3_347(.a(output_4_347), .b(output_4_12), .y(output_3_347));
wire output_5_347, output_5_12, output_4_347;
mixer gate_output_4_347(.a(output_5_347), .b(output_5_12), .y(output_4_347));
wire output_6_347, output_6_12, output_5_347;
mixer gate_output_5_347(.a(output_6_347), .b(output_6_12), .y(output_5_347));
wire output_7_347, output_7_12, output_6_347;
mixer gate_output_6_347(.a(output_7_347), .b(output_7_12), .y(output_6_347));
wire output_8_347, output_8_12, output_7_347;
mixer gate_output_7_347(.a(output_8_347), .b(output_8_12), .y(output_7_347));
wire output_9_347, output_9_12, output_8_347;
mixer gate_output_8_347(.a(output_9_347), .b(output_9_12), .y(output_8_347));
wire output_10_347, output_10_12, output_9_347;
mixer gate_output_9_347(.a(output_10_347), .b(output_10_12), .y(output_9_347));
wire output_11_347, output_11_12, output_10_347;
mixer gate_output_10_347(.a(output_11_347), .b(output_11_12), .y(output_10_347));
wire output_12_347, output_12_12, output_11_347;
mixer gate_output_11_347(.a(output_12_347), .b(output_12_12), .y(output_11_347));
wire output_13_347, output_13_12, output_12_347;
mixer gate_output_12_347(.a(output_13_347), .b(output_13_12), .y(output_12_347));
wire output_14_347, output_14_12, output_13_347;
mixer gate_output_13_347(.a(output_14_347), .b(output_14_12), .y(output_13_347));
wire output_15_347, output_15_12, output_14_347;
mixer gate_output_14_347(.a(output_15_347), .b(output_15_12), .y(output_14_347));
wire output_16_347, output_16_12, output_15_347;
mixer gate_output_15_347(.a(output_16_347), .b(output_16_12), .y(output_15_347));
wire output_1_348, output_1_13, output_0_348;
mixer gate_output_0_348(.a(output_1_348), .b(output_1_13), .y(output_0_348));
wire output_2_348, output_2_13, output_1_348;
mixer gate_output_1_348(.a(output_2_348), .b(output_2_13), .y(output_1_348));
wire output_3_348, output_3_13, output_2_348;
mixer gate_output_2_348(.a(output_3_348), .b(output_3_13), .y(output_2_348));
wire output_4_348, output_4_13, output_3_348;
mixer gate_output_3_348(.a(output_4_348), .b(output_4_13), .y(output_3_348));
wire output_5_348, output_5_13, output_4_348;
mixer gate_output_4_348(.a(output_5_348), .b(output_5_13), .y(output_4_348));
wire output_6_348, output_6_13, output_5_348;
mixer gate_output_5_348(.a(output_6_348), .b(output_6_13), .y(output_5_348));
wire output_7_348, output_7_13, output_6_348;
mixer gate_output_6_348(.a(output_7_348), .b(output_7_13), .y(output_6_348));
wire output_8_348, output_8_13, output_7_348;
mixer gate_output_7_348(.a(output_8_348), .b(output_8_13), .y(output_7_348));
wire output_9_348, output_9_13, output_8_348;
mixer gate_output_8_348(.a(output_9_348), .b(output_9_13), .y(output_8_348));
wire output_10_348, output_10_13, output_9_348;
mixer gate_output_9_348(.a(output_10_348), .b(output_10_13), .y(output_9_348));
wire output_11_348, output_11_13, output_10_348;
mixer gate_output_10_348(.a(output_11_348), .b(output_11_13), .y(output_10_348));
wire output_12_348, output_12_13, output_11_348;
mixer gate_output_11_348(.a(output_12_348), .b(output_12_13), .y(output_11_348));
wire output_13_348, output_13_13, output_12_348;
mixer gate_output_12_348(.a(output_13_348), .b(output_13_13), .y(output_12_348));
wire output_14_348, output_14_13, output_13_348;
mixer gate_output_13_348(.a(output_14_348), .b(output_14_13), .y(output_13_348));
wire output_15_348, output_15_13, output_14_348;
mixer gate_output_14_348(.a(output_15_348), .b(output_15_13), .y(output_14_348));
wire output_16_348, output_16_13, output_15_348;
mixer gate_output_15_348(.a(output_16_348), .b(output_16_13), .y(output_15_348));
wire output_1_349, output_1_14, output_0_349;
mixer gate_output_0_349(.a(output_1_349), .b(output_1_14), .y(output_0_349));
wire output_2_349, output_2_14, output_1_349;
mixer gate_output_1_349(.a(output_2_349), .b(output_2_14), .y(output_1_349));
wire output_3_349, output_3_14, output_2_349;
mixer gate_output_2_349(.a(output_3_349), .b(output_3_14), .y(output_2_349));
wire output_4_349, output_4_14, output_3_349;
mixer gate_output_3_349(.a(output_4_349), .b(output_4_14), .y(output_3_349));
wire output_5_349, output_5_14, output_4_349;
mixer gate_output_4_349(.a(output_5_349), .b(output_5_14), .y(output_4_349));
wire output_6_349, output_6_14, output_5_349;
mixer gate_output_5_349(.a(output_6_349), .b(output_6_14), .y(output_5_349));
wire output_7_349, output_7_14, output_6_349;
mixer gate_output_6_349(.a(output_7_349), .b(output_7_14), .y(output_6_349));
wire output_8_349, output_8_14, output_7_349;
mixer gate_output_7_349(.a(output_8_349), .b(output_8_14), .y(output_7_349));
wire output_9_349, output_9_14, output_8_349;
mixer gate_output_8_349(.a(output_9_349), .b(output_9_14), .y(output_8_349));
wire output_10_349, output_10_14, output_9_349;
mixer gate_output_9_349(.a(output_10_349), .b(output_10_14), .y(output_9_349));
wire output_11_349, output_11_14, output_10_349;
mixer gate_output_10_349(.a(output_11_349), .b(output_11_14), .y(output_10_349));
wire output_12_349, output_12_14, output_11_349;
mixer gate_output_11_349(.a(output_12_349), .b(output_12_14), .y(output_11_349));
wire output_13_349, output_13_14, output_12_349;
mixer gate_output_12_349(.a(output_13_349), .b(output_13_14), .y(output_12_349));
wire output_14_349, output_14_14, output_13_349;
mixer gate_output_13_349(.a(output_14_349), .b(output_14_14), .y(output_13_349));
wire output_15_349, output_15_14, output_14_349;
mixer gate_output_14_349(.a(output_15_349), .b(output_15_14), .y(output_14_349));
wire output_16_349, output_16_14, output_15_349;
mixer gate_output_15_349(.a(output_16_349), .b(output_16_14), .y(output_15_349));
wire output_1_350, output_1_15, output_0_350;
mixer gate_output_0_350(.a(output_1_350), .b(output_1_15), .y(output_0_350));
wire output_2_350, output_2_15, output_1_350;
mixer gate_output_1_350(.a(output_2_350), .b(output_2_15), .y(output_1_350));
wire output_3_350, output_3_15, output_2_350;
mixer gate_output_2_350(.a(output_3_350), .b(output_3_15), .y(output_2_350));
wire output_4_350, output_4_15, output_3_350;
mixer gate_output_3_350(.a(output_4_350), .b(output_4_15), .y(output_3_350));
wire output_5_350, output_5_15, output_4_350;
mixer gate_output_4_350(.a(output_5_350), .b(output_5_15), .y(output_4_350));
wire output_6_350, output_6_15, output_5_350;
mixer gate_output_5_350(.a(output_6_350), .b(output_6_15), .y(output_5_350));
wire output_7_350, output_7_15, output_6_350;
mixer gate_output_6_350(.a(output_7_350), .b(output_7_15), .y(output_6_350));
wire output_8_350, output_8_15, output_7_350;
mixer gate_output_7_350(.a(output_8_350), .b(output_8_15), .y(output_7_350));
wire output_9_350, output_9_15, output_8_350;
mixer gate_output_8_350(.a(output_9_350), .b(output_9_15), .y(output_8_350));
wire output_10_350, output_10_15, output_9_350;
mixer gate_output_9_350(.a(output_10_350), .b(output_10_15), .y(output_9_350));
wire output_11_350, output_11_15, output_10_350;
mixer gate_output_10_350(.a(output_11_350), .b(output_11_15), .y(output_10_350));
wire output_12_350, output_12_15, output_11_350;
mixer gate_output_11_350(.a(output_12_350), .b(output_12_15), .y(output_11_350));
wire output_13_350, output_13_15, output_12_350;
mixer gate_output_12_350(.a(output_13_350), .b(output_13_15), .y(output_12_350));
wire output_14_350, output_14_15, output_13_350;
mixer gate_output_13_350(.a(output_14_350), .b(output_14_15), .y(output_13_350));
wire output_15_350, output_15_15, output_14_350;
mixer gate_output_14_350(.a(output_15_350), .b(output_15_15), .y(output_14_350));
wire output_16_350, output_16_15, output_15_350;
mixer gate_output_15_350(.a(output_16_350), .b(output_16_15), .y(output_15_350));
wire output_1_351, output_1_0, output_0_351;
mixer gate_output_0_351(.a(output_1_351), .b(output_1_0), .y(output_0_351));
wire output_2_351, output_2_0, output_1_351;
mixer gate_output_1_351(.a(output_2_351), .b(output_2_0), .y(output_1_351));
wire output_3_351, output_3_0, output_2_351;
mixer gate_output_2_351(.a(output_3_351), .b(output_3_0), .y(output_2_351));
wire output_4_351, output_4_0, output_3_351;
mixer gate_output_3_351(.a(output_4_351), .b(output_4_0), .y(output_3_351));
wire output_5_351, output_5_0, output_4_351;
mixer gate_output_4_351(.a(output_5_351), .b(output_5_0), .y(output_4_351));
wire output_6_351, output_6_0, output_5_351;
mixer gate_output_5_351(.a(output_6_351), .b(output_6_0), .y(output_5_351));
wire output_7_351, output_7_0, output_6_351;
mixer gate_output_6_351(.a(output_7_351), .b(output_7_0), .y(output_6_351));
wire output_8_351, output_8_0, output_7_351;
mixer gate_output_7_351(.a(output_8_351), .b(output_8_0), .y(output_7_351));
wire output_9_351, output_9_0, output_8_351;
mixer gate_output_8_351(.a(output_9_351), .b(output_9_0), .y(output_8_351));
wire output_10_351, output_10_0, output_9_351;
mixer gate_output_9_351(.a(output_10_351), .b(output_10_0), .y(output_9_351));
wire output_11_351, output_11_0, output_10_351;
mixer gate_output_10_351(.a(output_11_351), .b(output_11_0), .y(output_10_351));
wire output_12_351, output_12_0, output_11_351;
mixer gate_output_11_351(.a(output_12_351), .b(output_12_0), .y(output_11_351));
wire output_13_351, output_13_0, output_12_351;
mixer gate_output_12_351(.a(output_13_351), .b(output_13_0), .y(output_12_351));
wire output_14_351, output_14_0, output_13_351;
mixer gate_output_13_351(.a(output_14_351), .b(output_14_0), .y(output_13_351));
wire output_15_351, output_15_0, output_14_351;
mixer gate_output_14_351(.a(output_15_351), .b(output_15_0), .y(output_14_351));
wire output_16_351, output_16_0, output_15_351;
mixer gate_output_15_351(.a(output_16_351), .b(output_16_0), .y(output_15_351));
wire output_1_352, output_1_1, output_0_352;
mixer gate_output_0_352(.a(output_1_352), .b(output_1_1), .y(output_0_352));
wire output_2_352, output_2_1, output_1_352;
mixer gate_output_1_352(.a(output_2_352), .b(output_2_1), .y(output_1_352));
wire output_3_352, output_3_1, output_2_352;
mixer gate_output_2_352(.a(output_3_352), .b(output_3_1), .y(output_2_352));
wire output_4_352, output_4_1, output_3_352;
mixer gate_output_3_352(.a(output_4_352), .b(output_4_1), .y(output_3_352));
wire output_5_352, output_5_1, output_4_352;
mixer gate_output_4_352(.a(output_5_352), .b(output_5_1), .y(output_4_352));
wire output_6_352, output_6_1, output_5_352;
mixer gate_output_5_352(.a(output_6_352), .b(output_6_1), .y(output_5_352));
wire output_7_352, output_7_1, output_6_352;
mixer gate_output_6_352(.a(output_7_352), .b(output_7_1), .y(output_6_352));
wire output_8_352, output_8_1, output_7_352;
mixer gate_output_7_352(.a(output_8_352), .b(output_8_1), .y(output_7_352));
wire output_9_352, output_9_1, output_8_352;
mixer gate_output_8_352(.a(output_9_352), .b(output_9_1), .y(output_8_352));
wire output_10_352, output_10_1, output_9_352;
mixer gate_output_9_352(.a(output_10_352), .b(output_10_1), .y(output_9_352));
wire output_11_352, output_11_1, output_10_352;
mixer gate_output_10_352(.a(output_11_352), .b(output_11_1), .y(output_10_352));
wire output_12_352, output_12_1, output_11_352;
mixer gate_output_11_352(.a(output_12_352), .b(output_12_1), .y(output_11_352));
wire output_13_352, output_13_1, output_12_352;
mixer gate_output_12_352(.a(output_13_352), .b(output_13_1), .y(output_12_352));
wire output_14_352, output_14_1, output_13_352;
mixer gate_output_13_352(.a(output_14_352), .b(output_14_1), .y(output_13_352));
wire output_15_352, output_15_1, output_14_352;
mixer gate_output_14_352(.a(output_15_352), .b(output_15_1), .y(output_14_352));
wire output_16_352, output_16_1, output_15_352;
mixer gate_output_15_352(.a(output_16_352), .b(output_16_1), .y(output_15_352));
wire output_1_353, output_1_2, output_0_353;
mixer gate_output_0_353(.a(output_1_353), .b(output_1_2), .y(output_0_353));
wire output_2_353, output_2_2, output_1_353;
mixer gate_output_1_353(.a(output_2_353), .b(output_2_2), .y(output_1_353));
wire output_3_353, output_3_2, output_2_353;
mixer gate_output_2_353(.a(output_3_353), .b(output_3_2), .y(output_2_353));
wire output_4_353, output_4_2, output_3_353;
mixer gate_output_3_353(.a(output_4_353), .b(output_4_2), .y(output_3_353));
wire output_5_353, output_5_2, output_4_353;
mixer gate_output_4_353(.a(output_5_353), .b(output_5_2), .y(output_4_353));
wire output_6_353, output_6_2, output_5_353;
mixer gate_output_5_353(.a(output_6_353), .b(output_6_2), .y(output_5_353));
wire output_7_353, output_7_2, output_6_353;
mixer gate_output_6_353(.a(output_7_353), .b(output_7_2), .y(output_6_353));
wire output_8_353, output_8_2, output_7_353;
mixer gate_output_7_353(.a(output_8_353), .b(output_8_2), .y(output_7_353));
wire output_9_353, output_9_2, output_8_353;
mixer gate_output_8_353(.a(output_9_353), .b(output_9_2), .y(output_8_353));
wire output_10_353, output_10_2, output_9_353;
mixer gate_output_9_353(.a(output_10_353), .b(output_10_2), .y(output_9_353));
wire output_11_353, output_11_2, output_10_353;
mixer gate_output_10_353(.a(output_11_353), .b(output_11_2), .y(output_10_353));
wire output_12_353, output_12_2, output_11_353;
mixer gate_output_11_353(.a(output_12_353), .b(output_12_2), .y(output_11_353));
wire output_13_353, output_13_2, output_12_353;
mixer gate_output_12_353(.a(output_13_353), .b(output_13_2), .y(output_12_353));
wire output_14_353, output_14_2, output_13_353;
mixer gate_output_13_353(.a(output_14_353), .b(output_14_2), .y(output_13_353));
wire output_15_353, output_15_2, output_14_353;
mixer gate_output_14_353(.a(output_15_353), .b(output_15_2), .y(output_14_353));
wire output_16_353, output_16_2, output_15_353;
mixer gate_output_15_353(.a(output_16_353), .b(output_16_2), .y(output_15_353));
wire output_1_354, output_1_3, output_0_354;
mixer gate_output_0_354(.a(output_1_354), .b(output_1_3), .y(output_0_354));
wire output_2_354, output_2_3, output_1_354;
mixer gate_output_1_354(.a(output_2_354), .b(output_2_3), .y(output_1_354));
wire output_3_354, output_3_3, output_2_354;
mixer gate_output_2_354(.a(output_3_354), .b(output_3_3), .y(output_2_354));
wire output_4_354, output_4_3, output_3_354;
mixer gate_output_3_354(.a(output_4_354), .b(output_4_3), .y(output_3_354));
wire output_5_354, output_5_3, output_4_354;
mixer gate_output_4_354(.a(output_5_354), .b(output_5_3), .y(output_4_354));
wire output_6_354, output_6_3, output_5_354;
mixer gate_output_5_354(.a(output_6_354), .b(output_6_3), .y(output_5_354));
wire output_7_354, output_7_3, output_6_354;
mixer gate_output_6_354(.a(output_7_354), .b(output_7_3), .y(output_6_354));
wire output_8_354, output_8_3, output_7_354;
mixer gate_output_7_354(.a(output_8_354), .b(output_8_3), .y(output_7_354));
wire output_9_354, output_9_3, output_8_354;
mixer gate_output_8_354(.a(output_9_354), .b(output_9_3), .y(output_8_354));
wire output_10_354, output_10_3, output_9_354;
mixer gate_output_9_354(.a(output_10_354), .b(output_10_3), .y(output_9_354));
wire output_11_354, output_11_3, output_10_354;
mixer gate_output_10_354(.a(output_11_354), .b(output_11_3), .y(output_10_354));
wire output_12_354, output_12_3, output_11_354;
mixer gate_output_11_354(.a(output_12_354), .b(output_12_3), .y(output_11_354));
wire output_13_354, output_13_3, output_12_354;
mixer gate_output_12_354(.a(output_13_354), .b(output_13_3), .y(output_12_354));
wire output_14_354, output_14_3, output_13_354;
mixer gate_output_13_354(.a(output_14_354), .b(output_14_3), .y(output_13_354));
wire output_15_354, output_15_3, output_14_354;
mixer gate_output_14_354(.a(output_15_354), .b(output_15_3), .y(output_14_354));
wire output_16_354, output_16_3, output_15_354;
mixer gate_output_15_354(.a(output_16_354), .b(output_16_3), .y(output_15_354));
wire output_1_355, output_1_4, output_0_355;
mixer gate_output_0_355(.a(output_1_355), .b(output_1_4), .y(output_0_355));
wire output_2_355, output_2_4, output_1_355;
mixer gate_output_1_355(.a(output_2_355), .b(output_2_4), .y(output_1_355));
wire output_3_355, output_3_4, output_2_355;
mixer gate_output_2_355(.a(output_3_355), .b(output_3_4), .y(output_2_355));
wire output_4_355, output_4_4, output_3_355;
mixer gate_output_3_355(.a(output_4_355), .b(output_4_4), .y(output_3_355));
wire output_5_355, output_5_4, output_4_355;
mixer gate_output_4_355(.a(output_5_355), .b(output_5_4), .y(output_4_355));
wire output_6_355, output_6_4, output_5_355;
mixer gate_output_5_355(.a(output_6_355), .b(output_6_4), .y(output_5_355));
wire output_7_355, output_7_4, output_6_355;
mixer gate_output_6_355(.a(output_7_355), .b(output_7_4), .y(output_6_355));
wire output_8_355, output_8_4, output_7_355;
mixer gate_output_7_355(.a(output_8_355), .b(output_8_4), .y(output_7_355));
wire output_9_355, output_9_4, output_8_355;
mixer gate_output_8_355(.a(output_9_355), .b(output_9_4), .y(output_8_355));
wire output_10_355, output_10_4, output_9_355;
mixer gate_output_9_355(.a(output_10_355), .b(output_10_4), .y(output_9_355));
wire output_11_355, output_11_4, output_10_355;
mixer gate_output_10_355(.a(output_11_355), .b(output_11_4), .y(output_10_355));
wire output_12_355, output_12_4, output_11_355;
mixer gate_output_11_355(.a(output_12_355), .b(output_12_4), .y(output_11_355));
wire output_13_355, output_13_4, output_12_355;
mixer gate_output_12_355(.a(output_13_355), .b(output_13_4), .y(output_12_355));
wire output_14_355, output_14_4, output_13_355;
mixer gate_output_13_355(.a(output_14_355), .b(output_14_4), .y(output_13_355));
wire output_15_355, output_15_4, output_14_355;
mixer gate_output_14_355(.a(output_15_355), .b(output_15_4), .y(output_14_355));
wire output_16_355, output_16_4, output_15_355;
mixer gate_output_15_355(.a(output_16_355), .b(output_16_4), .y(output_15_355));
wire output_1_356, output_1_5, output_0_356;
mixer gate_output_0_356(.a(output_1_356), .b(output_1_5), .y(output_0_356));
wire output_2_356, output_2_5, output_1_356;
mixer gate_output_1_356(.a(output_2_356), .b(output_2_5), .y(output_1_356));
wire output_3_356, output_3_5, output_2_356;
mixer gate_output_2_356(.a(output_3_356), .b(output_3_5), .y(output_2_356));
wire output_4_356, output_4_5, output_3_356;
mixer gate_output_3_356(.a(output_4_356), .b(output_4_5), .y(output_3_356));
wire output_5_356, output_5_5, output_4_356;
mixer gate_output_4_356(.a(output_5_356), .b(output_5_5), .y(output_4_356));
wire output_6_356, output_6_5, output_5_356;
mixer gate_output_5_356(.a(output_6_356), .b(output_6_5), .y(output_5_356));
wire output_7_356, output_7_5, output_6_356;
mixer gate_output_6_356(.a(output_7_356), .b(output_7_5), .y(output_6_356));
wire output_8_356, output_8_5, output_7_356;
mixer gate_output_7_356(.a(output_8_356), .b(output_8_5), .y(output_7_356));
wire output_9_356, output_9_5, output_8_356;
mixer gate_output_8_356(.a(output_9_356), .b(output_9_5), .y(output_8_356));
wire output_10_356, output_10_5, output_9_356;
mixer gate_output_9_356(.a(output_10_356), .b(output_10_5), .y(output_9_356));
wire output_11_356, output_11_5, output_10_356;
mixer gate_output_10_356(.a(output_11_356), .b(output_11_5), .y(output_10_356));
wire output_12_356, output_12_5, output_11_356;
mixer gate_output_11_356(.a(output_12_356), .b(output_12_5), .y(output_11_356));
wire output_13_356, output_13_5, output_12_356;
mixer gate_output_12_356(.a(output_13_356), .b(output_13_5), .y(output_12_356));
wire output_14_356, output_14_5, output_13_356;
mixer gate_output_13_356(.a(output_14_356), .b(output_14_5), .y(output_13_356));
wire output_15_356, output_15_5, output_14_356;
mixer gate_output_14_356(.a(output_15_356), .b(output_15_5), .y(output_14_356));
wire output_16_356, output_16_5, output_15_356;
mixer gate_output_15_356(.a(output_16_356), .b(output_16_5), .y(output_15_356));
wire output_1_357, output_1_6, output_0_357;
mixer gate_output_0_357(.a(output_1_357), .b(output_1_6), .y(output_0_357));
wire output_2_357, output_2_6, output_1_357;
mixer gate_output_1_357(.a(output_2_357), .b(output_2_6), .y(output_1_357));
wire output_3_357, output_3_6, output_2_357;
mixer gate_output_2_357(.a(output_3_357), .b(output_3_6), .y(output_2_357));
wire output_4_357, output_4_6, output_3_357;
mixer gate_output_3_357(.a(output_4_357), .b(output_4_6), .y(output_3_357));
wire output_5_357, output_5_6, output_4_357;
mixer gate_output_4_357(.a(output_5_357), .b(output_5_6), .y(output_4_357));
wire output_6_357, output_6_6, output_5_357;
mixer gate_output_5_357(.a(output_6_357), .b(output_6_6), .y(output_5_357));
wire output_7_357, output_7_6, output_6_357;
mixer gate_output_6_357(.a(output_7_357), .b(output_7_6), .y(output_6_357));
wire output_8_357, output_8_6, output_7_357;
mixer gate_output_7_357(.a(output_8_357), .b(output_8_6), .y(output_7_357));
wire output_9_357, output_9_6, output_8_357;
mixer gate_output_8_357(.a(output_9_357), .b(output_9_6), .y(output_8_357));
wire output_10_357, output_10_6, output_9_357;
mixer gate_output_9_357(.a(output_10_357), .b(output_10_6), .y(output_9_357));
wire output_11_357, output_11_6, output_10_357;
mixer gate_output_10_357(.a(output_11_357), .b(output_11_6), .y(output_10_357));
wire output_12_357, output_12_6, output_11_357;
mixer gate_output_11_357(.a(output_12_357), .b(output_12_6), .y(output_11_357));
wire output_13_357, output_13_6, output_12_357;
mixer gate_output_12_357(.a(output_13_357), .b(output_13_6), .y(output_12_357));
wire output_14_357, output_14_6, output_13_357;
mixer gate_output_13_357(.a(output_14_357), .b(output_14_6), .y(output_13_357));
wire output_15_357, output_15_6, output_14_357;
mixer gate_output_14_357(.a(output_15_357), .b(output_15_6), .y(output_14_357));
wire output_16_357, output_16_6, output_15_357;
mixer gate_output_15_357(.a(output_16_357), .b(output_16_6), .y(output_15_357));
wire output_1_358, output_1_7, output_0_358;
mixer gate_output_0_358(.a(output_1_358), .b(output_1_7), .y(output_0_358));
wire output_2_358, output_2_7, output_1_358;
mixer gate_output_1_358(.a(output_2_358), .b(output_2_7), .y(output_1_358));
wire output_3_358, output_3_7, output_2_358;
mixer gate_output_2_358(.a(output_3_358), .b(output_3_7), .y(output_2_358));
wire output_4_358, output_4_7, output_3_358;
mixer gate_output_3_358(.a(output_4_358), .b(output_4_7), .y(output_3_358));
wire output_5_358, output_5_7, output_4_358;
mixer gate_output_4_358(.a(output_5_358), .b(output_5_7), .y(output_4_358));
wire output_6_358, output_6_7, output_5_358;
mixer gate_output_5_358(.a(output_6_358), .b(output_6_7), .y(output_5_358));
wire output_7_358, output_7_7, output_6_358;
mixer gate_output_6_358(.a(output_7_358), .b(output_7_7), .y(output_6_358));
wire output_8_358, output_8_7, output_7_358;
mixer gate_output_7_358(.a(output_8_358), .b(output_8_7), .y(output_7_358));
wire output_9_358, output_9_7, output_8_358;
mixer gate_output_8_358(.a(output_9_358), .b(output_9_7), .y(output_8_358));
wire output_10_358, output_10_7, output_9_358;
mixer gate_output_9_358(.a(output_10_358), .b(output_10_7), .y(output_9_358));
wire output_11_358, output_11_7, output_10_358;
mixer gate_output_10_358(.a(output_11_358), .b(output_11_7), .y(output_10_358));
wire output_12_358, output_12_7, output_11_358;
mixer gate_output_11_358(.a(output_12_358), .b(output_12_7), .y(output_11_358));
wire output_13_358, output_13_7, output_12_358;
mixer gate_output_12_358(.a(output_13_358), .b(output_13_7), .y(output_12_358));
wire output_14_358, output_14_7, output_13_358;
mixer gate_output_13_358(.a(output_14_358), .b(output_14_7), .y(output_13_358));
wire output_15_358, output_15_7, output_14_358;
mixer gate_output_14_358(.a(output_15_358), .b(output_15_7), .y(output_14_358));
wire output_16_358, output_16_7, output_15_358;
mixer gate_output_15_358(.a(output_16_358), .b(output_16_7), .y(output_15_358));
wire output_1_359, output_1_8, output_0_359;
mixer gate_output_0_359(.a(output_1_359), .b(output_1_8), .y(output_0_359));
wire output_2_359, output_2_8, output_1_359;
mixer gate_output_1_359(.a(output_2_359), .b(output_2_8), .y(output_1_359));
wire output_3_359, output_3_8, output_2_359;
mixer gate_output_2_359(.a(output_3_359), .b(output_3_8), .y(output_2_359));
wire output_4_359, output_4_8, output_3_359;
mixer gate_output_3_359(.a(output_4_359), .b(output_4_8), .y(output_3_359));
wire output_5_359, output_5_8, output_4_359;
mixer gate_output_4_359(.a(output_5_359), .b(output_5_8), .y(output_4_359));
wire output_6_359, output_6_8, output_5_359;
mixer gate_output_5_359(.a(output_6_359), .b(output_6_8), .y(output_5_359));
wire output_7_359, output_7_8, output_6_359;
mixer gate_output_6_359(.a(output_7_359), .b(output_7_8), .y(output_6_359));
wire output_8_359, output_8_8, output_7_359;
mixer gate_output_7_359(.a(output_8_359), .b(output_8_8), .y(output_7_359));
wire output_9_359, output_9_8, output_8_359;
mixer gate_output_8_359(.a(output_9_359), .b(output_9_8), .y(output_8_359));
wire output_10_359, output_10_8, output_9_359;
mixer gate_output_9_359(.a(output_10_359), .b(output_10_8), .y(output_9_359));
wire output_11_359, output_11_8, output_10_359;
mixer gate_output_10_359(.a(output_11_359), .b(output_11_8), .y(output_10_359));
wire output_12_359, output_12_8, output_11_359;
mixer gate_output_11_359(.a(output_12_359), .b(output_12_8), .y(output_11_359));
wire output_13_359, output_13_8, output_12_359;
mixer gate_output_12_359(.a(output_13_359), .b(output_13_8), .y(output_12_359));
wire output_14_359, output_14_8, output_13_359;
mixer gate_output_13_359(.a(output_14_359), .b(output_14_8), .y(output_13_359));
wire output_15_359, output_15_8, output_14_359;
mixer gate_output_14_359(.a(output_15_359), .b(output_15_8), .y(output_14_359));
wire output_16_359, output_16_8, output_15_359;
mixer gate_output_15_359(.a(output_16_359), .b(output_16_8), .y(output_15_359));
wire output_1_360, output_1_9, output_0_360;
mixer gate_output_0_360(.a(output_1_360), .b(output_1_9), .y(output_0_360));
wire output_2_360, output_2_9, output_1_360;
mixer gate_output_1_360(.a(output_2_360), .b(output_2_9), .y(output_1_360));
wire output_3_360, output_3_9, output_2_360;
mixer gate_output_2_360(.a(output_3_360), .b(output_3_9), .y(output_2_360));
wire output_4_360, output_4_9, output_3_360;
mixer gate_output_3_360(.a(output_4_360), .b(output_4_9), .y(output_3_360));
wire output_5_360, output_5_9, output_4_360;
mixer gate_output_4_360(.a(output_5_360), .b(output_5_9), .y(output_4_360));
wire output_6_360, output_6_9, output_5_360;
mixer gate_output_5_360(.a(output_6_360), .b(output_6_9), .y(output_5_360));
wire output_7_360, output_7_9, output_6_360;
mixer gate_output_6_360(.a(output_7_360), .b(output_7_9), .y(output_6_360));
wire output_8_360, output_8_9, output_7_360;
mixer gate_output_7_360(.a(output_8_360), .b(output_8_9), .y(output_7_360));
wire output_9_360, output_9_9, output_8_360;
mixer gate_output_8_360(.a(output_9_360), .b(output_9_9), .y(output_8_360));
wire output_10_360, output_10_9, output_9_360;
mixer gate_output_9_360(.a(output_10_360), .b(output_10_9), .y(output_9_360));
wire output_11_360, output_11_9, output_10_360;
mixer gate_output_10_360(.a(output_11_360), .b(output_11_9), .y(output_10_360));
wire output_12_360, output_12_9, output_11_360;
mixer gate_output_11_360(.a(output_12_360), .b(output_12_9), .y(output_11_360));
wire output_13_360, output_13_9, output_12_360;
mixer gate_output_12_360(.a(output_13_360), .b(output_13_9), .y(output_12_360));
wire output_14_360, output_14_9, output_13_360;
mixer gate_output_13_360(.a(output_14_360), .b(output_14_9), .y(output_13_360));
wire output_15_360, output_15_9, output_14_360;
mixer gate_output_14_360(.a(output_15_360), .b(output_15_9), .y(output_14_360));
wire output_16_360, output_16_9, output_15_360;
mixer gate_output_15_360(.a(output_16_360), .b(output_16_9), .y(output_15_360));
wire output_1_361, output_1_10, output_0_361;
mixer gate_output_0_361(.a(output_1_361), .b(output_1_10), .y(output_0_361));
wire output_2_361, output_2_10, output_1_361;
mixer gate_output_1_361(.a(output_2_361), .b(output_2_10), .y(output_1_361));
wire output_3_361, output_3_10, output_2_361;
mixer gate_output_2_361(.a(output_3_361), .b(output_3_10), .y(output_2_361));
wire output_4_361, output_4_10, output_3_361;
mixer gate_output_3_361(.a(output_4_361), .b(output_4_10), .y(output_3_361));
wire output_5_361, output_5_10, output_4_361;
mixer gate_output_4_361(.a(output_5_361), .b(output_5_10), .y(output_4_361));
wire output_6_361, output_6_10, output_5_361;
mixer gate_output_5_361(.a(output_6_361), .b(output_6_10), .y(output_5_361));
wire output_7_361, output_7_10, output_6_361;
mixer gate_output_6_361(.a(output_7_361), .b(output_7_10), .y(output_6_361));
wire output_8_361, output_8_10, output_7_361;
mixer gate_output_7_361(.a(output_8_361), .b(output_8_10), .y(output_7_361));
wire output_9_361, output_9_10, output_8_361;
mixer gate_output_8_361(.a(output_9_361), .b(output_9_10), .y(output_8_361));
wire output_10_361, output_10_10, output_9_361;
mixer gate_output_9_361(.a(output_10_361), .b(output_10_10), .y(output_9_361));
wire output_11_361, output_11_10, output_10_361;
mixer gate_output_10_361(.a(output_11_361), .b(output_11_10), .y(output_10_361));
wire output_12_361, output_12_10, output_11_361;
mixer gate_output_11_361(.a(output_12_361), .b(output_12_10), .y(output_11_361));
wire output_13_361, output_13_10, output_12_361;
mixer gate_output_12_361(.a(output_13_361), .b(output_13_10), .y(output_12_361));
wire output_14_361, output_14_10, output_13_361;
mixer gate_output_13_361(.a(output_14_361), .b(output_14_10), .y(output_13_361));
wire output_15_361, output_15_10, output_14_361;
mixer gate_output_14_361(.a(output_15_361), .b(output_15_10), .y(output_14_361));
wire output_16_361, output_16_10, output_15_361;
mixer gate_output_15_361(.a(output_16_361), .b(output_16_10), .y(output_15_361));
wire output_1_362, output_1_11, output_0_362;
mixer gate_output_0_362(.a(output_1_362), .b(output_1_11), .y(output_0_362));
wire output_2_362, output_2_11, output_1_362;
mixer gate_output_1_362(.a(output_2_362), .b(output_2_11), .y(output_1_362));
wire output_3_362, output_3_11, output_2_362;
mixer gate_output_2_362(.a(output_3_362), .b(output_3_11), .y(output_2_362));
wire output_4_362, output_4_11, output_3_362;
mixer gate_output_3_362(.a(output_4_362), .b(output_4_11), .y(output_3_362));
wire output_5_362, output_5_11, output_4_362;
mixer gate_output_4_362(.a(output_5_362), .b(output_5_11), .y(output_4_362));
wire output_6_362, output_6_11, output_5_362;
mixer gate_output_5_362(.a(output_6_362), .b(output_6_11), .y(output_5_362));
wire output_7_362, output_7_11, output_6_362;
mixer gate_output_6_362(.a(output_7_362), .b(output_7_11), .y(output_6_362));
wire output_8_362, output_8_11, output_7_362;
mixer gate_output_7_362(.a(output_8_362), .b(output_8_11), .y(output_7_362));
wire output_9_362, output_9_11, output_8_362;
mixer gate_output_8_362(.a(output_9_362), .b(output_9_11), .y(output_8_362));
wire output_10_362, output_10_11, output_9_362;
mixer gate_output_9_362(.a(output_10_362), .b(output_10_11), .y(output_9_362));
wire output_11_362, output_11_11, output_10_362;
mixer gate_output_10_362(.a(output_11_362), .b(output_11_11), .y(output_10_362));
wire output_12_362, output_12_11, output_11_362;
mixer gate_output_11_362(.a(output_12_362), .b(output_12_11), .y(output_11_362));
wire output_13_362, output_13_11, output_12_362;
mixer gate_output_12_362(.a(output_13_362), .b(output_13_11), .y(output_12_362));
wire output_14_362, output_14_11, output_13_362;
mixer gate_output_13_362(.a(output_14_362), .b(output_14_11), .y(output_13_362));
wire output_15_362, output_15_11, output_14_362;
mixer gate_output_14_362(.a(output_15_362), .b(output_15_11), .y(output_14_362));
wire output_16_362, output_16_11, output_15_362;
mixer gate_output_15_362(.a(output_16_362), .b(output_16_11), .y(output_15_362));
wire output_1_363, output_1_12, output_0_363;
mixer gate_output_0_363(.a(output_1_363), .b(output_1_12), .y(output_0_363));
wire output_2_363, output_2_12, output_1_363;
mixer gate_output_1_363(.a(output_2_363), .b(output_2_12), .y(output_1_363));
wire output_3_363, output_3_12, output_2_363;
mixer gate_output_2_363(.a(output_3_363), .b(output_3_12), .y(output_2_363));
wire output_4_363, output_4_12, output_3_363;
mixer gate_output_3_363(.a(output_4_363), .b(output_4_12), .y(output_3_363));
wire output_5_363, output_5_12, output_4_363;
mixer gate_output_4_363(.a(output_5_363), .b(output_5_12), .y(output_4_363));
wire output_6_363, output_6_12, output_5_363;
mixer gate_output_5_363(.a(output_6_363), .b(output_6_12), .y(output_5_363));
wire output_7_363, output_7_12, output_6_363;
mixer gate_output_6_363(.a(output_7_363), .b(output_7_12), .y(output_6_363));
wire output_8_363, output_8_12, output_7_363;
mixer gate_output_7_363(.a(output_8_363), .b(output_8_12), .y(output_7_363));
wire output_9_363, output_9_12, output_8_363;
mixer gate_output_8_363(.a(output_9_363), .b(output_9_12), .y(output_8_363));
wire output_10_363, output_10_12, output_9_363;
mixer gate_output_9_363(.a(output_10_363), .b(output_10_12), .y(output_9_363));
wire output_11_363, output_11_12, output_10_363;
mixer gate_output_10_363(.a(output_11_363), .b(output_11_12), .y(output_10_363));
wire output_12_363, output_12_12, output_11_363;
mixer gate_output_11_363(.a(output_12_363), .b(output_12_12), .y(output_11_363));
wire output_13_363, output_13_12, output_12_363;
mixer gate_output_12_363(.a(output_13_363), .b(output_13_12), .y(output_12_363));
wire output_14_363, output_14_12, output_13_363;
mixer gate_output_13_363(.a(output_14_363), .b(output_14_12), .y(output_13_363));
wire output_15_363, output_15_12, output_14_363;
mixer gate_output_14_363(.a(output_15_363), .b(output_15_12), .y(output_14_363));
wire output_16_363, output_16_12, output_15_363;
mixer gate_output_15_363(.a(output_16_363), .b(output_16_12), .y(output_15_363));
wire output_1_364, output_1_13, output_0_364;
mixer gate_output_0_364(.a(output_1_364), .b(output_1_13), .y(output_0_364));
wire output_2_364, output_2_13, output_1_364;
mixer gate_output_1_364(.a(output_2_364), .b(output_2_13), .y(output_1_364));
wire output_3_364, output_3_13, output_2_364;
mixer gate_output_2_364(.a(output_3_364), .b(output_3_13), .y(output_2_364));
wire output_4_364, output_4_13, output_3_364;
mixer gate_output_3_364(.a(output_4_364), .b(output_4_13), .y(output_3_364));
wire output_5_364, output_5_13, output_4_364;
mixer gate_output_4_364(.a(output_5_364), .b(output_5_13), .y(output_4_364));
wire output_6_364, output_6_13, output_5_364;
mixer gate_output_5_364(.a(output_6_364), .b(output_6_13), .y(output_5_364));
wire output_7_364, output_7_13, output_6_364;
mixer gate_output_6_364(.a(output_7_364), .b(output_7_13), .y(output_6_364));
wire output_8_364, output_8_13, output_7_364;
mixer gate_output_7_364(.a(output_8_364), .b(output_8_13), .y(output_7_364));
wire output_9_364, output_9_13, output_8_364;
mixer gate_output_8_364(.a(output_9_364), .b(output_9_13), .y(output_8_364));
wire output_10_364, output_10_13, output_9_364;
mixer gate_output_9_364(.a(output_10_364), .b(output_10_13), .y(output_9_364));
wire output_11_364, output_11_13, output_10_364;
mixer gate_output_10_364(.a(output_11_364), .b(output_11_13), .y(output_10_364));
wire output_12_364, output_12_13, output_11_364;
mixer gate_output_11_364(.a(output_12_364), .b(output_12_13), .y(output_11_364));
wire output_13_364, output_13_13, output_12_364;
mixer gate_output_12_364(.a(output_13_364), .b(output_13_13), .y(output_12_364));
wire output_14_364, output_14_13, output_13_364;
mixer gate_output_13_364(.a(output_14_364), .b(output_14_13), .y(output_13_364));
wire output_15_364, output_15_13, output_14_364;
mixer gate_output_14_364(.a(output_15_364), .b(output_15_13), .y(output_14_364));
wire output_16_364, output_16_13, output_15_364;
mixer gate_output_15_364(.a(output_16_364), .b(output_16_13), .y(output_15_364));
wire output_1_365, output_1_14, output_0_365;
mixer gate_output_0_365(.a(output_1_365), .b(output_1_14), .y(output_0_365));
wire output_2_365, output_2_14, output_1_365;
mixer gate_output_1_365(.a(output_2_365), .b(output_2_14), .y(output_1_365));
wire output_3_365, output_3_14, output_2_365;
mixer gate_output_2_365(.a(output_3_365), .b(output_3_14), .y(output_2_365));
wire output_4_365, output_4_14, output_3_365;
mixer gate_output_3_365(.a(output_4_365), .b(output_4_14), .y(output_3_365));
wire output_5_365, output_5_14, output_4_365;
mixer gate_output_4_365(.a(output_5_365), .b(output_5_14), .y(output_4_365));
wire output_6_365, output_6_14, output_5_365;
mixer gate_output_5_365(.a(output_6_365), .b(output_6_14), .y(output_5_365));
wire output_7_365, output_7_14, output_6_365;
mixer gate_output_6_365(.a(output_7_365), .b(output_7_14), .y(output_6_365));
wire output_8_365, output_8_14, output_7_365;
mixer gate_output_7_365(.a(output_8_365), .b(output_8_14), .y(output_7_365));
wire output_9_365, output_9_14, output_8_365;
mixer gate_output_8_365(.a(output_9_365), .b(output_9_14), .y(output_8_365));
wire output_10_365, output_10_14, output_9_365;
mixer gate_output_9_365(.a(output_10_365), .b(output_10_14), .y(output_9_365));
wire output_11_365, output_11_14, output_10_365;
mixer gate_output_10_365(.a(output_11_365), .b(output_11_14), .y(output_10_365));
wire output_12_365, output_12_14, output_11_365;
mixer gate_output_11_365(.a(output_12_365), .b(output_12_14), .y(output_11_365));
wire output_13_365, output_13_14, output_12_365;
mixer gate_output_12_365(.a(output_13_365), .b(output_13_14), .y(output_12_365));
wire output_14_365, output_14_14, output_13_365;
mixer gate_output_13_365(.a(output_14_365), .b(output_14_14), .y(output_13_365));
wire output_15_365, output_15_14, output_14_365;
mixer gate_output_14_365(.a(output_15_365), .b(output_15_14), .y(output_14_365));
wire output_16_365, output_16_14, output_15_365;
mixer gate_output_15_365(.a(output_16_365), .b(output_16_14), .y(output_15_365));
wire output_1_366, output_1_15, output_0_366;
mixer gate_output_0_366(.a(output_1_366), .b(output_1_15), .y(output_0_366));
wire output_2_366, output_2_15, output_1_366;
mixer gate_output_1_366(.a(output_2_366), .b(output_2_15), .y(output_1_366));
wire output_3_366, output_3_15, output_2_366;
mixer gate_output_2_366(.a(output_3_366), .b(output_3_15), .y(output_2_366));
wire output_4_366, output_4_15, output_3_366;
mixer gate_output_3_366(.a(output_4_366), .b(output_4_15), .y(output_3_366));
wire output_5_366, output_5_15, output_4_366;
mixer gate_output_4_366(.a(output_5_366), .b(output_5_15), .y(output_4_366));
wire output_6_366, output_6_15, output_5_366;
mixer gate_output_5_366(.a(output_6_366), .b(output_6_15), .y(output_5_366));
wire output_7_366, output_7_15, output_6_366;
mixer gate_output_6_366(.a(output_7_366), .b(output_7_15), .y(output_6_366));
wire output_8_366, output_8_15, output_7_366;
mixer gate_output_7_366(.a(output_8_366), .b(output_8_15), .y(output_7_366));
wire output_9_366, output_9_15, output_8_366;
mixer gate_output_8_366(.a(output_9_366), .b(output_9_15), .y(output_8_366));
wire output_10_366, output_10_15, output_9_366;
mixer gate_output_9_366(.a(output_10_366), .b(output_10_15), .y(output_9_366));
wire output_11_366, output_11_15, output_10_366;
mixer gate_output_10_366(.a(output_11_366), .b(output_11_15), .y(output_10_366));
wire output_12_366, output_12_15, output_11_366;
mixer gate_output_11_366(.a(output_12_366), .b(output_12_15), .y(output_11_366));
wire output_13_366, output_13_15, output_12_366;
mixer gate_output_12_366(.a(output_13_366), .b(output_13_15), .y(output_12_366));
wire output_14_366, output_14_15, output_13_366;
mixer gate_output_13_366(.a(output_14_366), .b(output_14_15), .y(output_13_366));
wire output_15_366, output_15_15, output_14_366;
mixer gate_output_14_366(.a(output_15_366), .b(output_15_15), .y(output_14_366));
wire output_16_366, output_16_15, output_15_366;
mixer gate_output_15_366(.a(output_16_366), .b(output_16_15), .y(output_15_366));
wire output_1_367, output_1_0, output_0_367;
mixer gate_output_0_367(.a(output_1_367), .b(output_1_0), .y(output_0_367));
wire output_2_367, output_2_0, output_1_367;
mixer gate_output_1_367(.a(output_2_367), .b(output_2_0), .y(output_1_367));
wire output_3_367, output_3_0, output_2_367;
mixer gate_output_2_367(.a(output_3_367), .b(output_3_0), .y(output_2_367));
wire output_4_367, output_4_0, output_3_367;
mixer gate_output_3_367(.a(output_4_367), .b(output_4_0), .y(output_3_367));
wire output_5_367, output_5_0, output_4_367;
mixer gate_output_4_367(.a(output_5_367), .b(output_5_0), .y(output_4_367));
wire output_6_367, output_6_0, output_5_367;
mixer gate_output_5_367(.a(output_6_367), .b(output_6_0), .y(output_5_367));
wire output_7_367, output_7_0, output_6_367;
mixer gate_output_6_367(.a(output_7_367), .b(output_7_0), .y(output_6_367));
wire output_8_367, output_8_0, output_7_367;
mixer gate_output_7_367(.a(output_8_367), .b(output_8_0), .y(output_7_367));
wire output_9_367, output_9_0, output_8_367;
mixer gate_output_8_367(.a(output_9_367), .b(output_9_0), .y(output_8_367));
wire output_10_367, output_10_0, output_9_367;
mixer gate_output_9_367(.a(output_10_367), .b(output_10_0), .y(output_9_367));
wire output_11_367, output_11_0, output_10_367;
mixer gate_output_10_367(.a(output_11_367), .b(output_11_0), .y(output_10_367));
wire output_12_367, output_12_0, output_11_367;
mixer gate_output_11_367(.a(output_12_367), .b(output_12_0), .y(output_11_367));
wire output_13_367, output_13_0, output_12_367;
mixer gate_output_12_367(.a(output_13_367), .b(output_13_0), .y(output_12_367));
wire output_14_367, output_14_0, output_13_367;
mixer gate_output_13_367(.a(output_14_367), .b(output_14_0), .y(output_13_367));
wire output_15_367, output_15_0, output_14_367;
mixer gate_output_14_367(.a(output_15_367), .b(output_15_0), .y(output_14_367));
wire output_16_367, output_16_0, output_15_367;
mixer gate_output_15_367(.a(output_16_367), .b(output_16_0), .y(output_15_367));
wire output_1_368, output_1_1, output_0_368;
mixer gate_output_0_368(.a(output_1_368), .b(output_1_1), .y(output_0_368));
wire output_2_368, output_2_1, output_1_368;
mixer gate_output_1_368(.a(output_2_368), .b(output_2_1), .y(output_1_368));
wire output_3_368, output_3_1, output_2_368;
mixer gate_output_2_368(.a(output_3_368), .b(output_3_1), .y(output_2_368));
wire output_4_368, output_4_1, output_3_368;
mixer gate_output_3_368(.a(output_4_368), .b(output_4_1), .y(output_3_368));
wire output_5_368, output_5_1, output_4_368;
mixer gate_output_4_368(.a(output_5_368), .b(output_5_1), .y(output_4_368));
wire output_6_368, output_6_1, output_5_368;
mixer gate_output_5_368(.a(output_6_368), .b(output_6_1), .y(output_5_368));
wire output_7_368, output_7_1, output_6_368;
mixer gate_output_6_368(.a(output_7_368), .b(output_7_1), .y(output_6_368));
wire output_8_368, output_8_1, output_7_368;
mixer gate_output_7_368(.a(output_8_368), .b(output_8_1), .y(output_7_368));
wire output_9_368, output_9_1, output_8_368;
mixer gate_output_8_368(.a(output_9_368), .b(output_9_1), .y(output_8_368));
wire output_10_368, output_10_1, output_9_368;
mixer gate_output_9_368(.a(output_10_368), .b(output_10_1), .y(output_9_368));
wire output_11_368, output_11_1, output_10_368;
mixer gate_output_10_368(.a(output_11_368), .b(output_11_1), .y(output_10_368));
wire output_12_368, output_12_1, output_11_368;
mixer gate_output_11_368(.a(output_12_368), .b(output_12_1), .y(output_11_368));
wire output_13_368, output_13_1, output_12_368;
mixer gate_output_12_368(.a(output_13_368), .b(output_13_1), .y(output_12_368));
wire output_14_368, output_14_1, output_13_368;
mixer gate_output_13_368(.a(output_14_368), .b(output_14_1), .y(output_13_368));
wire output_15_368, output_15_1, output_14_368;
mixer gate_output_14_368(.a(output_15_368), .b(output_15_1), .y(output_14_368));
wire output_16_368, output_16_1, output_15_368;
mixer gate_output_15_368(.a(output_16_368), .b(output_16_1), .y(output_15_368));
wire output_1_369, output_1_2, output_0_369;
mixer gate_output_0_369(.a(output_1_369), .b(output_1_2), .y(output_0_369));
wire output_2_369, output_2_2, output_1_369;
mixer gate_output_1_369(.a(output_2_369), .b(output_2_2), .y(output_1_369));
wire output_3_369, output_3_2, output_2_369;
mixer gate_output_2_369(.a(output_3_369), .b(output_3_2), .y(output_2_369));
wire output_4_369, output_4_2, output_3_369;
mixer gate_output_3_369(.a(output_4_369), .b(output_4_2), .y(output_3_369));
wire output_5_369, output_5_2, output_4_369;
mixer gate_output_4_369(.a(output_5_369), .b(output_5_2), .y(output_4_369));
wire output_6_369, output_6_2, output_5_369;
mixer gate_output_5_369(.a(output_6_369), .b(output_6_2), .y(output_5_369));
wire output_7_369, output_7_2, output_6_369;
mixer gate_output_6_369(.a(output_7_369), .b(output_7_2), .y(output_6_369));
wire output_8_369, output_8_2, output_7_369;
mixer gate_output_7_369(.a(output_8_369), .b(output_8_2), .y(output_7_369));
wire output_9_369, output_9_2, output_8_369;
mixer gate_output_8_369(.a(output_9_369), .b(output_9_2), .y(output_8_369));
wire output_10_369, output_10_2, output_9_369;
mixer gate_output_9_369(.a(output_10_369), .b(output_10_2), .y(output_9_369));
wire output_11_369, output_11_2, output_10_369;
mixer gate_output_10_369(.a(output_11_369), .b(output_11_2), .y(output_10_369));
wire output_12_369, output_12_2, output_11_369;
mixer gate_output_11_369(.a(output_12_369), .b(output_12_2), .y(output_11_369));
wire output_13_369, output_13_2, output_12_369;
mixer gate_output_12_369(.a(output_13_369), .b(output_13_2), .y(output_12_369));
wire output_14_369, output_14_2, output_13_369;
mixer gate_output_13_369(.a(output_14_369), .b(output_14_2), .y(output_13_369));
wire output_15_369, output_15_2, output_14_369;
mixer gate_output_14_369(.a(output_15_369), .b(output_15_2), .y(output_14_369));
wire output_16_369, output_16_2, output_15_369;
mixer gate_output_15_369(.a(output_16_369), .b(output_16_2), .y(output_15_369));
wire output_1_370, output_1_3, output_0_370;
mixer gate_output_0_370(.a(output_1_370), .b(output_1_3), .y(output_0_370));
wire output_2_370, output_2_3, output_1_370;
mixer gate_output_1_370(.a(output_2_370), .b(output_2_3), .y(output_1_370));
wire output_3_370, output_3_3, output_2_370;
mixer gate_output_2_370(.a(output_3_370), .b(output_3_3), .y(output_2_370));
wire output_4_370, output_4_3, output_3_370;
mixer gate_output_3_370(.a(output_4_370), .b(output_4_3), .y(output_3_370));
wire output_5_370, output_5_3, output_4_370;
mixer gate_output_4_370(.a(output_5_370), .b(output_5_3), .y(output_4_370));
wire output_6_370, output_6_3, output_5_370;
mixer gate_output_5_370(.a(output_6_370), .b(output_6_3), .y(output_5_370));
wire output_7_370, output_7_3, output_6_370;
mixer gate_output_6_370(.a(output_7_370), .b(output_7_3), .y(output_6_370));
wire output_8_370, output_8_3, output_7_370;
mixer gate_output_7_370(.a(output_8_370), .b(output_8_3), .y(output_7_370));
wire output_9_370, output_9_3, output_8_370;
mixer gate_output_8_370(.a(output_9_370), .b(output_9_3), .y(output_8_370));
wire output_10_370, output_10_3, output_9_370;
mixer gate_output_9_370(.a(output_10_370), .b(output_10_3), .y(output_9_370));
wire output_11_370, output_11_3, output_10_370;
mixer gate_output_10_370(.a(output_11_370), .b(output_11_3), .y(output_10_370));
wire output_12_370, output_12_3, output_11_370;
mixer gate_output_11_370(.a(output_12_370), .b(output_12_3), .y(output_11_370));
wire output_13_370, output_13_3, output_12_370;
mixer gate_output_12_370(.a(output_13_370), .b(output_13_3), .y(output_12_370));
wire output_14_370, output_14_3, output_13_370;
mixer gate_output_13_370(.a(output_14_370), .b(output_14_3), .y(output_13_370));
wire output_15_370, output_15_3, output_14_370;
mixer gate_output_14_370(.a(output_15_370), .b(output_15_3), .y(output_14_370));
wire output_16_370, output_16_3, output_15_370;
mixer gate_output_15_370(.a(output_16_370), .b(output_16_3), .y(output_15_370));
wire output_1_371, output_1_4, output_0_371;
mixer gate_output_0_371(.a(output_1_371), .b(output_1_4), .y(output_0_371));
wire output_2_371, output_2_4, output_1_371;
mixer gate_output_1_371(.a(output_2_371), .b(output_2_4), .y(output_1_371));
wire output_3_371, output_3_4, output_2_371;
mixer gate_output_2_371(.a(output_3_371), .b(output_3_4), .y(output_2_371));
wire output_4_371, output_4_4, output_3_371;
mixer gate_output_3_371(.a(output_4_371), .b(output_4_4), .y(output_3_371));
wire output_5_371, output_5_4, output_4_371;
mixer gate_output_4_371(.a(output_5_371), .b(output_5_4), .y(output_4_371));
wire output_6_371, output_6_4, output_5_371;
mixer gate_output_5_371(.a(output_6_371), .b(output_6_4), .y(output_5_371));
wire output_7_371, output_7_4, output_6_371;
mixer gate_output_6_371(.a(output_7_371), .b(output_7_4), .y(output_6_371));
wire output_8_371, output_8_4, output_7_371;
mixer gate_output_7_371(.a(output_8_371), .b(output_8_4), .y(output_7_371));
wire output_9_371, output_9_4, output_8_371;
mixer gate_output_8_371(.a(output_9_371), .b(output_9_4), .y(output_8_371));
wire output_10_371, output_10_4, output_9_371;
mixer gate_output_9_371(.a(output_10_371), .b(output_10_4), .y(output_9_371));
wire output_11_371, output_11_4, output_10_371;
mixer gate_output_10_371(.a(output_11_371), .b(output_11_4), .y(output_10_371));
wire output_12_371, output_12_4, output_11_371;
mixer gate_output_11_371(.a(output_12_371), .b(output_12_4), .y(output_11_371));
wire output_13_371, output_13_4, output_12_371;
mixer gate_output_12_371(.a(output_13_371), .b(output_13_4), .y(output_12_371));
wire output_14_371, output_14_4, output_13_371;
mixer gate_output_13_371(.a(output_14_371), .b(output_14_4), .y(output_13_371));
wire output_15_371, output_15_4, output_14_371;
mixer gate_output_14_371(.a(output_15_371), .b(output_15_4), .y(output_14_371));
wire output_16_371, output_16_4, output_15_371;
mixer gate_output_15_371(.a(output_16_371), .b(output_16_4), .y(output_15_371));
wire output_1_372, output_1_5, output_0_372;
mixer gate_output_0_372(.a(output_1_372), .b(output_1_5), .y(output_0_372));
wire output_2_372, output_2_5, output_1_372;
mixer gate_output_1_372(.a(output_2_372), .b(output_2_5), .y(output_1_372));
wire output_3_372, output_3_5, output_2_372;
mixer gate_output_2_372(.a(output_3_372), .b(output_3_5), .y(output_2_372));
wire output_4_372, output_4_5, output_3_372;
mixer gate_output_3_372(.a(output_4_372), .b(output_4_5), .y(output_3_372));
wire output_5_372, output_5_5, output_4_372;
mixer gate_output_4_372(.a(output_5_372), .b(output_5_5), .y(output_4_372));
wire output_6_372, output_6_5, output_5_372;
mixer gate_output_5_372(.a(output_6_372), .b(output_6_5), .y(output_5_372));
wire output_7_372, output_7_5, output_6_372;
mixer gate_output_6_372(.a(output_7_372), .b(output_7_5), .y(output_6_372));
wire output_8_372, output_8_5, output_7_372;
mixer gate_output_7_372(.a(output_8_372), .b(output_8_5), .y(output_7_372));
wire output_9_372, output_9_5, output_8_372;
mixer gate_output_8_372(.a(output_9_372), .b(output_9_5), .y(output_8_372));
wire output_10_372, output_10_5, output_9_372;
mixer gate_output_9_372(.a(output_10_372), .b(output_10_5), .y(output_9_372));
wire output_11_372, output_11_5, output_10_372;
mixer gate_output_10_372(.a(output_11_372), .b(output_11_5), .y(output_10_372));
wire output_12_372, output_12_5, output_11_372;
mixer gate_output_11_372(.a(output_12_372), .b(output_12_5), .y(output_11_372));
wire output_13_372, output_13_5, output_12_372;
mixer gate_output_12_372(.a(output_13_372), .b(output_13_5), .y(output_12_372));
wire output_14_372, output_14_5, output_13_372;
mixer gate_output_13_372(.a(output_14_372), .b(output_14_5), .y(output_13_372));
wire output_15_372, output_15_5, output_14_372;
mixer gate_output_14_372(.a(output_15_372), .b(output_15_5), .y(output_14_372));
wire output_16_372, output_16_5, output_15_372;
mixer gate_output_15_372(.a(output_16_372), .b(output_16_5), .y(output_15_372));
wire output_1_373, output_1_6, output_0_373;
mixer gate_output_0_373(.a(output_1_373), .b(output_1_6), .y(output_0_373));
wire output_2_373, output_2_6, output_1_373;
mixer gate_output_1_373(.a(output_2_373), .b(output_2_6), .y(output_1_373));
wire output_3_373, output_3_6, output_2_373;
mixer gate_output_2_373(.a(output_3_373), .b(output_3_6), .y(output_2_373));
wire output_4_373, output_4_6, output_3_373;
mixer gate_output_3_373(.a(output_4_373), .b(output_4_6), .y(output_3_373));
wire output_5_373, output_5_6, output_4_373;
mixer gate_output_4_373(.a(output_5_373), .b(output_5_6), .y(output_4_373));
wire output_6_373, output_6_6, output_5_373;
mixer gate_output_5_373(.a(output_6_373), .b(output_6_6), .y(output_5_373));
wire output_7_373, output_7_6, output_6_373;
mixer gate_output_6_373(.a(output_7_373), .b(output_7_6), .y(output_6_373));
wire output_8_373, output_8_6, output_7_373;
mixer gate_output_7_373(.a(output_8_373), .b(output_8_6), .y(output_7_373));
wire output_9_373, output_9_6, output_8_373;
mixer gate_output_8_373(.a(output_9_373), .b(output_9_6), .y(output_8_373));
wire output_10_373, output_10_6, output_9_373;
mixer gate_output_9_373(.a(output_10_373), .b(output_10_6), .y(output_9_373));
wire output_11_373, output_11_6, output_10_373;
mixer gate_output_10_373(.a(output_11_373), .b(output_11_6), .y(output_10_373));
wire output_12_373, output_12_6, output_11_373;
mixer gate_output_11_373(.a(output_12_373), .b(output_12_6), .y(output_11_373));
wire output_13_373, output_13_6, output_12_373;
mixer gate_output_12_373(.a(output_13_373), .b(output_13_6), .y(output_12_373));
wire output_14_373, output_14_6, output_13_373;
mixer gate_output_13_373(.a(output_14_373), .b(output_14_6), .y(output_13_373));
wire output_15_373, output_15_6, output_14_373;
mixer gate_output_14_373(.a(output_15_373), .b(output_15_6), .y(output_14_373));
wire output_16_373, output_16_6, output_15_373;
mixer gate_output_15_373(.a(output_16_373), .b(output_16_6), .y(output_15_373));
wire output_1_374, output_1_7, output_0_374;
mixer gate_output_0_374(.a(output_1_374), .b(output_1_7), .y(output_0_374));
wire output_2_374, output_2_7, output_1_374;
mixer gate_output_1_374(.a(output_2_374), .b(output_2_7), .y(output_1_374));
wire output_3_374, output_3_7, output_2_374;
mixer gate_output_2_374(.a(output_3_374), .b(output_3_7), .y(output_2_374));
wire output_4_374, output_4_7, output_3_374;
mixer gate_output_3_374(.a(output_4_374), .b(output_4_7), .y(output_3_374));
wire output_5_374, output_5_7, output_4_374;
mixer gate_output_4_374(.a(output_5_374), .b(output_5_7), .y(output_4_374));
wire output_6_374, output_6_7, output_5_374;
mixer gate_output_5_374(.a(output_6_374), .b(output_6_7), .y(output_5_374));
wire output_7_374, output_7_7, output_6_374;
mixer gate_output_6_374(.a(output_7_374), .b(output_7_7), .y(output_6_374));
wire output_8_374, output_8_7, output_7_374;
mixer gate_output_7_374(.a(output_8_374), .b(output_8_7), .y(output_7_374));
wire output_9_374, output_9_7, output_8_374;
mixer gate_output_8_374(.a(output_9_374), .b(output_9_7), .y(output_8_374));
wire output_10_374, output_10_7, output_9_374;
mixer gate_output_9_374(.a(output_10_374), .b(output_10_7), .y(output_9_374));
wire output_11_374, output_11_7, output_10_374;
mixer gate_output_10_374(.a(output_11_374), .b(output_11_7), .y(output_10_374));
wire output_12_374, output_12_7, output_11_374;
mixer gate_output_11_374(.a(output_12_374), .b(output_12_7), .y(output_11_374));
wire output_13_374, output_13_7, output_12_374;
mixer gate_output_12_374(.a(output_13_374), .b(output_13_7), .y(output_12_374));
wire output_14_374, output_14_7, output_13_374;
mixer gate_output_13_374(.a(output_14_374), .b(output_14_7), .y(output_13_374));
wire output_15_374, output_15_7, output_14_374;
mixer gate_output_14_374(.a(output_15_374), .b(output_15_7), .y(output_14_374));
wire output_16_374, output_16_7, output_15_374;
mixer gate_output_15_374(.a(output_16_374), .b(output_16_7), .y(output_15_374));
wire output_1_375, output_1_8, output_0_375;
mixer gate_output_0_375(.a(output_1_375), .b(output_1_8), .y(output_0_375));
wire output_2_375, output_2_8, output_1_375;
mixer gate_output_1_375(.a(output_2_375), .b(output_2_8), .y(output_1_375));
wire output_3_375, output_3_8, output_2_375;
mixer gate_output_2_375(.a(output_3_375), .b(output_3_8), .y(output_2_375));
wire output_4_375, output_4_8, output_3_375;
mixer gate_output_3_375(.a(output_4_375), .b(output_4_8), .y(output_3_375));
wire output_5_375, output_5_8, output_4_375;
mixer gate_output_4_375(.a(output_5_375), .b(output_5_8), .y(output_4_375));
wire output_6_375, output_6_8, output_5_375;
mixer gate_output_5_375(.a(output_6_375), .b(output_6_8), .y(output_5_375));
wire output_7_375, output_7_8, output_6_375;
mixer gate_output_6_375(.a(output_7_375), .b(output_7_8), .y(output_6_375));
wire output_8_375, output_8_8, output_7_375;
mixer gate_output_7_375(.a(output_8_375), .b(output_8_8), .y(output_7_375));
wire output_9_375, output_9_8, output_8_375;
mixer gate_output_8_375(.a(output_9_375), .b(output_9_8), .y(output_8_375));
wire output_10_375, output_10_8, output_9_375;
mixer gate_output_9_375(.a(output_10_375), .b(output_10_8), .y(output_9_375));
wire output_11_375, output_11_8, output_10_375;
mixer gate_output_10_375(.a(output_11_375), .b(output_11_8), .y(output_10_375));
wire output_12_375, output_12_8, output_11_375;
mixer gate_output_11_375(.a(output_12_375), .b(output_12_8), .y(output_11_375));
wire output_13_375, output_13_8, output_12_375;
mixer gate_output_12_375(.a(output_13_375), .b(output_13_8), .y(output_12_375));
wire output_14_375, output_14_8, output_13_375;
mixer gate_output_13_375(.a(output_14_375), .b(output_14_8), .y(output_13_375));
wire output_15_375, output_15_8, output_14_375;
mixer gate_output_14_375(.a(output_15_375), .b(output_15_8), .y(output_14_375));
wire output_16_375, output_16_8, output_15_375;
mixer gate_output_15_375(.a(output_16_375), .b(output_16_8), .y(output_15_375));
wire output_1_376, output_1_9, output_0_376;
mixer gate_output_0_376(.a(output_1_376), .b(output_1_9), .y(output_0_376));
wire output_2_376, output_2_9, output_1_376;
mixer gate_output_1_376(.a(output_2_376), .b(output_2_9), .y(output_1_376));
wire output_3_376, output_3_9, output_2_376;
mixer gate_output_2_376(.a(output_3_376), .b(output_3_9), .y(output_2_376));
wire output_4_376, output_4_9, output_3_376;
mixer gate_output_3_376(.a(output_4_376), .b(output_4_9), .y(output_3_376));
wire output_5_376, output_5_9, output_4_376;
mixer gate_output_4_376(.a(output_5_376), .b(output_5_9), .y(output_4_376));
wire output_6_376, output_6_9, output_5_376;
mixer gate_output_5_376(.a(output_6_376), .b(output_6_9), .y(output_5_376));
wire output_7_376, output_7_9, output_6_376;
mixer gate_output_6_376(.a(output_7_376), .b(output_7_9), .y(output_6_376));
wire output_8_376, output_8_9, output_7_376;
mixer gate_output_7_376(.a(output_8_376), .b(output_8_9), .y(output_7_376));
wire output_9_376, output_9_9, output_8_376;
mixer gate_output_8_376(.a(output_9_376), .b(output_9_9), .y(output_8_376));
wire output_10_376, output_10_9, output_9_376;
mixer gate_output_9_376(.a(output_10_376), .b(output_10_9), .y(output_9_376));
wire output_11_376, output_11_9, output_10_376;
mixer gate_output_10_376(.a(output_11_376), .b(output_11_9), .y(output_10_376));
wire output_12_376, output_12_9, output_11_376;
mixer gate_output_11_376(.a(output_12_376), .b(output_12_9), .y(output_11_376));
wire output_13_376, output_13_9, output_12_376;
mixer gate_output_12_376(.a(output_13_376), .b(output_13_9), .y(output_12_376));
wire output_14_376, output_14_9, output_13_376;
mixer gate_output_13_376(.a(output_14_376), .b(output_14_9), .y(output_13_376));
wire output_15_376, output_15_9, output_14_376;
mixer gate_output_14_376(.a(output_15_376), .b(output_15_9), .y(output_14_376));
wire output_16_376, output_16_9, output_15_376;
mixer gate_output_15_376(.a(output_16_376), .b(output_16_9), .y(output_15_376));
wire output_1_377, output_1_10, output_0_377;
mixer gate_output_0_377(.a(output_1_377), .b(output_1_10), .y(output_0_377));
wire output_2_377, output_2_10, output_1_377;
mixer gate_output_1_377(.a(output_2_377), .b(output_2_10), .y(output_1_377));
wire output_3_377, output_3_10, output_2_377;
mixer gate_output_2_377(.a(output_3_377), .b(output_3_10), .y(output_2_377));
wire output_4_377, output_4_10, output_3_377;
mixer gate_output_3_377(.a(output_4_377), .b(output_4_10), .y(output_3_377));
wire output_5_377, output_5_10, output_4_377;
mixer gate_output_4_377(.a(output_5_377), .b(output_5_10), .y(output_4_377));
wire output_6_377, output_6_10, output_5_377;
mixer gate_output_5_377(.a(output_6_377), .b(output_6_10), .y(output_5_377));
wire output_7_377, output_7_10, output_6_377;
mixer gate_output_6_377(.a(output_7_377), .b(output_7_10), .y(output_6_377));
wire output_8_377, output_8_10, output_7_377;
mixer gate_output_7_377(.a(output_8_377), .b(output_8_10), .y(output_7_377));
wire output_9_377, output_9_10, output_8_377;
mixer gate_output_8_377(.a(output_9_377), .b(output_9_10), .y(output_8_377));
wire output_10_377, output_10_10, output_9_377;
mixer gate_output_9_377(.a(output_10_377), .b(output_10_10), .y(output_9_377));
wire output_11_377, output_11_10, output_10_377;
mixer gate_output_10_377(.a(output_11_377), .b(output_11_10), .y(output_10_377));
wire output_12_377, output_12_10, output_11_377;
mixer gate_output_11_377(.a(output_12_377), .b(output_12_10), .y(output_11_377));
wire output_13_377, output_13_10, output_12_377;
mixer gate_output_12_377(.a(output_13_377), .b(output_13_10), .y(output_12_377));
wire output_14_377, output_14_10, output_13_377;
mixer gate_output_13_377(.a(output_14_377), .b(output_14_10), .y(output_13_377));
wire output_15_377, output_15_10, output_14_377;
mixer gate_output_14_377(.a(output_15_377), .b(output_15_10), .y(output_14_377));
wire output_16_377, output_16_10, output_15_377;
mixer gate_output_15_377(.a(output_16_377), .b(output_16_10), .y(output_15_377));
wire output_1_378, output_1_11, output_0_378;
mixer gate_output_0_378(.a(output_1_378), .b(output_1_11), .y(output_0_378));
wire output_2_378, output_2_11, output_1_378;
mixer gate_output_1_378(.a(output_2_378), .b(output_2_11), .y(output_1_378));
wire output_3_378, output_3_11, output_2_378;
mixer gate_output_2_378(.a(output_3_378), .b(output_3_11), .y(output_2_378));
wire output_4_378, output_4_11, output_3_378;
mixer gate_output_3_378(.a(output_4_378), .b(output_4_11), .y(output_3_378));
wire output_5_378, output_5_11, output_4_378;
mixer gate_output_4_378(.a(output_5_378), .b(output_5_11), .y(output_4_378));
wire output_6_378, output_6_11, output_5_378;
mixer gate_output_5_378(.a(output_6_378), .b(output_6_11), .y(output_5_378));
wire output_7_378, output_7_11, output_6_378;
mixer gate_output_6_378(.a(output_7_378), .b(output_7_11), .y(output_6_378));
wire output_8_378, output_8_11, output_7_378;
mixer gate_output_7_378(.a(output_8_378), .b(output_8_11), .y(output_7_378));
wire output_9_378, output_9_11, output_8_378;
mixer gate_output_8_378(.a(output_9_378), .b(output_9_11), .y(output_8_378));
wire output_10_378, output_10_11, output_9_378;
mixer gate_output_9_378(.a(output_10_378), .b(output_10_11), .y(output_9_378));
wire output_11_378, output_11_11, output_10_378;
mixer gate_output_10_378(.a(output_11_378), .b(output_11_11), .y(output_10_378));
wire output_12_378, output_12_11, output_11_378;
mixer gate_output_11_378(.a(output_12_378), .b(output_12_11), .y(output_11_378));
wire output_13_378, output_13_11, output_12_378;
mixer gate_output_12_378(.a(output_13_378), .b(output_13_11), .y(output_12_378));
wire output_14_378, output_14_11, output_13_378;
mixer gate_output_13_378(.a(output_14_378), .b(output_14_11), .y(output_13_378));
wire output_15_378, output_15_11, output_14_378;
mixer gate_output_14_378(.a(output_15_378), .b(output_15_11), .y(output_14_378));
wire output_16_378, output_16_11, output_15_378;
mixer gate_output_15_378(.a(output_16_378), .b(output_16_11), .y(output_15_378));
wire output_1_379, output_1_12, output_0_379;
mixer gate_output_0_379(.a(output_1_379), .b(output_1_12), .y(output_0_379));
wire output_2_379, output_2_12, output_1_379;
mixer gate_output_1_379(.a(output_2_379), .b(output_2_12), .y(output_1_379));
wire output_3_379, output_3_12, output_2_379;
mixer gate_output_2_379(.a(output_3_379), .b(output_3_12), .y(output_2_379));
wire output_4_379, output_4_12, output_3_379;
mixer gate_output_3_379(.a(output_4_379), .b(output_4_12), .y(output_3_379));
wire output_5_379, output_5_12, output_4_379;
mixer gate_output_4_379(.a(output_5_379), .b(output_5_12), .y(output_4_379));
wire output_6_379, output_6_12, output_5_379;
mixer gate_output_5_379(.a(output_6_379), .b(output_6_12), .y(output_5_379));
wire output_7_379, output_7_12, output_6_379;
mixer gate_output_6_379(.a(output_7_379), .b(output_7_12), .y(output_6_379));
wire output_8_379, output_8_12, output_7_379;
mixer gate_output_7_379(.a(output_8_379), .b(output_8_12), .y(output_7_379));
wire output_9_379, output_9_12, output_8_379;
mixer gate_output_8_379(.a(output_9_379), .b(output_9_12), .y(output_8_379));
wire output_10_379, output_10_12, output_9_379;
mixer gate_output_9_379(.a(output_10_379), .b(output_10_12), .y(output_9_379));
wire output_11_379, output_11_12, output_10_379;
mixer gate_output_10_379(.a(output_11_379), .b(output_11_12), .y(output_10_379));
wire output_12_379, output_12_12, output_11_379;
mixer gate_output_11_379(.a(output_12_379), .b(output_12_12), .y(output_11_379));
wire output_13_379, output_13_12, output_12_379;
mixer gate_output_12_379(.a(output_13_379), .b(output_13_12), .y(output_12_379));
wire output_14_379, output_14_12, output_13_379;
mixer gate_output_13_379(.a(output_14_379), .b(output_14_12), .y(output_13_379));
wire output_15_379, output_15_12, output_14_379;
mixer gate_output_14_379(.a(output_15_379), .b(output_15_12), .y(output_14_379));
wire output_16_379, output_16_12, output_15_379;
mixer gate_output_15_379(.a(output_16_379), .b(output_16_12), .y(output_15_379));
wire output_1_380, output_1_13, output_0_380;
mixer gate_output_0_380(.a(output_1_380), .b(output_1_13), .y(output_0_380));
wire output_2_380, output_2_13, output_1_380;
mixer gate_output_1_380(.a(output_2_380), .b(output_2_13), .y(output_1_380));
wire output_3_380, output_3_13, output_2_380;
mixer gate_output_2_380(.a(output_3_380), .b(output_3_13), .y(output_2_380));
wire output_4_380, output_4_13, output_3_380;
mixer gate_output_3_380(.a(output_4_380), .b(output_4_13), .y(output_3_380));
wire output_5_380, output_5_13, output_4_380;
mixer gate_output_4_380(.a(output_5_380), .b(output_5_13), .y(output_4_380));
wire output_6_380, output_6_13, output_5_380;
mixer gate_output_5_380(.a(output_6_380), .b(output_6_13), .y(output_5_380));
wire output_7_380, output_7_13, output_6_380;
mixer gate_output_6_380(.a(output_7_380), .b(output_7_13), .y(output_6_380));
wire output_8_380, output_8_13, output_7_380;
mixer gate_output_7_380(.a(output_8_380), .b(output_8_13), .y(output_7_380));
wire output_9_380, output_9_13, output_8_380;
mixer gate_output_8_380(.a(output_9_380), .b(output_9_13), .y(output_8_380));
wire output_10_380, output_10_13, output_9_380;
mixer gate_output_9_380(.a(output_10_380), .b(output_10_13), .y(output_9_380));
wire output_11_380, output_11_13, output_10_380;
mixer gate_output_10_380(.a(output_11_380), .b(output_11_13), .y(output_10_380));
wire output_12_380, output_12_13, output_11_380;
mixer gate_output_11_380(.a(output_12_380), .b(output_12_13), .y(output_11_380));
wire output_13_380, output_13_13, output_12_380;
mixer gate_output_12_380(.a(output_13_380), .b(output_13_13), .y(output_12_380));
wire output_14_380, output_14_13, output_13_380;
mixer gate_output_13_380(.a(output_14_380), .b(output_14_13), .y(output_13_380));
wire output_15_380, output_15_13, output_14_380;
mixer gate_output_14_380(.a(output_15_380), .b(output_15_13), .y(output_14_380));
wire output_16_380, output_16_13, output_15_380;
mixer gate_output_15_380(.a(output_16_380), .b(output_16_13), .y(output_15_380));
wire output_1_381, output_1_14, output_0_381;
mixer gate_output_0_381(.a(output_1_381), .b(output_1_14), .y(output_0_381));
wire output_2_381, output_2_14, output_1_381;
mixer gate_output_1_381(.a(output_2_381), .b(output_2_14), .y(output_1_381));
wire output_3_381, output_3_14, output_2_381;
mixer gate_output_2_381(.a(output_3_381), .b(output_3_14), .y(output_2_381));
wire output_4_381, output_4_14, output_3_381;
mixer gate_output_3_381(.a(output_4_381), .b(output_4_14), .y(output_3_381));
wire output_5_381, output_5_14, output_4_381;
mixer gate_output_4_381(.a(output_5_381), .b(output_5_14), .y(output_4_381));
wire output_6_381, output_6_14, output_5_381;
mixer gate_output_5_381(.a(output_6_381), .b(output_6_14), .y(output_5_381));
wire output_7_381, output_7_14, output_6_381;
mixer gate_output_6_381(.a(output_7_381), .b(output_7_14), .y(output_6_381));
wire output_8_381, output_8_14, output_7_381;
mixer gate_output_7_381(.a(output_8_381), .b(output_8_14), .y(output_7_381));
wire output_9_381, output_9_14, output_8_381;
mixer gate_output_8_381(.a(output_9_381), .b(output_9_14), .y(output_8_381));
wire output_10_381, output_10_14, output_9_381;
mixer gate_output_9_381(.a(output_10_381), .b(output_10_14), .y(output_9_381));
wire output_11_381, output_11_14, output_10_381;
mixer gate_output_10_381(.a(output_11_381), .b(output_11_14), .y(output_10_381));
wire output_12_381, output_12_14, output_11_381;
mixer gate_output_11_381(.a(output_12_381), .b(output_12_14), .y(output_11_381));
wire output_13_381, output_13_14, output_12_381;
mixer gate_output_12_381(.a(output_13_381), .b(output_13_14), .y(output_12_381));
wire output_14_381, output_14_14, output_13_381;
mixer gate_output_13_381(.a(output_14_381), .b(output_14_14), .y(output_13_381));
wire output_15_381, output_15_14, output_14_381;
mixer gate_output_14_381(.a(output_15_381), .b(output_15_14), .y(output_14_381));
wire output_16_381, output_16_14, output_15_381;
mixer gate_output_15_381(.a(output_16_381), .b(output_16_14), .y(output_15_381));
wire output_1_382, output_1_15, output_0_382;
mixer gate_output_0_382(.a(output_1_382), .b(output_1_15), .y(output_0_382));
wire output_2_382, output_2_15, output_1_382;
mixer gate_output_1_382(.a(output_2_382), .b(output_2_15), .y(output_1_382));
wire output_3_382, output_3_15, output_2_382;
mixer gate_output_2_382(.a(output_3_382), .b(output_3_15), .y(output_2_382));
wire output_4_382, output_4_15, output_3_382;
mixer gate_output_3_382(.a(output_4_382), .b(output_4_15), .y(output_3_382));
wire output_5_382, output_5_15, output_4_382;
mixer gate_output_4_382(.a(output_5_382), .b(output_5_15), .y(output_4_382));
wire output_6_382, output_6_15, output_5_382;
mixer gate_output_5_382(.a(output_6_382), .b(output_6_15), .y(output_5_382));
wire output_7_382, output_7_15, output_6_382;
mixer gate_output_6_382(.a(output_7_382), .b(output_7_15), .y(output_6_382));
wire output_8_382, output_8_15, output_7_382;
mixer gate_output_7_382(.a(output_8_382), .b(output_8_15), .y(output_7_382));
wire output_9_382, output_9_15, output_8_382;
mixer gate_output_8_382(.a(output_9_382), .b(output_9_15), .y(output_8_382));
wire output_10_382, output_10_15, output_9_382;
mixer gate_output_9_382(.a(output_10_382), .b(output_10_15), .y(output_9_382));
wire output_11_382, output_11_15, output_10_382;
mixer gate_output_10_382(.a(output_11_382), .b(output_11_15), .y(output_10_382));
wire output_12_382, output_12_15, output_11_382;
mixer gate_output_11_382(.a(output_12_382), .b(output_12_15), .y(output_11_382));
wire output_13_382, output_13_15, output_12_382;
mixer gate_output_12_382(.a(output_13_382), .b(output_13_15), .y(output_12_382));
wire output_14_382, output_14_15, output_13_382;
mixer gate_output_13_382(.a(output_14_382), .b(output_14_15), .y(output_13_382));
wire output_15_382, output_15_15, output_14_382;
mixer gate_output_14_382(.a(output_15_382), .b(output_15_15), .y(output_14_382));
wire output_16_382, output_16_15, output_15_382;
mixer gate_output_15_382(.a(output_16_382), .b(output_16_15), .y(output_15_382));
wire output_1_383, output_1_0, output_0_383;
mixer gate_output_0_383(.a(output_1_383), .b(output_1_0), .y(output_0_383));
wire output_2_383, output_2_0, output_1_383;
mixer gate_output_1_383(.a(output_2_383), .b(output_2_0), .y(output_1_383));
wire output_3_383, output_3_0, output_2_383;
mixer gate_output_2_383(.a(output_3_383), .b(output_3_0), .y(output_2_383));
wire output_4_383, output_4_0, output_3_383;
mixer gate_output_3_383(.a(output_4_383), .b(output_4_0), .y(output_3_383));
wire output_5_383, output_5_0, output_4_383;
mixer gate_output_4_383(.a(output_5_383), .b(output_5_0), .y(output_4_383));
wire output_6_383, output_6_0, output_5_383;
mixer gate_output_5_383(.a(output_6_383), .b(output_6_0), .y(output_5_383));
wire output_7_383, output_7_0, output_6_383;
mixer gate_output_6_383(.a(output_7_383), .b(output_7_0), .y(output_6_383));
wire output_8_383, output_8_0, output_7_383;
mixer gate_output_7_383(.a(output_8_383), .b(output_8_0), .y(output_7_383));
wire output_9_383, output_9_0, output_8_383;
mixer gate_output_8_383(.a(output_9_383), .b(output_9_0), .y(output_8_383));
wire output_10_383, output_10_0, output_9_383;
mixer gate_output_9_383(.a(output_10_383), .b(output_10_0), .y(output_9_383));
wire output_11_383, output_11_0, output_10_383;
mixer gate_output_10_383(.a(output_11_383), .b(output_11_0), .y(output_10_383));
wire output_12_383, output_12_0, output_11_383;
mixer gate_output_11_383(.a(output_12_383), .b(output_12_0), .y(output_11_383));
wire output_13_383, output_13_0, output_12_383;
mixer gate_output_12_383(.a(output_13_383), .b(output_13_0), .y(output_12_383));
wire output_14_383, output_14_0, output_13_383;
mixer gate_output_13_383(.a(output_14_383), .b(output_14_0), .y(output_13_383));
wire output_15_383, output_15_0, output_14_383;
mixer gate_output_14_383(.a(output_15_383), .b(output_15_0), .y(output_14_383));
wire output_16_383, output_16_0, output_15_383;
mixer gate_output_15_383(.a(output_16_383), .b(output_16_0), .y(output_15_383));
wire output_1_384, output_1_1, output_0_384;
mixer gate_output_0_384(.a(output_1_384), .b(output_1_1), .y(output_0_384));
wire output_2_384, output_2_1, output_1_384;
mixer gate_output_1_384(.a(output_2_384), .b(output_2_1), .y(output_1_384));
wire output_3_384, output_3_1, output_2_384;
mixer gate_output_2_384(.a(output_3_384), .b(output_3_1), .y(output_2_384));
wire output_4_384, output_4_1, output_3_384;
mixer gate_output_3_384(.a(output_4_384), .b(output_4_1), .y(output_3_384));
wire output_5_384, output_5_1, output_4_384;
mixer gate_output_4_384(.a(output_5_384), .b(output_5_1), .y(output_4_384));
wire output_6_384, output_6_1, output_5_384;
mixer gate_output_5_384(.a(output_6_384), .b(output_6_1), .y(output_5_384));
wire output_7_384, output_7_1, output_6_384;
mixer gate_output_6_384(.a(output_7_384), .b(output_7_1), .y(output_6_384));
wire output_8_384, output_8_1, output_7_384;
mixer gate_output_7_384(.a(output_8_384), .b(output_8_1), .y(output_7_384));
wire output_9_384, output_9_1, output_8_384;
mixer gate_output_8_384(.a(output_9_384), .b(output_9_1), .y(output_8_384));
wire output_10_384, output_10_1, output_9_384;
mixer gate_output_9_384(.a(output_10_384), .b(output_10_1), .y(output_9_384));
wire output_11_384, output_11_1, output_10_384;
mixer gate_output_10_384(.a(output_11_384), .b(output_11_1), .y(output_10_384));
wire output_12_384, output_12_1, output_11_384;
mixer gate_output_11_384(.a(output_12_384), .b(output_12_1), .y(output_11_384));
wire output_13_384, output_13_1, output_12_384;
mixer gate_output_12_384(.a(output_13_384), .b(output_13_1), .y(output_12_384));
wire output_14_384, output_14_1, output_13_384;
mixer gate_output_13_384(.a(output_14_384), .b(output_14_1), .y(output_13_384));
wire output_15_384, output_15_1, output_14_384;
mixer gate_output_14_384(.a(output_15_384), .b(output_15_1), .y(output_14_384));
wire output_16_384, output_16_1, output_15_384;
mixer gate_output_15_384(.a(output_16_384), .b(output_16_1), .y(output_15_384));
wire output_1_385, output_1_2, output_0_385;
mixer gate_output_0_385(.a(output_1_385), .b(output_1_2), .y(output_0_385));
wire output_2_385, output_2_2, output_1_385;
mixer gate_output_1_385(.a(output_2_385), .b(output_2_2), .y(output_1_385));
wire output_3_385, output_3_2, output_2_385;
mixer gate_output_2_385(.a(output_3_385), .b(output_3_2), .y(output_2_385));
wire output_4_385, output_4_2, output_3_385;
mixer gate_output_3_385(.a(output_4_385), .b(output_4_2), .y(output_3_385));
wire output_5_385, output_5_2, output_4_385;
mixer gate_output_4_385(.a(output_5_385), .b(output_5_2), .y(output_4_385));
wire output_6_385, output_6_2, output_5_385;
mixer gate_output_5_385(.a(output_6_385), .b(output_6_2), .y(output_5_385));
wire output_7_385, output_7_2, output_6_385;
mixer gate_output_6_385(.a(output_7_385), .b(output_7_2), .y(output_6_385));
wire output_8_385, output_8_2, output_7_385;
mixer gate_output_7_385(.a(output_8_385), .b(output_8_2), .y(output_7_385));
wire output_9_385, output_9_2, output_8_385;
mixer gate_output_8_385(.a(output_9_385), .b(output_9_2), .y(output_8_385));
wire output_10_385, output_10_2, output_9_385;
mixer gate_output_9_385(.a(output_10_385), .b(output_10_2), .y(output_9_385));
wire output_11_385, output_11_2, output_10_385;
mixer gate_output_10_385(.a(output_11_385), .b(output_11_2), .y(output_10_385));
wire output_12_385, output_12_2, output_11_385;
mixer gate_output_11_385(.a(output_12_385), .b(output_12_2), .y(output_11_385));
wire output_13_385, output_13_2, output_12_385;
mixer gate_output_12_385(.a(output_13_385), .b(output_13_2), .y(output_12_385));
wire output_14_385, output_14_2, output_13_385;
mixer gate_output_13_385(.a(output_14_385), .b(output_14_2), .y(output_13_385));
wire output_15_385, output_15_2, output_14_385;
mixer gate_output_14_385(.a(output_15_385), .b(output_15_2), .y(output_14_385));
wire output_16_385, output_16_2, output_15_385;
mixer gate_output_15_385(.a(output_16_385), .b(output_16_2), .y(output_15_385));
wire output_1_386, output_1_3, output_0_386;
mixer gate_output_0_386(.a(output_1_386), .b(output_1_3), .y(output_0_386));
wire output_2_386, output_2_3, output_1_386;
mixer gate_output_1_386(.a(output_2_386), .b(output_2_3), .y(output_1_386));
wire output_3_386, output_3_3, output_2_386;
mixer gate_output_2_386(.a(output_3_386), .b(output_3_3), .y(output_2_386));
wire output_4_386, output_4_3, output_3_386;
mixer gate_output_3_386(.a(output_4_386), .b(output_4_3), .y(output_3_386));
wire output_5_386, output_5_3, output_4_386;
mixer gate_output_4_386(.a(output_5_386), .b(output_5_3), .y(output_4_386));
wire output_6_386, output_6_3, output_5_386;
mixer gate_output_5_386(.a(output_6_386), .b(output_6_3), .y(output_5_386));
wire output_7_386, output_7_3, output_6_386;
mixer gate_output_6_386(.a(output_7_386), .b(output_7_3), .y(output_6_386));
wire output_8_386, output_8_3, output_7_386;
mixer gate_output_7_386(.a(output_8_386), .b(output_8_3), .y(output_7_386));
wire output_9_386, output_9_3, output_8_386;
mixer gate_output_8_386(.a(output_9_386), .b(output_9_3), .y(output_8_386));
wire output_10_386, output_10_3, output_9_386;
mixer gate_output_9_386(.a(output_10_386), .b(output_10_3), .y(output_9_386));
wire output_11_386, output_11_3, output_10_386;
mixer gate_output_10_386(.a(output_11_386), .b(output_11_3), .y(output_10_386));
wire output_12_386, output_12_3, output_11_386;
mixer gate_output_11_386(.a(output_12_386), .b(output_12_3), .y(output_11_386));
wire output_13_386, output_13_3, output_12_386;
mixer gate_output_12_386(.a(output_13_386), .b(output_13_3), .y(output_12_386));
wire output_14_386, output_14_3, output_13_386;
mixer gate_output_13_386(.a(output_14_386), .b(output_14_3), .y(output_13_386));
wire output_15_386, output_15_3, output_14_386;
mixer gate_output_14_386(.a(output_15_386), .b(output_15_3), .y(output_14_386));
wire output_16_386, output_16_3, output_15_386;
mixer gate_output_15_386(.a(output_16_386), .b(output_16_3), .y(output_15_386));
wire output_1_387, output_1_4, output_0_387;
mixer gate_output_0_387(.a(output_1_387), .b(output_1_4), .y(output_0_387));
wire output_2_387, output_2_4, output_1_387;
mixer gate_output_1_387(.a(output_2_387), .b(output_2_4), .y(output_1_387));
wire output_3_387, output_3_4, output_2_387;
mixer gate_output_2_387(.a(output_3_387), .b(output_3_4), .y(output_2_387));
wire output_4_387, output_4_4, output_3_387;
mixer gate_output_3_387(.a(output_4_387), .b(output_4_4), .y(output_3_387));
wire output_5_387, output_5_4, output_4_387;
mixer gate_output_4_387(.a(output_5_387), .b(output_5_4), .y(output_4_387));
wire output_6_387, output_6_4, output_5_387;
mixer gate_output_5_387(.a(output_6_387), .b(output_6_4), .y(output_5_387));
wire output_7_387, output_7_4, output_6_387;
mixer gate_output_6_387(.a(output_7_387), .b(output_7_4), .y(output_6_387));
wire output_8_387, output_8_4, output_7_387;
mixer gate_output_7_387(.a(output_8_387), .b(output_8_4), .y(output_7_387));
wire output_9_387, output_9_4, output_8_387;
mixer gate_output_8_387(.a(output_9_387), .b(output_9_4), .y(output_8_387));
wire output_10_387, output_10_4, output_9_387;
mixer gate_output_9_387(.a(output_10_387), .b(output_10_4), .y(output_9_387));
wire output_11_387, output_11_4, output_10_387;
mixer gate_output_10_387(.a(output_11_387), .b(output_11_4), .y(output_10_387));
wire output_12_387, output_12_4, output_11_387;
mixer gate_output_11_387(.a(output_12_387), .b(output_12_4), .y(output_11_387));
wire output_13_387, output_13_4, output_12_387;
mixer gate_output_12_387(.a(output_13_387), .b(output_13_4), .y(output_12_387));
wire output_14_387, output_14_4, output_13_387;
mixer gate_output_13_387(.a(output_14_387), .b(output_14_4), .y(output_13_387));
wire output_15_387, output_15_4, output_14_387;
mixer gate_output_14_387(.a(output_15_387), .b(output_15_4), .y(output_14_387));
wire output_16_387, output_16_4, output_15_387;
mixer gate_output_15_387(.a(output_16_387), .b(output_16_4), .y(output_15_387));
wire output_1_388, output_1_5, output_0_388;
mixer gate_output_0_388(.a(output_1_388), .b(output_1_5), .y(output_0_388));
wire output_2_388, output_2_5, output_1_388;
mixer gate_output_1_388(.a(output_2_388), .b(output_2_5), .y(output_1_388));
wire output_3_388, output_3_5, output_2_388;
mixer gate_output_2_388(.a(output_3_388), .b(output_3_5), .y(output_2_388));
wire output_4_388, output_4_5, output_3_388;
mixer gate_output_3_388(.a(output_4_388), .b(output_4_5), .y(output_3_388));
wire output_5_388, output_5_5, output_4_388;
mixer gate_output_4_388(.a(output_5_388), .b(output_5_5), .y(output_4_388));
wire output_6_388, output_6_5, output_5_388;
mixer gate_output_5_388(.a(output_6_388), .b(output_6_5), .y(output_5_388));
wire output_7_388, output_7_5, output_6_388;
mixer gate_output_6_388(.a(output_7_388), .b(output_7_5), .y(output_6_388));
wire output_8_388, output_8_5, output_7_388;
mixer gate_output_7_388(.a(output_8_388), .b(output_8_5), .y(output_7_388));
wire output_9_388, output_9_5, output_8_388;
mixer gate_output_8_388(.a(output_9_388), .b(output_9_5), .y(output_8_388));
wire output_10_388, output_10_5, output_9_388;
mixer gate_output_9_388(.a(output_10_388), .b(output_10_5), .y(output_9_388));
wire output_11_388, output_11_5, output_10_388;
mixer gate_output_10_388(.a(output_11_388), .b(output_11_5), .y(output_10_388));
wire output_12_388, output_12_5, output_11_388;
mixer gate_output_11_388(.a(output_12_388), .b(output_12_5), .y(output_11_388));
wire output_13_388, output_13_5, output_12_388;
mixer gate_output_12_388(.a(output_13_388), .b(output_13_5), .y(output_12_388));
wire output_14_388, output_14_5, output_13_388;
mixer gate_output_13_388(.a(output_14_388), .b(output_14_5), .y(output_13_388));
wire output_15_388, output_15_5, output_14_388;
mixer gate_output_14_388(.a(output_15_388), .b(output_15_5), .y(output_14_388));
wire output_16_388, output_16_5, output_15_388;
mixer gate_output_15_388(.a(output_16_388), .b(output_16_5), .y(output_15_388));
wire output_1_389, output_1_6, output_0_389;
mixer gate_output_0_389(.a(output_1_389), .b(output_1_6), .y(output_0_389));
wire output_2_389, output_2_6, output_1_389;
mixer gate_output_1_389(.a(output_2_389), .b(output_2_6), .y(output_1_389));
wire output_3_389, output_3_6, output_2_389;
mixer gate_output_2_389(.a(output_3_389), .b(output_3_6), .y(output_2_389));
wire output_4_389, output_4_6, output_3_389;
mixer gate_output_3_389(.a(output_4_389), .b(output_4_6), .y(output_3_389));
wire output_5_389, output_5_6, output_4_389;
mixer gate_output_4_389(.a(output_5_389), .b(output_5_6), .y(output_4_389));
wire output_6_389, output_6_6, output_5_389;
mixer gate_output_5_389(.a(output_6_389), .b(output_6_6), .y(output_5_389));
wire output_7_389, output_7_6, output_6_389;
mixer gate_output_6_389(.a(output_7_389), .b(output_7_6), .y(output_6_389));
wire output_8_389, output_8_6, output_7_389;
mixer gate_output_7_389(.a(output_8_389), .b(output_8_6), .y(output_7_389));
wire output_9_389, output_9_6, output_8_389;
mixer gate_output_8_389(.a(output_9_389), .b(output_9_6), .y(output_8_389));
wire output_10_389, output_10_6, output_9_389;
mixer gate_output_9_389(.a(output_10_389), .b(output_10_6), .y(output_9_389));
wire output_11_389, output_11_6, output_10_389;
mixer gate_output_10_389(.a(output_11_389), .b(output_11_6), .y(output_10_389));
wire output_12_389, output_12_6, output_11_389;
mixer gate_output_11_389(.a(output_12_389), .b(output_12_6), .y(output_11_389));
wire output_13_389, output_13_6, output_12_389;
mixer gate_output_12_389(.a(output_13_389), .b(output_13_6), .y(output_12_389));
wire output_14_389, output_14_6, output_13_389;
mixer gate_output_13_389(.a(output_14_389), .b(output_14_6), .y(output_13_389));
wire output_15_389, output_15_6, output_14_389;
mixer gate_output_14_389(.a(output_15_389), .b(output_15_6), .y(output_14_389));
wire output_16_389, output_16_6, output_15_389;
mixer gate_output_15_389(.a(output_16_389), .b(output_16_6), .y(output_15_389));
wire output_1_390, output_1_7, output_0_390;
mixer gate_output_0_390(.a(output_1_390), .b(output_1_7), .y(output_0_390));
wire output_2_390, output_2_7, output_1_390;
mixer gate_output_1_390(.a(output_2_390), .b(output_2_7), .y(output_1_390));
wire output_3_390, output_3_7, output_2_390;
mixer gate_output_2_390(.a(output_3_390), .b(output_3_7), .y(output_2_390));
wire output_4_390, output_4_7, output_3_390;
mixer gate_output_3_390(.a(output_4_390), .b(output_4_7), .y(output_3_390));
wire output_5_390, output_5_7, output_4_390;
mixer gate_output_4_390(.a(output_5_390), .b(output_5_7), .y(output_4_390));
wire output_6_390, output_6_7, output_5_390;
mixer gate_output_5_390(.a(output_6_390), .b(output_6_7), .y(output_5_390));
wire output_7_390, output_7_7, output_6_390;
mixer gate_output_6_390(.a(output_7_390), .b(output_7_7), .y(output_6_390));
wire output_8_390, output_8_7, output_7_390;
mixer gate_output_7_390(.a(output_8_390), .b(output_8_7), .y(output_7_390));
wire output_9_390, output_9_7, output_8_390;
mixer gate_output_8_390(.a(output_9_390), .b(output_9_7), .y(output_8_390));
wire output_10_390, output_10_7, output_9_390;
mixer gate_output_9_390(.a(output_10_390), .b(output_10_7), .y(output_9_390));
wire output_11_390, output_11_7, output_10_390;
mixer gate_output_10_390(.a(output_11_390), .b(output_11_7), .y(output_10_390));
wire output_12_390, output_12_7, output_11_390;
mixer gate_output_11_390(.a(output_12_390), .b(output_12_7), .y(output_11_390));
wire output_13_390, output_13_7, output_12_390;
mixer gate_output_12_390(.a(output_13_390), .b(output_13_7), .y(output_12_390));
wire output_14_390, output_14_7, output_13_390;
mixer gate_output_13_390(.a(output_14_390), .b(output_14_7), .y(output_13_390));
wire output_15_390, output_15_7, output_14_390;
mixer gate_output_14_390(.a(output_15_390), .b(output_15_7), .y(output_14_390));
wire output_16_390, output_16_7, output_15_390;
mixer gate_output_15_390(.a(output_16_390), .b(output_16_7), .y(output_15_390));
wire output_1_391, output_1_8, output_0_391;
mixer gate_output_0_391(.a(output_1_391), .b(output_1_8), .y(output_0_391));
wire output_2_391, output_2_8, output_1_391;
mixer gate_output_1_391(.a(output_2_391), .b(output_2_8), .y(output_1_391));
wire output_3_391, output_3_8, output_2_391;
mixer gate_output_2_391(.a(output_3_391), .b(output_3_8), .y(output_2_391));
wire output_4_391, output_4_8, output_3_391;
mixer gate_output_3_391(.a(output_4_391), .b(output_4_8), .y(output_3_391));
wire output_5_391, output_5_8, output_4_391;
mixer gate_output_4_391(.a(output_5_391), .b(output_5_8), .y(output_4_391));
wire output_6_391, output_6_8, output_5_391;
mixer gate_output_5_391(.a(output_6_391), .b(output_6_8), .y(output_5_391));
wire output_7_391, output_7_8, output_6_391;
mixer gate_output_6_391(.a(output_7_391), .b(output_7_8), .y(output_6_391));
wire output_8_391, output_8_8, output_7_391;
mixer gate_output_7_391(.a(output_8_391), .b(output_8_8), .y(output_7_391));
wire output_9_391, output_9_8, output_8_391;
mixer gate_output_8_391(.a(output_9_391), .b(output_9_8), .y(output_8_391));
wire output_10_391, output_10_8, output_9_391;
mixer gate_output_9_391(.a(output_10_391), .b(output_10_8), .y(output_9_391));
wire output_11_391, output_11_8, output_10_391;
mixer gate_output_10_391(.a(output_11_391), .b(output_11_8), .y(output_10_391));
wire output_12_391, output_12_8, output_11_391;
mixer gate_output_11_391(.a(output_12_391), .b(output_12_8), .y(output_11_391));
wire output_13_391, output_13_8, output_12_391;
mixer gate_output_12_391(.a(output_13_391), .b(output_13_8), .y(output_12_391));
wire output_14_391, output_14_8, output_13_391;
mixer gate_output_13_391(.a(output_14_391), .b(output_14_8), .y(output_13_391));
wire output_15_391, output_15_8, output_14_391;
mixer gate_output_14_391(.a(output_15_391), .b(output_15_8), .y(output_14_391));
wire output_16_391, output_16_8, output_15_391;
mixer gate_output_15_391(.a(output_16_391), .b(output_16_8), .y(output_15_391));
wire output_1_392, output_1_9, output_0_392;
mixer gate_output_0_392(.a(output_1_392), .b(output_1_9), .y(output_0_392));
wire output_2_392, output_2_9, output_1_392;
mixer gate_output_1_392(.a(output_2_392), .b(output_2_9), .y(output_1_392));
wire output_3_392, output_3_9, output_2_392;
mixer gate_output_2_392(.a(output_3_392), .b(output_3_9), .y(output_2_392));
wire output_4_392, output_4_9, output_3_392;
mixer gate_output_3_392(.a(output_4_392), .b(output_4_9), .y(output_3_392));
wire output_5_392, output_5_9, output_4_392;
mixer gate_output_4_392(.a(output_5_392), .b(output_5_9), .y(output_4_392));
wire output_6_392, output_6_9, output_5_392;
mixer gate_output_5_392(.a(output_6_392), .b(output_6_9), .y(output_5_392));
wire output_7_392, output_7_9, output_6_392;
mixer gate_output_6_392(.a(output_7_392), .b(output_7_9), .y(output_6_392));
wire output_8_392, output_8_9, output_7_392;
mixer gate_output_7_392(.a(output_8_392), .b(output_8_9), .y(output_7_392));
wire output_9_392, output_9_9, output_8_392;
mixer gate_output_8_392(.a(output_9_392), .b(output_9_9), .y(output_8_392));
wire output_10_392, output_10_9, output_9_392;
mixer gate_output_9_392(.a(output_10_392), .b(output_10_9), .y(output_9_392));
wire output_11_392, output_11_9, output_10_392;
mixer gate_output_10_392(.a(output_11_392), .b(output_11_9), .y(output_10_392));
wire output_12_392, output_12_9, output_11_392;
mixer gate_output_11_392(.a(output_12_392), .b(output_12_9), .y(output_11_392));
wire output_13_392, output_13_9, output_12_392;
mixer gate_output_12_392(.a(output_13_392), .b(output_13_9), .y(output_12_392));
wire output_14_392, output_14_9, output_13_392;
mixer gate_output_13_392(.a(output_14_392), .b(output_14_9), .y(output_13_392));
wire output_15_392, output_15_9, output_14_392;
mixer gate_output_14_392(.a(output_15_392), .b(output_15_9), .y(output_14_392));
wire output_16_392, output_16_9, output_15_392;
mixer gate_output_15_392(.a(output_16_392), .b(output_16_9), .y(output_15_392));
wire output_1_393, output_1_10, output_0_393;
mixer gate_output_0_393(.a(output_1_393), .b(output_1_10), .y(output_0_393));
wire output_2_393, output_2_10, output_1_393;
mixer gate_output_1_393(.a(output_2_393), .b(output_2_10), .y(output_1_393));
wire output_3_393, output_3_10, output_2_393;
mixer gate_output_2_393(.a(output_3_393), .b(output_3_10), .y(output_2_393));
wire output_4_393, output_4_10, output_3_393;
mixer gate_output_3_393(.a(output_4_393), .b(output_4_10), .y(output_3_393));
wire output_5_393, output_5_10, output_4_393;
mixer gate_output_4_393(.a(output_5_393), .b(output_5_10), .y(output_4_393));
wire output_6_393, output_6_10, output_5_393;
mixer gate_output_5_393(.a(output_6_393), .b(output_6_10), .y(output_5_393));
wire output_7_393, output_7_10, output_6_393;
mixer gate_output_6_393(.a(output_7_393), .b(output_7_10), .y(output_6_393));
wire output_8_393, output_8_10, output_7_393;
mixer gate_output_7_393(.a(output_8_393), .b(output_8_10), .y(output_7_393));
wire output_9_393, output_9_10, output_8_393;
mixer gate_output_8_393(.a(output_9_393), .b(output_9_10), .y(output_8_393));
wire output_10_393, output_10_10, output_9_393;
mixer gate_output_9_393(.a(output_10_393), .b(output_10_10), .y(output_9_393));
wire output_11_393, output_11_10, output_10_393;
mixer gate_output_10_393(.a(output_11_393), .b(output_11_10), .y(output_10_393));
wire output_12_393, output_12_10, output_11_393;
mixer gate_output_11_393(.a(output_12_393), .b(output_12_10), .y(output_11_393));
wire output_13_393, output_13_10, output_12_393;
mixer gate_output_12_393(.a(output_13_393), .b(output_13_10), .y(output_12_393));
wire output_14_393, output_14_10, output_13_393;
mixer gate_output_13_393(.a(output_14_393), .b(output_14_10), .y(output_13_393));
wire output_15_393, output_15_10, output_14_393;
mixer gate_output_14_393(.a(output_15_393), .b(output_15_10), .y(output_14_393));
wire output_16_393, output_16_10, output_15_393;
mixer gate_output_15_393(.a(output_16_393), .b(output_16_10), .y(output_15_393));
wire output_1_394, output_1_11, output_0_394;
mixer gate_output_0_394(.a(output_1_394), .b(output_1_11), .y(output_0_394));
wire output_2_394, output_2_11, output_1_394;
mixer gate_output_1_394(.a(output_2_394), .b(output_2_11), .y(output_1_394));
wire output_3_394, output_3_11, output_2_394;
mixer gate_output_2_394(.a(output_3_394), .b(output_3_11), .y(output_2_394));
wire output_4_394, output_4_11, output_3_394;
mixer gate_output_3_394(.a(output_4_394), .b(output_4_11), .y(output_3_394));
wire output_5_394, output_5_11, output_4_394;
mixer gate_output_4_394(.a(output_5_394), .b(output_5_11), .y(output_4_394));
wire output_6_394, output_6_11, output_5_394;
mixer gate_output_5_394(.a(output_6_394), .b(output_6_11), .y(output_5_394));
wire output_7_394, output_7_11, output_6_394;
mixer gate_output_6_394(.a(output_7_394), .b(output_7_11), .y(output_6_394));
wire output_8_394, output_8_11, output_7_394;
mixer gate_output_7_394(.a(output_8_394), .b(output_8_11), .y(output_7_394));
wire output_9_394, output_9_11, output_8_394;
mixer gate_output_8_394(.a(output_9_394), .b(output_9_11), .y(output_8_394));
wire output_10_394, output_10_11, output_9_394;
mixer gate_output_9_394(.a(output_10_394), .b(output_10_11), .y(output_9_394));
wire output_11_394, output_11_11, output_10_394;
mixer gate_output_10_394(.a(output_11_394), .b(output_11_11), .y(output_10_394));
wire output_12_394, output_12_11, output_11_394;
mixer gate_output_11_394(.a(output_12_394), .b(output_12_11), .y(output_11_394));
wire output_13_394, output_13_11, output_12_394;
mixer gate_output_12_394(.a(output_13_394), .b(output_13_11), .y(output_12_394));
wire output_14_394, output_14_11, output_13_394;
mixer gate_output_13_394(.a(output_14_394), .b(output_14_11), .y(output_13_394));
wire output_15_394, output_15_11, output_14_394;
mixer gate_output_14_394(.a(output_15_394), .b(output_15_11), .y(output_14_394));
wire output_16_394, output_16_11, output_15_394;
mixer gate_output_15_394(.a(output_16_394), .b(output_16_11), .y(output_15_394));
wire output_1_395, output_1_12, output_0_395;
mixer gate_output_0_395(.a(output_1_395), .b(output_1_12), .y(output_0_395));
wire output_2_395, output_2_12, output_1_395;
mixer gate_output_1_395(.a(output_2_395), .b(output_2_12), .y(output_1_395));
wire output_3_395, output_3_12, output_2_395;
mixer gate_output_2_395(.a(output_3_395), .b(output_3_12), .y(output_2_395));
wire output_4_395, output_4_12, output_3_395;
mixer gate_output_3_395(.a(output_4_395), .b(output_4_12), .y(output_3_395));
wire output_5_395, output_5_12, output_4_395;
mixer gate_output_4_395(.a(output_5_395), .b(output_5_12), .y(output_4_395));
wire output_6_395, output_6_12, output_5_395;
mixer gate_output_5_395(.a(output_6_395), .b(output_6_12), .y(output_5_395));
wire output_7_395, output_7_12, output_6_395;
mixer gate_output_6_395(.a(output_7_395), .b(output_7_12), .y(output_6_395));
wire output_8_395, output_8_12, output_7_395;
mixer gate_output_7_395(.a(output_8_395), .b(output_8_12), .y(output_7_395));
wire output_9_395, output_9_12, output_8_395;
mixer gate_output_8_395(.a(output_9_395), .b(output_9_12), .y(output_8_395));
wire output_10_395, output_10_12, output_9_395;
mixer gate_output_9_395(.a(output_10_395), .b(output_10_12), .y(output_9_395));
wire output_11_395, output_11_12, output_10_395;
mixer gate_output_10_395(.a(output_11_395), .b(output_11_12), .y(output_10_395));
wire output_12_395, output_12_12, output_11_395;
mixer gate_output_11_395(.a(output_12_395), .b(output_12_12), .y(output_11_395));
wire output_13_395, output_13_12, output_12_395;
mixer gate_output_12_395(.a(output_13_395), .b(output_13_12), .y(output_12_395));
wire output_14_395, output_14_12, output_13_395;
mixer gate_output_13_395(.a(output_14_395), .b(output_14_12), .y(output_13_395));
wire output_15_395, output_15_12, output_14_395;
mixer gate_output_14_395(.a(output_15_395), .b(output_15_12), .y(output_14_395));
wire output_16_395, output_16_12, output_15_395;
mixer gate_output_15_395(.a(output_16_395), .b(output_16_12), .y(output_15_395));
wire output_1_396, output_1_13, output_0_396;
mixer gate_output_0_396(.a(output_1_396), .b(output_1_13), .y(output_0_396));
wire output_2_396, output_2_13, output_1_396;
mixer gate_output_1_396(.a(output_2_396), .b(output_2_13), .y(output_1_396));
wire output_3_396, output_3_13, output_2_396;
mixer gate_output_2_396(.a(output_3_396), .b(output_3_13), .y(output_2_396));
wire output_4_396, output_4_13, output_3_396;
mixer gate_output_3_396(.a(output_4_396), .b(output_4_13), .y(output_3_396));
wire output_5_396, output_5_13, output_4_396;
mixer gate_output_4_396(.a(output_5_396), .b(output_5_13), .y(output_4_396));
wire output_6_396, output_6_13, output_5_396;
mixer gate_output_5_396(.a(output_6_396), .b(output_6_13), .y(output_5_396));
wire output_7_396, output_7_13, output_6_396;
mixer gate_output_6_396(.a(output_7_396), .b(output_7_13), .y(output_6_396));
wire output_8_396, output_8_13, output_7_396;
mixer gate_output_7_396(.a(output_8_396), .b(output_8_13), .y(output_7_396));
wire output_9_396, output_9_13, output_8_396;
mixer gate_output_8_396(.a(output_9_396), .b(output_9_13), .y(output_8_396));
wire output_10_396, output_10_13, output_9_396;
mixer gate_output_9_396(.a(output_10_396), .b(output_10_13), .y(output_9_396));
wire output_11_396, output_11_13, output_10_396;
mixer gate_output_10_396(.a(output_11_396), .b(output_11_13), .y(output_10_396));
wire output_12_396, output_12_13, output_11_396;
mixer gate_output_11_396(.a(output_12_396), .b(output_12_13), .y(output_11_396));
wire output_13_396, output_13_13, output_12_396;
mixer gate_output_12_396(.a(output_13_396), .b(output_13_13), .y(output_12_396));
wire output_14_396, output_14_13, output_13_396;
mixer gate_output_13_396(.a(output_14_396), .b(output_14_13), .y(output_13_396));
wire output_15_396, output_15_13, output_14_396;
mixer gate_output_14_396(.a(output_15_396), .b(output_15_13), .y(output_14_396));
wire output_16_396, output_16_13, output_15_396;
mixer gate_output_15_396(.a(output_16_396), .b(output_16_13), .y(output_15_396));
wire output_1_397, output_1_14, output_0_397;
mixer gate_output_0_397(.a(output_1_397), .b(output_1_14), .y(output_0_397));
wire output_2_397, output_2_14, output_1_397;
mixer gate_output_1_397(.a(output_2_397), .b(output_2_14), .y(output_1_397));
wire output_3_397, output_3_14, output_2_397;
mixer gate_output_2_397(.a(output_3_397), .b(output_3_14), .y(output_2_397));
wire output_4_397, output_4_14, output_3_397;
mixer gate_output_3_397(.a(output_4_397), .b(output_4_14), .y(output_3_397));
wire output_5_397, output_5_14, output_4_397;
mixer gate_output_4_397(.a(output_5_397), .b(output_5_14), .y(output_4_397));
wire output_6_397, output_6_14, output_5_397;
mixer gate_output_5_397(.a(output_6_397), .b(output_6_14), .y(output_5_397));
wire output_7_397, output_7_14, output_6_397;
mixer gate_output_6_397(.a(output_7_397), .b(output_7_14), .y(output_6_397));
wire output_8_397, output_8_14, output_7_397;
mixer gate_output_7_397(.a(output_8_397), .b(output_8_14), .y(output_7_397));
wire output_9_397, output_9_14, output_8_397;
mixer gate_output_8_397(.a(output_9_397), .b(output_9_14), .y(output_8_397));
wire output_10_397, output_10_14, output_9_397;
mixer gate_output_9_397(.a(output_10_397), .b(output_10_14), .y(output_9_397));
wire output_11_397, output_11_14, output_10_397;
mixer gate_output_10_397(.a(output_11_397), .b(output_11_14), .y(output_10_397));
wire output_12_397, output_12_14, output_11_397;
mixer gate_output_11_397(.a(output_12_397), .b(output_12_14), .y(output_11_397));
wire output_13_397, output_13_14, output_12_397;
mixer gate_output_12_397(.a(output_13_397), .b(output_13_14), .y(output_12_397));
wire output_14_397, output_14_14, output_13_397;
mixer gate_output_13_397(.a(output_14_397), .b(output_14_14), .y(output_13_397));
wire output_15_397, output_15_14, output_14_397;
mixer gate_output_14_397(.a(output_15_397), .b(output_15_14), .y(output_14_397));
wire output_16_397, output_16_14, output_15_397;
mixer gate_output_15_397(.a(output_16_397), .b(output_16_14), .y(output_15_397));
wire output_1_398, output_1_15, output_0_398;
mixer gate_output_0_398(.a(output_1_398), .b(output_1_15), .y(output_0_398));
wire output_2_398, output_2_15, output_1_398;
mixer gate_output_1_398(.a(output_2_398), .b(output_2_15), .y(output_1_398));
wire output_3_398, output_3_15, output_2_398;
mixer gate_output_2_398(.a(output_3_398), .b(output_3_15), .y(output_2_398));
wire output_4_398, output_4_15, output_3_398;
mixer gate_output_3_398(.a(output_4_398), .b(output_4_15), .y(output_3_398));
wire output_5_398, output_5_15, output_4_398;
mixer gate_output_4_398(.a(output_5_398), .b(output_5_15), .y(output_4_398));
wire output_6_398, output_6_15, output_5_398;
mixer gate_output_5_398(.a(output_6_398), .b(output_6_15), .y(output_5_398));
wire output_7_398, output_7_15, output_6_398;
mixer gate_output_6_398(.a(output_7_398), .b(output_7_15), .y(output_6_398));
wire output_8_398, output_8_15, output_7_398;
mixer gate_output_7_398(.a(output_8_398), .b(output_8_15), .y(output_7_398));
wire output_9_398, output_9_15, output_8_398;
mixer gate_output_8_398(.a(output_9_398), .b(output_9_15), .y(output_8_398));
wire output_10_398, output_10_15, output_9_398;
mixer gate_output_9_398(.a(output_10_398), .b(output_10_15), .y(output_9_398));
wire output_11_398, output_11_15, output_10_398;
mixer gate_output_10_398(.a(output_11_398), .b(output_11_15), .y(output_10_398));
wire output_12_398, output_12_15, output_11_398;
mixer gate_output_11_398(.a(output_12_398), .b(output_12_15), .y(output_11_398));
wire output_13_398, output_13_15, output_12_398;
mixer gate_output_12_398(.a(output_13_398), .b(output_13_15), .y(output_12_398));
wire output_14_398, output_14_15, output_13_398;
mixer gate_output_13_398(.a(output_14_398), .b(output_14_15), .y(output_13_398));
wire output_15_398, output_15_15, output_14_398;
mixer gate_output_14_398(.a(output_15_398), .b(output_15_15), .y(output_14_398));
wire output_16_398, output_16_15, output_15_398;
mixer gate_output_15_398(.a(output_16_398), .b(output_16_15), .y(output_15_398));
wire output_1_399, output_1_0, output_0_399;
mixer gate_output_0_399(.a(output_1_399), .b(output_1_0), .y(output_0_399));
wire output_2_399, output_2_0, output_1_399;
mixer gate_output_1_399(.a(output_2_399), .b(output_2_0), .y(output_1_399));
wire output_3_399, output_3_0, output_2_399;
mixer gate_output_2_399(.a(output_3_399), .b(output_3_0), .y(output_2_399));
wire output_4_399, output_4_0, output_3_399;
mixer gate_output_3_399(.a(output_4_399), .b(output_4_0), .y(output_3_399));
wire output_5_399, output_5_0, output_4_399;
mixer gate_output_4_399(.a(output_5_399), .b(output_5_0), .y(output_4_399));
wire output_6_399, output_6_0, output_5_399;
mixer gate_output_5_399(.a(output_6_399), .b(output_6_0), .y(output_5_399));
wire output_7_399, output_7_0, output_6_399;
mixer gate_output_6_399(.a(output_7_399), .b(output_7_0), .y(output_6_399));
wire output_8_399, output_8_0, output_7_399;
mixer gate_output_7_399(.a(output_8_399), .b(output_8_0), .y(output_7_399));
wire output_9_399, output_9_0, output_8_399;
mixer gate_output_8_399(.a(output_9_399), .b(output_9_0), .y(output_8_399));
wire output_10_399, output_10_0, output_9_399;
mixer gate_output_9_399(.a(output_10_399), .b(output_10_0), .y(output_9_399));
wire output_11_399, output_11_0, output_10_399;
mixer gate_output_10_399(.a(output_11_399), .b(output_11_0), .y(output_10_399));
wire output_12_399, output_12_0, output_11_399;
mixer gate_output_11_399(.a(output_12_399), .b(output_12_0), .y(output_11_399));
wire output_13_399, output_13_0, output_12_399;
mixer gate_output_12_399(.a(output_13_399), .b(output_13_0), .y(output_12_399));
wire output_14_399, output_14_0, output_13_399;
mixer gate_output_13_399(.a(output_14_399), .b(output_14_0), .y(output_13_399));
wire output_15_399, output_15_0, output_14_399;
mixer gate_output_14_399(.a(output_15_399), .b(output_15_0), .y(output_14_399));
wire output_16_399, output_16_0, output_15_399;
mixer gate_output_15_399(.a(output_16_399), .b(output_16_0), .y(output_15_399));
wire output_1_400, output_1_1, output_0_400;
mixer gate_output_0_400(.a(output_1_400), .b(output_1_1), .y(output_0_400));
wire output_2_400, output_2_1, output_1_400;
mixer gate_output_1_400(.a(output_2_400), .b(output_2_1), .y(output_1_400));
wire output_3_400, output_3_1, output_2_400;
mixer gate_output_2_400(.a(output_3_400), .b(output_3_1), .y(output_2_400));
wire output_4_400, output_4_1, output_3_400;
mixer gate_output_3_400(.a(output_4_400), .b(output_4_1), .y(output_3_400));
wire output_5_400, output_5_1, output_4_400;
mixer gate_output_4_400(.a(output_5_400), .b(output_5_1), .y(output_4_400));
wire output_6_400, output_6_1, output_5_400;
mixer gate_output_5_400(.a(output_6_400), .b(output_6_1), .y(output_5_400));
wire output_7_400, output_7_1, output_6_400;
mixer gate_output_6_400(.a(output_7_400), .b(output_7_1), .y(output_6_400));
wire output_8_400, output_8_1, output_7_400;
mixer gate_output_7_400(.a(output_8_400), .b(output_8_1), .y(output_7_400));
wire output_9_400, output_9_1, output_8_400;
mixer gate_output_8_400(.a(output_9_400), .b(output_9_1), .y(output_8_400));
wire output_10_400, output_10_1, output_9_400;
mixer gate_output_9_400(.a(output_10_400), .b(output_10_1), .y(output_9_400));
wire output_11_400, output_11_1, output_10_400;
mixer gate_output_10_400(.a(output_11_400), .b(output_11_1), .y(output_10_400));
wire output_12_400, output_12_1, output_11_400;
mixer gate_output_11_400(.a(output_12_400), .b(output_12_1), .y(output_11_400));
wire output_13_400, output_13_1, output_12_400;
mixer gate_output_12_400(.a(output_13_400), .b(output_13_1), .y(output_12_400));
wire output_14_400, output_14_1, output_13_400;
mixer gate_output_13_400(.a(output_14_400), .b(output_14_1), .y(output_13_400));
wire output_15_400, output_15_1, output_14_400;
mixer gate_output_14_400(.a(output_15_400), .b(output_15_1), .y(output_14_400));
wire output_16_400, output_16_1, output_15_400;
mixer gate_output_15_400(.a(output_16_400), .b(output_16_1), .y(output_15_400));
wire output_1_401, output_1_2, output_0_401;
mixer gate_output_0_401(.a(output_1_401), .b(output_1_2), .y(output_0_401));
wire output_2_401, output_2_2, output_1_401;
mixer gate_output_1_401(.a(output_2_401), .b(output_2_2), .y(output_1_401));
wire output_3_401, output_3_2, output_2_401;
mixer gate_output_2_401(.a(output_3_401), .b(output_3_2), .y(output_2_401));
wire output_4_401, output_4_2, output_3_401;
mixer gate_output_3_401(.a(output_4_401), .b(output_4_2), .y(output_3_401));
wire output_5_401, output_5_2, output_4_401;
mixer gate_output_4_401(.a(output_5_401), .b(output_5_2), .y(output_4_401));
wire output_6_401, output_6_2, output_5_401;
mixer gate_output_5_401(.a(output_6_401), .b(output_6_2), .y(output_5_401));
wire output_7_401, output_7_2, output_6_401;
mixer gate_output_6_401(.a(output_7_401), .b(output_7_2), .y(output_6_401));
wire output_8_401, output_8_2, output_7_401;
mixer gate_output_7_401(.a(output_8_401), .b(output_8_2), .y(output_7_401));
wire output_9_401, output_9_2, output_8_401;
mixer gate_output_8_401(.a(output_9_401), .b(output_9_2), .y(output_8_401));
wire output_10_401, output_10_2, output_9_401;
mixer gate_output_9_401(.a(output_10_401), .b(output_10_2), .y(output_9_401));
wire output_11_401, output_11_2, output_10_401;
mixer gate_output_10_401(.a(output_11_401), .b(output_11_2), .y(output_10_401));
wire output_12_401, output_12_2, output_11_401;
mixer gate_output_11_401(.a(output_12_401), .b(output_12_2), .y(output_11_401));
wire output_13_401, output_13_2, output_12_401;
mixer gate_output_12_401(.a(output_13_401), .b(output_13_2), .y(output_12_401));
wire output_14_401, output_14_2, output_13_401;
mixer gate_output_13_401(.a(output_14_401), .b(output_14_2), .y(output_13_401));
wire output_15_401, output_15_2, output_14_401;
mixer gate_output_14_401(.a(output_15_401), .b(output_15_2), .y(output_14_401));
wire output_16_401, output_16_2, output_15_401;
mixer gate_output_15_401(.a(output_16_401), .b(output_16_2), .y(output_15_401));
wire output_1_402, output_1_3, output_0_402;
mixer gate_output_0_402(.a(output_1_402), .b(output_1_3), .y(output_0_402));
wire output_2_402, output_2_3, output_1_402;
mixer gate_output_1_402(.a(output_2_402), .b(output_2_3), .y(output_1_402));
wire output_3_402, output_3_3, output_2_402;
mixer gate_output_2_402(.a(output_3_402), .b(output_3_3), .y(output_2_402));
wire output_4_402, output_4_3, output_3_402;
mixer gate_output_3_402(.a(output_4_402), .b(output_4_3), .y(output_3_402));
wire output_5_402, output_5_3, output_4_402;
mixer gate_output_4_402(.a(output_5_402), .b(output_5_3), .y(output_4_402));
wire output_6_402, output_6_3, output_5_402;
mixer gate_output_5_402(.a(output_6_402), .b(output_6_3), .y(output_5_402));
wire output_7_402, output_7_3, output_6_402;
mixer gate_output_6_402(.a(output_7_402), .b(output_7_3), .y(output_6_402));
wire output_8_402, output_8_3, output_7_402;
mixer gate_output_7_402(.a(output_8_402), .b(output_8_3), .y(output_7_402));
wire output_9_402, output_9_3, output_8_402;
mixer gate_output_8_402(.a(output_9_402), .b(output_9_3), .y(output_8_402));
wire output_10_402, output_10_3, output_9_402;
mixer gate_output_9_402(.a(output_10_402), .b(output_10_3), .y(output_9_402));
wire output_11_402, output_11_3, output_10_402;
mixer gate_output_10_402(.a(output_11_402), .b(output_11_3), .y(output_10_402));
wire output_12_402, output_12_3, output_11_402;
mixer gate_output_11_402(.a(output_12_402), .b(output_12_3), .y(output_11_402));
wire output_13_402, output_13_3, output_12_402;
mixer gate_output_12_402(.a(output_13_402), .b(output_13_3), .y(output_12_402));
wire output_14_402, output_14_3, output_13_402;
mixer gate_output_13_402(.a(output_14_402), .b(output_14_3), .y(output_13_402));
wire output_15_402, output_15_3, output_14_402;
mixer gate_output_14_402(.a(output_15_402), .b(output_15_3), .y(output_14_402));
wire output_16_402, output_16_3, output_15_402;
mixer gate_output_15_402(.a(output_16_402), .b(output_16_3), .y(output_15_402));
wire output_1_403, output_1_4, output_0_403;
mixer gate_output_0_403(.a(output_1_403), .b(output_1_4), .y(output_0_403));
wire output_2_403, output_2_4, output_1_403;
mixer gate_output_1_403(.a(output_2_403), .b(output_2_4), .y(output_1_403));
wire output_3_403, output_3_4, output_2_403;
mixer gate_output_2_403(.a(output_3_403), .b(output_3_4), .y(output_2_403));
wire output_4_403, output_4_4, output_3_403;
mixer gate_output_3_403(.a(output_4_403), .b(output_4_4), .y(output_3_403));
wire output_5_403, output_5_4, output_4_403;
mixer gate_output_4_403(.a(output_5_403), .b(output_5_4), .y(output_4_403));
wire output_6_403, output_6_4, output_5_403;
mixer gate_output_5_403(.a(output_6_403), .b(output_6_4), .y(output_5_403));
wire output_7_403, output_7_4, output_6_403;
mixer gate_output_6_403(.a(output_7_403), .b(output_7_4), .y(output_6_403));
wire output_8_403, output_8_4, output_7_403;
mixer gate_output_7_403(.a(output_8_403), .b(output_8_4), .y(output_7_403));
wire output_9_403, output_9_4, output_8_403;
mixer gate_output_8_403(.a(output_9_403), .b(output_9_4), .y(output_8_403));
wire output_10_403, output_10_4, output_9_403;
mixer gate_output_9_403(.a(output_10_403), .b(output_10_4), .y(output_9_403));
wire output_11_403, output_11_4, output_10_403;
mixer gate_output_10_403(.a(output_11_403), .b(output_11_4), .y(output_10_403));
wire output_12_403, output_12_4, output_11_403;
mixer gate_output_11_403(.a(output_12_403), .b(output_12_4), .y(output_11_403));
wire output_13_403, output_13_4, output_12_403;
mixer gate_output_12_403(.a(output_13_403), .b(output_13_4), .y(output_12_403));
wire output_14_403, output_14_4, output_13_403;
mixer gate_output_13_403(.a(output_14_403), .b(output_14_4), .y(output_13_403));
wire output_15_403, output_15_4, output_14_403;
mixer gate_output_14_403(.a(output_15_403), .b(output_15_4), .y(output_14_403));
wire output_16_403, output_16_4, output_15_403;
mixer gate_output_15_403(.a(output_16_403), .b(output_16_4), .y(output_15_403));
wire output_1_404, output_1_5, output_0_404;
mixer gate_output_0_404(.a(output_1_404), .b(output_1_5), .y(output_0_404));
wire output_2_404, output_2_5, output_1_404;
mixer gate_output_1_404(.a(output_2_404), .b(output_2_5), .y(output_1_404));
wire output_3_404, output_3_5, output_2_404;
mixer gate_output_2_404(.a(output_3_404), .b(output_3_5), .y(output_2_404));
wire output_4_404, output_4_5, output_3_404;
mixer gate_output_3_404(.a(output_4_404), .b(output_4_5), .y(output_3_404));
wire output_5_404, output_5_5, output_4_404;
mixer gate_output_4_404(.a(output_5_404), .b(output_5_5), .y(output_4_404));
wire output_6_404, output_6_5, output_5_404;
mixer gate_output_5_404(.a(output_6_404), .b(output_6_5), .y(output_5_404));
wire output_7_404, output_7_5, output_6_404;
mixer gate_output_6_404(.a(output_7_404), .b(output_7_5), .y(output_6_404));
wire output_8_404, output_8_5, output_7_404;
mixer gate_output_7_404(.a(output_8_404), .b(output_8_5), .y(output_7_404));
wire output_9_404, output_9_5, output_8_404;
mixer gate_output_8_404(.a(output_9_404), .b(output_9_5), .y(output_8_404));
wire output_10_404, output_10_5, output_9_404;
mixer gate_output_9_404(.a(output_10_404), .b(output_10_5), .y(output_9_404));
wire output_11_404, output_11_5, output_10_404;
mixer gate_output_10_404(.a(output_11_404), .b(output_11_5), .y(output_10_404));
wire output_12_404, output_12_5, output_11_404;
mixer gate_output_11_404(.a(output_12_404), .b(output_12_5), .y(output_11_404));
wire output_13_404, output_13_5, output_12_404;
mixer gate_output_12_404(.a(output_13_404), .b(output_13_5), .y(output_12_404));
wire output_14_404, output_14_5, output_13_404;
mixer gate_output_13_404(.a(output_14_404), .b(output_14_5), .y(output_13_404));
wire output_15_404, output_15_5, output_14_404;
mixer gate_output_14_404(.a(output_15_404), .b(output_15_5), .y(output_14_404));
wire output_16_404, output_16_5, output_15_404;
mixer gate_output_15_404(.a(output_16_404), .b(output_16_5), .y(output_15_404));
wire output_1_405, output_1_6, output_0_405;
mixer gate_output_0_405(.a(output_1_405), .b(output_1_6), .y(output_0_405));
wire output_2_405, output_2_6, output_1_405;
mixer gate_output_1_405(.a(output_2_405), .b(output_2_6), .y(output_1_405));
wire output_3_405, output_3_6, output_2_405;
mixer gate_output_2_405(.a(output_3_405), .b(output_3_6), .y(output_2_405));
wire output_4_405, output_4_6, output_3_405;
mixer gate_output_3_405(.a(output_4_405), .b(output_4_6), .y(output_3_405));
wire output_5_405, output_5_6, output_4_405;
mixer gate_output_4_405(.a(output_5_405), .b(output_5_6), .y(output_4_405));
wire output_6_405, output_6_6, output_5_405;
mixer gate_output_5_405(.a(output_6_405), .b(output_6_6), .y(output_5_405));
wire output_7_405, output_7_6, output_6_405;
mixer gate_output_6_405(.a(output_7_405), .b(output_7_6), .y(output_6_405));
wire output_8_405, output_8_6, output_7_405;
mixer gate_output_7_405(.a(output_8_405), .b(output_8_6), .y(output_7_405));
wire output_9_405, output_9_6, output_8_405;
mixer gate_output_8_405(.a(output_9_405), .b(output_9_6), .y(output_8_405));
wire output_10_405, output_10_6, output_9_405;
mixer gate_output_9_405(.a(output_10_405), .b(output_10_6), .y(output_9_405));
wire output_11_405, output_11_6, output_10_405;
mixer gate_output_10_405(.a(output_11_405), .b(output_11_6), .y(output_10_405));
wire output_12_405, output_12_6, output_11_405;
mixer gate_output_11_405(.a(output_12_405), .b(output_12_6), .y(output_11_405));
wire output_13_405, output_13_6, output_12_405;
mixer gate_output_12_405(.a(output_13_405), .b(output_13_6), .y(output_12_405));
wire output_14_405, output_14_6, output_13_405;
mixer gate_output_13_405(.a(output_14_405), .b(output_14_6), .y(output_13_405));
wire output_15_405, output_15_6, output_14_405;
mixer gate_output_14_405(.a(output_15_405), .b(output_15_6), .y(output_14_405));
wire output_16_405, output_16_6, output_15_405;
mixer gate_output_15_405(.a(output_16_405), .b(output_16_6), .y(output_15_405));
wire output_1_406, output_1_7, output_0_406;
mixer gate_output_0_406(.a(output_1_406), .b(output_1_7), .y(output_0_406));
wire output_2_406, output_2_7, output_1_406;
mixer gate_output_1_406(.a(output_2_406), .b(output_2_7), .y(output_1_406));
wire output_3_406, output_3_7, output_2_406;
mixer gate_output_2_406(.a(output_3_406), .b(output_3_7), .y(output_2_406));
wire output_4_406, output_4_7, output_3_406;
mixer gate_output_3_406(.a(output_4_406), .b(output_4_7), .y(output_3_406));
wire output_5_406, output_5_7, output_4_406;
mixer gate_output_4_406(.a(output_5_406), .b(output_5_7), .y(output_4_406));
wire output_6_406, output_6_7, output_5_406;
mixer gate_output_5_406(.a(output_6_406), .b(output_6_7), .y(output_5_406));
wire output_7_406, output_7_7, output_6_406;
mixer gate_output_6_406(.a(output_7_406), .b(output_7_7), .y(output_6_406));
wire output_8_406, output_8_7, output_7_406;
mixer gate_output_7_406(.a(output_8_406), .b(output_8_7), .y(output_7_406));
wire output_9_406, output_9_7, output_8_406;
mixer gate_output_8_406(.a(output_9_406), .b(output_9_7), .y(output_8_406));
wire output_10_406, output_10_7, output_9_406;
mixer gate_output_9_406(.a(output_10_406), .b(output_10_7), .y(output_9_406));
wire output_11_406, output_11_7, output_10_406;
mixer gate_output_10_406(.a(output_11_406), .b(output_11_7), .y(output_10_406));
wire output_12_406, output_12_7, output_11_406;
mixer gate_output_11_406(.a(output_12_406), .b(output_12_7), .y(output_11_406));
wire output_13_406, output_13_7, output_12_406;
mixer gate_output_12_406(.a(output_13_406), .b(output_13_7), .y(output_12_406));
wire output_14_406, output_14_7, output_13_406;
mixer gate_output_13_406(.a(output_14_406), .b(output_14_7), .y(output_13_406));
wire output_15_406, output_15_7, output_14_406;
mixer gate_output_14_406(.a(output_15_406), .b(output_15_7), .y(output_14_406));
wire output_16_406, output_16_7, output_15_406;
mixer gate_output_15_406(.a(output_16_406), .b(output_16_7), .y(output_15_406));
wire output_1_407, output_1_8, output_0_407;
mixer gate_output_0_407(.a(output_1_407), .b(output_1_8), .y(output_0_407));
wire output_2_407, output_2_8, output_1_407;
mixer gate_output_1_407(.a(output_2_407), .b(output_2_8), .y(output_1_407));
wire output_3_407, output_3_8, output_2_407;
mixer gate_output_2_407(.a(output_3_407), .b(output_3_8), .y(output_2_407));
wire output_4_407, output_4_8, output_3_407;
mixer gate_output_3_407(.a(output_4_407), .b(output_4_8), .y(output_3_407));
wire output_5_407, output_5_8, output_4_407;
mixer gate_output_4_407(.a(output_5_407), .b(output_5_8), .y(output_4_407));
wire output_6_407, output_6_8, output_5_407;
mixer gate_output_5_407(.a(output_6_407), .b(output_6_8), .y(output_5_407));
wire output_7_407, output_7_8, output_6_407;
mixer gate_output_6_407(.a(output_7_407), .b(output_7_8), .y(output_6_407));
wire output_8_407, output_8_8, output_7_407;
mixer gate_output_7_407(.a(output_8_407), .b(output_8_8), .y(output_7_407));
wire output_9_407, output_9_8, output_8_407;
mixer gate_output_8_407(.a(output_9_407), .b(output_9_8), .y(output_8_407));
wire output_10_407, output_10_8, output_9_407;
mixer gate_output_9_407(.a(output_10_407), .b(output_10_8), .y(output_9_407));
wire output_11_407, output_11_8, output_10_407;
mixer gate_output_10_407(.a(output_11_407), .b(output_11_8), .y(output_10_407));
wire output_12_407, output_12_8, output_11_407;
mixer gate_output_11_407(.a(output_12_407), .b(output_12_8), .y(output_11_407));
wire output_13_407, output_13_8, output_12_407;
mixer gate_output_12_407(.a(output_13_407), .b(output_13_8), .y(output_12_407));
wire output_14_407, output_14_8, output_13_407;
mixer gate_output_13_407(.a(output_14_407), .b(output_14_8), .y(output_13_407));
wire output_15_407, output_15_8, output_14_407;
mixer gate_output_14_407(.a(output_15_407), .b(output_15_8), .y(output_14_407));
wire output_16_407, output_16_8, output_15_407;
mixer gate_output_15_407(.a(output_16_407), .b(output_16_8), .y(output_15_407));
wire output_1_408, output_1_9, output_0_408;
mixer gate_output_0_408(.a(output_1_408), .b(output_1_9), .y(output_0_408));
wire output_2_408, output_2_9, output_1_408;
mixer gate_output_1_408(.a(output_2_408), .b(output_2_9), .y(output_1_408));
wire output_3_408, output_3_9, output_2_408;
mixer gate_output_2_408(.a(output_3_408), .b(output_3_9), .y(output_2_408));
wire output_4_408, output_4_9, output_3_408;
mixer gate_output_3_408(.a(output_4_408), .b(output_4_9), .y(output_3_408));
wire output_5_408, output_5_9, output_4_408;
mixer gate_output_4_408(.a(output_5_408), .b(output_5_9), .y(output_4_408));
wire output_6_408, output_6_9, output_5_408;
mixer gate_output_5_408(.a(output_6_408), .b(output_6_9), .y(output_5_408));
wire output_7_408, output_7_9, output_6_408;
mixer gate_output_6_408(.a(output_7_408), .b(output_7_9), .y(output_6_408));
wire output_8_408, output_8_9, output_7_408;
mixer gate_output_7_408(.a(output_8_408), .b(output_8_9), .y(output_7_408));
wire output_9_408, output_9_9, output_8_408;
mixer gate_output_8_408(.a(output_9_408), .b(output_9_9), .y(output_8_408));
wire output_10_408, output_10_9, output_9_408;
mixer gate_output_9_408(.a(output_10_408), .b(output_10_9), .y(output_9_408));
wire output_11_408, output_11_9, output_10_408;
mixer gate_output_10_408(.a(output_11_408), .b(output_11_9), .y(output_10_408));
wire output_12_408, output_12_9, output_11_408;
mixer gate_output_11_408(.a(output_12_408), .b(output_12_9), .y(output_11_408));
wire output_13_408, output_13_9, output_12_408;
mixer gate_output_12_408(.a(output_13_408), .b(output_13_9), .y(output_12_408));
wire output_14_408, output_14_9, output_13_408;
mixer gate_output_13_408(.a(output_14_408), .b(output_14_9), .y(output_13_408));
wire output_15_408, output_15_9, output_14_408;
mixer gate_output_14_408(.a(output_15_408), .b(output_15_9), .y(output_14_408));
wire output_16_408, output_16_9, output_15_408;
mixer gate_output_15_408(.a(output_16_408), .b(output_16_9), .y(output_15_408));
wire output_1_409, output_1_10, output_0_409;
mixer gate_output_0_409(.a(output_1_409), .b(output_1_10), .y(output_0_409));
wire output_2_409, output_2_10, output_1_409;
mixer gate_output_1_409(.a(output_2_409), .b(output_2_10), .y(output_1_409));
wire output_3_409, output_3_10, output_2_409;
mixer gate_output_2_409(.a(output_3_409), .b(output_3_10), .y(output_2_409));
wire output_4_409, output_4_10, output_3_409;
mixer gate_output_3_409(.a(output_4_409), .b(output_4_10), .y(output_3_409));
wire output_5_409, output_5_10, output_4_409;
mixer gate_output_4_409(.a(output_5_409), .b(output_5_10), .y(output_4_409));
wire output_6_409, output_6_10, output_5_409;
mixer gate_output_5_409(.a(output_6_409), .b(output_6_10), .y(output_5_409));
wire output_7_409, output_7_10, output_6_409;
mixer gate_output_6_409(.a(output_7_409), .b(output_7_10), .y(output_6_409));
wire output_8_409, output_8_10, output_7_409;
mixer gate_output_7_409(.a(output_8_409), .b(output_8_10), .y(output_7_409));
wire output_9_409, output_9_10, output_8_409;
mixer gate_output_8_409(.a(output_9_409), .b(output_9_10), .y(output_8_409));
wire output_10_409, output_10_10, output_9_409;
mixer gate_output_9_409(.a(output_10_409), .b(output_10_10), .y(output_9_409));
wire output_11_409, output_11_10, output_10_409;
mixer gate_output_10_409(.a(output_11_409), .b(output_11_10), .y(output_10_409));
wire output_12_409, output_12_10, output_11_409;
mixer gate_output_11_409(.a(output_12_409), .b(output_12_10), .y(output_11_409));
wire output_13_409, output_13_10, output_12_409;
mixer gate_output_12_409(.a(output_13_409), .b(output_13_10), .y(output_12_409));
wire output_14_409, output_14_10, output_13_409;
mixer gate_output_13_409(.a(output_14_409), .b(output_14_10), .y(output_13_409));
wire output_15_409, output_15_10, output_14_409;
mixer gate_output_14_409(.a(output_15_409), .b(output_15_10), .y(output_14_409));
wire output_16_409, output_16_10, output_15_409;
mixer gate_output_15_409(.a(output_16_409), .b(output_16_10), .y(output_15_409));
wire output_1_410, output_1_11, output_0_410;
mixer gate_output_0_410(.a(output_1_410), .b(output_1_11), .y(output_0_410));
wire output_2_410, output_2_11, output_1_410;
mixer gate_output_1_410(.a(output_2_410), .b(output_2_11), .y(output_1_410));
wire output_3_410, output_3_11, output_2_410;
mixer gate_output_2_410(.a(output_3_410), .b(output_3_11), .y(output_2_410));
wire output_4_410, output_4_11, output_3_410;
mixer gate_output_3_410(.a(output_4_410), .b(output_4_11), .y(output_3_410));
wire output_5_410, output_5_11, output_4_410;
mixer gate_output_4_410(.a(output_5_410), .b(output_5_11), .y(output_4_410));
wire output_6_410, output_6_11, output_5_410;
mixer gate_output_5_410(.a(output_6_410), .b(output_6_11), .y(output_5_410));
wire output_7_410, output_7_11, output_6_410;
mixer gate_output_6_410(.a(output_7_410), .b(output_7_11), .y(output_6_410));
wire output_8_410, output_8_11, output_7_410;
mixer gate_output_7_410(.a(output_8_410), .b(output_8_11), .y(output_7_410));
wire output_9_410, output_9_11, output_8_410;
mixer gate_output_8_410(.a(output_9_410), .b(output_9_11), .y(output_8_410));
wire output_10_410, output_10_11, output_9_410;
mixer gate_output_9_410(.a(output_10_410), .b(output_10_11), .y(output_9_410));
wire output_11_410, output_11_11, output_10_410;
mixer gate_output_10_410(.a(output_11_410), .b(output_11_11), .y(output_10_410));
wire output_12_410, output_12_11, output_11_410;
mixer gate_output_11_410(.a(output_12_410), .b(output_12_11), .y(output_11_410));
wire output_13_410, output_13_11, output_12_410;
mixer gate_output_12_410(.a(output_13_410), .b(output_13_11), .y(output_12_410));
wire output_14_410, output_14_11, output_13_410;
mixer gate_output_13_410(.a(output_14_410), .b(output_14_11), .y(output_13_410));
wire output_15_410, output_15_11, output_14_410;
mixer gate_output_14_410(.a(output_15_410), .b(output_15_11), .y(output_14_410));
wire output_16_410, output_16_11, output_15_410;
mixer gate_output_15_410(.a(output_16_410), .b(output_16_11), .y(output_15_410));
wire output_1_411, output_1_12, output_0_411;
mixer gate_output_0_411(.a(output_1_411), .b(output_1_12), .y(output_0_411));
wire output_2_411, output_2_12, output_1_411;
mixer gate_output_1_411(.a(output_2_411), .b(output_2_12), .y(output_1_411));
wire output_3_411, output_3_12, output_2_411;
mixer gate_output_2_411(.a(output_3_411), .b(output_3_12), .y(output_2_411));
wire output_4_411, output_4_12, output_3_411;
mixer gate_output_3_411(.a(output_4_411), .b(output_4_12), .y(output_3_411));
wire output_5_411, output_5_12, output_4_411;
mixer gate_output_4_411(.a(output_5_411), .b(output_5_12), .y(output_4_411));
wire output_6_411, output_6_12, output_5_411;
mixer gate_output_5_411(.a(output_6_411), .b(output_6_12), .y(output_5_411));
wire output_7_411, output_7_12, output_6_411;
mixer gate_output_6_411(.a(output_7_411), .b(output_7_12), .y(output_6_411));
wire output_8_411, output_8_12, output_7_411;
mixer gate_output_7_411(.a(output_8_411), .b(output_8_12), .y(output_7_411));
wire output_9_411, output_9_12, output_8_411;
mixer gate_output_8_411(.a(output_9_411), .b(output_9_12), .y(output_8_411));
wire output_10_411, output_10_12, output_9_411;
mixer gate_output_9_411(.a(output_10_411), .b(output_10_12), .y(output_9_411));
wire output_11_411, output_11_12, output_10_411;
mixer gate_output_10_411(.a(output_11_411), .b(output_11_12), .y(output_10_411));
wire output_12_411, output_12_12, output_11_411;
mixer gate_output_11_411(.a(output_12_411), .b(output_12_12), .y(output_11_411));
wire output_13_411, output_13_12, output_12_411;
mixer gate_output_12_411(.a(output_13_411), .b(output_13_12), .y(output_12_411));
wire output_14_411, output_14_12, output_13_411;
mixer gate_output_13_411(.a(output_14_411), .b(output_14_12), .y(output_13_411));
wire output_15_411, output_15_12, output_14_411;
mixer gate_output_14_411(.a(output_15_411), .b(output_15_12), .y(output_14_411));
wire output_16_411, output_16_12, output_15_411;
mixer gate_output_15_411(.a(output_16_411), .b(output_16_12), .y(output_15_411));
wire output_1_412, output_1_13, output_0_412;
mixer gate_output_0_412(.a(output_1_412), .b(output_1_13), .y(output_0_412));
wire output_2_412, output_2_13, output_1_412;
mixer gate_output_1_412(.a(output_2_412), .b(output_2_13), .y(output_1_412));
wire output_3_412, output_3_13, output_2_412;
mixer gate_output_2_412(.a(output_3_412), .b(output_3_13), .y(output_2_412));
wire output_4_412, output_4_13, output_3_412;
mixer gate_output_3_412(.a(output_4_412), .b(output_4_13), .y(output_3_412));
wire output_5_412, output_5_13, output_4_412;
mixer gate_output_4_412(.a(output_5_412), .b(output_5_13), .y(output_4_412));
wire output_6_412, output_6_13, output_5_412;
mixer gate_output_5_412(.a(output_6_412), .b(output_6_13), .y(output_5_412));
wire output_7_412, output_7_13, output_6_412;
mixer gate_output_6_412(.a(output_7_412), .b(output_7_13), .y(output_6_412));
wire output_8_412, output_8_13, output_7_412;
mixer gate_output_7_412(.a(output_8_412), .b(output_8_13), .y(output_7_412));
wire output_9_412, output_9_13, output_8_412;
mixer gate_output_8_412(.a(output_9_412), .b(output_9_13), .y(output_8_412));
wire output_10_412, output_10_13, output_9_412;
mixer gate_output_9_412(.a(output_10_412), .b(output_10_13), .y(output_9_412));
wire output_11_412, output_11_13, output_10_412;
mixer gate_output_10_412(.a(output_11_412), .b(output_11_13), .y(output_10_412));
wire output_12_412, output_12_13, output_11_412;
mixer gate_output_11_412(.a(output_12_412), .b(output_12_13), .y(output_11_412));
wire output_13_412, output_13_13, output_12_412;
mixer gate_output_12_412(.a(output_13_412), .b(output_13_13), .y(output_12_412));
wire output_14_412, output_14_13, output_13_412;
mixer gate_output_13_412(.a(output_14_412), .b(output_14_13), .y(output_13_412));
wire output_15_412, output_15_13, output_14_412;
mixer gate_output_14_412(.a(output_15_412), .b(output_15_13), .y(output_14_412));
wire output_16_412, output_16_13, output_15_412;
mixer gate_output_15_412(.a(output_16_412), .b(output_16_13), .y(output_15_412));
wire output_1_413, output_1_14, output_0_413;
mixer gate_output_0_413(.a(output_1_413), .b(output_1_14), .y(output_0_413));
wire output_2_413, output_2_14, output_1_413;
mixer gate_output_1_413(.a(output_2_413), .b(output_2_14), .y(output_1_413));
wire output_3_413, output_3_14, output_2_413;
mixer gate_output_2_413(.a(output_3_413), .b(output_3_14), .y(output_2_413));
wire output_4_413, output_4_14, output_3_413;
mixer gate_output_3_413(.a(output_4_413), .b(output_4_14), .y(output_3_413));
wire output_5_413, output_5_14, output_4_413;
mixer gate_output_4_413(.a(output_5_413), .b(output_5_14), .y(output_4_413));
wire output_6_413, output_6_14, output_5_413;
mixer gate_output_5_413(.a(output_6_413), .b(output_6_14), .y(output_5_413));
wire output_7_413, output_7_14, output_6_413;
mixer gate_output_6_413(.a(output_7_413), .b(output_7_14), .y(output_6_413));
wire output_8_413, output_8_14, output_7_413;
mixer gate_output_7_413(.a(output_8_413), .b(output_8_14), .y(output_7_413));
wire output_9_413, output_9_14, output_8_413;
mixer gate_output_8_413(.a(output_9_413), .b(output_9_14), .y(output_8_413));
wire output_10_413, output_10_14, output_9_413;
mixer gate_output_9_413(.a(output_10_413), .b(output_10_14), .y(output_9_413));
wire output_11_413, output_11_14, output_10_413;
mixer gate_output_10_413(.a(output_11_413), .b(output_11_14), .y(output_10_413));
wire output_12_413, output_12_14, output_11_413;
mixer gate_output_11_413(.a(output_12_413), .b(output_12_14), .y(output_11_413));
wire output_13_413, output_13_14, output_12_413;
mixer gate_output_12_413(.a(output_13_413), .b(output_13_14), .y(output_12_413));
wire output_14_413, output_14_14, output_13_413;
mixer gate_output_13_413(.a(output_14_413), .b(output_14_14), .y(output_13_413));
wire output_15_413, output_15_14, output_14_413;
mixer gate_output_14_413(.a(output_15_413), .b(output_15_14), .y(output_14_413));
wire output_16_413, output_16_14, output_15_413;
mixer gate_output_15_413(.a(output_16_413), .b(output_16_14), .y(output_15_413));
wire output_1_414, output_1_15, output_0_414;
mixer gate_output_0_414(.a(output_1_414), .b(output_1_15), .y(output_0_414));
wire output_2_414, output_2_15, output_1_414;
mixer gate_output_1_414(.a(output_2_414), .b(output_2_15), .y(output_1_414));
wire output_3_414, output_3_15, output_2_414;
mixer gate_output_2_414(.a(output_3_414), .b(output_3_15), .y(output_2_414));
wire output_4_414, output_4_15, output_3_414;
mixer gate_output_3_414(.a(output_4_414), .b(output_4_15), .y(output_3_414));
wire output_5_414, output_5_15, output_4_414;
mixer gate_output_4_414(.a(output_5_414), .b(output_5_15), .y(output_4_414));
wire output_6_414, output_6_15, output_5_414;
mixer gate_output_5_414(.a(output_6_414), .b(output_6_15), .y(output_5_414));
wire output_7_414, output_7_15, output_6_414;
mixer gate_output_6_414(.a(output_7_414), .b(output_7_15), .y(output_6_414));
wire output_8_414, output_8_15, output_7_414;
mixer gate_output_7_414(.a(output_8_414), .b(output_8_15), .y(output_7_414));
wire output_9_414, output_9_15, output_8_414;
mixer gate_output_8_414(.a(output_9_414), .b(output_9_15), .y(output_8_414));
wire output_10_414, output_10_15, output_9_414;
mixer gate_output_9_414(.a(output_10_414), .b(output_10_15), .y(output_9_414));
wire output_11_414, output_11_15, output_10_414;
mixer gate_output_10_414(.a(output_11_414), .b(output_11_15), .y(output_10_414));
wire output_12_414, output_12_15, output_11_414;
mixer gate_output_11_414(.a(output_12_414), .b(output_12_15), .y(output_11_414));
wire output_13_414, output_13_15, output_12_414;
mixer gate_output_12_414(.a(output_13_414), .b(output_13_15), .y(output_12_414));
wire output_14_414, output_14_15, output_13_414;
mixer gate_output_13_414(.a(output_14_414), .b(output_14_15), .y(output_13_414));
wire output_15_414, output_15_15, output_14_414;
mixer gate_output_14_414(.a(output_15_414), .b(output_15_15), .y(output_14_414));
wire output_16_414, output_16_15, output_15_414;
mixer gate_output_15_414(.a(output_16_414), .b(output_16_15), .y(output_15_414));
wire output_1_415, output_1_0, output_0_415;
mixer gate_output_0_415(.a(output_1_415), .b(output_1_0), .y(output_0_415));
wire output_2_415, output_2_0, output_1_415;
mixer gate_output_1_415(.a(output_2_415), .b(output_2_0), .y(output_1_415));
wire output_3_415, output_3_0, output_2_415;
mixer gate_output_2_415(.a(output_3_415), .b(output_3_0), .y(output_2_415));
wire output_4_415, output_4_0, output_3_415;
mixer gate_output_3_415(.a(output_4_415), .b(output_4_0), .y(output_3_415));
wire output_5_415, output_5_0, output_4_415;
mixer gate_output_4_415(.a(output_5_415), .b(output_5_0), .y(output_4_415));
wire output_6_415, output_6_0, output_5_415;
mixer gate_output_5_415(.a(output_6_415), .b(output_6_0), .y(output_5_415));
wire output_7_415, output_7_0, output_6_415;
mixer gate_output_6_415(.a(output_7_415), .b(output_7_0), .y(output_6_415));
wire output_8_415, output_8_0, output_7_415;
mixer gate_output_7_415(.a(output_8_415), .b(output_8_0), .y(output_7_415));
wire output_9_415, output_9_0, output_8_415;
mixer gate_output_8_415(.a(output_9_415), .b(output_9_0), .y(output_8_415));
wire output_10_415, output_10_0, output_9_415;
mixer gate_output_9_415(.a(output_10_415), .b(output_10_0), .y(output_9_415));
wire output_11_415, output_11_0, output_10_415;
mixer gate_output_10_415(.a(output_11_415), .b(output_11_0), .y(output_10_415));
wire output_12_415, output_12_0, output_11_415;
mixer gate_output_11_415(.a(output_12_415), .b(output_12_0), .y(output_11_415));
wire output_13_415, output_13_0, output_12_415;
mixer gate_output_12_415(.a(output_13_415), .b(output_13_0), .y(output_12_415));
wire output_14_415, output_14_0, output_13_415;
mixer gate_output_13_415(.a(output_14_415), .b(output_14_0), .y(output_13_415));
wire output_15_415, output_15_0, output_14_415;
mixer gate_output_14_415(.a(output_15_415), .b(output_15_0), .y(output_14_415));
wire output_16_415, output_16_0, output_15_415;
mixer gate_output_15_415(.a(output_16_415), .b(output_16_0), .y(output_15_415));
wire output_1_416, output_1_1, output_0_416;
mixer gate_output_0_416(.a(output_1_416), .b(output_1_1), .y(output_0_416));
wire output_2_416, output_2_1, output_1_416;
mixer gate_output_1_416(.a(output_2_416), .b(output_2_1), .y(output_1_416));
wire output_3_416, output_3_1, output_2_416;
mixer gate_output_2_416(.a(output_3_416), .b(output_3_1), .y(output_2_416));
wire output_4_416, output_4_1, output_3_416;
mixer gate_output_3_416(.a(output_4_416), .b(output_4_1), .y(output_3_416));
wire output_5_416, output_5_1, output_4_416;
mixer gate_output_4_416(.a(output_5_416), .b(output_5_1), .y(output_4_416));
wire output_6_416, output_6_1, output_5_416;
mixer gate_output_5_416(.a(output_6_416), .b(output_6_1), .y(output_5_416));
wire output_7_416, output_7_1, output_6_416;
mixer gate_output_6_416(.a(output_7_416), .b(output_7_1), .y(output_6_416));
wire output_8_416, output_8_1, output_7_416;
mixer gate_output_7_416(.a(output_8_416), .b(output_8_1), .y(output_7_416));
wire output_9_416, output_9_1, output_8_416;
mixer gate_output_8_416(.a(output_9_416), .b(output_9_1), .y(output_8_416));
wire output_10_416, output_10_1, output_9_416;
mixer gate_output_9_416(.a(output_10_416), .b(output_10_1), .y(output_9_416));
wire output_11_416, output_11_1, output_10_416;
mixer gate_output_10_416(.a(output_11_416), .b(output_11_1), .y(output_10_416));
wire output_12_416, output_12_1, output_11_416;
mixer gate_output_11_416(.a(output_12_416), .b(output_12_1), .y(output_11_416));
wire output_13_416, output_13_1, output_12_416;
mixer gate_output_12_416(.a(output_13_416), .b(output_13_1), .y(output_12_416));
wire output_14_416, output_14_1, output_13_416;
mixer gate_output_13_416(.a(output_14_416), .b(output_14_1), .y(output_13_416));
wire output_15_416, output_15_1, output_14_416;
mixer gate_output_14_416(.a(output_15_416), .b(output_15_1), .y(output_14_416));
wire output_16_416, output_16_1, output_15_416;
mixer gate_output_15_416(.a(output_16_416), .b(output_16_1), .y(output_15_416));
wire output_1_417, output_1_2, output_0_417;
mixer gate_output_0_417(.a(output_1_417), .b(output_1_2), .y(output_0_417));
wire output_2_417, output_2_2, output_1_417;
mixer gate_output_1_417(.a(output_2_417), .b(output_2_2), .y(output_1_417));
wire output_3_417, output_3_2, output_2_417;
mixer gate_output_2_417(.a(output_3_417), .b(output_3_2), .y(output_2_417));
wire output_4_417, output_4_2, output_3_417;
mixer gate_output_3_417(.a(output_4_417), .b(output_4_2), .y(output_3_417));
wire output_5_417, output_5_2, output_4_417;
mixer gate_output_4_417(.a(output_5_417), .b(output_5_2), .y(output_4_417));
wire output_6_417, output_6_2, output_5_417;
mixer gate_output_5_417(.a(output_6_417), .b(output_6_2), .y(output_5_417));
wire output_7_417, output_7_2, output_6_417;
mixer gate_output_6_417(.a(output_7_417), .b(output_7_2), .y(output_6_417));
wire output_8_417, output_8_2, output_7_417;
mixer gate_output_7_417(.a(output_8_417), .b(output_8_2), .y(output_7_417));
wire output_9_417, output_9_2, output_8_417;
mixer gate_output_8_417(.a(output_9_417), .b(output_9_2), .y(output_8_417));
wire output_10_417, output_10_2, output_9_417;
mixer gate_output_9_417(.a(output_10_417), .b(output_10_2), .y(output_9_417));
wire output_11_417, output_11_2, output_10_417;
mixer gate_output_10_417(.a(output_11_417), .b(output_11_2), .y(output_10_417));
wire output_12_417, output_12_2, output_11_417;
mixer gate_output_11_417(.a(output_12_417), .b(output_12_2), .y(output_11_417));
wire output_13_417, output_13_2, output_12_417;
mixer gate_output_12_417(.a(output_13_417), .b(output_13_2), .y(output_12_417));
wire output_14_417, output_14_2, output_13_417;
mixer gate_output_13_417(.a(output_14_417), .b(output_14_2), .y(output_13_417));
wire output_15_417, output_15_2, output_14_417;
mixer gate_output_14_417(.a(output_15_417), .b(output_15_2), .y(output_14_417));
wire output_16_417, output_16_2, output_15_417;
mixer gate_output_15_417(.a(output_16_417), .b(output_16_2), .y(output_15_417));
wire output_1_418, output_1_3, output_0_418;
mixer gate_output_0_418(.a(output_1_418), .b(output_1_3), .y(output_0_418));
wire output_2_418, output_2_3, output_1_418;
mixer gate_output_1_418(.a(output_2_418), .b(output_2_3), .y(output_1_418));
wire output_3_418, output_3_3, output_2_418;
mixer gate_output_2_418(.a(output_3_418), .b(output_3_3), .y(output_2_418));
wire output_4_418, output_4_3, output_3_418;
mixer gate_output_3_418(.a(output_4_418), .b(output_4_3), .y(output_3_418));
wire output_5_418, output_5_3, output_4_418;
mixer gate_output_4_418(.a(output_5_418), .b(output_5_3), .y(output_4_418));
wire output_6_418, output_6_3, output_5_418;
mixer gate_output_5_418(.a(output_6_418), .b(output_6_3), .y(output_5_418));
wire output_7_418, output_7_3, output_6_418;
mixer gate_output_6_418(.a(output_7_418), .b(output_7_3), .y(output_6_418));
wire output_8_418, output_8_3, output_7_418;
mixer gate_output_7_418(.a(output_8_418), .b(output_8_3), .y(output_7_418));
wire output_9_418, output_9_3, output_8_418;
mixer gate_output_8_418(.a(output_9_418), .b(output_9_3), .y(output_8_418));
wire output_10_418, output_10_3, output_9_418;
mixer gate_output_9_418(.a(output_10_418), .b(output_10_3), .y(output_9_418));
wire output_11_418, output_11_3, output_10_418;
mixer gate_output_10_418(.a(output_11_418), .b(output_11_3), .y(output_10_418));
wire output_12_418, output_12_3, output_11_418;
mixer gate_output_11_418(.a(output_12_418), .b(output_12_3), .y(output_11_418));
wire output_13_418, output_13_3, output_12_418;
mixer gate_output_12_418(.a(output_13_418), .b(output_13_3), .y(output_12_418));
wire output_14_418, output_14_3, output_13_418;
mixer gate_output_13_418(.a(output_14_418), .b(output_14_3), .y(output_13_418));
wire output_15_418, output_15_3, output_14_418;
mixer gate_output_14_418(.a(output_15_418), .b(output_15_3), .y(output_14_418));
wire output_16_418, output_16_3, output_15_418;
mixer gate_output_15_418(.a(output_16_418), .b(output_16_3), .y(output_15_418));
wire output_1_419, output_1_4, output_0_419;
mixer gate_output_0_419(.a(output_1_419), .b(output_1_4), .y(output_0_419));
wire output_2_419, output_2_4, output_1_419;
mixer gate_output_1_419(.a(output_2_419), .b(output_2_4), .y(output_1_419));
wire output_3_419, output_3_4, output_2_419;
mixer gate_output_2_419(.a(output_3_419), .b(output_3_4), .y(output_2_419));
wire output_4_419, output_4_4, output_3_419;
mixer gate_output_3_419(.a(output_4_419), .b(output_4_4), .y(output_3_419));
wire output_5_419, output_5_4, output_4_419;
mixer gate_output_4_419(.a(output_5_419), .b(output_5_4), .y(output_4_419));
wire output_6_419, output_6_4, output_5_419;
mixer gate_output_5_419(.a(output_6_419), .b(output_6_4), .y(output_5_419));
wire output_7_419, output_7_4, output_6_419;
mixer gate_output_6_419(.a(output_7_419), .b(output_7_4), .y(output_6_419));
wire output_8_419, output_8_4, output_7_419;
mixer gate_output_7_419(.a(output_8_419), .b(output_8_4), .y(output_7_419));
wire output_9_419, output_9_4, output_8_419;
mixer gate_output_8_419(.a(output_9_419), .b(output_9_4), .y(output_8_419));
wire output_10_419, output_10_4, output_9_419;
mixer gate_output_9_419(.a(output_10_419), .b(output_10_4), .y(output_9_419));
wire output_11_419, output_11_4, output_10_419;
mixer gate_output_10_419(.a(output_11_419), .b(output_11_4), .y(output_10_419));
wire output_12_419, output_12_4, output_11_419;
mixer gate_output_11_419(.a(output_12_419), .b(output_12_4), .y(output_11_419));
wire output_13_419, output_13_4, output_12_419;
mixer gate_output_12_419(.a(output_13_419), .b(output_13_4), .y(output_12_419));
wire output_14_419, output_14_4, output_13_419;
mixer gate_output_13_419(.a(output_14_419), .b(output_14_4), .y(output_13_419));
wire output_15_419, output_15_4, output_14_419;
mixer gate_output_14_419(.a(output_15_419), .b(output_15_4), .y(output_14_419));
wire output_16_419, output_16_4, output_15_419;
mixer gate_output_15_419(.a(output_16_419), .b(output_16_4), .y(output_15_419));
wire output_1_420, output_1_5, output_0_420;
mixer gate_output_0_420(.a(output_1_420), .b(output_1_5), .y(output_0_420));
wire output_2_420, output_2_5, output_1_420;
mixer gate_output_1_420(.a(output_2_420), .b(output_2_5), .y(output_1_420));
wire output_3_420, output_3_5, output_2_420;
mixer gate_output_2_420(.a(output_3_420), .b(output_3_5), .y(output_2_420));
wire output_4_420, output_4_5, output_3_420;
mixer gate_output_3_420(.a(output_4_420), .b(output_4_5), .y(output_3_420));
wire output_5_420, output_5_5, output_4_420;
mixer gate_output_4_420(.a(output_5_420), .b(output_5_5), .y(output_4_420));
wire output_6_420, output_6_5, output_5_420;
mixer gate_output_5_420(.a(output_6_420), .b(output_6_5), .y(output_5_420));
wire output_7_420, output_7_5, output_6_420;
mixer gate_output_6_420(.a(output_7_420), .b(output_7_5), .y(output_6_420));
wire output_8_420, output_8_5, output_7_420;
mixer gate_output_7_420(.a(output_8_420), .b(output_8_5), .y(output_7_420));
wire output_9_420, output_9_5, output_8_420;
mixer gate_output_8_420(.a(output_9_420), .b(output_9_5), .y(output_8_420));
wire output_10_420, output_10_5, output_9_420;
mixer gate_output_9_420(.a(output_10_420), .b(output_10_5), .y(output_9_420));
wire output_11_420, output_11_5, output_10_420;
mixer gate_output_10_420(.a(output_11_420), .b(output_11_5), .y(output_10_420));
wire output_12_420, output_12_5, output_11_420;
mixer gate_output_11_420(.a(output_12_420), .b(output_12_5), .y(output_11_420));
wire output_13_420, output_13_5, output_12_420;
mixer gate_output_12_420(.a(output_13_420), .b(output_13_5), .y(output_12_420));
wire output_14_420, output_14_5, output_13_420;
mixer gate_output_13_420(.a(output_14_420), .b(output_14_5), .y(output_13_420));
wire output_15_420, output_15_5, output_14_420;
mixer gate_output_14_420(.a(output_15_420), .b(output_15_5), .y(output_14_420));
wire output_16_420, output_16_5, output_15_420;
mixer gate_output_15_420(.a(output_16_420), .b(output_16_5), .y(output_15_420));
wire output_1_421, output_1_6, output_0_421;
mixer gate_output_0_421(.a(output_1_421), .b(output_1_6), .y(output_0_421));
wire output_2_421, output_2_6, output_1_421;
mixer gate_output_1_421(.a(output_2_421), .b(output_2_6), .y(output_1_421));
wire output_3_421, output_3_6, output_2_421;
mixer gate_output_2_421(.a(output_3_421), .b(output_3_6), .y(output_2_421));
wire output_4_421, output_4_6, output_3_421;
mixer gate_output_3_421(.a(output_4_421), .b(output_4_6), .y(output_3_421));
wire output_5_421, output_5_6, output_4_421;
mixer gate_output_4_421(.a(output_5_421), .b(output_5_6), .y(output_4_421));
wire output_6_421, output_6_6, output_5_421;
mixer gate_output_5_421(.a(output_6_421), .b(output_6_6), .y(output_5_421));
wire output_7_421, output_7_6, output_6_421;
mixer gate_output_6_421(.a(output_7_421), .b(output_7_6), .y(output_6_421));
wire output_8_421, output_8_6, output_7_421;
mixer gate_output_7_421(.a(output_8_421), .b(output_8_6), .y(output_7_421));
wire output_9_421, output_9_6, output_8_421;
mixer gate_output_8_421(.a(output_9_421), .b(output_9_6), .y(output_8_421));
wire output_10_421, output_10_6, output_9_421;
mixer gate_output_9_421(.a(output_10_421), .b(output_10_6), .y(output_9_421));
wire output_11_421, output_11_6, output_10_421;
mixer gate_output_10_421(.a(output_11_421), .b(output_11_6), .y(output_10_421));
wire output_12_421, output_12_6, output_11_421;
mixer gate_output_11_421(.a(output_12_421), .b(output_12_6), .y(output_11_421));
wire output_13_421, output_13_6, output_12_421;
mixer gate_output_12_421(.a(output_13_421), .b(output_13_6), .y(output_12_421));
wire output_14_421, output_14_6, output_13_421;
mixer gate_output_13_421(.a(output_14_421), .b(output_14_6), .y(output_13_421));
wire output_15_421, output_15_6, output_14_421;
mixer gate_output_14_421(.a(output_15_421), .b(output_15_6), .y(output_14_421));
wire output_16_421, output_16_6, output_15_421;
mixer gate_output_15_421(.a(output_16_421), .b(output_16_6), .y(output_15_421));
wire output_1_422, output_1_7, output_0_422;
mixer gate_output_0_422(.a(output_1_422), .b(output_1_7), .y(output_0_422));
wire output_2_422, output_2_7, output_1_422;
mixer gate_output_1_422(.a(output_2_422), .b(output_2_7), .y(output_1_422));
wire output_3_422, output_3_7, output_2_422;
mixer gate_output_2_422(.a(output_3_422), .b(output_3_7), .y(output_2_422));
wire output_4_422, output_4_7, output_3_422;
mixer gate_output_3_422(.a(output_4_422), .b(output_4_7), .y(output_3_422));
wire output_5_422, output_5_7, output_4_422;
mixer gate_output_4_422(.a(output_5_422), .b(output_5_7), .y(output_4_422));
wire output_6_422, output_6_7, output_5_422;
mixer gate_output_5_422(.a(output_6_422), .b(output_6_7), .y(output_5_422));
wire output_7_422, output_7_7, output_6_422;
mixer gate_output_6_422(.a(output_7_422), .b(output_7_7), .y(output_6_422));
wire output_8_422, output_8_7, output_7_422;
mixer gate_output_7_422(.a(output_8_422), .b(output_8_7), .y(output_7_422));
wire output_9_422, output_9_7, output_8_422;
mixer gate_output_8_422(.a(output_9_422), .b(output_9_7), .y(output_8_422));
wire output_10_422, output_10_7, output_9_422;
mixer gate_output_9_422(.a(output_10_422), .b(output_10_7), .y(output_9_422));
wire output_11_422, output_11_7, output_10_422;
mixer gate_output_10_422(.a(output_11_422), .b(output_11_7), .y(output_10_422));
wire output_12_422, output_12_7, output_11_422;
mixer gate_output_11_422(.a(output_12_422), .b(output_12_7), .y(output_11_422));
wire output_13_422, output_13_7, output_12_422;
mixer gate_output_12_422(.a(output_13_422), .b(output_13_7), .y(output_12_422));
wire output_14_422, output_14_7, output_13_422;
mixer gate_output_13_422(.a(output_14_422), .b(output_14_7), .y(output_13_422));
wire output_15_422, output_15_7, output_14_422;
mixer gate_output_14_422(.a(output_15_422), .b(output_15_7), .y(output_14_422));
wire output_16_422, output_16_7, output_15_422;
mixer gate_output_15_422(.a(output_16_422), .b(output_16_7), .y(output_15_422));
wire output_1_423, output_1_8, output_0_423;
mixer gate_output_0_423(.a(output_1_423), .b(output_1_8), .y(output_0_423));
wire output_2_423, output_2_8, output_1_423;
mixer gate_output_1_423(.a(output_2_423), .b(output_2_8), .y(output_1_423));
wire output_3_423, output_3_8, output_2_423;
mixer gate_output_2_423(.a(output_3_423), .b(output_3_8), .y(output_2_423));
wire output_4_423, output_4_8, output_3_423;
mixer gate_output_3_423(.a(output_4_423), .b(output_4_8), .y(output_3_423));
wire output_5_423, output_5_8, output_4_423;
mixer gate_output_4_423(.a(output_5_423), .b(output_5_8), .y(output_4_423));
wire output_6_423, output_6_8, output_5_423;
mixer gate_output_5_423(.a(output_6_423), .b(output_6_8), .y(output_5_423));
wire output_7_423, output_7_8, output_6_423;
mixer gate_output_6_423(.a(output_7_423), .b(output_7_8), .y(output_6_423));
wire output_8_423, output_8_8, output_7_423;
mixer gate_output_7_423(.a(output_8_423), .b(output_8_8), .y(output_7_423));
wire output_9_423, output_9_8, output_8_423;
mixer gate_output_8_423(.a(output_9_423), .b(output_9_8), .y(output_8_423));
wire output_10_423, output_10_8, output_9_423;
mixer gate_output_9_423(.a(output_10_423), .b(output_10_8), .y(output_9_423));
wire output_11_423, output_11_8, output_10_423;
mixer gate_output_10_423(.a(output_11_423), .b(output_11_8), .y(output_10_423));
wire output_12_423, output_12_8, output_11_423;
mixer gate_output_11_423(.a(output_12_423), .b(output_12_8), .y(output_11_423));
wire output_13_423, output_13_8, output_12_423;
mixer gate_output_12_423(.a(output_13_423), .b(output_13_8), .y(output_12_423));
wire output_14_423, output_14_8, output_13_423;
mixer gate_output_13_423(.a(output_14_423), .b(output_14_8), .y(output_13_423));
wire output_15_423, output_15_8, output_14_423;
mixer gate_output_14_423(.a(output_15_423), .b(output_15_8), .y(output_14_423));
wire output_16_423, output_16_8, output_15_423;
mixer gate_output_15_423(.a(output_16_423), .b(output_16_8), .y(output_15_423));
wire output_1_424, output_1_9, output_0_424;
mixer gate_output_0_424(.a(output_1_424), .b(output_1_9), .y(output_0_424));
wire output_2_424, output_2_9, output_1_424;
mixer gate_output_1_424(.a(output_2_424), .b(output_2_9), .y(output_1_424));
wire output_3_424, output_3_9, output_2_424;
mixer gate_output_2_424(.a(output_3_424), .b(output_3_9), .y(output_2_424));
wire output_4_424, output_4_9, output_3_424;
mixer gate_output_3_424(.a(output_4_424), .b(output_4_9), .y(output_3_424));
wire output_5_424, output_5_9, output_4_424;
mixer gate_output_4_424(.a(output_5_424), .b(output_5_9), .y(output_4_424));
wire output_6_424, output_6_9, output_5_424;
mixer gate_output_5_424(.a(output_6_424), .b(output_6_9), .y(output_5_424));
wire output_7_424, output_7_9, output_6_424;
mixer gate_output_6_424(.a(output_7_424), .b(output_7_9), .y(output_6_424));
wire output_8_424, output_8_9, output_7_424;
mixer gate_output_7_424(.a(output_8_424), .b(output_8_9), .y(output_7_424));
wire output_9_424, output_9_9, output_8_424;
mixer gate_output_8_424(.a(output_9_424), .b(output_9_9), .y(output_8_424));
wire output_10_424, output_10_9, output_9_424;
mixer gate_output_9_424(.a(output_10_424), .b(output_10_9), .y(output_9_424));
wire output_11_424, output_11_9, output_10_424;
mixer gate_output_10_424(.a(output_11_424), .b(output_11_9), .y(output_10_424));
wire output_12_424, output_12_9, output_11_424;
mixer gate_output_11_424(.a(output_12_424), .b(output_12_9), .y(output_11_424));
wire output_13_424, output_13_9, output_12_424;
mixer gate_output_12_424(.a(output_13_424), .b(output_13_9), .y(output_12_424));
wire output_14_424, output_14_9, output_13_424;
mixer gate_output_13_424(.a(output_14_424), .b(output_14_9), .y(output_13_424));
wire output_15_424, output_15_9, output_14_424;
mixer gate_output_14_424(.a(output_15_424), .b(output_15_9), .y(output_14_424));
wire output_16_424, output_16_9, output_15_424;
mixer gate_output_15_424(.a(output_16_424), .b(output_16_9), .y(output_15_424));
wire output_1_425, output_1_10, output_0_425;
mixer gate_output_0_425(.a(output_1_425), .b(output_1_10), .y(output_0_425));
wire output_2_425, output_2_10, output_1_425;
mixer gate_output_1_425(.a(output_2_425), .b(output_2_10), .y(output_1_425));
wire output_3_425, output_3_10, output_2_425;
mixer gate_output_2_425(.a(output_3_425), .b(output_3_10), .y(output_2_425));
wire output_4_425, output_4_10, output_3_425;
mixer gate_output_3_425(.a(output_4_425), .b(output_4_10), .y(output_3_425));
wire output_5_425, output_5_10, output_4_425;
mixer gate_output_4_425(.a(output_5_425), .b(output_5_10), .y(output_4_425));
wire output_6_425, output_6_10, output_5_425;
mixer gate_output_5_425(.a(output_6_425), .b(output_6_10), .y(output_5_425));
wire output_7_425, output_7_10, output_6_425;
mixer gate_output_6_425(.a(output_7_425), .b(output_7_10), .y(output_6_425));
wire output_8_425, output_8_10, output_7_425;
mixer gate_output_7_425(.a(output_8_425), .b(output_8_10), .y(output_7_425));
wire output_9_425, output_9_10, output_8_425;
mixer gate_output_8_425(.a(output_9_425), .b(output_9_10), .y(output_8_425));
wire output_10_425, output_10_10, output_9_425;
mixer gate_output_9_425(.a(output_10_425), .b(output_10_10), .y(output_9_425));
wire output_11_425, output_11_10, output_10_425;
mixer gate_output_10_425(.a(output_11_425), .b(output_11_10), .y(output_10_425));
wire output_12_425, output_12_10, output_11_425;
mixer gate_output_11_425(.a(output_12_425), .b(output_12_10), .y(output_11_425));
wire output_13_425, output_13_10, output_12_425;
mixer gate_output_12_425(.a(output_13_425), .b(output_13_10), .y(output_12_425));
wire output_14_425, output_14_10, output_13_425;
mixer gate_output_13_425(.a(output_14_425), .b(output_14_10), .y(output_13_425));
wire output_15_425, output_15_10, output_14_425;
mixer gate_output_14_425(.a(output_15_425), .b(output_15_10), .y(output_14_425));
wire output_16_425, output_16_10, output_15_425;
mixer gate_output_15_425(.a(output_16_425), .b(output_16_10), .y(output_15_425));
wire output_1_426, output_1_11, output_0_426;
mixer gate_output_0_426(.a(output_1_426), .b(output_1_11), .y(output_0_426));
wire output_2_426, output_2_11, output_1_426;
mixer gate_output_1_426(.a(output_2_426), .b(output_2_11), .y(output_1_426));
wire output_3_426, output_3_11, output_2_426;
mixer gate_output_2_426(.a(output_3_426), .b(output_3_11), .y(output_2_426));
wire output_4_426, output_4_11, output_3_426;
mixer gate_output_3_426(.a(output_4_426), .b(output_4_11), .y(output_3_426));
wire output_5_426, output_5_11, output_4_426;
mixer gate_output_4_426(.a(output_5_426), .b(output_5_11), .y(output_4_426));
wire output_6_426, output_6_11, output_5_426;
mixer gate_output_5_426(.a(output_6_426), .b(output_6_11), .y(output_5_426));
wire output_7_426, output_7_11, output_6_426;
mixer gate_output_6_426(.a(output_7_426), .b(output_7_11), .y(output_6_426));
wire output_8_426, output_8_11, output_7_426;
mixer gate_output_7_426(.a(output_8_426), .b(output_8_11), .y(output_7_426));
wire output_9_426, output_9_11, output_8_426;
mixer gate_output_8_426(.a(output_9_426), .b(output_9_11), .y(output_8_426));
wire output_10_426, output_10_11, output_9_426;
mixer gate_output_9_426(.a(output_10_426), .b(output_10_11), .y(output_9_426));
wire output_11_426, output_11_11, output_10_426;
mixer gate_output_10_426(.a(output_11_426), .b(output_11_11), .y(output_10_426));
wire output_12_426, output_12_11, output_11_426;
mixer gate_output_11_426(.a(output_12_426), .b(output_12_11), .y(output_11_426));
wire output_13_426, output_13_11, output_12_426;
mixer gate_output_12_426(.a(output_13_426), .b(output_13_11), .y(output_12_426));
wire output_14_426, output_14_11, output_13_426;
mixer gate_output_13_426(.a(output_14_426), .b(output_14_11), .y(output_13_426));
wire output_15_426, output_15_11, output_14_426;
mixer gate_output_14_426(.a(output_15_426), .b(output_15_11), .y(output_14_426));
wire output_16_426, output_16_11, output_15_426;
mixer gate_output_15_426(.a(output_16_426), .b(output_16_11), .y(output_15_426));
wire output_1_427, output_1_12, output_0_427;
mixer gate_output_0_427(.a(output_1_427), .b(output_1_12), .y(output_0_427));
wire output_2_427, output_2_12, output_1_427;
mixer gate_output_1_427(.a(output_2_427), .b(output_2_12), .y(output_1_427));
wire output_3_427, output_3_12, output_2_427;
mixer gate_output_2_427(.a(output_3_427), .b(output_3_12), .y(output_2_427));
wire output_4_427, output_4_12, output_3_427;
mixer gate_output_3_427(.a(output_4_427), .b(output_4_12), .y(output_3_427));
wire output_5_427, output_5_12, output_4_427;
mixer gate_output_4_427(.a(output_5_427), .b(output_5_12), .y(output_4_427));
wire output_6_427, output_6_12, output_5_427;
mixer gate_output_5_427(.a(output_6_427), .b(output_6_12), .y(output_5_427));
wire output_7_427, output_7_12, output_6_427;
mixer gate_output_6_427(.a(output_7_427), .b(output_7_12), .y(output_6_427));
wire output_8_427, output_8_12, output_7_427;
mixer gate_output_7_427(.a(output_8_427), .b(output_8_12), .y(output_7_427));
wire output_9_427, output_9_12, output_8_427;
mixer gate_output_8_427(.a(output_9_427), .b(output_9_12), .y(output_8_427));
wire output_10_427, output_10_12, output_9_427;
mixer gate_output_9_427(.a(output_10_427), .b(output_10_12), .y(output_9_427));
wire output_11_427, output_11_12, output_10_427;
mixer gate_output_10_427(.a(output_11_427), .b(output_11_12), .y(output_10_427));
wire output_12_427, output_12_12, output_11_427;
mixer gate_output_11_427(.a(output_12_427), .b(output_12_12), .y(output_11_427));
wire output_13_427, output_13_12, output_12_427;
mixer gate_output_12_427(.a(output_13_427), .b(output_13_12), .y(output_12_427));
wire output_14_427, output_14_12, output_13_427;
mixer gate_output_13_427(.a(output_14_427), .b(output_14_12), .y(output_13_427));
wire output_15_427, output_15_12, output_14_427;
mixer gate_output_14_427(.a(output_15_427), .b(output_15_12), .y(output_14_427));
wire output_16_427, output_16_12, output_15_427;
mixer gate_output_15_427(.a(output_16_427), .b(output_16_12), .y(output_15_427));
wire output_1_428, output_1_13, output_0_428;
mixer gate_output_0_428(.a(output_1_428), .b(output_1_13), .y(output_0_428));
wire output_2_428, output_2_13, output_1_428;
mixer gate_output_1_428(.a(output_2_428), .b(output_2_13), .y(output_1_428));
wire output_3_428, output_3_13, output_2_428;
mixer gate_output_2_428(.a(output_3_428), .b(output_3_13), .y(output_2_428));
wire output_4_428, output_4_13, output_3_428;
mixer gate_output_3_428(.a(output_4_428), .b(output_4_13), .y(output_3_428));
wire output_5_428, output_5_13, output_4_428;
mixer gate_output_4_428(.a(output_5_428), .b(output_5_13), .y(output_4_428));
wire output_6_428, output_6_13, output_5_428;
mixer gate_output_5_428(.a(output_6_428), .b(output_6_13), .y(output_5_428));
wire output_7_428, output_7_13, output_6_428;
mixer gate_output_6_428(.a(output_7_428), .b(output_7_13), .y(output_6_428));
wire output_8_428, output_8_13, output_7_428;
mixer gate_output_7_428(.a(output_8_428), .b(output_8_13), .y(output_7_428));
wire output_9_428, output_9_13, output_8_428;
mixer gate_output_8_428(.a(output_9_428), .b(output_9_13), .y(output_8_428));
wire output_10_428, output_10_13, output_9_428;
mixer gate_output_9_428(.a(output_10_428), .b(output_10_13), .y(output_9_428));
wire output_11_428, output_11_13, output_10_428;
mixer gate_output_10_428(.a(output_11_428), .b(output_11_13), .y(output_10_428));
wire output_12_428, output_12_13, output_11_428;
mixer gate_output_11_428(.a(output_12_428), .b(output_12_13), .y(output_11_428));
wire output_13_428, output_13_13, output_12_428;
mixer gate_output_12_428(.a(output_13_428), .b(output_13_13), .y(output_12_428));
wire output_14_428, output_14_13, output_13_428;
mixer gate_output_13_428(.a(output_14_428), .b(output_14_13), .y(output_13_428));
wire output_15_428, output_15_13, output_14_428;
mixer gate_output_14_428(.a(output_15_428), .b(output_15_13), .y(output_14_428));
wire output_16_428, output_16_13, output_15_428;
mixer gate_output_15_428(.a(output_16_428), .b(output_16_13), .y(output_15_428));
wire output_1_429, output_1_14, output_0_429;
mixer gate_output_0_429(.a(output_1_429), .b(output_1_14), .y(output_0_429));
wire output_2_429, output_2_14, output_1_429;
mixer gate_output_1_429(.a(output_2_429), .b(output_2_14), .y(output_1_429));
wire output_3_429, output_3_14, output_2_429;
mixer gate_output_2_429(.a(output_3_429), .b(output_3_14), .y(output_2_429));
wire output_4_429, output_4_14, output_3_429;
mixer gate_output_3_429(.a(output_4_429), .b(output_4_14), .y(output_3_429));
wire output_5_429, output_5_14, output_4_429;
mixer gate_output_4_429(.a(output_5_429), .b(output_5_14), .y(output_4_429));
wire output_6_429, output_6_14, output_5_429;
mixer gate_output_5_429(.a(output_6_429), .b(output_6_14), .y(output_5_429));
wire output_7_429, output_7_14, output_6_429;
mixer gate_output_6_429(.a(output_7_429), .b(output_7_14), .y(output_6_429));
wire output_8_429, output_8_14, output_7_429;
mixer gate_output_7_429(.a(output_8_429), .b(output_8_14), .y(output_7_429));
wire output_9_429, output_9_14, output_8_429;
mixer gate_output_8_429(.a(output_9_429), .b(output_9_14), .y(output_8_429));
wire output_10_429, output_10_14, output_9_429;
mixer gate_output_9_429(.a(output_10_429), .b(output_10_14), .y(output_9_429));
wire output_11_429, output_11_14, output_10_429;
mixer gate_output_10_429(.a(output_11_429), .b(output_11_14), .y(output_10_429));
wire output_12_429, output_12_14, output_11_429;
mixer gate_output_11_429(.a(output_12_429), .b(output_12_14), .y(output_11_429));
wire output_13_429, output_13_14, output_12_429;
mixer gate_output_12_429(.a(output_13_429), .b(output_13_14), .y(output_12_429));
wire output_14_429, output_14_14, output_13_429;
mixer gate_output_13_429(.a(output_14_429), .b(output_14_14), .y(output_13_429));
wire output_15_429, output_15_14, output_14_429;
mixer gate_output_14_429(.a(output_15_429), .b(output_15_14), .y(output_14_429));
wire output_16_429, output_16_14, output_15_429;
mixer gate_output_15_429(.a(output_16_429), .b(output_16_14), .y(output_15_429));
wire output_1_430, output_1_15, output_0_430;
mixer gate_output_0_430(.a(output_1_430), .b(output_1_15), .y(output_0_430));
wire output_2_430, output_2_15, output_1_430;
mixer gate_output_1_430(.a(output_2_430), .b(output_2_15), .y(output_1_430));
wire output_3_430, output_3_15, output_2_430;
mixer gate_output_2_430(.a(output_3_430), .b(output_3_15), .y(output_2_430));
wire output_4_430, output_4_15, output_3_430;
mixer gate_output_3_430(.a(output_4_430), .b(output_4_15), .y(output_3_430));
wire output_5_430, output_5_15, output_4_430;
mixer gate_output_4_430(.a(output_5_430), .b(output_5_15), .y(output_4_430));
wire output_6_430, output_6_15, output_5_430;
mixer gate_output_5_430(.a(output_6_430), .b(output_6_15), .y(output_5_430));
wire output_7_430, output_7_15, output_6_430;
mixer gate_output_6_430(.a(output_7_430), .b(output_7_15), .y(output_6_430));
wire output_8_430, output_8_15, output_7_430;
mixer gate_output_7_430(.a(output_8_430), .b(output_8_15), .y(output_7_430));
wire output_9_430, output_9_15, output_8_430;
mixer gate_output_8_430(.a(output_9_430), .b(output_9_15), .y(output_8_430));
wire output_10_430, output_10_15, output_9_430;
mixer gate_output_9_430(.a(output_10_430), .b(output_10_15), .y(output_9_430));
wire output_11_430, output_11_15, output_10_430;
mixer gate_output_10_430(.a(output_11_430), .b(output_11_15), .y(output_10_430));
wire output_12_430, output_12_15, output_11_430;
mixer gate_output_11_430(.a(output_12_430), .b(output_12_15), .y(output_11_430));
wire output_13_430, output_13_15, output_12_430;
mixer gate_output_12_430(.a(output_13_430), .b(output_13_15), .y(output_12_430));
wire output_14_430, output_14_15, output_13_430;
mixer gate_output_13_430(.a(output_14_430), .b(output_14_15), .y(output_13_430));
wire output_15_430, output_15_15, output_14_430;
mixer gate_output_14_430(.a(output_15_430), .b(output_15_15), .y(output_14_430));
wire output_16_430, output_16_15, output_15_430;
mixer gate_output_15_430(.a(output_16_430), .b(output_16_15), .y(output_15_430));
wire output_1_431, output_1_0, output_0_431;
mixer gate_output_0_431(.a(output_1_431), .b(output_1_0), .y(output_0_431));
wire output_2_431, output_2_0, output_1_431;
mixer gate_output_1_431(.a(output_2_431), .b(output_2_0), .y(output_1_431));
wire output_3_431, output_3_0, output_2_431;
mixer gate_output_2_431(.a(output_3_431), .b(output_3_0), .y(output_2_431));
wire output_4_431, output_4_0, output_3_431;
mixer gate_output_3_431(.a(output_4_431), .b(output_4_0), .y(output_3_431));
wire output_5_431, output_5_0, output_4_431;
mixer gate_output_4_431(.a(output_5_431), .b(output_5_0), .y(output_4_431));
wire output_6_431, output_6_0, output_5_431;
mixer gate_output_5_431(.a(output_6_431), .b(output_6_0), .y(output_5_431));
wire output_7_431, output_7_0, output_6_431;
mixer gate_output_6_431(.a(output_7_431), .b(output_7_0), .y(output_6_431));
wire output_8_431, output_8_0, output_7_431;
mixer gate_output_7_431(.a(output_8_431), .b(output_8_0), .y(output_7_431));
wire output_9_431, output_9_0, output_8_431;
mixer gate_output_8_431(.a(output_9_431), .b(output_9_0), .y(output_8_431));
wire output_10_431, output_10_0, output_9_431;
mixer gate_output_9_431(.a(output_10_431), .b(output_10_0), .y(output_9_431));
wire output_11_431, output_11_0, output_10_431;
mixer gate_output_10_431(.a(output_11_431), .b(output_11_0), .y(output_10_431));
wire output_12_431, output_12_0, output_11_431;
mixer gate_output_11_431(.a(output_12_431), .b(output_12_0), .y(output_11_431));
wire output_13_431, output_13_0, output_12_431;
mixer gate_output_12_431(.a(output_13_431), .b(output_13_0), .y(output_12_431));
wire output_14_431, output_14_0, output_13_431;
mixer gate_output_13_431(.a(output_14_431), .b(output_14_0), .y(output_13_431));
wire output_15_431, output_15_0, output_14_431;
mixer gate_output_14_431(.a(output_15_431), .b(output_15_0), .y(output_14_431));
wire output_16_431, output_16_0, output_15_431;
mixer gate_output_15_431(.a(output_16_431), .b(output_16_0), .y(output_15_431));
wire output_1_432, output_1_1, output_0_432;
mixer gate_output_0_432(.a(output_1_432), .b(output_1_1), .y(output_0_432));
wire output_2_432, output_2_1, output_1_432;
mixer gate_output_1_432(.a(output_2_432), .b(output_2_1), .y(output_1_432));
wire output_3_432, output_3_1, output_2_432;
mixer gate_output_2_432(.a(output_3_432), .b(output_3_1), .y(output_2_432));
wire output_4_432, output_4_1, output_3_432;
mixer gate_output_3_432(.a(output_4_432), .b(output_4_1), .y(output_3_432));
wire output_5_432, output_5_1, output_4_432;
mixer gate_output_4_432(.a(output_5_432), .b(output_5_1), .y(output_4_432));
wire output_6_432, output_6_1, output_5_432;
mixer gate_output_5_432(.a(output_6_432), .b(output_6_1), .y(output_5_432));
wire output_7_432, output_7_1, output_6_432;
mixer gate_output_6_432(.a(output_7_432), .b(output_7_1), .y(output_6_432));
wire output_8_432, output_8_1, output_7_432;
mixer gate_output_7_432(.a(output_8_432), .b(output_8_1), .y(output_7_432));
wire output_9_432, output_9_1, output_8_432;
mixer gate_output_8_432(.a(output_9_432), .b(output_9_1), .y(output_8_432));
wire output_10_432, output_10_1, output_9_432;
mixer gate_output_9_432(.a(output_10_432), .b(output_10_1), .y(output_9_432));
wire output_11_432, output_11_1, output_10_432;
mixer gate_output_10_432(.a(output_11_432), .b(output_11_1), .y(output_10_432));
wire output_12_432, output_12_1, output_11_432;
mixer gate_output_11_432(.a(output_12_432), .b(output_12_1), .y(output_11_432));
wire output_13_432, output_13_1, output_12_432;
mixer gate_output_12_432(.a(output_13_432), .b(output_13_1), .y(output_12_432));
wire output_14_432, output_14_1, output_13_432;
mixer gate_output_13_432(.a(output_14_432), .b(output_14_1), .y(output_13_432));
wire output_15_432, output_15_1, output_14_432;
mixer gate_output_14_432(.a(output_15_432), .b(output_15_1), .y(output_14_432));
wire output_16_432, output_16_1, output_15_432;
mixer gate_output_15_432(.a(output_16_432), .b(output_16_1), .y(output_15_432));
wire output_1_433, output_1_2, output_0_433;
mixer gate_output_0_433(.a(output_1_433), .b(output_1_2), .y(output_0_433));
wire output_2_433, output_2_2, output_1_433;
mixer gate_output_1_433(.a(output_2_433), .b(output_2_2), .y(output_1_433));
wire output_3_433, output_3_2, output_2_433;
mixer gate_output_2_433(.a(output_3_433), .b(output_3_2), .y(output_2_433));
wire output_4_433, output_4_2, output_3_433;
mixer gate_output_3_433(.a(output_4_433), .b(output_4_2), .y(output_3_433));
wire output_5_433, output_5_2, output_4_433;
mixer gate_output_4_433(.a(output_5_433), .b(output_5_2), .y(output_4_433));
wire output_6_433, output_6_2, output_5_433;
mixer gate_output_5_433(.a(output_6_433), .b(output_6_2), .y(output_5_433));
wire output_7_433, output_7_2, output_6_433;
mixer gate_output_6_433(.a(output_7_433), .b(output_7_2), .y(output_6_433));
wire output_8_433, output_8_2, output_7_433;
mixer gate_output_7_433(.a(output_8_433), .b(output_8_2), .y(output_7_433));
wire output_9_433, output_9_2, output_8_433;
mixer gate_output_8_433(.a(output_9_433), .b(output_9_2), .y(output_8_433));
wire output_10_433, output_10_2, output_9_433;
mixer gate_output_9_433(.a(output_10_433), .b(output_10_2), .y(output_9_433));
wire output_11_433, output_11_2, output_10_433;
mixer gate_output_10_433(.a(output_11_433), .b(output_11_2), .y(output_10_433));
wire output_12_433, output_12_2, output_11_433;
mixer gate_output_11_433(.a(output_12_433), .b(output_12_2), .y(output_11_433));
wire output_13_433, output_13_2, output_12_433;
mixer gate_output_12_433(.a(output_13_433), .b(output_13_2), .y(output_12_433));
wire output_14_433, output_14_2, output_13_433;
mixer gate_output_13_433(.a(output_14_433), .b(output_14_2), .y(output_13_433));
wire output_15_433, output_15_2, output_14_433;
mixer gate_output_14_433(.a(output_15_433), .b(output_15_2), .y(output_14_433));
wire output_16_433, output_16_2, output_15_433;
mixer gate_output_15_433(.a(output_16_433), .b(output_16_2), .y(output_15_433));
wire output_1_434, output_1_3, output_0_434;
mixer gate_output_0_434(.a(output_1_434), .b(output_1_3), .y(output_0_434));
wire output_2_434, output_2_3, output_1_434;
mixer gate_output_1_434(.a(output_2_434), .b(output_2_3), .y(output_1_434));
wire output_3_434, output_3_3, output_2_434;
mixer gate_output_2_434(.a(output_3_434), .b(output_3_3), .y(output_2_434));
wire output_4_434, output_4_3, output_3_434;
mixer gate_output_3_434(.a(output_4_434), .b(output_4_3), .y(output_3_434));
wire output_5_434, output_5_3, output_4_434;
mixer gate_output_4_434(.a(output_5_434), .b(output_5_3), .y(output_4_434));
wire output_6_434, output_6_3, output_5_434;
mixer gate_output_5_434(.a(output_6_434), .b(output_6_3), .y(output_5_434));
wire output_7_434, output_7_3, output_6_434;
mixer gate_output_6_434(.a(output_7_434), .b(output_7_3), .y(output_6_434));
wire output_8_434, output_8_3, output_7_434;
mixer gate_output_7_434(.a(output_8_434), .b(output_8_3), .y(output_7_434));
wire output_9_434, output_9_3, output_8_434;
mixer gate_output_8_434(.a(output_9_434), .b(output_9_3), .y(output_8_434));
wire output_10_434, output_10_3, output_9_434;
mixer gate_output_9_434(.a(output_10_434), .b(output_10_3), .y(output_9_434));
wire output_11_434, output_11_3, output_10_434;
mixer gate_output_10_434(.a(output_11_434), .b(output_11_3), .y(output_10_434));
wire output_12_434, output_12_3, output_11_434;
mixer gate_output_11_434(.a(output_12_434), .b(output_12_3), .y(output_11_434));
wire output_13_434, output_13_3, output_12_434;
mixer gate_output_12_434(.a(output_13_434), .b(output_13_3), .y(output_12_434));
wire output_14_434, output_14_3, output_13_434;
mixer gate_output_13_434(.a(output_14_434), .b(output_14_3), .y(output_13_434));
wire output_15_434, output_15_3, output_14_434;
mixer gate_output_14_434(.a(output_15_434), .b(output_15_3), .y(output_14_434));
wire output_16_434, output_16_3, output_15_434;
mixer gate_output_15_434(.a(output_16_434), .b(output_16_3), .y(output_15_434));
wire output_1_435, output_1_4, output_0_435;
mixer gate_output_0_435(.a(output_1_435), .b(output_1_4), .y(output_0_435));
wire output_2_435, output_2_4, output_1_435;
mixer gate_output_1_435(.a(output_2_435), .b(output_2_4), .y(output_1_435));
wire output_3_435, output_3_4, output_2_435;
mixer gate_output_2_435(.a(output_3_435), .b(output_3_4), .y(output_2_435));
wire output_4_435, output_4_4, output_3_435;
mixer gate_output_3_435(.a(output_4_435), .b(output_4_4), .y(output_3_435));
wire output_5_435, output_5_4, output_4_435;
mixer gate_output_4_435(.a(output_5_435), .b(output_5_4), .y(output_4_435));
wire output_6_435, output_6_4, output_5_435;
mixer gate_output_5_435(.a(output_6_435), .b(output_6_4), .y(output_5_435));
wire output_7_435, output_7_4, output_6_435;
mixer gate_output_6_435(.a(output_7_435), .b(output_7_4), .y(output_6_435));
wire output_8_435, output_8_4, output_7_435;
mixer gate_output_7_435(.a(output_8_435), .b(output_8_4), .y(output_7_435));
wire output_9_435, output_9_4, output_8_435;
mixer gate_output_8_435(.a(output_9_435), .b(output_9_4), .y(output_8_435));
wire output_10_435, output_10_4, output_9_435;
mixer gate_output_9_435(.a(output_10_435), .b(output_10_4), .y(output_9_435));
wire output_11_435, output_11_4, output_10_435;
mixer gate_output_10_435(.a(output_11_435), .b(output_11_4), .y(output_10_435));
wire output_12_435, output_12_4, output_11_435;
mixer gate_output_11_435(.a(output_12_435), .b(output_12_4), .y(output_11_435));
wire output_13_435, output_13_4, output_12_435;
mixer gate_output_12_435(.a(output_13_435), .b(output_13_4), .y(output_12_435));
wire output_14_435, output_14_4, output_13_435;
mixer gate_output_13_435(.a(output_14_435), .b(output_14_4), .y(output_13_435));
wire output_15_435, output_15_4, output_14_435;
mixer gate_output_14_435(.a(output_15_435), .b(output_15_4), .y(output_14_435));
wire output_16_435, output_16_4, output_15_435;
mixer gate_output_15_435(.a(output_16_435), .b(output_16_4), .y(output_15_435));
wire output_1_436, output_1_5, output_0_436;
mixer gate_output_0_436(.a(output_1_436), .b(output_1_5), .y(output_0_436));
wire output_2_436, output_2_5, output_1_436;
mixer gate_output_1_436(.a(output_2_436), .b(output_2_5), .y(output_1_436));
wire output_3_436, output_3_5, output_2_436;
mixer gate_output_2_436(.a(output_3_436), .b(output_3_5), .y(output_2_436));
wire output_4_436, output_4_5, output_3_436;
mixer gate_output_3_436(.a(output_4_436), .b(output_4_5), .y(output_3_436));
wire output_5_436, output_5_5, output_4_436;
mixer gate_output_4_436(.a(output_5_436), .b(output_5_5), .y(output_4_436));
wire output_6_436, output_6_5, output_5_436;
mixer gate_output_5_436(.a(output_6_436), .b(output_6_5), .y(output_5_436));
wire output_7_436, output_7_5, output_6_436;
mixer gate_output_6_436(.a(output_7_436), .b(output_7_5), .y(output_6_436));
wire output_8_436, output_8_5, output_7_436;
mixer gate_output_7_436(.a(output_8_436), .b(output_8_5), .y(output_7_436));
wire output_9_436, output_9_5, output_8_436;
mixer gate_output_8_436(.a(output_9_436), .b(output_9_5), .y(output_8_436));
wire output_10_436, output_10_5, output_9_436;
mixer gate_output_9_436(.a(output_10_436), .b(output_10_5), .y(output_9_436));
wire output_11_436, output_11_5, output_10_436;
mixer gate_output_10_436(.a(output_11_436), .b(output_11_5), .y(output_10_436));
wire output_12_436, output_12_5, output_11_436;
mixer gate_output_11_436(.a(output_12_436), .b(output_12_5), .y(output_11_436));
wire output_13_436, output_13_5, output_12_436;
mixer gate_output_12_436(.a(output_13_436), .b(output_13_5), .y(output_12_436));
wire output_14_436, output_14_5, output_13_436;
mixer gate_output_13_436(.a(output_14_436), .b(output_14_5), .y(output_13_436));
wire output_15_436, output_15_5, output_14_436;
mixer gate_output_14_436(.a(output_15_436), .b(output_15_5), .y(output_14_436));
wire output_16_436, output_16_5, output_15_436;
mixer gate_output_15_436(.a(output_16_436), .b(output_16_5), .y(output_15_436));
wire output_1_437, output_1_6, output_0_437;
mixer gate_output_0_437(.a(output_1_437), .b(output_1_6), .y(output_0_437));
wire output_2_437, output_2_6, output_1_437;
mixer gate_output_1_437(.a(output_2_437), .b(output_2_6), .y(output_1_437));
wire output_3_437, output_3_6, output_2_437;
mixer gate_output_2_437(.a(output_3_437), .b(output_3_6), .y(output_2_437));
wire output_4_437, output_4_6, output_3_437;
mixer gate_output_3_437(.a(output_4_437), .b(output_4_6), .y(output_3_437));
wire output_5_437, output_5_6, output_4_437;
mixer gate_output_4_437(.a(output_5_437), .b(output_5_6), .y(output_4_437));
wire output_6_437, output_6_6, output_5_437;
mixer gate_output_5_437(.a(output_6_437), .b(output_6_6), .y(output_5_437));
wire output_7_437, output_7_6, output_6_437;
mixer gate_output_6_437(.a(output_7_437), .b(output_7_6), .y(output_6_437));
wire output_8_437, output_8_6, output_7_437;
mixer gate_output_7_437(.a(output_8_437), .b(output_8_6), .y(output_7_437));
wire output_9_437, output_9_6, output_8_437;
mixer gate_output_8_437(.a(output_9_437), .b(output_9_6), .y(output_8_437));
wire output_10_437, output_10_6, output_9_437;
mixer gate_output_9_437(.a(output_10_437), .b(output_10_6), .y(output_9_437));
wire output_11_437, output_11_6, output_10_437;
mixer gate_output_10_437(.a(output_11_437), .b(output_11_6), .y(output_10_437));
wire output_12_437, output_12_6, output_11_437;
mixer gate_output_11_437(.a(output_12_437), .b(output_12_6), .y(output_11_437));
wire output_13_437, output_13_6, output_12_437;
mixer gate_output_12_437(.a(output_13_437), .b(output_13_6), .y(output_12_437));
wire output_14_437, output_14_6, output_13_437;
mixer gate_output_13_437(.a(output_14_437), .b(output_14_6), .y(output_13_437));
wire output_15_437, output_15_6, output_14_437;
mixer gate_output_14_437(.a(output_15_437), .b(output_15_6), .y(output_14_437));
wire output_16_437, output_16_6, output_15_437;
mixer gate_output_15_437(.a(output_16_437), .b(output_16_6), .y(output_15_437));
wire output_1_438, output_1_7, output_0_438;
mixer gate_output_0_438(.a(output_1_438), .b(output_1_7), .y(output_0_438));
wire output_2_438, output_2_7, output_1_438;
mixer gate_output_1_438(.a(output_2_438), .b(output_2_7), .y(output_1_438));
wire output_3_438, output_3_7, output_2_438;
mixer gate_output_2_438(.a(output_3_438), .b(output_3_7), .y(output_2_438));
wire output_4_438, output_4_7, output_3_438;
mixer gate_output_3_438(.a(output_4_438), .b(output_4_7), .y(output_3_438));
wire output_5_438, output_5_7, output_4_438;
mixer gate_output_4_438(.a(output_5_438), .b(output_5_7), .y(output_4_438));
wire output_6_438, output_6_7, output_5_438;
mixer gate_output_5_438(.a(output_6_438), .b(output_6_7), .y(output_5_438));
wire output_7_438, output_7_7, output_6_438;
mixer gate_output_6_438(.a(output_7_438), .b(output_7_7), .y(output_6_438));
wire output_8_438, output_8_7, output_7_438;
mixer gate_output_7_438(.a(output_8_438), .b(output_8_7), .y(output_7_438));
wire output_9_438, output_9_7, output_8_438;
mixer gate_output_8_438(.a(output_9_438), .b(output_9_7), .y(output_8_438));
wire output_10_438, output_10_7, output_9_438;
mixer gate_output_9_438(.a(output_10_438), .b(output_10_7), .y(output_9_438));
wire output_11_438, output_11_7, output_10_438;
mixer gate_output_10_438(.a(output_11_438), .b(output_11_7), .y(output_10_438));
wire output_12_438, output_12_7, output_11_438;
mixer gate_output_11_438(.a(output_12_438), .b(output_12_7), .y(output_11_438));
wire output_13_438, output_13_7, output_12_438;
mixer gate_output_12_438(.a(output_13_438), .b(output_13_7), .y(output_12_438));
wire output_14_438, output_14_7, output_13_438;
mixer gate_output_13_438(.a(output_14_438), .b(output_14_7), .y(output_13_438));
wire output_15_438, output_15_7, output_14_438;
mixer gate_output_14_438(.a(output_15_438), .b(output_15_7), .y(output_14_438));
wire output_16_438, output_16_7, output_15_438;
mixer gate_output_15_438(.a(output_16_438), .b(output_16_7), .y(output_15_438));
wire output_1_439, output_1_8, output_0_439;
mixer gate_output_0_439(.a(output_1_439), .b(output_1_8), .y(output_0_439));
wire output_2_439, output_2_8, output_1_439;
mixer gate_output_1_439(.a(output_2_439), .b(output_2_8), .y(output_1_439));
wire output_3_439, output_3_8, output_2_439;
mixer gate_output_2_439(.a(output_3_439), .b(output_3_8), .y(output_2_439));
wire output_4_439, output_4_8, output_3_439;
mixer gate_output_3_439(.a(output_4_439), .b(output_4_8), .y(output_3_439));
wire output_5_439, output_5_8, output_4_439;
mixer gate_output_4_439(.a(output_5_439), .b(output_5_8), .y(output_4_439));
wire output_6_439, output_6_8, output_5_439;
mixer gate_output_5_439(.a(output_6_439), .b(output_6_8), .y(output_5_439));
wire output_7_439, output_7_8, output_6_439;
mixer gate_output_6_439(.a(output_7_439), .b(output_7_8), .y(output_6_439));
wire output_8_439, output_8_8, output_7_439;
mixer gate_output_7_439(.a(output_8_439), .b(output_8_8), .y(output_7_439));
wire output_9_439, output_9_8, output_8_439;
mixer gate_output_8_439(.a(output_9_439), .b(output_9_8), .y(output_8_439));
wire output_10_439, output_10_8, output_9_439;
mixer gate_output_9_439(.a(output_10_439), .b(output_10_8), .y(output_9_439));
wire output_11_439, output_11_8, output_10_439;
mixer gate_output_10_439(.a(output_11_439), .b(output_11_8), .y(output_10_439));
wire output_12_439, output_12_8, output_11_439;
mixer gate_output_11_439(.a(output_12_439), .b(output_12_8), .y(output_11_439));
wire output_13_439, output_13_8, output_12_439;
mixer gate_output_12_439(.a(output_13_439), .b(output_13_8), .y(output_12_439));
wire output_14_439, output_14_8, output_13_439;
mixer gate_output_13_439(.a(output_14_439), .b(output_14_8), .y(output_13_439));
wire output_15_439, output_15_8, output_14_439;
mixer gate_output_14_439(.a(output_15_439), .b(output_15_8), .y(output_14_439));
wire output_16_439, output_16_8, output_15_439;
mixer gate_output_15_439(.a(output_16_439), .b(output_16_8), .y(output_15_439));
wire output_1_440, output_1_9, output_0_440;
mixer gate_output_0_440(.a(output_1_440), .b(output_1_9), .y(output_0_440));
wire output_2_440, output_2_9, output_1_440;
mixer gate_output_1_440(.a(output_2_440), .b(output_2_9), .y(output_1_440));
wire output_3_440, output_3_9, output_2_440;
mixer gate_output_2_440(.a(output_3_440), .b(output_3_9), .y(output_2_440));
wire output_4_440, output_4_9, output_3_440;
mixer gate_output_3_440(.a(output_4_440), .b(output_4_9), .y(output_3_440));
wire output_5_440, output_5_9, output_4_440;
mixer gate_output_4_440(.a(output_5_440), .b(output_5_9), .y(output_4_440));
wire output_6_440, output_6_9, output_5_440;
mixer gate_output_5_440(.a(output_6_440), .b(output_6_9), .y(output_5_440));
wire output_7_440, output_7_9, output_6_440;
mixer gate_output_6_440(.a(output_7_440), .b(output_7_9), .y(output_6_440));
wire output_8_440, output_8_9, output_7_440;
mixer gate_output_7_440(.a(output_8_440), .b(output_8_9), .y(output_7_440));
wire output_9_440, output_9_9, output_8_440;
mixer gate_output_8_440(.a(output_9_440), .b(output_9_9), .y(output_8_440));
wire output_10_440, output_10_9, output_9_440;
mixer gate_output_9_440(.a(output_10_440), .b(output_10_9), .y(output_9_440));
wire output_11_440, output_11_9, output_10_440;
mixer gate_output_10_440(.a(output_11_440), .b(output_11_9), .y(output_10_440));
wire output_12_440, output_12_9, output_11_440;
mixer gate_output_11_440(.a(output_12_440), .b(output_12_9), .y(output_11_440));
wire output_13_440, output_13_9, output_12_440;
mixer gate_output_12_440(.a(output_13_440), .b(output_13_9), .y(output_12_440));
wire output_14_440, output_14_9, output_13_440;
mixer gate_output_13_440(.a(output_14_440), .b(output_14_9), .y(output_13_440));
wire output_15_440, output_15_9, output_14_440;
mixer gate_output_14_440(.a(output_15_440), .b(output_15_9), .y(output_14_440));
wire output_16_440, output_16_9, output_15_440;
mixer gate_output_15_440(.a(output_16_440), .b(output_16_9), .y(output_15_440));
wire output_1_441, output_1_10, output_0_441;
mixer gate_output_0_441(.a(output_1_441), .b(output_1_10), .y(output_0_441));
wire output_2_441, output_2_10, output_1_441;
mixer gate_output_1_441(.a(output_2_441), .b(output_2_10), .y(output_1_441));
wire output_3_441, output_3_10, output_2_441;
mixer gate_output_2_441(.a(output_3_441), .b(output_3_10), .y(output_2_441));
wire output_4_441, output_4_10, output_3_441;
mixer gate_output_3_441(.a(output_4_441), .b(output_4_10), .y(output_3_441));
wire output_5_441, output_5_10, output_4_441;
mixer gate_output_4_441(.a(output_5_441), .b(output_5_10), .y(output_4_441));
wire output_6_441, output_6_10, output_5_441;
mixer gate_output_5_441(.a(output_6_441), .b(output_6_10), .y(output_5_441));
wire output_7_441, output_7_10, output_6_441;
mixer gate_output_6_441(.a(output_7_441), .b(output_7_10), .y(output_6_441));
wire output_8_441, output_8_10, output_7_441;
mixer gate_output_7_441(.a(output_8_441), .b(output_8_10), .y(output_7_441));
wire output_9_441, output_9_10, output_8_441;
mixer gate_output_8_441(.a(output_9_441), .b(output_9_10), .y(output_8_441));
wire output_10_441, output_10_10, output_9_441;
mixer gate_output_9_441(.a(output_10_441), .b(output_10_10), .y(output_9_441));
wire output_11_441, output_11_10, output_10_441;
mixer gate_output_10_441(.a(output_11_441), .b(output_11_10), .y(output_10_441));
wire output_12_441, output_12_10, output_11_441;
mixer gate_output_11_441(.a(output_12_441), .b(output_12_10), .y(output_11_441));
wire output_13_441, output_13_10, output_12_441;
mixer gate_output_12_441(.a(output_13_441), .b(output_13_10), .y(output_12_441));
wire output_14_441, output_14_10, output_13_441;
mixer gate_output_13_441(.a(output_14_441), .b(output_14_10), .y(output_13_441));
wire output_15_441, output_15_10, output_14_441;
mixer gate_output_14_441(.a(output_15_441), .b(output_15_10), .y(output_14_441));
wire output_16_441, output_16_10, output_15_441;
mixer gate_output_15_441(.a(output_16_441), .b(output_16_10), .y(output_15_441));
wire output_1_442, output_1_11, output_0_442;
mixer gate_output_0_442(.a(output_1_442), .b(output_1_11), .y(output_0_442));
wire output_2_442, output_2_11, output_1_442;
mixer gate_output_1_442(.a(output_2_442), .b(output_2_11), .y(output_1_442));
wire output_3_442, output_3_11, output_2_442;
mixer gate_output_2_442(.a(output_3_442), .b(output_3_11), .y(output_2_442));
wire output_4_442, output_4_11, output_3_442;
mixer gate_output_3_442(.a(output_4_442), .b(output_4_11), .y(output_3_442));
wire output_5_442, output_5_11, output_4_442;
mixer gate_output_4_442(.a(output_5_442), .b(output_5_11), .y(output_4_442));
wire output_6_442, output_6_11, output_5_442;
mixer gate_output_5_442(.a(output_6_442), .b(output_6_11), .y(output_5_442));
wire output_7_442, output_7_11, output_6_442;
mixer gate_output_6_442(.a(output_7_442), .b(output_7_11), .y(output_6_442));
wire output_8_442, output_8_11, output_7_442;
mixer gate_output_7_442(.a(output_8_442), .b(output_8_11), .y(output_7_442));
wire output_9_442, output_9_11, output_8_442;
mixer gate_output_8_442(.a(output_9_442), .b(output_9_11), .y(output_8_442));
wire output_10_442, output_10_11, output_9_442;
mixer gate_output_9_442(.a(output_10_442), .b(output_10_11), .y(output_9_442));
wire output_11_442, output_11_11, output_10_442;
mixer gate_output_10_442(.a(output_11_442), .b(output_11_11), .y(output_10_442));
wire output_12_442, output_12_11, output_11_442;
mixer gate_output_11_442(.a(output_12_442), .b(output_12_11), .y(output_11_442));
wire output_13_442, output_13_11, output_12_442;
mixer gate_output_12_442(.a(output_13_442), .b(output_13_11), .y(output_12_442));
wire output_14_442, output_14_11, output_13_442;
mixer gate_output_13_442(.a(output_14_442), .b(output_14_11), .y(output_13_442));
wire output_15_442, output_15_11, output_14_442;
mixer gate_output_14_442(.a(output_15_442), .b(output_15_11), .y(output_14_442));
wire output_16_442, output_16_11, output_15_442;
mixer gate_output_15_442(.a(output_16_442), .b(output_16_11), .y(output_15_442));
wire output_1_443, output_1_12, output_0_443;
mixer gate_output_0_443(.a(output_1_443), .b(output_1_12), .y(output_0_443));
wire output_2_443, output_2_12, output_1_443;
mixer gate_output_1_443(.a(output_2_443), .b(output_2_12), .y(output_1_443));
wire output_3_443, output_3_12, output_2_443;
mixer gate_output_2_443(.a(output_3_443), .b(output_3_12), .y(output_2_443));
wire output_4_443, output_4_12, output_3_443;
mixer gate_output_3_443(.a(output_4_443), .b(output_4_12), .y(output_3_443));
wire output_5_443, output_5_12, output_4_443;
mixer gate_output_4_443(.a(output_5_443), .b(output_5_12), .y(output_4_443));
wire output_6_443, output_6_12, output_5_443;
mixer gate_output_5_443(.a(output_6_443), .b(output_6_12), .y(output_5_443));
wire output_7_443, output_7_12, output_6_443;
mixer gate_output_6_443(.a(output_7_443), .b(output_7_12), .y(output_6_443));
wire output_8_443, output_8_12, output_7_443;
mixer gate_output_7_443(.a(output_8_443), .b(output_8_12), .y(output_7_443));
wire output_9_443, output_9_12, output_8_443;
mixer gate_output_8_443(.a(output_9_443), .b(output_9_12), .y(output_8_443));
wire output_10_443, output_10_12, output_9_443;
mixer gate_output_9_443(.a(output_10_443), .b(output_10_12), .y(output_9_443));
wire output_11_443, output_11_12, output_10_443;
mixer gate_output_10_443(.a(output_11_443), .b(output_11_12), .y(output_10_443));
wire output_12_443, output_12_12, output_11_443;
mixer gate_output_11_443(.a(output_12_443), .b(output_12_12), .y(output_11_443));
wire output_13_443, output_13_12, output_12_443;
mixer gate_output_12_443(.a(output_13_443), .b(output_13_12), .y(output_12_443));
wire output_14_443, output_14_12, output_13_443;
mixer gate_output_13_443(.a(output_14_443), .b(output_14_12), .y(output_13_443));
wire output_15_443, output_15_12, output_14_443;
mixer gate_output_14_443(.a(output_15_443), .b(output_15_12), .y(output_14_443));
wire output_16_443, output_16_12, output_15_443;
mixer gate_output_15_443(.a(output_16_443), .b(output_16_12), .y(output_15_443));
wire output_1_444, output_1_13, output_0_444;
mixer gate_output_0_444(.a(output_1_444), .b(output_1_13), .y(output_0_444));
wire output_2_444, output_2_13, output_1_444;
mixer gate_output_1_444(.a(output_2_444), .b(output_2_13), .y(output_1_444));
wire output_3_444, output_3_13, output_2_444;
mixer gate_output_2_444(.a(output_3_444), .b(output_3_13), .y(output_2_444));
wire output_4_444, output_4_13, output_3_444;
mixer gate_output_3_444(.a(output_4_444), .b(output_4_13), .y(output_3_444));
wire output_5_444, output_5_13, output_4_444;
mixer gate_output_4_444(.a(output_5_444), .b(output_5_13), .y(output_4_444));
wire output_6_444, output_6_13, output_5_444;
mixer gate_output_5_444(.a(output_6_444), .b(output_6_13), .y(output_5_444));
wire output_7_444, output_7_13, output_6_444;
mixer gate_output_6_444(.a(output_7_444), .b(output_7_13), .y(output_6_444));
wire output_8_444, output_8_13, output_7_444;
mixer gate_output_7_444(.a(output_8_444), .b(output_8_13), .y(output_7_444));
wire output_9_444, output_9_13, output_8_444;
mixer gate_output_8_444(.a(output_9_444), .b(output_9_13), .y(output_8_444));
wire output_10_444, output_10_13, output_9_444;
mixer gate_output_9_444(.a(output_10_444), .b(output_10_13), .y(output_9_444));
wire output_11_444, output_11_13, output_10_444;
mixer gate_output_10_444(.a(output_11_444), .b(output_11_13), .y(output_10_444));
wire output_12_444, output_12_13, output_11_444;
mixer gate_output_11_444(.a(output_12_444), .b(output_12_13), .y(output_11_444));
wire output_13_444, output_13_13, output_12_444;
mixer gate_output_12_444(.a(output_13_444), .b(output_13_13), .y(output_12_444));
wire output_14_444, output_14_13, output_13_444;
mixer gate_output_13_444(.a(output_14_444), .b(output_14_13), .y(output_13_444));
wire output_15_444, output_15_13, output_14_444;
mixer gate_output_14_444(.a(output_15_444), .b(output_15_13), .y(output_14_444));
wire output_16_444, output_16_13, output_15_444;
mixer gate_output_15_444(.a(output_16_444), .b(output_16_13), .y(output_15_444));
wire output_1_445, output_1_14, output_0_445;
mixer gate_output_0_445(.a(output_1_445), .b(output_1_14), .y(output_0_445));
wire output_2_445, output_2_14, output_1_445;
mixer gate_output_1_445(.a(output_2_445), .b(output_2_14), .y(output_1_445));
wire output_3_445, output_3_14, output_2_445;
mixer gate_output_2_445(.a(output_3_445), .b(output_3_14), .y(output_2_445));
wire output_4_445, output_4_14, output_3_445;
mixer gate_output_3_445(.a(output_4_445), .b(output_4_14), .y(output_3_445));
wire output_5_445, output_5_14, output_4_445;
mixer gate_output_4_445(.a(output_5_445), .b(output_5_14), .y(output_4_445));
wire output_6_445, output_6_14, output_5_445;
mixer gate_output_5_445(.a(output_6_445), .b(output_6_14), .y(output_5_445));
wire output_7_445, output_7_14, output_6_445;
mixer gate_output_6_445(.a(output_7_445), .b(output_7_14), .y(output_6_445));
wire output_8_445, output_8_14, output_7_445;
mixer gate_output_7_445(.a(output_8_445), .b(output_8_14), .y(output_7_445));
wire output_9_445, output_9_14, output_8_445;
mixer gate_output_8_445(.a(output_9_445), .b(output_9_14), .y(output_8_445));
wire output_10_445, output_10_14, output_9_445;
mixer gate_output_9_445(.a(output_10_445), .b(output_10_14), .y(output_9_445));
wire output_11_445, output_11_14, output_10_445;
mixer gate_output_10_445(.a(output_11_445), .b(output_11_14), .y(output_10_445));
wire output_12_445, output_12_14, output_11_445;
mixer gate_output_11_445(.a(output_12_445), .b(output_12_14), .y(output_11_445));
wire output_13_445, output_13_14, output_12_445;
mixer gate_output_12_445(.a(output_13_445), .b(output_13_14), .y(output_12_445));
wire output_14_445, output_14_14, output_13_445;
mixer gate_output_13_445(.a(output_14_445), .b(output_14_14), .y(output_13_445));
wire output_15_445, output_15_14, output_14_445;
mixer gate_output_14_445(.a(output_15_445), .b(output_15_14), .y(output_14_445));
wire output_16_445, output_16_14, output_15_445;
mixer gate_output_15_445(.a(output_16_445), .b(output_16_14), .y(output_15_445));
wire output_1_446, output_1_15, output_0_446;
mixer gate_output_0_446(.a(output_1_446), .b(output_1_15), .y(output_0_446));
wire output_2_446, output_2_15, output_1_446;
mixer gate_output_1_446(.a(output_2_446), .b(output_2_15), .y(output_1_446));
wire output_3_446, output_3_15, output_2_446;
mixer gate_output_2_446(.a(output_3_446), .b(output_3_15), .y(output_2_446));
wire output_4_446, output_4_15, output_3_446;
mixer gate_output_3_446(.a(output_4_446), .b(output_4_15), .y(output_3_446));
wire output_5_446, output_5_15, output_4_446;
mixer gate_output_4_446(.a(output_5_446), .b(output_5_15), .y(output_4_446));
wire output_6_446, output_6_15, output_5_446;
mixer gate_output_5_446(.a(output_6_446), .b(output_6_15), .y(output_5_446));
wire output_7_446, output_7_15, output_6_446;
mixer gate_output_6_446(.a(output_7_446), .b(output_7_15), .y(output_6_446));
wire output_8_446, output_8_15, output_7_446;
mixer gate_output_7_446(.a(output_8_446), .b(output_8_15), .y(output_7_446));
wire output_9_446, output_9_15, output_8_446;
mixer gate_output_8_446(.a(output_9_446), .b(output_9_15), .y(output_8_446));
wire output_10_446, output_10_15, output_9_446;
mixer gate_output_9_446(.a(output_10_446), .b(output_10_15), .y(output_9_446));
wire output_11_446, output_11_15, output_10_446;
mixer gate_output_10_446(.a(output_11_446), .b(output_11_15), .y(output_10_446));
wire output_12_446, output_12_15, output_11_446;
mixer gate_output_11_446(.a(output_12_446), .b(output_12_15), .y(output_11_446));
wire output_13_446, output_13_15, output_12_446;
mixer gate_output_12_446(.a(output_13_446), .b(output_13_15), .y(output_12_446));
wire output_14_446, output_14_15, output_13_446;
mixer gate_output_13_446(.a(output_14_446), .b(output_14_15), .y(output_13_446));
wire output_15_446, output_15_15, output_14_446;
mixer gate_output_14_446(.a(output_15_446), .b(output_15_15), .y(output_14_446));
wire output_16_446, output_16_15, output_15_446;
mixer gate_output_15_446(.a(output_16_446), .b(output_16_15), .y(output_15_446));
wire output_1_447, output_1_0, output_0_447;
mixer gate_output_0_447(.a(output_1_447), .b(output_1_0), .y(output_0_447));
wire output_2_447, output_2_0, output_1_447;
mixer gate_output_1_447(.a(output_2_447), .b(output_2_0), .y(output_1_447));
wire output_3_447, output_3_0, output_2_447;
mixer gate_output_2_447(.a(output_3_447), .b(output_3_0), .y(output_2_447));
wire output_4_447, output_4_0, output_3_447;
mixer gate_output_3_447(.a(output_4_447), .b(output_4_0), .y(output_3_447));
wire output_5_447, output_5_0, output_4_447;
mixer gate_output_4_447(.a(output_5_447), .b(output_5_0), .y(output_4_447));
wire output_6_447, output_6_0, output_5_447;
mixer gate_output_5_447(.a(output_6_447), .b(output_6_0), .y(output_5_447));
wire output_7_447, output_7_0, output_6_447;
mixer gate_output_6_447(.a(output_7_447), .b(output_7_0), .y(output_6_447));
wire output_8_447, output_8_0, output_7_447;
mixer gate_output_7_447(.a(output_8_447), .b(output_8_0), .y(output_7_447));
wire output_9_447, output_9_0, output_8_447;
mixer gate_output_8_447(.a(output_9_447), .b(output_9_0), .y(output_8_447));
wire output_10_447, output_10_0, output_9_447;
mixer gate_output_9_447(.a(output_10_447), .b(output_10_0), .y(output_9_447));
wire output_11_447, output_11_0, output_10_447;
mixer gate_output_10_447(.a(output_11_447), .b(output_11_0), .y(output_10_447));
wire output_12_447, output_12_0, output_11_447;
mixer gate_output_11_447(.a(output_12_447), .b(output_12_0), .y(output_11_447));
wire output_13_447, output_13_0, output_12_447;
mixer gate_output_12_447(.a(output_13_447), .b(output_13_0), .y(output_12_447));
wire output_14_447, output_14_0, output_13_447;
mixer gate_output_13_447(.a(output_14_447), .b(output_14_0), .y(output_13_447));
wire output_15_447, output_15_0, output_14_447;
mixer gate_output_14_447(.a(output_15_447), .b(output_15_0), .y(output_14_447));
wire output_16_447, output_16_0, output_15_447;
mixer gate_output_15_447(.a(output_16_447), .b(output_16_0), .y(output_15_447));
wire output_1_448, output_1_1, output_0_448;
mixer gate_output_0_448(.a(output_1_448), .b(output_1_1), .y(output_0_448));
wire output_2_448, output_2_1, output_1_448;
mixer gate_output_1_448(.a(output_2_448), .b(output_2_1), .y(output_1_448));
wire output_3_448, output_3_1, output_2_448;
mixer gate_output_2_448(.a(output_3_448), .b(output_3_1), .y(output_2_448));
wire output_4_448, output_4_1, output_3_448;
mixer gate_output_3_448(.a(output_4_448), .b(output_4_1), .y(output_3_448));
wire output_5_448, output_5_1, output_4_448;
mixer gate_output_4_448(.a(output_5_448), .b(output_5_1), .y(output_4_448));
wire output_6_448, output_6_1, output_5_448;
mixer gate_output_5_448(.a(output_6_448), .b(output_6_1), .y(output_5_448));
wire output_7_448, output_7_1, output_6_448;
mixer gate_output_6_448(.a(output_7_448), .b(output_7_1), .y(output_6_448));
wire output_8_448, output_8_1, output_7_448;
mixer gate_output_7_448(.a(output_8_448), .b(output_8_1), .y(output_7_448));
wire output_9_448, output_9_1, output_8_448;
mixer gate_output_8_448(.a(output_9_448), .b(output_9_1), .y(output_8_448));
wire output_10_448, output_10_1, output_9_448;
mixer gate_output_9_448(.a(output_10_448), .b(output_10_1), .y(output_9_448));
wire output_11_448, output_11_1, output_10_448;
mixer gate_output_10_448(.a(output_11_448), .b(output_11_1), .y(output_10_448));
wire output_12_448, output_12_1, output_11_448;
mixer gate_output_11_448(.a(output_12_448), .b(output_12_1), .y(output_11_448));
wire output_13_448, output_13_1, output_12_448;
mixer gate_output_12_448(.a(output_13_448), .b(output_13_1), .y(output_12_448));
wire output_14_448, output_14_1, output_13_448;
mixer gate_output_13_448(.a(output_14_448), .b(output_14_1), .y(output_13_448));
wire output_15_448, output_15_1, output_14_448;
mixer gate_output_14_448(.a(output_15_448), .b(output_15_1), .y(output_14_448));
wire output_16_448, output_16_1, output_15_448;
mixer gate_output_15_448(.a(output_16_448), .b(output_16_1), .y(output_15_448));
wire output_1_449, output_1_2, output_0_449;
mixer gate_output_0_449(.a(output_1_449), .b(output_1_2), .y(output_0_449));
wire output_2_449, output_2_2, output_1_449;
mixer gate_output_1_449(.a(output_2_449), .b(output_2_2), .y(output_1_449));
wire output_3_449, output_3_2, output_2_449;
mixer gate_output_2_449(.a(output_3_449), .b(output_3_2), .y(output_2_449));
wire output_4_449, output_4_2, output_3_449;
mixer gate_output_3_449(.a(output_4_449), .b(output_4_2), .y(output_3_449));
wire output_5_449, output_5_2, output_4_449;
mixer gate_output_4_449(.a(output_5_449), .b(output_5_2), .y(output_4_449));
wire output_6_449, output_6_2, output_5_449;
mixer gate_output_5_449(.a(output_6_449), .b(output_6_2), .y(output_5_449));
wire output_7_449, output_7_2, output_6_449;
mixer gate_output_6_449(.a(output_7_449), .b(output_7_2), .y(output_6_449));
wire output_8_449, output_8_2, output_7_449;
mixer gate_output_7_449(.a(output_8_449), .b(output_8_2), .y(output_7_449));
wire output_9_449, output_9_2, output_8_449;
mixer gate_output_8_449(.a(output_9_449), .b(output_9_2), .y(output_8_449));
wire output_10_449, output_10_2, output_9_449;
mixer gate_output_9_449(.a(output_10_449), .b(output_10_2), .y(output_9_449));
wire output_11_449, output_11_2, output_10_449;
mixer gate_output_10_449(.a(output_11_449), .b(output_11_2), .y(output_10_449));
wire output_12_449, output_12_2, output_11_449;
mixer gate_output_11_449(.a(output_12_449), .b(output_12_2), .y(output_11_449));
wire output_13_449, output_13_2, output_12_449;
mixer gate_output_12_449(.a(output_13_449), .b(output_13_2), .y(output_12_449));
wire output_14_449, output_14_2, output_13_449;
mixer gate_output_13_449(.a(output_14_449), .b(output_14_2), .y(output_13_449));
wire output_15_449, output_15_2, output_14_449;
mixer gate_output_14_449(.a(output_15_449), .b(output_15_2), .y(output_14_449));
wire output_16_449, output_16_2, output_15_449;
mixer gate_output_15_449(.a(output_16_449), .b(output_16_2), .y(output_15_449));
wire output_1_450, output_1_3, output_0_450;
mixer gate_output_0_450(.a(output_1_450), .b(output_1_3), .y(output_0_450));
wire output_2_450, output_2_3, output_1_450;
mixer gate_output_1_450(.a(output_2_450), .b(output_2_3), .y(output_1_450));
wire output_3_450, output_3_3, output_2_450;
mixer gate_output_2_450(.a(output_3_450), .b(output_3_3), .y(output_2_450));
wire output_4_450, output_4_3, output_3_450;
mixer gate_output_3_450(.a(output_4_450), .b(output_4_3), .y(output_3_450));
wire output_5_450, output_5_3, output_4_450;
mixer gate_output_4_450(.a(output_5_450), .b(output_5_3), .y(output_4_450));
wire output_6_450, output_6_3, output_5_450;
mixer gate_output_5_450(.a(output_6_450), .b(output_6_3), .y(output_5_450));
wire output_7_450, output_7_3, output_6_450;
mixer gate_output_6_450(.a(output_7_450), .b(output_7_3), .y(output_6_450));
wire output_8_450, output_8_3, output_7_450;
mixer gate_output_7_450(.a(output_8_450), .b(output_8_3), .y(output_7_450));
wire output_9_450, output_9_3, output_8_450;
mixer gate_output_8_450(.a(output_9_450), .b(output_9_3), .y(output_8_450));
wire output_10_450, output_10_3, output_9_450;
mixer gate_output_9_450(.a(output_10_450), .b(output_10_3), .y(output_9_450));
wire output_11_450, output_11_3, output_10_450;
mixer gate_output_10_450(.a(output_11_450), .b(output_11_3), .y(output_10_450));
wire output_12_450, output_12_3, output_11_450;
mixer gate_output_11_450(.a(output_12_450), .b(output_12_3), .y(output_11_450));
wire output_13_450, output_13_3, output_12_450;
mixer gate_output_12_450(.a(output_13_450), .b(output_13_3), .y(output_12_450));
wire output_14_450, output_14_3, output_13_450;
mixer gate_output_13_450(.a(output_14_450), .b(output_14_3), .y(output_13_450));
wire output_15_450, output_15_3, output_14_450;
mixer gate_output_14_450(.a(output_15_450), .b(output_15_3), .y(output_14_450));
wire output_16_450, output_16_3, output_15_450;
mixer gate_output_15_450(.a(output_16_450), .b(output_16_3), .y(output_15_450));
wire output_1_451, output_1_4, output_0_451;
mixer gate_output_0_451(.a(output_1_451), .b(output_1_4), .y(output_0_451));
wire output_2_451, output_2_4, output_1_451;
mixer gate_output_1_451(.a(output_2_451), .b(output_2_4), .y(output_1_451));
wire output_3_451, output_3_4, output_2_451;
mixer gate_output_2_451(.a(output_3_451), .b(output_3_4), .y(output_2_451));
wire output_4_451, output_4_4, output_3_451;
mixer gate_output_3_451(.a(output_4_451), .b(output_4_4), .y(output_3_451));
wire output_5_451, output_5_4, output_4_451;
mixer gate_output_4_451(.a(output_5_451), .b(output_5_4), .y(output_4_451));
wire output_6_451, output_6_4, output_5_451;
mixer gate_output_5_451(.a(output_6_451), .b(output_6_4), .y(output_5_451));
wire output_7_451, output_7_4, output_6_451;
mixer gate_output_6_451(.a(output_7_451), .b(output_7_4), .y(output_6_451));
wire output_8_451, output_8_4, output_7_451;
mixer gate_output_7_451(.a(output_8_451), .b(output_8_4), .y(output_7_451));
wire output_9_451, output_9_4, output_8_451;
mixer gate_output_8_451(.a(output_9_451), .b(output_9_4), .y(output_8_451));
wire output_10_451, output_10_4, output_9_451;
mixer gate_output_9_451(.a(output_10_451), .b(output_10_4), .y(output_9_451));
wire output_11_451, output_11_4, output_10_451;
mixer gate_output_10_451(.a(output_11_451), .b(output_11_4), .y(output_10_451));
wire output_12_451, output_12_4, output_11_451;
mixer gate_output_11_451(.a(output_12_451), .b(output_12_4), .y(output_11_451));
wire output_13_451, output_13_4, output_12_451;
mixer gate_output_12_451(.a(output_13_451), .b(output_13_4), .y(output_12_451));
wire output_14_451, output_14_4, output_13_451;
mixer gate_output_13_451(.a(output_14_451), .b(output_14_4), .y(output_13_451));
wire output_15_451, output_15_4, output_14_451;
mixer gate_output_14_451(.a(output_15_451), .b(output_15_4), .y(output_14_451));
wire output_16_451, output_16_4, output_15_451;
mixer gate_output_15_451(.a(output_16_451), .b(output_16_4), .y(output_15_451));
wire output_1_452, output_1_5, output_0_452;
mixer gate_output_0_452(.a(output_1_452), .b(output_1_5), .y(output_0_452));
wire output_2_452, output_2_5, output_1_452;
mixer gate_output_1_452(.a(output_2_452), .b(output_2_5), .y(output_1_452));
wire output_3_452, output_3_5, output_2_452;
mixer gate_output_2_452(.a(output_3_452), .b(output_3_5), .y(output_2_452));
wire output_4_452, output_4_5, output_3_452;
mixer gate_output_3_452(.a(output_4_452), .b(output_4_5), .y(output_3_452));
wire output_5_452, output_5_5, output_4_452;
mixer gate_output_4_452(.a(output_5_452), .b(output_5_5), .y(output_4_452));
wire output_6_452, output_6_5, output_5_452;
mixer gate_output_5_452(.a(output_6_452), .b(output_6_5), .y(output_5_452));
wire output_7_452, output_7_5, output_6_452;
mixer gate_output_6_452(.a(output_7_452), .b(output_7_5), .y(output_6_452));
wire output_8_452, output_8_5, output_7_452;
mixer gate_output_7_452(.a(output_8_452), .b(output_8_5), .y(output_7_452));
wire output_9_452, output_9_5, output_8_452;
mixer gate_output_8_452(.a(output_9_452), .b(output_9_5), .y(output_8_452));
wire output_10_452, output_10_5, output_9_452;
mixer gate_output_9_452(.a(output_10_452), .b(output_10_5), .y(output_9_452));
wire output_11_452, output_11_5, output_10_452;
mixer gate_output_10_452(.a(output_11_452), .b(output_11_5), .y(output_10_452));
wire output_12_452, output_12_5, output_11_452;
mixer gate_output_11_452(.a(output_12_452), .b(output_12_5), .y(output_11_452));
wire output_13_452, output_13_5, output_12_452;
mixer gate_output_12_452(.a(output_13_452), .b(output_13_5), .y(output_12_452));
wire output_14_452, output_14_5, output_13_452;
mixer gate_output_13_452(.a(output_14_452), .b(output_14_5), .y(output_13_452));
wire output_15_452, output_15_5, output_14_452;
mixer gate_output_14_452(.a(output_15_452), .b(output_15_5), .y(output_14_452));
wire output_16_452, output_16_5, output_15_452;
mixer gate_output_15_452(.a(output_16_452), .b(output_16_5), .y(output_15_452));
wire output_1_453, output_1_6, output_0_453;
mixer gate_output_0_453(.a(output_1_453), .b(output_1_6), .y(output_0_453));
wire output_2_453, output_2_6, output_1_453;
mixer gate_output_1_453(.a(output_2_453), .b(output_2_6), .y(output_1_453));
wire output_3_453, output_3_6, output_2_453;
mixer gate_output_2_453(.a(output_3_453), .b(output_3_6), .y(output_2_453));
wire output_4_453, output_4_6, output_3_453;
mixer gate_output_3_453(.a(output_4_453), .b(output_4_6), .y(output_3_453));
wire output_5_453, output_5_6, output_4_453;
mixer gate_output_4_453(.a(output_5_453), .b(output_5_6), .y(output_4_453));
wire output_6_453, output_6_6, output_5_453;
mixer gate_output_5_453(.a(output_6_453), .b(output_6_6), .y(output_5_453));
wire output_7_453, output_7_6, output_6_453;
mixer gate_output_6_453(.a(output_7_453), .b(output_7_6), .y(output_6_453));
wire output_8_453, output_8_6, output_7_453;
mixer gate_output_7_453(.a(output_8_453), .b(output_8_6), .y(output_7_453));
wire output_9_453, output_9_6, output_8_453;
mixer gate_output_8_453(.a(output_9_453), .b(output_9_6), .y(output_8_453));
wire output_10_453, output_10_6, output_9_453;
mixer gate_output_9_453(.a(output_10_453), .b(output_10_6), .y(output_9_453));
wire output_11_453, output_11_6, output_10_453;
mixer gate_output_10_453(.a(output_11_453), .b(output_11_6), .y(output_10_453));
wire output_12_453, output_12_6, output_11_453;
mixer gate_output_11_453(.a(output_12_453), .b(output_12_6), .y(output_11_453));
wire output_13_453, output_13_6, output_12_453;
mixer gate_output_12_453(.a(output_13_453), .b(output_13_6), .y(output_12_453));
wire output_14_453, output_14_6, output_13_453;
mixer gate_output_13_453(.a(output_14_453), .b(output_14_6), .y(output_13_453));
wire output_15_453, output_15_6, output_14_453;
mixer gate_output_14_453(.a(output_15_453), .b(output_15_6), .y(output_14_453));
wire output_16_453, output_16_6, output_15_453;
mixer gate_output_15_453(.a(output_16_453), .b(output_16_6), .y(output_15_453));
wire output_1_454, output_1_7, output_0_454;
mixer gate_output_0_454(.a(output_1_454), .b(output_1_7), .y(output_0_454));
wire output_2_454, output_2_7, output_1_454;
mixer gate_output_1_454(.a(output_2_454), .b(output_2_7), .y(output_1_454));
wire output_3_454, output_3_7, output_2_454;
mixer gate_output_2_454(.a(output_3_454), .b(output_3_7), .y(output_2_454));
wire output_4_454, output_4_7, output_3_454;
mixer gate_output_3_454(.a(output_4_454), .b(output_4_7), .y(output_3_454));
wire output_5_454, output_5_7, output_4_454;
mixer gate_output_4_454(.a(output_5_454), .b(output_5_7), .y(output_4_454));
wire output_6_454, output_6_7, output_5_454;
mixer gate_output_5_454(.a(output_6_454), .b(output_6_7), .y(output_5_454));
wire output_7_454, output_7_7, output_6_454;
mixer gate_output_6_454(.a(output_7_454), .b(output_7_7), .y(output_6_454));
wire output_8_454, output_8_7, output_7_454;
mixer gate_output_7_454(.a(output_8_454), .b(output_8_7), .y(output_7_454));
wire output_9_454, output_9_7, output_8_454;
mixer gate_output_8_454(.a(output_9_454), .b(output_9_7), .y(output_8_454));
wire output_10_454, output_10_7, output_9_454;
mixer gate_output_9_454(.a(output_10_454), .b(output_10_7), .y(output_9_454));
wire output_11_454, output_11_7, output_10_454;
mixer gate_output_10_454(.a(output_11_454), .b(output_11_7), .y(output_10_454));
wire output_12_454, output_12_7, output_11_454;
mixer gate_output_11_454(.a(output_12_454), .b(output_12_7), .y(output_11_454));
wire output_13_454, output_13_7, output_12_454;
mixer gate_output_12_454(.a(output_13_454), .b(output_13_7), .y(output_12_454));
wire output_14_454, output_14_7, output_13_454;
mixer gate_output_13_454(.a(output_14_454), .b(output_14_7), .y(output_13_454));
wire output_15_454, output_15_7, output_14_454;
mixer gate_output_14_454(.a(output_15_454), .b(output_15_7), .y(output_14_454));
wire output_16_454, output_16_7, output_15_454;
mixer gate_output_15_454(.a(output_16_454), .b(output_16_7), .y(output_15_454));
wire output_1_455, output_1_8, output_0_455;
mixer gate_output_0_455(.a(output_1_455), .b(output_1_8), .y(output_0_455));
wire output_2_455, output_2_8, output_1_455;
mixer gate_output_1_455(.a(output_2_455), .b(output_2_8), .y(output_1_455));
wire output_3_455, output_3_8, output_2_455;
mixer gate_output_2_455(.a(output_3_455), .b(output_3_8), .y(output_2_455));
wire output_4_455, output_4_8, output_3_455;
mixer gate_output_3_455(.a(output_4_455), .b(output_4_8), .y(output_3_455));
wire output_5_455, output_5_8, output_4_455;
mixer gate_output_4_455(.a(output_5_455), .b(output_5_8), .y(output_4_455));
wire output_6_455, output_6_8, output_5_455;
mixer gate_output_5_455(.a(output_6_455), .b(output_6_8), .y(output_5_455));
wire output_7_455, output_7_8, output_6_455;
mixer gate_output_6_455(.a(output_7_455), .b(output_7_8), .y(output_6_455));
wire output_8_455, output_8_8, output_7_455;
mixer gate_output_7_455(.a(output_8_455), .b(output_8_8), .y(output_7_455));
wire output_9_455, output_9_8, output_8_455;
mixer gate_output_8_455(.a(output_9_455), .b(output_9_8), .y(output_8_455));
wire output_10_455, output_10_8, output_9_455;
mixer gate_output_9_455(.a(output_10_455), .b(output_10_8), .y(output_9_455));
wire output_11_455, output_11_8, output_10_455;
mixer gate_output_10_455(.a(output_11_455), .b(output_11_8), .y(output_10_455));
wire output_12_455, output_12_8, output_11_455;
mixer gate_output_11_455(.a(output_12_455), .b(output_12_8), .y(output_11_455));
wire output_13_455, output_13_8, output_12_455;
mixer gate_output_12_455(.a(output_13_455), .b(output_13_8), .y(output_12_455));
wire output_14_455, output_14_8, output_13_455;
mixer gate_output_13_455(.a(output_14_455), .b(output_14_8), .y(output_13_455));
wire output_15_455, output_15_8, output_14_455;
mixer gate_output_14_455(.a(output_15_455), .b(output_15_8), .y(output_14_455));
wire output_16_455, output_16_8, output_15_455;
mixer gate_output_15_455(.a(output_16_455), .b(output_16_8), .y(output_15_455));
wire output_1_456, output_1_9, output_0_456;
mixer gate_output_0_456(.a(output_1_456), .b(output_1_9), .y(output_0_456));
wire output_2_456, output_2_9, output_1_456;
mixer gate_output_1_456(.a(output_2_456), .b(output_2_9), .y(output_1_456));
wire output_3_456, output_3_9, output_2_456;
mixer gate_output_2_456(.a(output_3_456), .b(output_3_9), .y(output_2_456));
wire output_4_456, output_4_9, output_3_456;
mixer gate_output_3_456(.a(output_4_456), .b(output_4_9), .y(output_3_456));
wire output_5_456, output_5_9, output_4_456;
mixer gate_output_4_456(.a(output_5_456), .b(output_5_9), .y(output_4_456));
wire output_6_456, output_6_9, output_5_456;
mixer gate_output_5_456(.a(output_6_456), .b(output_6_9), .y(output_5_456));
wire output_7_456, output_7_9, output_6_456;
mixer gate_output_6_456(.a(output_7_456), .b(output_7_9), .y(output_6_456));
wire output_8_456, output_8_9, output_7_456;
mixer gate_output_7_456(.a(output_8_456), .b(output_8_9), .y(output_7_456));
wire output_9_456, output_9_9, output_8_456;
mixer gate_output_8_456(.a(output_9_456), .b(output_9_9), .y(output_8_456));
wire output_10_456, output_10_9, output_9_456;
mixer gate_output_9_456(.a(output_10_456), .b(output_10_9), .y(output_9_456));
wire output_11_456, output_11_9, output_10_456;
mixer gate_output_10_456(.a(output_11_456), .b(output_11_9), .y(output_10_456));
wire output_12_456, output_12_9, output_11_456;
mixer gate_output_11_456(.a(output_12_456), .b(output_12_9), .y(output_11_456));
wire output_13_456, output_13_9, output_12_456;
mixer gate_output_12_456(.a(output_13_456), .b(output_13_9), .y(output_12_456));
wire output_14_456, output_14_9, output_13_456;
mixer gate_output_13_456(.a(output_14_456), .b(output_14_9), .y(output_13_456));
wire output_15_456, output_15_9, output_14_456;
mixer gate_output_14_456(.a(output_15_456), .b(output_15_9), .y(output_14_456));
wire output_16_456, output_16_9, output_15_456;
mixer gate_output_15_456(.a(output_16_456), .b(output_16_9), .y(output_15_456));
wire output_1_457, output_1_10, output_0_457;
mixer gate_output_0_457(.a(output_1_457), .b(output_1_10), .y(output_0_457));
wire output_2_457, output_2_10, output_1_457;
mixer gate_output_1_457(.a(output_2_457), .b(output_2_10), .y(output_1_457));
wire output_3_457, output_3_10, output_2_457;
mixer gate_output_2_457(.a(output_3_457), .b(output_3_10), .y(output_2_457));
wire output_4_457, output_4_10, output_3_457;
mixer gate_output_3_457(.a(output_4_457), .b(output_4_10), .y(output_3_457));
wire output_5_457, output_5_10, output_4_457;
mixer gate_output_4_457(.a(output_5_457), .b(output_5_10), .y(output_4_457));
wire output_6_457, output_6_10, output_5_457;
mixer gate_output_5_457(.a(output_6_457), .b(output_6_10), .y(output_5_457));
wire output_7_457, output_7_10, output_6_457;
mixer gate_output_6_457(.a(output_7_457), .b(output_7_10), .y(output_6_457));
wire output_8_457, output_8_10, output_7_457;
mixer gate_output_7_457(.a(output_8_457), .b(output_8_10), .y(output_7_457));
wire output_9_457, output_9_10, output_8_457;
mixer gate_output_8_457(.a(output_9_457), .b(output_9_10), .y(output_8_457));
wire output_10_457, output_10_10, output_9_457;
mixer gate_output_9_457(.a(output_10_457), .b(output_10_10), .y(output_9_457));
wire output_11_457, output_11_10, output_10_457;
mixer gate_output_10_457(.a(output_11_457), .b(output_11_10), .y(output_10_457));
wire output_12_457, output_12_10, output_11_457;
mixer gate_output_11_457(.a(output_12_457), .b(output_12_10), .y(output_11_457));
wire output_13_457, output_13_10, output_12_457;
mixer gate_output_12_457(.a(output_13_457), .b(output_13_10), .y(output_12_457));
wire output_14_457, output_14_10, output_13_457;
mixer gate_output_13_457(.a(output_14_457), .b(output_14_10), .y(output_13_457));
wire output_15_457, output_15_10, output_14_457;
mixer gate_output_14_457(.a(output_15_457), .b(output_15_10), .y(output_14_457));
wire output_16_457, output_16_10, output_15_457;
mixer gate_output_15_457(.a(output_16_457), .b(output_16_10), .y(output_15_457));
wire output_1_458, output_1_11, output_0_458;
mixer gate_output_0_458(.a(output_1_458), .b(output_1_11), .y(output_0_458));
wire output_2_458, output_2_11, output_1_458;
mixer gate_output_1_458(.a(output_2_458), .b(output_2_11), .y(output_1_458));
wire output_3_458, output_3_11, output_2_458;
mixer gate_output_2_458(.a(output_3_458), .b(output_3_11), .y(output_2_458));
wire output_4_458, output_4_11, output_3_458;
mixer gate_output_3_458(.a(output_4_458), .b(output_4_11), .y(output_3_458));
wire output_5_458, output_5_11, output_4_458;
mixer gate_output_4_458(.a(output_5_458), .b(output_5_11), .y(output_4_458));
wire output_6_458, output_6_11, output_5_458;
mixer gate_output_5_458(.a(output_6_458), .b(output_6_11), .y(output_5_458));
wire output_7_458, output_7_11, output_6_458;
mixer gate_output_6_458(.a(output_7_458), .b(output_7_11), .y(output_6_458));
wire output_8_458, output_8_11, output_7_458;
mixer gate_output_7_458(.a(output_8_458), .b(output_8_11), .y(output_7_458));
wire output_9_458, output_9_11, output_8_458;
mixer gate_output_8_458(.a(output_9_458), .b(output_9_11), .y(output_8_458));
wire output_10_458, output_10_11, output_9_458;
mixer gate_output_9_458(.a(output_10_458), .b(output_10_11), .y(output_9_458));
wire output_11_458, output_11_11, output_10_458;
mixer gate_output_10_458(.a(output_11_458), .b(output_11_11), .y(output_10_458));
wire output_12_458, output_12_11, output_11_458;
mixer gate_output_11_458(.a(output_12_458), .b(output_12_11), .y(output_11_458));
wire output_13_458, output_13_11, output_12_458;
mixer gate_output_12_458(.a(output_13_458), .b(output_13_11), .y(output_12_458));
wire output_14_458, output_14_11, output_13_458;
mixer gate_output_13_458(.a(output_14_458), .b(output_14_11), .y(output_13_458));
wire output_15_458, output_15_11, output_14_458;
mixer gate_output_14_458(.a(output_15_458), .b(output_15_11), .y(output_14_458));
wire output_16_458, output_16_11, output_15_458;
mixer gate_output_15_458(.a(output_16_458), .b(output_16_11), .y(output_15_458));
wire output_1_459, output_1_12, output_0_459;
mixer gate_output_0_459(.a(output_1_459), .b(output_1_12), .y(output_0_459));
wire output_2_459, output_2_12, output_1_459;
mixer gate_output_1_459(.a(output_2_459), .b(output_2_12), .y(output_1_459));
wire output_3_459, output_3_12, output_2_459;
mixer gate_output_2_459(.a(output_3_459), .b(output_3_12), .y(output_2_459));
wire output_4_459, output_4_12, output_3_459;
mixer gate_output_3_459(.a(output_4_459), .b(output_4_12), .y(output_3_459));
wire output_5_459, output_5_12, output_4_459;
mixer gate_output_4_459(.a(output_5_459), .b(output_5_12), .y(output_4_459));
wire output_6_459, output_6_12, output_5_459;
mixer gate_output_5_459(.a(output_6_459), .b(output_6_12), .y(output_5_459));
wire output_7_459, output_7_12, output_6_459;
mixer gate_output_6_459(.a(output_7_459), .b(output_7_12), .y(output_6_459));
wire output_8_459, output_8_12, output_7_459;
mixer gate_output_7_459(.a(output_8_459), .b(output_8_12), .y(output_7_459));
wire output_9_459, output_9_12, output_8_459;
mixer gate_output_8_459(.a(output_9_459), .b(output_9_12), .y(output_8_459));
wire output_10_459, output_10_12, output_9_459;
mixer gate_output_9_459(.a(output_10_459), .b(output_10_12), .y(output_9_459));
wire output_11_459, output_11_12, output_10_459;
mixer gate_output_10_459(.a(output_11_459), .b(output_11_12), .y(output_10_459));
wire output_12_459, output_12_12, output_11_459;
mixer gate_output_11_459(.a(output_12_459), .b(output_12_12), .y(output_11_459));
wire output_13_459, output_13_12, output_12_459;
mixer gate_output_12_459(.a(output_13_459), .b(output_13_12), .y(output_12_459));
wire output_14_459, output_14_12, output_13_459;
mixer gate_output_13_459(.a(output_14_459), .b(output_14_12), .y(output_13_459));
wire output_15_459, output_15_12, output_14_459;
mixer gate_output_14_459(.a(output_15_459), .b(output_15_12), .y(output_14_459));
wire output_16_459, output_16_12, output_15_459;
mixer gate_output_15_459(.a(output_16_459), .b(output_16_12), .y(output_15_459));
wire output_1_460, output_1_13, output_0_460;
mixer gate_output_0_460(.a(output_1_460), .b(output_1_13), .y(output_0_460));
wire output_2_460, output_2_13, output_1_460;
mixer gate_output_1_460(.a(output_2_460), .b(output_2_13), .y(output_1_460));
wire output_3_460, output_3_13, output_2_460;
mixer gate_output_2_460(.a(output_3_460), .b(output_3_13), .y(output_2_460));
wire output_4_460, output_4_13, output_3_460;
mixer gate_output_3_460(.a(output_4_460), .b(output_4_13), .y(output_3_460));
wire output_5_460, output_5_13, output_4_460;
mixer gate_output_4_460(.a(output_5_460), .b(output_5_13), .y(output_4_460));
wire output_6_460, output_6_13, output_5_460;
mixer gate_output_5_460(.a(output_6_460), .b(output_6_13), .y(output_5_460));
wire output_7_460, output_7_13, output_6_460;
mixer gate_output_6_460(.a(output_7_460), .b(output_7_13), .y(output_6_460));
wire output_8_460, output_8_13, output_7_460;
mixer gate_output_7_460(.a(output_8_460), .b(output_8_13), .y(output_7_460));
wire output_9_460, output_9_13, output_8_460;
mixer gate_output_8_460(.a(output_9_460), .b(output_9_13), .y(output_8_460));
wire output_10_460, output_10_13, output_9_460;
mixer gate_output_9_460(.a(output_10_460), .b(output_10_13), .y(output_9_460));
wire output_11_460, output_11_13, output_10_460;
mixer gate_output_10_460(.a(output_11_460), .b(output_11_13), .y(output_10_460));
wire output_12_460, output_12_13, output_11_460;
mixer gate_output_11_460(.a(output_12_460), .b(output_12_13), .y(output_11_460));
wire output_13_460, output_13_13, output_12_460;
mixer gate_output_12_460(.a(output_13_460), .b(output_13_13), .y(output_12_460));
wire output_14_460, output_14_13, output_13_460;
mixer gate_output_13_460(.a(output_14_460), .b(output_14_13), .y(output_13_460));
wire output_15_460, output_15_13, output_14_460;
mixer gate_output_14_460(.a(output_15_460), .b(output_15_13), .y(output_14_460));
wire output_16_460, output_16_13, output_15_460;
mixer gate_output_15_460(.a(output_16_460), .b(output_16_13), .y(output_15_460));
wire output_1_461, output_1_14, output_0_461;
mixer gate_output_0_461(.a(output_1_461), .b(output_1_14), .y(output_0_461));
wire output_2_461, output_2_14, output_1_461;
mixer gate_output_1_461(.a(output_2_461), .b(output_2_14), .y(output_1_461));
wire output_3_461, output_3_14, output_2_461;
mixer gate_output_2_461(.a(output_3_461), .b(output_3_14), .y(output_2_461));
wire output_4_461, output_4_14, output_3_461;
mixer gate_output_3_461(.a(output_4_461), .b(output_4_14), .y(output_3_461));
wire output_5_461, output_5_14, output_4_461;
mixer gate_output_4_461(.a(output_5_461), .b(output_5_14), .y(output_4_461));
wire output_6_461, output_6_14, output_5_461;
mixer gate_output_5_461(.a(output_6_461), .b(output_6_14), .y(output_5_461));
wire output_7_461, output_7_14, output_6_461;
mixer gate_output_6_461(.a(output_7_461), .b(output_7_14), .y(output_6_461));
wire output_8_461, output_8_14, output_7_461;
mixer gate_output_7_461(.a(output_8_461), .b(output_8_14), .y(output_7_461));
wire output_9_461, output_9_14, output_8_461;
mixer gate_output_8_461(.a(output_9_461), .b(output_9_14), .y(output_8_461));
wire output_10_461, output_10_14, output_9_461;
mixer gate_output_9_461(.a(output_10_461), .b(output_10_14), .y(output_9_461));
wire output_11_461, output_11_14, output_10_461;
mixer gate_output_10_461(.a(output_11_461), .b(output_11_14), .y(output_10_461));
wire output_12_461, output_12_14, output_11_461;
mixer gate_output_11_461(.a(output_12_461), .b(output_12_14), .y(output_11_461));
wire output_13_461, output_13_14, output_12_461;
mixer gate_output_12_461(.a(output_13_461), .b(output_13_14), .y(output_12_461));
wire output_14_461, output_14_14, output_13_461;
mixer gate_output_13_461(.a(output_14_461), .b(output_14_14), .y(output_13_461));
wire output_15_461, output_15_14, output_14_461;
mixer gate_output_14_461(.a(output_15_461), .b(output_15_14), .y(output_14_461));
wire output_16_461, output_16_14, output_15_461;
mixer gate_output_15_461(.a(output_16_461), .b(output_16_14), .y(output_15_461));
wire output_1_462, output_1_15, output_0_462;
mixer gate_output_0_462(.a(output_1_462), .b(output_1_15), .y(output_0_462));
wire output_2_462, output_2_15, output_1_462;
mixer gate_output_1_462(.a(output_2_462), .b(output_2_15), .y(output_1_462));
wire output_3_462, output_3_15, output_2_462;
mixer gate_output_2_462(.a(output_3_462), .b(output_3_15), .y(output_2_462));
wire output_4_462, output_4_15, output_3_462;
mixer gate_output_3_462(.a(output_4_462), .b(output_4_15), .y(output_3_462));
wire output_5_462, output_5_15, output_4_462;
mixer gate_output_4_462(.a(output_5_462), .b(output_5_15), .y(output_4_462));
wire output_6_462, output_6_15, output_5_462;
mixer gate_output_5_462(.a(output_6_462), .b(output_6_15), .y(output_5_462));
wire output_7_462, output_7_15, output_6_462;
mixer gate_output_6_462(.a(output_7_462), .b(output_7_15), .y(output_6_462));
wire output_8_462, output_8_15, output_7_462;
mixer gate_output_7_462(.a(output_8_462), .b(output_8_15), .y(output_7_462));
wire output_9_462, output_9_15, output_8_462;
mixer gate_output_8_462(.a(output_9_462), .b(output_9_15), .y(output_8_462));
wire output_10_462, output_10_15, output_9_462;
mixer gate_output_9_462(.a(output_10_462), .b(output_10_15), .y(output_9_462));
wire output_11_462, output_11_15, output_10_462;
mixer gate_output_10_462(.a(output_11_462), .b(output_11_15), .y(output_10_462));
wire output_12_462, output_12_15, output_11_462;
mixer gate_output_11_462(.a(output_12_462), .b(output_12_15), .y(output_11_462));
wire output_13_462, output_13_15, output_12_462;
mixer gate_output_12_462(.a(output_13_462), .b(output_13_15), .y(output_12_462));
wire output_14_462, output_14_15, output_13_462;
mixer gate_output_13_462(.a(output_14_462), .b(output_14_15), .y(output_13_462));
wire output_15_462, output_15_15, output_14_462;
mixer gate_output_14_462(.a(output_15_462), .b(output_15_15), .y(output_14_462));
wire output_16_462, output_16_15, output_15_462;
mixer gate_output_15_462(.a(output_16_462), .b(output_16_15), .y(output_15_462));
wire output_1_463, output_1_0, output_0_463;
mixer gate_output_0_463(.a(output_1_463), .b(output_1_0), .y(output_0_463));
wire output_2_463, output_2_0, output_1_463;
mixer gate_output_1_463(.a(output_2_463), .b(output_2_0), .y(output_1_463));
wire output_3_463, output_3_0, output_2_463;
mixer gate_output_2_463(.a(output_3_463), .b(output_3_0), .y(output_2_463));
wire output_4_463, output_4_0, output_3_463;
mixer gate_output_3_463(.a(output_4_463), .b(output_4_0), .y(output_3_463));
wire output_5_463, output_5_0, output_4_463;
mixer gate_output_4_463(.a(output_5_463), .b(output_5_0), .y(output_4_463));
wire output_6_463, output_6_0, output_5_463;
mixer gate_output_5_463(.a(output_6_463), .b(output_6_0), .y(output_5_463));
wire output_7_463, output_7_0, output_6_463;
mixer gate_output_6_463(.a(output_7_463), .b(output_7_0), .y(output_6_463));
wire output_8_463, output_8_0, output_7_463;
mixer gate_output_7_463(.a(output_8_463), .b(output_8_0), .y(output_7_463));
wire output_9_463, output_9_0, output_8_463;
mixer gate_output_8_463(.a(output_9_463), .b(output_9_0), .y(output_8_463));
wire output_10_463, output_10_0, output_9_463;
mixer gate_output_9_463(.a(output_10_463), .b(output_10_0), .y(output_9_463));
wire output_11_463, output_11_0, output_10_463;
mixer gate_output_10_463(.a(output_11_463), .b(output_11_0), .y(output_10_463));
wire output_12_463, output_12_0, output_11_463;
mixer gate_output_11_463(.a(output_12_463), .b(output_12_0), .y(output_11_463));
wire output_13_463, output_13_0, output_12_463;
mixer gate_output_12_463(.a(output_13_463), .b(output_13_0), .y(output_12_463));
wire output_14_463, output_14_0, output_13_463;
mixer gate_output_13_463(.a(output_14_463), .b(output_14_0), .y(output_13_463));
wire output_15_463, output_15_0, output_14_463;
mixer gate_output_14_463(.a(output_15_463), .b(output_15_0), .y(output_14_463));
wire output_16_463, output_16_0, output_15_463;
mixer gate_output_15_463(.a(output_16_463), .b(output_16_0), .y(output_15_463));
wire output_1_464, output_1_1, output_0_464;
mixer gate_output_0_464(.a(output_1_464), .b(output_1_1), .y(output_0_464));
wire output_2_464, output_2_1, output_1_464;
mixer gate_output_1_464(.a(output_2_464), .b(output_2_1), .y(output_1_464));
wire output_3_464, output_3_1, output_2_464;
mixer gate_output_2_464(.a(output_3_464), .b(output_3_1), .y(output_2_464));
wire output_4_464, output_4_1, output_3_464;
mixer gate_output_3_464(.a(output_4_464), .b(output_4_1), .y(output_3_464));
wire output_5_464, output_5_1, output_4_464;
mixer gate_output_4_464(.a(output_5_464), .b(output_5_1), .y(output_4_464));
wire output_6_464, output_6_1, output_5_464;
mixer gate_output_5_464(.a(output_6_464), .b(output_6_1), .y(output_5_464));
wire output_7_464, output_7_1, output_6_464;
mixer gate_output_6_464(.a(output_7_464), .b(output_7_1), .y(output_6_464));
wire output_8_464, output_8_1, output_7_464;
mixer gate_output_7_464(.a(output_8_464), .b(output_8_1), .y(output_7_464));
wire output_9_464, output_9_1, output_8_464;
mixer gate_output_8_464(.a(output_9_464), .b(output_9_1), .y(output_8_464));
wire output_10_464, output_10_1, output_9_464;
mixer gate_output_9_464(.a(output_10_464), .b(output_10_1), .y(output_9_464));
wire output_11_464, output_11_1, output_10_464;
mixer gate_output_10_464(.a(output_11_464), .b(output_11_1), .y(output_10_464));
wire output_12_464, output_12_1, output_11_464;
mixer gate_output_11_464(.a(output_12_464), .b(output_12_1), .y(output_11_464));
wire output_13_464, output_13_1, output_12_464;
mixer gate_output_12_464(.a(output_13_464), .b(output_13_1), .y(output_12_464));
wire output_14_464, output_14_1, output_13_464;
mixer gate_output_13_464(.a(output_14_464), .b(output_14_1), .y(output_13_464));
wire output_15_464, output_15_1, output_14_464;
mixer gate_output_14_464(.a(output_15_464), .b(output_15_1), .y(output_14_464));
wire output_16_464, output_16_1, output_15_464;
mixer gate_output_15_464(.a(output_16_464), .b(output_16_1), .y(output_15_464));
wire output_1_465, output_1_2, output_0_465;
mixer gate_output_0_465(.a(output_1_465), .b(output_1_2), .y(output_0_465));
wire output_2_465, output_2_2, output_1_465;
mixer gate_output_1_465(.a(output_2_465), .b(output_2_2), .y(output_1_465));
wire output_3_465, output_3_2, output_2_465;
mixer gate_output_2_465(.a(output_3_465), .b(output_3_2), .y(output_2_465));
wire output_4_465, output_4_2, output_3_465;
mixer gate_output_3_465(.a(output_4_465), .b(output_4_2), .y(output_3_465));
wire output_5_465, output_5_2, output_4_465;
mixer gate_output_4_465(.a(output_5_465), .b(output_5_2), .y(output_4_465));
wire output_6_465, output_6_2, output_5_465;
mixer gate_output_5_465(.a(output_6_465), .b(output_6_2), .y(output_5_465));
wire output_7_465, output_7_2, output_6_465;
mixer gate_output_6_465(.a(output_7_465), .b(output_7_2), .y(output_6_465));
wire output_8_465, output_8_2, output_7_465;
mixer gate_output_7_465(.a(output_8_465), .b(output_8_2), .y(output_7_465));
wire output_9_465, output_9_2, output_8_465;
mixer gate_output_8_465(.a(output_9_465), .b(output_9_2), .y(output_8_465));
wire output_10_465, output_10_2, output_9_465;
mixer gate_output_9_465(.a(output_10_465), .b(output_10_2), .y(output_9_465));
wire output_11_465, output_11_2, output_10_465;
mixer gate_output_10_465(.a(output_11_465), .b(output_11_2), .y(output_10_465));
wire output_12_465, output_12_2, output_11_465;
mixer gate_output_11_465(.a(output_12_465), .b(output_12_2), .y(output_11_465));
wire output_13_465, output_13_2, output_12_465;
mixer gate_output_12_465(.a(output_13_465), .b(output_13_2), .y(output_12_465));
wire output_14_465, output_14_2, output_13_465;
mixer gate_output_13_465(.a(output_14_465), .b(output_14_2), .y(output_13_465));
wire output_15_465, output_15_2, output_14_465;
mixer gate_output_14_465(.a(output_15_465), .b(output_15_2), .y(output_14_465));
wire output_16_465, output_16_2, output_15_465;
mixer gate_output_15_465(.a(output_16_465), .b(output_16_2), .y(output_15_465));
wire output_1_466, output_1_3, output_0_466;
mixer gate_output_0_466(.a(output_1_466), .b(output_1_3), .y(output_0_466));
wire output_2_466, output_2_3, output_1_466;
mixer gate_output_1_466(.a(output_2_466), .b(output_2_3), .y(output_1_466));
wire output_3_466, output_3_3, output_2_466;
mixer gate_output_2_466(.a(output_3_466), .b(output_3_3), .y(output_2_466));
wire output_4_466, output_4_3, output_3_466;
mixer gate_output_3_466(.a(output_4_466), .b(output_4_3), .y(output_3_466));
wire output_5_466, output_5_3, output_4_466;
mixer gate_output_4_466(.a(output_5_466), .b(output_5_3), .y(output_4_466));
wire output_6_466, output_6_3, output_5_466;
mixer gate_output_5_466(.a(output_6_466), .b(output_6_3), .y(output_5_466));
wire output_7_466, output_7_3, output_6_466;
mixer gate_output_6_466(.a(output_7_466), .b(output_7_3), .y(output_6_466));
wire output_8_466, output_8_3, output_7_466;
mixer gate_output_7_466(.a(output_8_466), .b(output_8_3), .y(output_7_466));
wire output_9_466, output_9_3, output_8_466;
mixer gate_output_8_466(.a(output_9_466), .b(output_9_3), .y(output_8_466));
wire output_10_466, output_10_3, output_9_466;
mixer gate_output_9_466(.a(output_10_466), .b(output_10_3), .y(output_9_466));
wire output_11_466, output_11_3, output_10_466;
mixer gate_output_10_466(.a(output_11_466), .b(output_11_3), .y(output_10_466));
wire output_12_466, output_12_3, output_11_466;
mixer gate_output_11_466(.a(output_12_466), .b(output_12_3), .y(output_11_466));
wire output_13_466, output_13_3, output_12_466;
mixer gate_output_12_466(.a(output_13_466), .b(output_13_3), .y(output_12_466));
wire output_14_466, output_14_3, output_13_466;
mixer gate_output_13_466(.a(output_14_466), .b(output_14_3), .y(output_13_466));
wire output_15_466, output_15_3, output_14_466;
mixer gate_output_14_466(.a(output_15_466), .b(output_15_3), .y(output_14_466));
wire output_16_466, output_16_3, output_15_466;
mixer gate_output_15_466(.a(output_16_466), .b(output_16_3), .y(output_15_466));
wire output_1_467, output_1_4, output_0_467;
mixer gate_output_0_467(.a(output_1_467), .b(output_1_4), .y(output_0_467));
wire output_2_467, output_2_4, output_1_467;
mixer gate_output_1_467(.a(output_2_467), .b(output_2_4), .y(output_1_467));
wire output_3_467, output_3_4, output_2_467;
mixer gate_output_2_467(.a(output_3_467), .b(output_3_4), .y(output_2_467));
wire output_4_467, output_4_4, output_3_467;
mixer gate_output_3_467(.a(output_4_467), .b(output_4_4), .y(output_3_467));
wire output_5_467, output_5_4, output_4_467;
mixer gate_output_4_467(.a(output_5_467), .b(output_5_4), .y(output_4_467));
wire output_6_467, output_6_4, output_5_467;
mixer gate_output_5_467(.a(output_6_467), .b(output_6_4), .y(output_5_467));
wire output_7_467, output_7_4, output_6_467;
mixer gate_output_6_467(.a(output_7_467), .b(output_7_4), .y(output_6_467));
wire output_8_467, output_8_4, output_7_467;
mixer gate_output_7_467(.a(output_8_467), .b(output_8_4), .y(output_7_467));
wire output_9_467, output_9_4, output_8_467;
mixer gate_output_8_467(.a(output_9_467), .b(output_9_4), .y(output_8_467));
wire output_10_467, output_10_4, output_9_467;
mixer gate_output_9_467(.a(output_10_467), .b(output_10_4), .y(output_9_467));
wire output_11_467, output_11_4, output_10_467;
mixer gate_output_10_467(.a(output_11_467), .b(output_11_4), .y(output_10_467));
wire output_12_467, output_12_4, output_11_467;
mixer gate_output_11_467(.a(output_12_467), .b(output_12_4), .y(output_11_467));
wire output_13_467, output_13_4, output_12_467;
mixer gate_output_12_467(.a(output_13_467), .b(output_13_4), .y(output_12_467));
wire output_14_467, output_14_4, output_13_467;
mixer gate_output_13_467(.a(output_14_467), .b(output_14_4), .y(output_13_467));
wire output_15_467, output_15_4, output_14_467;
mixer gate_output_14_467(.a(output_15_467), .b(output_15_4), .y(output_14_467));
wire output_16_467, output_16_4, output_15_467;
mixer gate_output_15_467(.a(output_16_467), .b(output_16_4), .y(output_15_467));
wire output_1_468, output_1_5, output_0_468;
mixer gate_output_0_468(.a(output_1_468), .b(output_1_5), .y(output_0_468));
wire output_2_468, output_2_5, output_1_468;
mixer gate_output_1_468(.a(output_2_468), .b(output_2_5), .y(output_1_468));
wire output_3_468, output_3_5, output_2_468;
mixer gate_output_2_468(.a(output_3_468), .b(output_3_5), .y(output_2_468));
wire output_4_468, output_4_5, output_3_468;
mixer gate_output_3_468(.a(output_4_468), .b(output_4_5), .y(output_3_468));
wire output_5_468, output_5_5, output_4_468;
mixer gate_output_4_468(.a(output_5_468), .b(output_5_5), .y(output_4_468));
wire output_6_468, output_6_5, output_5_468;
mixer gate_output_5_468(.a(output_6_468), .b(output_6_5), .y(output_5_468));
wire output_7_468, output_7_5, output_6_468;
mixer gate_output_6_468(.a(output_7_468), .b(output_7_5), .y(output_6_468));
wire output_8_468, output_8_5, output_7_468;
mixer gate_output_7_468(.a(output_8_468), .b(output_8_5), .y(output_7_468));
wire output_9_468, output_9_5, output_8_468;
mixer gate_output_8_468(.a(output_9_468), .b(output_9_5), .y(output_8_468));
wire output_10_468, output_10_5, output_9_468;
mixer gate_output_9_468(.a(output_10_468), .b(output_10_5), .y(output_9_468));
wire output_11_468, output_11_5, output_10_468;
mixer gate_output_10_468(.a(output_11_468), .b(output_11_5), .y(output_10_468));
wire output_12_468, output_12_5, output_11_468;
mixer gate_output_11_468(.a(output_12_468), .b(output_12_5), .y(output_11_468));
wire output_13_468, output_13_5, output_12_468;
mixer gate_output_12_468(.a(output_13_468), .b(output_13_5), .y(output_12_468));
wire output_14_468, output_14_5, output_13_468;
mixer gate_output_13_468(.a(output_14_468), .b(output_14_5), .y(output_13_468));
wire output_15_468, output_15_5, output_14_468;
mixer gate_output_14_468(.a(output_15_468), .b(output_15_5), .y(output_14_468));
wire output_16_468, output_16_5, output_15_468;
mixer gate_output_15_468(.a(output_16_468), .b(output_16_5), .y(output_15_468));
wire output_1_469, output_1_6, output_0_469;
mixer gate_output_0_469(.a(output_1_469), .b(output_1_6), .y(output_0_469));
wire output_2_469, output_2_6, output_1_469;
mixer gate_output_1_469(.a(output_2_469), .b(output_2_6), .y(output_1_469));
wire output_3_469, output_3_6, output_2_469;
mixer gate_output_2_469(.a(output_3_469), .b(output_3_6), .y(output_2_469));
wire output_4_469, output_4_6, output_3_469;
mixer gate_output_3_469(.a(output_4_469), .b(output_4_6), .y(output_3_469));
wire output_5_469, output_5_6, output_4_469;
mixer gate_output_4_469(.a(output_5_469), .b(output_5_6), .y(output_4_469));
wire output_6_469, output_6_6, output_5_469;
mixer gate_output_5_469(.a(output_6_469), .b(output_6_6), .y(output_5_469));
wire output_7_469, output_7_6, output_6_469;
mixer gate_output_6_469(.a(output_7_469), .b(output_7_6), .y(output_6_469));
wire output_8_469, output_8_6, output_7_469;
mixer gate_output_7_469(.a(output_8_469), .b(output_8_6), .y(output_7_469));
wire output_9_469, output_9_6, output_8_469;
mixer gate_output_8_469(.a(output_9_469), .b(output_9_6), .y(output_8_469));
wire output_10_469, output_10_6, output_9_469;
mixer gate_output_9_469(.a(output_10_469), .b(output_10_6), .y(output_9_469));
wire output_11_469, output_11_6, output_10_469;
mixer gate_output_10_469(.a(output_11_469), .b(output_11_6), .y(output_10_469));
wire output_12_469, output_12_6, output_11_469;
mixer gate_output_11_469(.a(output_12_469), .b(output_12_6), .y(output_11_469));
wire output_13_469, output_13_6, output_12_469;
mixer gate_output_12_469(.a(output_13_469), .b(output_13_6), .y(output_12_469));
wire output_14_469, output_14_6, output_13_469;
mixer gate_output_13_469(.a(output_14_469), .b(output_14_6), .y(output_13_469));
wire output_15_469, output_15_6, output_14_469;
mixer gate_output_14_469(.a(output_15_469), .b(output_15_6), .y(output_14_469));
wire output_16_469, output_16_6, output_15_469;
mixer gate_output_15_469(.a(output_16_469), .b(output_16_6), .y(output_15_469));
wire output_1_470, output_1_7, output_0_470;
mixer gate_output_0_470(.a(output_1_470), .b(output_1_7), .y(output_0_470));
wire output_2_470, output_2_7, output_1_470;
mixer gate_output_1_470(.a(output_2_470), .b(output_2_7), .y(output_1_470));
wire output_3_470, output_3_7, output_2_470;
mixer gate_output_2_470(.a(output_3_470), .b(output_3_7), .y(output_2_470));
wire output_4_470, output_4_7, output_3_470;
mixer gate_output_3_470(.a(output_4_470), .b(output_4_7), .y(output_3_470));
wire output_5_470, output_5_7, output_4_470;
mixer gate_output_4_470(.a(output_5_470), .b(output_5_7), .y(output_4_470));
wire output_6_470, output_6_7, output_5_470;
mixer gate_output_5_470(.a(output_6_470), .b(output_6_7), .y(output_5_470));
wire output_7_470, output_7_7, output_6_470;
mixer gate_output_6_470(.a(output_7_470), .b(output_7_7), .y(output_6_470));
wire output_8_470, output_8_7, output_7_470;
mixer gate_output_7_470(.a(output_8_470), .b(output_8_7), .y(output_7_470));
wire output_9_470, output_9_7, output_8_470;
mixer gate_output_8_470(.a(output_9_470), .b(output_9_7), .y(output_8_470));
wire output_10_470, output_10_7, output_9_470;
mixer gate_output_9_470(.a(output_10_470), .b(output_10_7), .y(output_9_470));
wire output_11_470, output_11_7, output_10_470;
mixer gate_output_10_470(.a(output_11_470), .b(output_11_7), .y(output_10_470));
wire output_12_470, output_12_7, output_11_470;
mixer gate_output_11_470(.a(output_12_470), .b(output_12_7), .y(output_11_470));
wire output_13_470, output_13_7, output_12_470;
mixer gate_output_12_470(.a(output_13_470), .b(output_13_7), .y(output_12_470));
wire output_14_470, output_14_7, output_13_470;
mixer gate_output_13_470(.a(output_14_470), .b(output_14_7), .y(output_13_470));
wire output_15_470, output_15_7, output_14_470;
mixer gate_output_14_470(.a(output_15_470), .b(output_15_7), .y(output_14_470));
wire output_16_470, output_16_7, output_15_470;
mixer gate_output_15_470(.a(output_16_470), .b(output_16_7), .y(output_15_470));
wire output_1_471, output_1_8, output_0_471;
mixer gate_output_0_471(.a(output_1_471), .b(output_1_8), .y(output_0_471));
wire output_2_471, output_2_8, output_1_471;
mixer gate_output_1_471(.a(output_2_471), .b(output_2_8), .y(output_1_471));
wire output_3_471, output_3_8, output_2_471;
mixer gate_output_2_471(.a(output_3_471), .b(output_3_8), .y(output_2_471));
wire output_4_471, output_4_8, output_3_471;
mixer gate_output_3_471(.a(output_4_471), .b(output_4_8), .y(output_3_471));
wire output_5_471, output_5_8, output_4_471;
mixer gate_output_4_471(.a(output_5_471), .b(output_5_8), .y(output_4_471));
wire output_6_471, output_6_8, output_5_471;
mixer gate_output_5_471(.a(output_6_471), .b(output_6_8), .y(output_5_471));
wire output_7_471, output_7_8, output_6_471;
mixer gate_output_6_471(.a(output_7_471), .b(output_7_8), .y(output_6_471));
wire output_8_471, output_8_8, output_7_471;
mixer gate_output_7_471(.a(output_8_471), .b(output_8_8), .y(output_7_471));
wire output_9_471, output_9_8, output_8_471;
mixer gate_output_8_471(.a(output_9_471), .b(output_9_8), .y(output_8_471));
wire output_10_471, output_10_8, output_9_471;
mixer gate_output_9_471(.a(output_10_471), .b(output_10_8), .y(output_9_471));
wire output_11_471, output_11_8, output_10_471;
mixer gate_output_10_471(.a(output_11_471), .b(output_11_8), .y(output_10_471));
wire output_12_471, output_12_8, output_11_471;
mixer gate_output_11_471(.a(output_12_471), .b(output_12_8), .y(output_11_471));
wire output_13_471, output_13_8, output_12_471;
mixer gate_output_12_471(.a(output_13_471), .b(output_13_8), .y(output_12_471));
wire output_14_471, output_14_8, output_13_471;
mixer gate_output_13_471(.a(output_14_471), .b(output_14_8), .y(output_13_471));
wire output_15_471, output_15_8, output_14_471;
mixer gate_output_14_471(.a(output_15_471), .b(output_15_8), .y(output_14_471));
wire output_16_471, output_16_8, output_15_471;
mixer gate_output_15_471(.a(output_16_471), .b(output_16_8), .y(output_15_471));
wire output_1_472, output_1_9, output_0_472;
mixer gate_output_0_472(.a(output_1_472), .b(output_1_9), .y(output_0_472));
wire output_2_472, output_2_9, output_1_472;
mixer gate_output_1_472(.a(output_2_472), .b(output_2_9), .y(output_1_472));
wire output_3_472, output_3_9, output_2_472;
mixer gate_output_2_472(.a(output_3_472), .b(output_3_9), .y(output_2_472));
wire output_4_472, output_4_9, output_3_472;
mixer gate_output_3_472(.a(output_4_472), .b(output_4_9), .y(output_3_472));
wire output_5_472, output_5_9, output_4_472;
mixer gate_output_4_472(.a(output_5_472), .b(output_5_9), .y(output_4_472));
wire output_6_472, output_6_9, output_5_472;
mixer gate_output_5_472(.a(output_6_472), .b(output_6_9), .y(output_5_472));
wire output_7_472, output_7_9, output_6_472;
mixer gate_output_6_472(.a(output_7_472), .b(output_7_9), .y(output_6_472));
wire output_8_472, output_8_9, output_7_472;
mixer gate_output_7_472(.a(output_8_472), .b(output_8_9), .y(output_7_472));
wire output_9_472, output_9_9, output_8_472;
mixer gate_output_8_472(.a(output_9_472), .b(output_9_9), .y(output_8_472));
wire output_10_472, output_10_9, output_9_472;
mixer gate_output_9_472(.a(output_10_472), .b(output_10_9), .y(output_9_472));
wire output_11_472, output_11_9, output_10_472;
mixer gate_output_10_472(.a(output_11_472), .b(output_11_9), .y(output_10_472));
wire output_12_472, output_12_9, output_11_472;
mixer gate_output_11_472(.a(output_12_472), .b(output_12_9), .y(output_11_472));
wire output_13_472, output_13_9, output_12_472;
mixer gate_output_12_472(.a(output_13_472), .b(output_13_9), .y(output_12_472));
wire output_14_472, output_14_9, output_13_472;
mixer gate_output_13_472(.a(output_14_472), .b(output_14_9), .y(output_13_472));
wire output_15_472, output_15_9, output_14_472;
mixer gate_output_14_472(.a(output_15_472), .b(output_15_9), .y(output_14_472));
wire output_16_472, output_16_9, output_15_472;
mixer gate_output_15_472(.a(output_16_472), .b(output_16_9), .y(output_15_472));
wire output_1_473, output_1_10, output_0_473;
mixer gate_output_0_473(.a(output_1_473), .b(output_1_10), .y(output_0_473));
wire output_2_473, output_2_10, output_1_473;
mixer gate_output_1_473(.a(output_2_473), .b(output_2_10), .y(output_1_473));
wire output_3_473, output_3_10, output_2_473;
mixer gate_output_2_473(.a(output_3_473), .b(output_3_10), .y(output_2_473));
wire output_4_473, output_4_10, output_3_473;
mixer gate_output_3_473(.a(output_4_473), .b(output_4_10), .y(output_3_473));
wire output_5_473, output_5_10, output_4_473;
mixer gate_output_4_473(.a(output_5_473), .b(output_5_10), .y(output_4_473));
wire output_6_473, output_6_10, output_5_473;
mixer gate_output_5_473(.a(output_6_473), .b(output_6_10), .y(output_5_473));
wire output_7_473, output_7_10, output_6_473;
mixer gate_output_6_473(.a(output_7_473), .b(output_7_10), .y(output_6_473));
wire output_8_473, output_8_10, output_7_473;
mixer gate_output_7_473(.a(output_8_473), .b(output_8_10), .y(output_7_473));
wire output_9_473, output_9_10, output_8_473;
mixer gate_output_8_473(.a(output_9_473), .b(output_9_10), .y(output_8_473));
wire output_10_473, output_10_10, output_9_473;
mixer gate_output_9_473(.a(output_10_473), .b(output_10_10), .y(output_9_473));
wire output_11_473, output_11_10, output_10_473;
mixer gate_output_10_473(.a(output_11_473), .b(output_11_10), .y(output_10_473));
wire output_12_473, output_12_10, output_11_473;
mixer gate_output_11_473(.a(output_12_473), .b(output_12_10), .y(output_11_473));
wire output_13_473, output_13_10, output_12_473;
mixer gate_output_12_473(.a(output_13_473), .b(output_13_10), .y(output_12_473));
wire output_14_473, output_14_10, output_13_473;
mixer gate_output_13_473(.a(output_14_473), .b(output_14_10), .y(output_13_473));
wire output_15_473, output_15_10, output_14_473;
mixer gate_output_14_473(.a(output_15_473), .b(output_15_10), .y(output_14_473));
wire output_16_473, output_16_10, output_15_473;
mixer gate_output_15_473(.a(output_16_473), .b(output_16_10), .y(output_15_473));
wire output_1_474, output_1_11, output_0_474;
mixer gate_output_0_474(.a(output_1_474), .b(output_1_11), .y(output_0_474));
wire output_2_474, output_2_11, output_1_474;
mixer gate_output_1_474(.a(output_2_474), .b(output_2_11), .y(output_1_474));
wire output_3_474, output_3_11, output_2_474;
mixer gate_output_2_474(.a(output_3_474), .b(output_3_11), .y(output_2_474));
wire output_4_474, output_4_11, output_3_474;
mixer gate_output_3_474(.a(output_4_474), .b(output_4_11), .y(output_3_474));
wire output_5_474, output_5_11, output_4_474;
mixer gate_output_4_474(.a(output_5_474), .b(output_5_11), .y(output_4_474));
wire output_6_474, output_6_11, output_5_474;
mixer gate_output_5_474(.a(output_6_474), .b(output_6_11), .y(output_5_474));
wire output_7_474, output_7_11, output_6_474;
mixer gate_output_6_474(.a(output_7_474), .b(output_7_11), .y(output_6_474));
wire output_8_474, output_8_11, output_7_474;
mixer gate_output_7_474(.a(output_8_474), .b(output_8_11), .y(output_7_474));
wire output_9_474, output_9_11, output_8_474;
mixer gate_output_8_474(.a(output_9_474), .b(output_9_11), .y(output_8_474));
wire output_10_474, output_10_11, output_9_474;
mixer gate_output_9_474(.a(output_10_474), .b(output_10_11), .y(output_9_474));
wire output_11_474, output_11_11, output_10_474;
mixer gate_output_10_474(.a(output_11_474), .b(output_11_11), .y(output_10_474));
wire output_12_474, output_12_11, output_11_474;
mixer gate_output_11_474(.a(output_12_474), .b(output_12_11), .y(output_11_474));
wire output_13_474, output_13_11, output_12_474;
mixer gate_output_12_474(.a(output_13_474), .b(output_13_11), .y(output_12_474));
wire output_14_474, output_14_11, output_13_474;
mixer gate_output_13_474(.a(output_14_474), .b(output_14_11), .y(output_13_474));
wire output_15_474, output_15_11, output_14_474;
mixer gate_output_14_474(.a(output_15_474), .b(output_15_11), .y(output_14_474));
wire output_16_474, output_16_11, output_15_474;
mixer gate_output_15_474(.a(output_16_474), .b(output_16_11), .y(output_15_474));
wire output_1_475, output_1_12, output_0_475;
mixer gate_output_0_475(.a(output_1_475), .b(output_1_12), .y(output_0_475));
wire output_2_475, output_2_12, output_1_475;
mixer gate_output_1_475(.a(output_2_475), .b(output_2_12), .y(output_1_475));
wire output_3_475, output_3_12, output_2_475;
mixer gate_output_2_475(.a(output_3_475), .b(output_3_12), .y(output_2_475));
wire output_4_475, output_4_12, output_3_475;
mixer gate_output_3_475(.a(output_4_475), .b(output_4_12), .y(output_3_475));
wire output_5_475, output_5_12, output_4_475;
mixer gate_output_4_475(.a(output_5_475), .b(output_5_12), .y(output_4_475));
wire output_6_475, output_6_12, output_5_475;
mixer gate_output_5_475(.a(output_6_475), .b(output_6_12), .y(output_5_475));
wire output_7_475, output_7_12, output_6_475;
mixer gate_output_6_475(.a(output_7_475), .b(output_7_12), .y(output_6_475));
wire output_8_475, output_8_12, output_7_475;
mixer gate_output_7_475(.a(output_8_475), .b(output_8_12), .y(output_7_475));
wire output_9_475, output_9_12, output_8_475;
mixer gate_output_8_475(.a(output_9_475), .b(output_9_12), .y(output_8_475));
wire output_10_475, output_10_12, output_9_475;
mixer gate_output_9_475(.a(output_10_475), .b(output_10_12), .y(output_9_475));
wire output_11_475, output_11_12, output_10_475;
mixer gate_output_10_475(.a(output_11_475), .b(output_11_12), .y(output_10_475));
wire output_12_475, output_12_12, output_11_475;
mixer gate_output_11_475(.a(output_12_475), .b(output_12_12), .y(output_11_475));
wire output_13_475, output_13_12, output_12_475;
mixer gate_output_12_475(.a(output_13_475), .b(output_13_12), .y(output_12_475));
wire output_14_475, output_14_12, output_13_475;
mixer gate_output_13_475(.a(output_14_475), .b(output_14_12), .y(output_13_475));
wire output_15_475, output_15_12, output_14_475;
mixer gate_output_14_475(.a(output_15_475), .b(output_15_12), .y(output_14_475));
wire output_16_475, output_16_12, output_15_475;
mixer gate_output_15_475(.a(output_16_475), .b(output_16_12), .y(output_15_475));
wire output_1_476, output_1_13, output_0_476;
mixer gate_output_0_476(.a(output_1_476), .b(output_1_13), .y(output_0_476));
wire output_2_476, output_2_13, output_1_476;
mixer gate_output_1_476(.a(output_2_476), .b(output_2_13), .y(output_1_476));
wire output_3_476, output_3_13, output_2_476;
mixer gate_output_2_476(.a(output_3_476), .b(output_3_13), .y(output_2_476));
wire output_4_476, output_4_13, output_3_476;
mixer gate_output_3_476(.a(output_4_476), .b(output_4_13), .y(output_3_476));
wire output_5_476, output_5_13, output_4_476;
mixer gate_output_4_476(.a(output_5_476), .b(output_5_13), .y(output_4_476));
wire output_6_476, output_6_13, output_5_476;
mixer gate_output_5_476(.a(output_6_476), .b(output_6_13), .y(output_5_476));
wire output_7_476, output_7_13, output_6_476;
mixer gate_output_6_476(.a(output_7_476), .b(output_7_13), .y(output_6_476));
wire output_8_476, output_8_13, output_7_476;
mixer gate_output_7_476(.a(output_8_476), .b(output_8_13), .y(output_7_476));
wire output_9_476, output_9_13, output_8_476;
mixer gate_output_8_476(.a(output_9_476), .b(output_9_13), .y(output_8_476));
wire output_10_476, output_10_13, output_9_476;
mixer gate_output_9_476(.a(output_10_476), .b(output_10_13), .y(output_9_476));
wire output_11_476, output_11_13, output_10_476;
mixer gate_output_10_476(.a(output_11_476), .b(output_11_13), .y(output_10_476));
wire output_12_476, output_12_13, output_11_476;
mixer gate_output_11_476(.a(output_12_476), .b(output_12_13), .y(output_11_476));
wire output_13_476, output_13_13, output_12_476;
mixer gate_output_12_476(.a(output_13_476), .b(output_13_13), .y(output_12_476));
wire output_14_476, output_14_13, output_13_476;
mixer gate_output_13_476(.a(output_14_476), .b(output_14_13), .y(output_13_476));
wire output_15_476, output_15_13, output_14_476;
mixer gate_output_14_476(.a(output_15_476), .b(output_15_13), .y(output_14_476));
wire output_16_476, output_16_13, output_15_476;
mixer gate_output_15_476(.a(output_16_476), .b(output_16_13), .y(output_15_476));
wire output_1_477, output_1_14, output_0_477;
mixer gate_output_0_477(.a(output_1_477), .b(output_1_14), .y(output_0_477));
wire output_2_477, output_2_14, output_1_477;
mixer gate_output_1_477(.a(output_2_477), .b(output_2_14), .y(output_1_477));
wire output_3_477, output_3_14, output_2_477;
mixer gate_output_2_477(.a(output_3_477), .b(output_3_14), .y(output_2_477));
wire output_4_477, output_4_14, output_3_477;
mixer gate_output_3_477(.a(output_4_477), .b(output_4_14), .y(output_3_477));
wire output_5_477, output_5_14, output_4_477;
mixer gate_output_4_477(.a(output_5_477), .b(output_5_14), .y(output_4_477));
wire output_6_477, output_6_14, output_5_477;
mixer gate_output_5_477(.a(output_6_477), .b(output_6_14), .y(output_5_477));
wire output_7_477, output_7_14, output_6_477;
mixer gate_output_6_477(.a(output_7_477), .b(output_7_14), .y(output_6_477));
wire output_8_477, output_8_14, output_7_477;
mixer gate_output_7_477(.a(output_8_477), .b(output_8_14), .y(output_7_477));
wire output_9_477, output_9_14, output_8_477;
mixer gate_output_8_477(.a(output_9_477), .b(output_9_14), .y(output_8_477));
wire output_10_477, output_10_14, output_9_477;
mixer gate_output_9_477(.a(output_10_477), .b(output_10_14), .y(output_9_477));
wire output_11_477, output_11_14, output_10_477;
mixer gate_output_10_477(.a(output_11_477), .b(output_11_14), .y(output_10_477));
wire output_12_477, output_12_14, output_11_477;
mixer gate_output_11_477(.a(output_12_477), .b(output_12_14), .y(output_11_477));
wire output_13_477, output_13_14, output_12_477;
mixer gate_output_12_477(.a(output_13_477), .b(output_13_14), .y(output_12_477));
wire output_14_477, output_14_14, output_13_477;
mixer gate_output_13_477(.a(output_14_477), .b(output_14_14), .y(output_13_477));
wire output_15_477, output_15_14, output_14_477;
mixer gate_output_14_477(.a(output_15_477), .b(output_15_14), .y(output_14_477));
wire output_16_477, output_16_14, output_15_477;
mixer gate_output_15_477(.a(output_16_477), .b(output_16_14), .y(output_15_477));
wire output_1_478, output_1_15, output_0_478;
mixer gate_output_0_478(.a(output_1_478), .b(output_1_15), .y(output_0_478));
wire output_2_478, output_2_15, output_1_478;
mixer gate_output_1_478(.a(output_2_478), .b(output_2_15), .y(output_1_478));
wire output_3_478, output_3_15, output_2_478;
mixer gate_output_2_478(.a(output_3_478), .b(output_3_15), .y(output_2_478));
wire output_4_478, output_4_15, output_3_478;
mixer gate_output_3_478(.a(output_4_478), .b(output_4_15), .y(output_3_478));
wire output_5_478, output_5_15, output_4_478;
mixer gate_output_4_478(.a(output_5_478), .b(output_5_15), .y(output_4_478));
wire output_6_478, output_6_15, output_5_478;
mixer gate_output_5_478(.a(output_6_478), .b(output_6_15), .y(output_5_478));
wire output_7_478, output_7_15, output_6_478;
mixer gate_output_6_478(.a(output_7_478), .b(output_7_15), .y(output_6_478));
wire output_8_478, output_8_15, output_7_478;
mixer gate_output_7_478(.a(output_8_478), .b(output_8_15), .y(output_7_478));
wire output_9_478, output_9_15, output_8_478;
mixer gate_output_8_478(.a(output_9_478), .b(output_9_15), .y(output_8_478));
wire output_10_478, output_10_15, output_9_478;
mixer gate_output_9_478(.a(output_10_478), .b(output_10_15), .y(output_9_478));
wire output_11_478, output_11_15, output_10_478;
mixer gate_output_10_478(.a(output_11_478), .b(output_11_15), .y(output_10_478));
wire output_12_478, output_12_15, output_11_478;
mixer gate_output_11_478(.a(output_12_478), .b(output_12_15), .y(output_11_478));
wire output_13_478, output_13_15, output_12_478;
mixer gate_output_12_478(.a(output_13_478), .b(output_13_15), .y(output_12_478));
wire output_14_478, output_14_15, output_13_478;
mixer gate_output_13_478(.a(output_14_478), .b(output_14_15), .y(output_13_478));
wire output_15_478, output_15_15, output_14_478;
mixer gate_output_14_478(.a(output_15_478), .b(output_15_15), .y(output_14_478));
wire output_16_478, output_16_15, output_15_478;
mixer gate_output_15_478(.a(output_16_478), .b(output_16_15), .y(output_15_478));
wire output_1_479, output_1_0, output_0_479;
mixer gate_output_0_479(.a(output_1_479), .b(output_1_0), .y(output_0_479));
wire output_2_479, output_2_0, output_1_479;
mixer gate_output_1_479(.a(output_2_479), .b(output_2_0), .y(output_1_479));
wire output_3_479, output_3_0, output_2_479;
mixer gate_output_2_479(.a(output_3_479), .b(output_3_0), .y(output_2_479));
wire output_4_479, output_4_0, output_3_479;
mixer gate_output_3_479(.a(output_4_479), .b(output_4_0), .y(output_3_479));
wire output_5_479, output_5_0, output_4_479;
mixer gate_output_4_479(.a(output_5_479), .b(output_5_0), .y(output_4_479));
wire output_6_479, output_6_0, output_5_479;
mixer gate_output_5_479(.a(output_6_479), .b(output_6_0), .y(output_5_479));
wire output_7_479, output_7_0, output_6_479;
mixer gate_output_6_479(.a(output_7_479), .b(output_7_0), .y(output_6_479));
wire output_8_479, output_8_0, output_7_479;
mixer gate_output_7_479(.a(output_8_479), .b(output_8_0), .y(output_7_479));
wire output_9_479, output_9_0, output_8_479;
mixer gate_output_8_479(.a(output_9_479), .b(output_9_0), .y(output_8_479));
wire output_10_479, output_10_0, output_9_479;
mixer gate_output_9_479(.a(output_10_479), .b(output_10_0), .y(output_9_479));
wire output_11_479, output_11_0, output_10_479;
mixer gate_output_10_479(.a(output_11_479), .b(output_11_0), .y(output_10_479));
wire output_12_479, output_12_0, output_11_479;
mixer gate_output_11_479(.a(output_12_479), .b(output_12_0), .y(output_11_479));
wire output_13_479, output_13_0, output_12_479;
mixer gate_output_12_479(.a(output_13_479), .b(output_13_0), .y(output_12_479));
wire output_14_479, output_14_0, output_13_479;
mixer gate_output_13_479(.a(output_14_479), .b(output_14_0), .y(output_13_479));
wire output_15_479, output_15_0, output_14_479;
mixer gate_output_14_479(.a(output_15_479), .b(output_15_0), .y(output_14_479));
wire output_16_479, output_16_0, output_15_479;
mixer gate_output_15_479(.a(output_16_479), .b(output_16_0), .y(output_15_479));
wire output_1_480, output_1_1, output_0_480;
mixer gate_output_0_480(.a(output_1_480), .b(output_1_1), .y(output_0_480));
wire output_2_480, output_2_1, output_1_480;
mixer gate_output_1_480(.a(output_2_480), .b(output_2_1), .y(output_1_480));
wire output_3_480, output_3_1, output_2_480;
mixer gate_output_2_480(.a(output_3_480), .b(output_3_1), .y(output_2_480));
wire output_4_480, output_4_1, output_3_480;
mixer gate_output_3_480(.a(output_4_480), .b(output_4_1), .y(output_3_480));
wire output_5_480, output_5_1, output_4_480;
mixer gate_output_4_480(.a(output_5_480), .b(output_5_1), .y(output_4_480));
wire output_6_480, output_6_1, output_5_480;
mixer gate_output_5_480(.a(output_6_480), .b(output_6_1), .y(output_5_480));
wire output_7_480, output_7_1, output_6_480;
mixer gate_output_6_480(.a(output_7_480), .b(output_7_1), .y(output_6_480));
wire output_8_480, output_8_1, output_7_480;
mixer gate_output_7_480(.a(output_8_480), .b(output_8_1), .y(output_7_480));
wire output_9_480, output_9_1, output_8_480;
mixer gate_output_8_480(.a(output_9_480), .b(output_9_1), .y(output_8_480));
wire output_10_480, output_10_1, output_9_480;
mixer gate_output_9_480(.a(output_10_480), .b(output_10_1), .y(output_9_480));
wire output_11_480, output_11_1, output_10_480;
mixer gate_output_10_480(.a(output_11_480), .b(output_11_1), .y(output_10_480));
wire output_12_480, output_12_1, output_11_480;
mixer gate_output_11_480(.a(output_12_480), .b(output_12_1), .y(output_11_480));
wire output_13_480, output_13_1, output_12_480;
mixer gate_output_12_480(.a(output_13_480), .b(output_13_1), .y(output_12_480));
wire output_14_480, output_14_1, output_13_480;
mixer gate_output_13_480(.a(output_14_480), .b(output_14_1), .y(output_13_480));
wire output_15_480, output_15_1, output_14_480;
mixer gate_output_14_480(.a(output_15_480), .b(output_15_1), .y(output_14_480));
wire output_16_480, output_16_1, output_15_480;
mixer gate_output_15_480(.a(output_16_480), .b(output_16_1), .y(output_15_480));
wire output_1_481, output_1_2, output_0_481;
mixer gate_output_0_481(.a(output_1_481), .b(output_1_2), .y(output_0_481));
wire output_2_481, output_2_2, output_1_481;
mixer gate_output_1_481(.a(output_2_481), .b(output_2_2), .y(output_1_481));
wire output_3_481, output_3_2, output_2_481;
mixer gate_output_2_481(.a(output_3_481), .b(output_3_2), .y(output_2_481));
wire output_4_481, output_4_2, output_3_481;
mixer gate_output_3_481(.a(output_4_481), .b(output_4_2), .y(output_3_481));
wire output_5_481, output_5_2, output_4_481;
mixer gate_output_4_481(.a(output_5_481), .b(output_5_2), .y(output_4_481));
wire output_6_481, output_6_2, output_5_481;
mixer gate_output_5_481(.a(output_6_481), .b(output_6_2), .y(output_5_481));
wire output_7_481, output_7_2, output_6_481;
mixer gate_output_6_481(.a(output_7_481), .b(output_7_2), .y(output_6_481));
wire output_8_481, output_8_2, output_7_481;
mixer gate_output_7_481(.a(output_8_481), .b(output_8_2), .y(output_7_481));
wire output_9_481, output_9_2, output_8_481;
mixer gate_output_8_481(.a(output_9_481), .b(output_9_2), .y(output_8_481));
wire output_10_481, output_10_2, output_9_481;
mixer gate_output_9_481(.a(output_10_481), .b(output_10_2), .y(output_9_481));
wire output_11_481, output_11_2, output_10_481;
mixer gate_output_10_481(.a(output_11_481), .b(output_11_2), .y(output_10_481));
wire output_12_481, output_12_2, output_11_481;
mixer gate_output_11_481(.a(output_12_481), .b(output_12_2), .y(output_11_481));
wire output_13_481, output_13_2, output_12_481;
mixer gate_output_12_481(.a(output_13_481), .b(output_13_2), .y(output_12_481));
wire output_14_481, output_14_2, output_13_481;
mixer gate_output_13_481(.a(output_14_481), .b(output_14_2), .y(output_13_481));
wire output_15_481, output_15_2, output_14_481;
mixer gate_output_14_481(.a(output_15_481), .b(output_15_2), .y(output_14_481));
wire output_16_481, output_16_2, output_15_481;
mixer gate_output_15_481(.a(output_16_481), .b(output_16_2), .y(output_15_481));
wire output_1_482, output_1_3, output_0_482;
mixer gate_output_0_482(.a(output_1_482), .b(output_1_3), .y(output_0_482));
wire output_2_482, output_2_3, output_1_482;
mixer gate_output_1_482(.a(output_2_482), .b(output_2_3), .y(output_1_482));
wire output_3_482, output_3_3, output_2_482;
mixer gate_output_2_482(.a(output_3_482), .b(output_3_3), .y(output_2_482));
wire output_4_482, output_4_3, output_3_482;
mixer gate_output_3_482(.a(output_4_482), .b(output_4_3), .y(output_3_482));
wire output_5_482, output_5_3, output_4_482;
mixer gate_output_4_482(.a(output_5_482), .b(output_5_3), .y(output_4_482));
wire output_6_482, output_6_3, output_5_482;
mixer gate_output_5_482(.a(output_6_482), .b(output_6_3), .y(output_5_482));
wire output_7_482, output_7_3, output_6_482;
mixer gate_output_6_482(.a(output_7_482), .b(output_7_3), .y(output_6_482));
wire output_8_482, output_8_3, output_7_482;
mixer gate_output_7_482(.a(output_8_482), .b(output_8_3), .y(output_7_482));
wire output_9_482, output_9_3, output_8_482;
mixer gate_output_8_482(.a(output_9_482), .b(output_9_3), .y(output_8_482));
wire output_10_482, output_10_3, output_9_482;
mixer gate_output_9_482(.a(output_10_482), .b(output_10_3), .y(output_9_482));
wire output_11_482, output_11_3, output_10_482;
mixer gate_output_10_482(.a(output_11_482), .b(output_11_3), .y(output_10_482));
wire output_12_482, output_12_3, output_11_482;
mixer gate_output_11_482(.a(output_12_482), .b(output_12_3), .y(output_11_482));
wire output_13_482, output_13_3, output_12_482;
mixer gate_output_12_482(.a(output_13_482), .b(output_13_3), .y(output_12_482));
wire output_14_482, output_14_3, output_13_482;
mixer gate_output_13_482(.a(output_14_482), .b(output_14_3), .y(output_13_482));
wire output_15_482, output_15_3, output_14_482;
mixer gate_output_14_482(.a(output_15_482), .b(output_15_3), .y(output_14_482));
wire output_16_482, output_16_3, output_15_482;
mixer gate_output_15_482(.a(output_16_482), .b(output_16_3), .y(output_15_482));
wire output_1_483, output_1_4, output_0_483;
mixer gate_output_0_483(.a(output_1_483), .b(output_1_4), .y(output_0_483));
wire output_2_483, output_2_4, output_1_483;
mixer gate_output_1_483(.a(output_2_483), .b(output_2_4), .y(output_1_483));
wire output_3_483, output_3_4, output_2_483;
mixer gate_output_2_483(.a(output_3_483), .b(output_3_4), .y(output_2_483));
wire output_4_483, output_4_4, output_3_483;
mixer gate_output_3_483(.a(output_4_483), .b(output_4_4), .y(output_3_483));
wire output_5_483, output_5_4, output_4_483;
mixer gate_output_4_483(.a(output_5_483), .b(output_5_4), .y(output_4_483));
wire output_6_483, output_6_4, output_5_483;
mixer gate_output_5_483(.a(output_6_483), .b(output_6_4), .y(output_5_483));
wire output_7_483, output_7_4, output_6_483;
mixer gate_output_6_483(.a(output_7_483), .b(output_7_4), .y(output_6_483));
wire output_8_483, output_8_4, output_7_483;
mixer gate_output_7_483(.a(output_8_483), .b(output_8_4), .y(output_7_483));
wire output_9_483, output_9_4, output_8_483;
mixer gate_output_8_483(.a(output_9_483), .b(output_9_4), .y(output_8_483));
wire output_10_483, output_10_4, output_9_483;
mixer gate_output_9_483(.a(output_10_483), .b(output_10_4), .y(output_9_483));
wire output_11_483, output_11_4, output_10_483;
mixer gate_output_10_483(.a(output_11_483), .b(output_11_4), .y(output_10_483));
wire output_12_483, output_12_4, output_11_483;
mixer gate_output_11_483(.a(output_12_483), .b(output_12_4), .y(output_11_483));
wire output_13_483, output_13_4, output_12_483;
mixer gate_output_12_483(.a(output_13_483), .b(output_13_4), .y(output_12_483));
wire output_14_483, output_14_4, output_13_483;
mixer gate_output_13_483(.a(output_14_483), .b(output_14_4), .y(output_13_483));
wire output_15_483, output_15_4, output_14_483;
mixer gate_output_14_483(.a(output_15_483), .b(output_15_4), .y(output_14_483));
wire output_16_483, output_16_4, output_15_483;
mixer gate_output_15_483(.a(output_16_483), .b(output_16_4), .y(output_15_483));
wire output_1_484, output_1_5, output_0_484;
mixer gate_output_0_484(.a(output_1_484), .b(output_1_5), .y(output_0_484));
wire output_2_484, output_2_5, output_1_484;
mixer gate_output_1_484(.a(output_2_484), .b(output_2_5), .y(output_1_484));
wire output_3_484, output_3_5, output_2_484;
mixer gate_output_2_484(.a(output_3_484), .b(output_3_5), .y(output_2_484));
wire output_4_484, output_4_5, output_3_484;
mixer gate_output_3_484(.a(output_4_484), .b(output_4_5), .y(output_3_484));
wire output_5_484, output_5_5, output_4_484;
mixer gate_output_4_484(.a(output_5_484), .b(output_5_5), .y(output_4_484));
wire output_6_484, output_6_5, output_5_484;
mixer gate_output_5_484(.a(output_6_484), .b(output_6_5), .y(output_5_484));
wire output_7_484, output_7_5, output_6_484;
mixer gate_output_6_484(.a(output_7_484), .b(output_7_5), .y(output_6_484));
wire output_8_484, output_8_5, output_7_484;
mixer gate_output_7_484(.a(output_8_484), .b(output_8_5), .y(output_7_484));
wire output_9_484, output_9_5, output_8_484;
mixer gate_output_8_484(.a(output_9_484), .b(output_9_5), .y(output_8_484));
wire output_10_484, output_10_5, output_9_484;
mixer gate_output_9_484(.a(output_10_484), .b(output_10_5), .y(output_9_484));
wire output_11_484, output_11_5, output_10_484;
mixer gate_output_10_484(.a(output_11_484), .b(output_11_5), .y(output_10_484));
wire output_12_484, output_12_5, output_11_484;
mixer gate_output_11_484(.a(output_12_484), .b(output_12_5), .y(output_11_484));
wire output_13_484, output_13_5, output_12_484;
mixer gate_output_12_484(.a(output_13_484), .b(output_13_5), .y(output_12_484));
wire output_14_484, output_14_5, output_13_484;
mixer gate_output_13_484(.a(output_14_484), .b(output_14_5), .y(output_13_484));
wire output_15_484, output_15_5, output_14_484;
mixer gate_output_14_484(.a(output_15_484), .b(output_15_5), .y(output_14_484));
wire output_16_484, output_16_5, output_15_484;
mixer gate_output_15_484(.a(output_16_484), .b(output_16_5), .y(output_15_484));
wire output_1_485, output_1_6, output_0_485;
mixer gate_output_0_485(.a(output_1_485), .b(output_1_6), .y(output_0_485));
wire output_2_485, output_2_6, output_1_485;
mixer gate_output_1_485(.a(output_2_485), .b(output_2_6), .y(output_1_485));
wire output_3_485, output_3_6, output_2_485;
mixer gate_output_2_485(.a(output_3_485), .b(output_3_6), .y(output_2_485));
wire output_4_485, output_4_6, output_3_485;
mixer gate_output_3_485(.a(output_4_485), .b(output_4_6), .y(output_3_485));
wire output_5_485, output_5_6, output_4_485;
mixer gate_output_4_485(.a(output_5_485), .b(output_5_6), .y(output_4_485));
wire output_6_485, output_6_6, output_5_485;
mixer gate_output_5_485(.a(output_6_485), .b(output_6_6), .y(output_5_485));
wire output_7_485, output_7_6, output_6_485;
mixer gate_output_6_485(.a(output_7_485), .b(output_7_6), .y(output_6_485));
wire output_8_485, output_8_6, output_7_485;
mixer gate_output_7_485(.a(output_8_485), .b(output_8_6), .y(output_7_485));
wire output_9_485, output_9_6, output_8_485;
mixer gate_output_8_485(.a(output_9_485), .b(output_9_6), .y(output_8_485));
wire output_10_485, output_10_6, output_9_485;
mixer gate_output_9_485(.a(output_10_485), .b(output_10_6), .y(output_9_485));
wire output_11_485, output_11_6, output_10_485;
mixer gate_output_10_485(.a(output_11_485), .b(output_11_6), .y(output_10_485));
wire output_12_485, output_12_6, output_11_485;
mixer gate_output_11_485(.a(output_12_485), .b(output_12_6), .y(output_11_485));
wire output_13_485, output_13_6, output_12_485;
mixer gate_output_12_485(.a(output_13_485), .b(output_13_6), .y(output_12_485));
wire output_14_485, output_14_6, output_13_485;
mixer gate_output_13_485(.a(output_14_485), .b(output_14_6), .y(output_13_485));
wire output_15_485, output_15_6, output_14_485;
mixer gate_output_14_485(.a(output_15_485), .b(output_15_6), .y(output_14_485));
wire output_16_485, output_16_6, output_15_485;
mixer gate_output_15_485(.a(output_16_485), .b(output_16_6), .y(output_15_485));
wire output_1_486, output_1_7, output_0_486;
mixer gate_output_0_486(.a(output_1_486), .b(output_1_7), .y(output_0_486));
wire output_2_486, output_2_7, output_1_486;
mixer gate_output_1_486(.a(output_2_486), .b(output_2_7), .y(output_1_486));
wire output_3_486, output_3_7, output_2_486;
mixer gate_output_2_486(.a(output_3_486), .b(output_3_7), .y(output_2_486));
wire output_4_486, output_4_7, output_3_486;
mixer gate_output_3_486(.a(output_4_486), .b(output_4_7), .y(output_3_486));
wire output_5_486, output_5_7, output_4_486;
mixer gate_output_4_486(.a(output_5_486), .b(output_5_7), .y(output_4_486));
wire output_6_486, output_6_7, output_5_486;
mixer gate_output_5_486(.a(output_6_486), .b(output_6_7), .y(output_5_486));
wire output_7_486, output_7_7, output_6_486;
mixer gate_output_6_486(.a(output_7_486), .b(output_7_7), .y(output_6_486));
wire output_8_486, output_8_7, output_7_486;
mixer gate_output_7_486(.a(output_8_486), .b(output_8_7), .y(output_7_486));
wire output_9_486, output_9_7, output_8_486;
mixer gate_output_8_486(.a(output_9_486), .b(output_9_7), .y(output_8_486));
wire output_10_486, output_10_7, output_9_486;
mixer gate_output_9_486(.a(output_10_486), .b(output_10_7), .y(output_9_486));
wire output_11_486, output_11_7, output_10_486;
mixer gate_output_10_486(.a(output_11_486), .b(output_11_7), .y(output_10_486));
wire output_12_486, output_12_7, output_11_486;
mixer gate_output_11_486(.a(output_12_486), .b(output_12_7), .y(output_11_486));
wire output_13_486, output_13_7, output_12_486;
mixer gate_output_12_486(.a(output_13_486), .b(output_13_7), .y(output_12_486));
wire output_14_486, output_14_7, output_13_486;
mixer gate_output_13_486(.a(output_14_486), .b(output_14_7), .y(output_13_486));
wire output_15_486, output_15_7, output_14_486;
mixer gate_output_14_486(.a(output_15_486), .b(output_15_7), .y(output_14_486));
wire output_16_486, output_16_7, output_15_486;
mixer gate_output_15_486(.a(output_16_486), .b(output_16_7), .y(output_15_486));
wire output_1_487, output_1_8, output_0_487;
mixer gate_output_0_487(.a(output_1_487), .b(output_1_8), .y(output_0_487));
wire output_2_487, output_2_8, output_1_487;
mixer gate_output_1_487(.a(output_2_487), .b(output_2_8), .y(output_1_487));
wire output_3_487, output_3_8, output_2_487;
mixer gate_output_2_487(.a(output_3_487), .b(output_3_8), .y(output_2_487));
wire output_4_487, output_4_8, output_3_487;
mixer gate_output_3_487(.a(output_4_487), .b(output_4_8), .y(output_3_487));
wire output_5_487, output_5_8, output_4_487;
mixer gate_output_4_487(.a(output_5_487), .b(output_5_8), .y(output_4_487));
wire output_6_487, output_6_8, output_5_487;
mixer gate_output_5_487(.a(output_6_487), .b(output_6_8), .y(output_5_487));
wire output_7_487, output_7_8, output_6_487;
mixer gate_output_6_487(.a(output_7_487), .b(output_7_8), .y(output_6_487));
wire output_8_487, output_8_8, output_7_487;
mixer gate_output_7_487(.a(output_8_487), .b(output_8_8), .y(output_7_487));
wire output_9_487, output_9_8, output_8_487;
mixer gate_output_8_487(.a(output_9_487), .b(output_9_8), .y(output_8_487));
wire output_10_487, output_10_8, output_9_487;
mixer gate_output_9_487(.a(output_10_487), .b(output_10_8), .y(output_9_487));
wire output_11_487, output_11_8, output_10_487;
mixer gate_output_10_487(.a(output_11_487), .b(output_11_8), .y(output_10_487));
wire output_12_487, output_12_8, output_11_487;
mixer gate_output_11_487(.a(output_12_487), .b(output_12_8), .y(output_11_487));
wire output_13_487, output_13_8, output_12_487;
mixer gate_output_12_487(.a(output_13_487), .b(output_13_8), .y(output_12_487));
wire output_14_487, output_14_8, output_13_487;
mixer gate_output_13_487(.a(output_14_487), .b(output_14_8), .y(output_13_487));
wire output_15_487, output_15_8, output_14_487;
mixer gate_output_14_487(.a(output_15_487), .b(output_15_8), .y(output_14_487));
wire output_16_487, output_16_8, output_15_487;
mixer gate_output_15_487(.a(output_16_487), .b(output_16_8), .y(output_15_487));
wire output_1_488, output_1_9, output_0_488;
mixer gate_output_0_488(.a(output_1_488), .b(output_1_9), .y(output_0_488));
wire output_2_488, output_2_9, output_1_488;
mixer gate_output_1_488(.a(output_2_488), .b(output_2_9), .y(output_1_488));
wire output_3_488, output_3_9, output_2_488;
mixer gate_output_2_488(.a(output_3_488), .b(output_3_9), .y(output_2_488));
wire output_4_488, output_4_9, output_3_488;
mixer gate_output_3_488(.a(output_4_488), .b(output_4_9), .y(output_3_488));
wire output_5_488, output_5_9, output_4_488;
mixer gate_output_4_488(.a(output_5_488), .b(output_5_9), .y(output_4_488));
wire output_6_488, output_6_9, output_5_488;
mixer gate_output_5_488(.a(output_6_488), .b(output_6_9), .y(output_5_488));
wire output_7_488, output_7_9, output_6_488;
mixer gate_output_6_488(.a(output_7_488), .b(output_7_9), .y(output_6_488));
wire output_8_488, output_8_9, output_7_488;
mixer gate_output_7_488(.a(output_8_488), .b(output_8_9), .y(output_7_488));
wire output_9_488, output_9_9, output_8_488;
mixer gate_output_8_488(.a(output_9_488), .b(output_9_9), .y(output_8_488));
wire output_10_488, output_10_9, output_9_488;
mixer gate_output_9_488(.a(output_10_488), .b(output_10_9), .y(output_9_488));
wire output_11_488, output_11_9, output_10_488;
mixer gate_output_10_488(.a(output_11_488), .b(output_11_9), .y(output_10_488));
wire output_12_488, output_12_9, output_11_488;
mixer gate_output_11_488(.a(output_12_488), .b(output_12_9), .y(output_11_488));
wire output_13_488, output_13_9, output_12_488;
mixer gate_output_12_488(.a(output_13_488), .b(output_13_9), .y(output_12_488));
wire output_14_488, output_14_9, output_13_488;
mixer gate_output_13_488(.a(output_14_488), .b(output_14_9), .y(output_13_488));
wire output_15_488, output_15_9, output_14_488;
mixer gate_output_14_488(.a(output_15_488), .b(output_15_9), .y(output_14_488));
wire output_16_488, output_16_9, output_15_488;
mixer gate_output_15_488(.a(output_16_488), .b(output_16_9), .y(output_15_488));
wire output_1_489, output_1_10, output_0_489;
mixer gate_output_0_489(.a(output_1_489), .b(output_1_10), .y(output_0_489));
wire output_2_489, output_2_10, output_1_489;
mixer gate_output_1_489(.a(output_2_489), .b(output_2_10), .y(output_1_489));
wire output_3_489, output_3_10, output_2_489;
mixer gate_output_2_489(.a(output_3_489), .b(output_3_10), .y(output_2_489));
wire output_4_489, output_4_10, output_3_489;
mixer gate_output_3_489(.a(output_4_489), .b(output_4_10), .y(output_3_489));
wire output_5_489, output_5_10, output_4_489;
mixer gate_output_4_489(.a(output_5_489), .b(output_5_10), .y(output_4_489));
wire output_6_489, output_6_10, output_5_489;
mixer gate_output_5_489(.a(output_6_489), .b(output_6_10), .y(output_5_489));
wire output_7_489, output_7_10, output_6_489;
mixer gate_output_6_489(.a(output_7_489), .b(output_7_10), .y(output_6_489));
wire output_8_489, output_8_10, output_7_489;
mixer gate_output_7_489(.a(output_8_489), .b(output_8_10), .y(output_7_489));
wire output_9_489, output_9_10, output_8_489;
mixer gate_output_8_489(.a(output_9_489), .b(output_9_10), .y(output_8_489));
wire output_10_489, output_10_10, output_9_489;
mixer gate_output_9_489(.a(output_10_489), .b(output_10_10), .y(output_9_489));
wire output_11_489, output_11_10, output_10_489;
mixer gate_output_10_489(.a(output_11_489), .b(output_11_10), .y(output_10_489));
wire output_12_489, output_12_10, output_11_489;
mixer gate_output_11_489(.a(output_12_489), .b(output_12_10), .y(output_11_489));
wire output_13_489, output_13_10, output_12_489;
mixer gate_output_12_489(.a(output_13_489), .b(output_13_10), .y(output_12_489));
wire output_14_489, output_14_10, output_13_489;
mixer gate_output_13_489(.a(output_14_489), .b(output_14_10), .y(output_13_489));
wire output_15_489, output_15_10, output_14_489;
mixer gate_output_14_489(.a(output_15_489), .b(output_15_10), .y(output_14_489));
wire output_16_489, output_16_10, output_15_489;
mixer gate_output_15_489(.a(output_16_489), .b(output_16_10), .y(output_15_489));
wire output_1_490, output_1_11, output_0_490;
mixer gate_output_0_490(.a(output_1_490), .b(output_1_11), .y(output_0_490));
wire output_2_490, output_2_11, output_1_490;
mixer gate_output_1_490(.a(output_2_490), .b(output_2_11), .y(output_1_490));
wire output_3_490, output_3_11, output_2_490;
mixer gate_output_2_490(.a(output_3_490), .b(output_3_11), .y(output_2_490));
wire output_4_490, output_4_11, output_3_490;
mixer gate_output_3_490(.a(output_4_490), .b(output_4_11), .y(output_3_490));
wire output_5_490, output_5_11, output_4_490;
mixer gate_output_4_490(.a(output_5_490), .b(output_5_11), .y(output_4_490));
wire output_6_490, output_6_11, output_5_490;
mixer gate_output_5_490(.a(output_6_490), .b(output_6_11), .y(output_5_490));
wire output_7_490, output_7_11, output_6_490;
mixer gate_output_6_490(.a(output_7_490), .b(output_7_11), .y(output_6_490));
wire output_8_490, output_8_11, output_7_490;
mixer gate_output_7_490(.a(output_8_490), .b(output_8_11), .y(output_7_490));
wire output_9_490, output_9_11, output_8_490;
mixer gate_output_8_490(.a(output_9_490), .b(output_9_11), .y(output_8_490));
wire output_10_490, output_10_11, output_9_490;
mixer gate_output_9_490(.a(output_10_490), .b(output_10_11), .y(output_9_490));
wire output_11_490, output_11_11, output_10_490;
mixer gate_output_10_490(.a(output_11_490), .b(output_11_11), .y(output_10_490));
wire output_12_490, output_12_11, output_11_490;
mixer gate_output_11_490(.a(output_12_490), .b(output_12_11), .y(output_11_490));
wire output_13_490, output_13_11, output_12_490;
mixer gate_output_12_490(.a(output_13_490), .b(output_13_11), .y(output_12_490));
wire output_14_490, output_14_11, output_13_490;
mixer gate_output_13_490(.a(output_14_490), .b(output_14_11), .y(output_13_490));
wire output_15_490, output_15_11, output_14_490;
mixer gate_output_14_490(.a(output_15_490), .b(output_15_11), .y(output_14_490));
wire output_16_490, output_16_11, output_15_490;
mixer gate_output_15_490(.a(output_16_490), .b(output_16_11), .y(output_15_490));
wire output_1_491, output_1_12, output_0_491;
mixer gate_output_0_491(.a(output_1_491), .b(output_1_12), .y(output_0_491));
wire output_2_491, output_2_12, output_1_491;
mixer gate_output_1_491(.a(output_2_491), .b(output_2_12), .y(output_1_491));
wire output_3_491, output_3_12, output_2_491;
mixer gate_output_2_491(.a(output_3_491), .b(output_3_12), .y(output_2_491));
wire output_4_491, output_4_12, output_3_491;
mixer gate_output_3_491(.a(output_4_491), .b(output_4_12), .y(output_3_491));
wire output_5_491, output_5_12, output_4_491;
mixer gate_output_4_491(.a(output_5_491), .b(output_5_12), .y(output_4_491));
wire output_6_491, output_6_12, output_5_491;
mixer gate_output_5_491(.a(output_6_491), .b(output_6_12), .y(output_5_491));
wire output_7_491, output_7_12, output_6_491;
mixer gate_output_6_491(.a(output_7_491), .b(output_7_12), .y(output_6_491));
wire output_8_491, output_8_12, output_7_491;
mixer gate_output_7_491(.a(output_8_491), .b(output_8_12), .y(output_7_491));
wire output_9_491, output_9_12, output_8_491;
mixer gate_output_8_491(.a(output_9_491), .b(output_9_12), .y(output_8_491));
wire output_10_491, output_10_12, output_9_491;
mixer gate_output_9_491(.a(output_10_491), .b(output_10_12), .y(output_9_491));
wire output_11_491, output_11_12, output_10_491;
mixer gate_output_10_491(.a(output_11_491), .b(output_11_12), .y(output_10_491));
wire output_12_491, output_12_12, output_11_491;
mixer gate_output_11_491(.a(output_12_491), .b(output_12_12), .y(output_11_491));
wire output_13_491, output_13_12, output_12_491;
mixer gate_output_12_491(.a(output_13_491), .b(output_13_12), .y(output_12_491));
wire output_14_491, output_14_12, output_13_491;
mixer gate_output_13_491(.a(output_14_491), .b(output_14_12), .y(output_13_491));
wire output_15_491, output_15_12, output_14_491;
mixer gate_output_14_491(.a(output_15_491), .b(output_15_12), .y(output_14_491));
wire output_16_491, output_16_12, output_15_491;
mixer gate_output_15_491(.a(output_16_491), .b(output_16_12), .y(output_15_491));
wire output_1_492, output_1_13, output_0_492;
mixer gate_output_0_492(.a(output_1_492), .b(output_1_13), .y(output_0_492));
wire output_2_492, output_2_13, output_1_492;
mixer gate_output_1_492(.a(output_2_492), .b(output_2_13), .y(output_1_492));
wire output_3_492, output_3_13, output_2_492;
mixer gate_output_2_492(.a(output_3_492), .b(output_3_13), .y(output_2_492));
wire output_4_492, output_4_13, output_3_492;
mixer gate_output_3_492(.a(output_4_492), .b(output_4_13), .y(output_3_492));
wire output_5_492, output_5_13, output_4_492;
mixer gate_output_4_492(.a(output_5_492), .b(output_5_13), .y(output_4_492));
wire output_6_492, output_6_13, output_5_492;
mixer gate_output_5_492(.a(output_6_492), .b(output_6_13), .y(output_5_492));
wire output_7_492, output_7_13, output_6_492;
mixer gate_output_6_492(.a(output_7_492), .b(output_7_13), .y(output_6_492));
wire output_8_492, output_8_13, output_7_492;
mixer gate_output_7_492(.a(output_8_492), .b(output_8_13), .y(output_7_492));
wire output_9_492, output_9_13, output_8_492;
mixer gate_output_8_492(.a(output_9_492), .b(output_9_13), .y(output_8_492));
wire output_10_492, output_10_13, output_9_492;
mixer gate_output_9_492(.a(output_10_492), .b(output_10_13), .y(output_9_492));
wire output_11_492, output_11_13, output_10_492;
mixer gate_output_10_492(.a(output_11_492), .b(output_11_13), .y(output_10_492));
wire output_12_492, output_12_13, output_11_492;
mixer gate_output_11_492(.a(output_12_492), .b(output_12_13), .y(output_11_492));
wire output_13_492, output_13_13, output_12_492;
mixer gate_output_12_492(.a(output_13_492), .b(output_13_13), .y(output_12_492));
wire output_14_492, output_14_13, output_13_492;
mixer gate_output_13_492(.a(output_14_492), .b(output_14_13), .y(output_13_492));
wire output_15_492, output_15_13, output_14_492;
mixer gate_output_14_492(.a(output_15_492), .b(output_15_13), .y(output_14_492));
wire output_16_492, output_16_13, output_15_492;
mixer gate_output_15_492(.a(output_16_492), .b(output_16_13), .y(output_15_492));
wire output_1_493, output_1_14, output_0_493;
mixer gate_output_0_493(.a(output_1_493), .b(output_1_14), .y(output_0_493));
wire output_2_493, output_2_14, output_1_493;
mixer gate_output_1_493(.a(output_2_493), .b(output_2_14), .y(output_1_493));
wire output_3_493, output_3_14, output_2_493;
mixer gate_output_2_493(.a(output_3_493), .b(output_3_14), .y(output_2_493));
wire output_4_493, output_4_14, output_3_493;
mixer gate_output_3_493(.a(output_4_493), .b(output_4_14), .y(output_3_493));
wire output_5_493, output_5_14, output_4_493;
mixer gate_output_4_493(.a(output_5_493), .b(output_5_14), .y(output_4_493));
wire output_6_493, output_6_14, output_5_493;
mixer gate_output_5_493(.a(output_6_493), .b(output_6_14), .y(output_5_493));
wire output_7_493, output_7_14, output_6_493;
mixer gate_output_6_493(.a(output_7_493), .b(output_7_14), .y(output_6_493));
wire output_8_493, output_8_14, output_7_493;
mixer gate_output_7_493(.a(output_8_493), .b(output_8_14), .y(output_7_493));
wire output_9_493, output_9_14, output_8_493;
mixer gate_output_8_493(.a(output_9_493), .b(output_9_14), .y(output_8_493));
wire output_10_493, output_10_14, output_9_493;
mixer gate_output_9_493(.a(output_10_493), .b(output_10_14), .y(output_9_493));
wire output_11_493, output_11_14, output_10_493;
mixer gate_output_10_493(.a(output_11_493), .b(output_11_14), .y(output_10_493));
wire output_12_493, output_12_14, output_11_493;
mixer gate_output_11_493(.a(output_12_493), .b(output_12_14), .y(output_11_493));
wire output_13_493, output_13_14, output_12_493;
mixer gate_output_12_493(.a(output_13_493), .b(output_13_14), .y(output_12_493));
wire output_14_493, output_14_14, output_13_493;
mixer gate_output_13_493(.a(output_14_493), .b(output_14_14), .y(output_13_493));
wire output_15_493, output_15_14, output_14_493;
mixer gate_output_14_493(.a(output_15_493), .b(output_15_14), .y(output_14_493));
wire output_16_493, output_16_14, output_15_493;
mixer gate_output_15_493(.a(output_16_493), .b(output_16_14), .y(output_15_493));
wire output_1_494, output_1_15, output_0_494;
mixer gate_output_0_494(.a(output_1_494), .b(output_1_15), .y(output_0_494));
wire output_2_494, output_2_15, output_1_494;
mixer gate_output_1_494(.a(output_2_494), .b(output_2_15), .y(output_1_494));
wire output_3_494, output_3_15, output_2_494;
mixer gate_output_2_494(.a(output_3_494), .b(output_3_15), .y(output_2_494));
wire output_4_494, output_4_15, output_3_494;
mixer gate_output_3_494(.a(output_4_494), .b(output_4_15), .y(output_3_494));
wire output_5_494, output_5_15, output_4_494;
mixer gate_output_4_494(.a(output_5_494), .b(output_5_15), .y(output_4_494));
wire output_6_494, output_6_15, output_5_494;
mixer gate_output_5_494(.a(output_6_494), .b(output_6_15), .y(output_5_494));
wire output_7_494, output_7_15, output_6_494;
mixer gate_output_6_494(.a(output_7_494), .b(output_7_15), .y(output_6_494));
wire output_8_494, output_8_15, output_7_494;
mixer gate_output_7_494(.a(output_8_494), .b(output_8_15), .y(output_7_494));
wire output_9_494, output_9_15, output_8_494;
mixer gate_output_8_494(.a(output_9_494), .b(output_9_15), .y(output_8_494));
wire output_10_494, output_10_15, output_9_494;
mixer gate_output_9_494(.a(output_10_494), .b(output_10_15), .y(output_9_494));
wire output_11_494, output_11_15, output_10_494;
mixer gate_output_10_494(.a(output_11_494), .b(output_11_15), .y(output_10_494));
wire output_12_494, output_12_15, output_11_494;
mixer gate_output_11_494(.a(output_12_494), .b(output_12_15), .y(output_11_494));
wire output_13_494, output_13_15, output_12_494;
mixer gate_output_12_494(.a(output_13_494), .b(output_13_15), .y(output_12_494));
wire output_14_494, output_14_15, output_13_494;
mixer gate_output_13_494(.a(output_14_494), .b(output_14_15), .y(output_13_494));
wire output_15_494, output_15_15, output_14_494;
mixer gate_output_14_494(.a(output_15_494), .b(output_15_15), .y(output_14_494));
wire output_16_494, output_16_15, output_15_494;
mixer gate_output_15_494(.a(output_16_494), .b(output_16_15), .y(output_15_494));
wire output_1_495, output_1_0, output_0_495;
mixer gate_output_0_495(.a(output_1_495), .b(output_1_0), .y(output_0_495));
wire output_2_495, output_2_0, output_1_495;
mixer gate_output_1_495(.a(output_2_495), .b(output_2_0), .y(output_1_495));
wire output_3_495, output_3_0, output_2_495;
mixer gate_output_2_495(.a(output_3_495), .b(output_3_0), .y(output_2_495));
wire output_4_495, output_4_0, output_3_495;
mixer gate_output_3_495(.a(output_4_495), .b(output_4_0), .y(output_3_495));
wire output_5_495, output_5_0, output_4_495;
mixer gate_output_4_495(.a(output_5_495), .b(output_5_0), .y(output_4_495));
wire output_6_495, output_6_0, output_5_495;
mixer gate_output_5_495(.a(output_6_495), .b(output_6_0), .y(output_5_495));
wire output_7_495, output_7_0, output_6_495;
mixer gate_output_6_495(.a(output_7_495), .b(output_7_0), .y(output_6_495));
wire output_8_495, output_8_0, output_7_495;
mixer gate_output_7_495(.a(output_8_495), .b(output_8_0), .y(output_7_495));
wire output_9_495, output_9_0, output_8_495;
mixer gate_output_8_495(.a(output_9_495), .b(output_9_0), .y(output_8_495));
wire output_10_495, output_10_0, output_9_495;
mixer gate_output_9_495(.a(output_10_495), .b(output_10_0), .y(output_9_495));
wire output_11_495, output_11_0, output_10_495;
mixer gate_output_10_495(.a(output_11_495), .b(output_11_0), .y(output_10_495));
wire output_12_495, output_12_0, output_11_495;
mixer gate_output_11_495(.a(output_12_495), .b(output_12_0), .y(output_11_495));
wire output_13_495, output_13_0, output_12_495;
mixer gate_output_12_495(.a(output_13_495), .b(output_13_0), .y(output_12_495));
wire output_14_495, output_14_0, output_13_495;
mixer gate_output_13_495(.a(output_14_495), .b(output_14_0), .y(output_13_495));
wire output_15_495, output_15_0, output_14_495;
mixer gate_output_14_495(.a(output_15_495), .b(output_15_0), .y(output_14_495));
wire output_16_495, output_16_0, output_15_495;
mixer gate_output_15_495(.a(output_16_495), .b(output_16_0), .y(output_15_495));
wire output_1_496, output_1_1, output_0_496;
mixer gate_output_0_496(.a(output_1_496), .b(output_1_1), .y(output_0_496));
wire output_2_496, output_2_1, output_1_496;
mixer gate_output_1_496(.a(output_2_496), .b(output_2_1), .y(output_1_496));
wire output_3_496, output_3_1, output_2_496;
mixer gate_output_2_496(.a(output_3_496), .b(output_3_1), .y(output_2_496));
wire output_4_496, output_4_1, output_3_496;
mixer gate_output_3_496(.a(output_4_496), .b(output_4_1), .y(output_3_496));
wire output_5_496, output_5_1, output_4_496;
mixer gate_output_4_496(.a(output_5_496), .b(output_5_1), .y(output_4_496));
wire output_6_496, output_6_1, output_5_496;
mixer gate_output_5_496(.a(output_6_496), .b(output_6_1), .y(output_5_496));
wire output_7_496, output_7_1, output_6_496;
mixer gate_output_6_496(.a(output_7_496), .b(output_7_1), .y(output_6_496));
wire output_8_496, output_8_1, output_7_496;
mixer gate_output_7_496(.a(output_8_496), .b(output_8_1), .y(output_7_496));
wire output_9_496, output_9_1, output_8_496;
mixer gate_output_8_496(.a(output_9_496), .b(output_9_1), .y(output_8_496));
wire output_10_496, output_10_1, output_9_496;
mixer gate_output_9_496(.a(output_10_496), .b(output_10_1), .y(output_9_496));
wire output_11_496, output_11_1, output_10_496;
mixer gate_output_10_496(.a(output_11_496), .b(output_11_1), .y(output_10_496));
wire output_12_496, output_12_1, output_11_496;
mixer gate_output_11_496(.a(output_12_496), .b(output_12_1), .y(output_11_496));
wire output_13_496, output_13_1, output_12_496;
mixer gate_output_12_496(.a(output_13_496), .b(output_13_1), .y(output_12_496));
wire output_14_496, output_14_1, output_13_496;
mixer gate_output_13_496(.a(output_14_496), .b(output_14_1), .y(output_13_496));
wire output_15_496, output_15_1, output_14_496;
mixer gate_output_14_496(.a(output_15_496), .b(output_15_1), .y(output_14_496));
wire output_16_496, output_16_1, output_15_496;
mixer gate_output_15_496(.a(output_16_496), .b(output_16_1), .y(output_15_496));
wire output_1_497, output_1_2, output_0_497;
mixer gate_output_0_497(.a(output_1_497), .b(output_1_2), .y(output_0_497));
wire output_2_497, output_2_2, output_1_497;
mixer gate_output_1_497(.a(output_2_497), .b(output_2_2), .y(output_1_497));
wire output_3_497, output_3_2, output_2_497;
mixer gate_output_2_497(.a(output_3_497), .b(output_3_2), .y(output_2_497));
wire output_4_497, output_4_2, output_3_497;
mixer gate_output_3_497(.a(output_4_497), .b(output_4_2), .y(output_3_497));
wire output_5_497, output_5_2, output_4_497;
mixer gate_output_4_497(.a(output_5_497), .b(output_5_2), .y(output_4_497));
wire output_6_497, output_6_2, output_5_497;
mixer gate_output_5_497(.a(output_6_497), .b(output_6_2), .y(output_5_497));
wire output_7_497, output_7_2, output_6_497;
mixer gate_output_6_497(.a(output_7_497), .b(output_7_2), .y(output_6_497));
wire output_8_497, output_8_2, output_7_497;
mixer gate_output_7_497(.a(output_8_497), .b(output_8_2), .y(output_7_497));
wire output_9_497, output_9_2, output_8_497;
mixer gate_output_8_497(.a(output_9_497), .b(output_9_2), .y(output_8_497));
wire output_10_497, output_10_2, output_9_497;
mixer gate_output_9_497(.a(output_10_497), .b(output_10_2), .y(output_9_497));
wire output_11_497, output_11_2, output_10_497;
mixer gate_output_10_497(.a(output_11_497), .b(output_11_2), .y(output_10_497));
wire output_12_497, output_12_2, output_11_497;
mixer gate_output_11_497(.a(output_12_497), .b(output_12_2), .y(output_11_497));
wire output_13_497, output_13_2, output_12_497;
mixer gate_output_12_497(.a(output_13_497), .b(output_13_2), .y(output_12_497));
wire output_14_497, output_14_2, output_13_497;
mixer gate_output_13_497(.a(output_14_497), .b(output_14_2), .y(output_13_497));
wire output_15_497, output_15_2, output_14_497;
mixer gate_output_14_497(.a(output_15_497), .b(output_15_2), .y(output_14_497));
wire output_16_497, output_16_2, output_15_497;
mixer gate_output_15_497(.a(output_16_497), .b(output_16_2), .y(output_15_497));
wire output_1_498, output_1_3, output_0_498;
mixer gate_output_0_498(.a(output_1_498), .b(output_1_3), .y(output_0_498));
wire output_2_498, output_2_3, output_1_498;
mixer gate_output_1_498(.a(output_2_498), .b(output_2_3), .y(output_1_498));
wire output_3_498, output_3_3, output_2_498;
mixer gate_output_2_498(.a(output_3_498), .b(output_3_3), .y(output_2_498));
wire output_4_498, output_4_3, output_3_498;
mixer gate_output_3_498(.a(output_4_498), .b(output_4_3), .y(output_3_498));
wire output_5_498, output_5_3, output_4_498;
mixer gate_output_4_498(.a(output_5_498), .b(output_5_3), .y(output_4_498));
wire output_6_498, output_6_3, output_5_498;
mixer gate_output_5_498(.a(output_6_498), .b(output_6_3), .y(output_5_498));
wire output_7_498, output_7_3, output_6_498;
mixer gate_output_6_498(.a(output_7_498), .b(output_7_3), .y(output_6_498));
wire output_8_498, output_8_3, output_7_498;
mixer gate_output_7_498(.a(output_8_498), .b(output_8_3), .y(output_7_498));
wire output_9_498, output_9_3, output_8_498;
mixer gate_output_8_498(.a(output_9_498), .b(output_9_3), .y(output_8_498));
wire output_10_498, output_10_3, output_9_498;
mixer gate_output_9_498(.a(output_10_498), .b(output_10_3), .y(output_9_498));
wire output_11_498, output_11_3, output_10_498;
mixer gate_output_10_498(.a(output_11_498), .b(output_11_3), .y(output_10_498));
wire output_12_498, output_12_3, output_11_498;
mixer gate_output_11_498(.a(output_12_498), .b(output_12_3), .y(output_11_498));
wire output_13_498, output_13_3, output_12_498;
mixer gate_output_12_498(.a(output_13_498), .b(output_13_3), .y(output_12_498));
wire output_14_498, output_14_3, output_13_498;
mixer gate_output_13_498(.a(output_14_498), .b(output_14_3), .y(output_13_498));
wire output_15_498, output_15_3, output_14_498;
mixer gate_output_14_498(.a(output_15_498), .b(output_15_3), .y(output_14_498));
wire output_16_498, output_16_3, output_15_498;
mixer gate_output_15_498(.a(output_16_498), .b(output_16_3), .y(output_15_498));
wire output_1_499, output_1_4, output_0_499;
mixer gate_output_0_499(.a(output_1_499), .b(output_1_4), .y(output_0_499));
wire output_2_499, output_2_4, output_1_499;
mixer gate_output_1_499(.a(output_2_499), .b(output_2_4), .y(output_1_499));
wire output_3_499, output_3_4, output_2_499;
mixer gate_output_2_499(.a(output_3_499), .b(output_3_4), .y(output_2_499));
wire output_4_499, output_4_4, output_3_499;
mixer gate_output_3_499(.a(output_4_499), .b(output_4_4), .y(output_3_499));
wire output_5_499, output_5_4, output_4_499;
mixer gate_output_4_499(.a(output_5_499), .b(output_5_4), .y(output_4_499));
wire output_6_499, output_6_4, output_5_499;
mixer gate_output_5_499(.a(output_6_499), .b(output_6_4), .y(output_5_499));
wire output_7_499, output_7_4, output_6_499;
mixer gate_output_6_499(.a(output_7_499), .b(output_7_4), .y(output_6_499));
wire output_8_499, output_8_4, output_7_499;
mixer gate_output_7_499(.a(output_8_499), .b(output_8_4), .y(output_7_499));
wire output_9_499, output_9_4, output_8_499;
mixer gate_output_8_499(.a(output_9_499), .b(output_9_4), .y(output_8_499));
wire output_10_499, output_10_4, output_9_499;
mixer gate_output_9_499(.a(output_10_499), .b(output_10_4), .y(output_9_499));
wire output_11_499, output_11_4, output_10_499;
mixer gate_output_10_499(.a(output_11_499), .b(output_11_4), .y(output_10_499));
wire output_12_499, output_12_4, output_11_499;
mixer gate_output_11_499(.a(output_12_499), .b(output_12_4), .y(output_11_499));
wire output_13_499, output_13_4, output_12_499;
mixer gate_output_12_499(.a(output_13_499), .b(output_13_4), .y(output_12_499));
wire output_14_499, output_14_4, output_13_499;
mixer gate_output_13_499(.a(output_14_499), .b(output_14_4), .y(output_13_499));
wire output_15_499, output_15_4, output_14_499;
mixer gate_output_14_499(.a(output_15_499), .b(output_15_4), .y(output_14_499));
wire output_16_499, output_16_4, output_15_499;
mixer gate_output_15_499(.a(output_16_499), .b(output_16_4), .y(output_15_499));
wire output_1_500, output_1_5, output_0_500;
mixer gate_output_0_500(.a(output_1_500), .b(output_1_5), .y(output_0_500));
wire output_2_500, output_2_5, output_1_500;
mixer gate_output_1_500(.a(output_2_500), .b(output_2_5), .y(output_1_500));
wire output_3_500, output_3_5, output_2_500;
mixer gate_output_2_500(.a(output_3_500), .b(output_3_5), .y(output_2_500));
wire output_4_500, output_4_5, output_3_500;
mixer gate_output_3_500(.a(output_4_500), .b(output_4_5), .y(output_3_500));
wire output_5_500, output_5_5, output_4_500;
mixer gate_output_4_500(.a(output_5_500), .b(output_5_5), .y(output_4_500));
wire output_6_500, output_6_5, output_5_500;
mixer gate_output_5_500(.a(output_6_500), .b(output_6_5), .y(output_5_500));
wire output_7_500, output_7_5, output_6_500;
mixer gate_output_6_500(.a(output_7_500), .b(output_7_5), .y(output_6_500));
wire output_8_500, output_8_5, output_7_500;
mixer gate_output_7_500(.a(output_8_500), .b(output_8_5), .y(output_7_500));
wire output_9_500, output_9_5, output_8_500;
mixer gate_output_8_500(.a(output_9_500), .b(output_9_5), .y(output_8_500));
wire output_10_500, output_10_5, output_9_500;
mixer gate_output_9_500(.a(output_10_500), .b(output_10_5), .y(output_9_500));
wire output_11_500, output_11_5, output_10_500;
mixer gate_output_10_500(.a(output_11_500), .b(output_11_5), .y(output_10_500));
wire output_12_500, output_12_5, output_11_500;
mixer gate_output_11_500(.a(output_12_500), .b(output_12_5), .y(output_11_500));
wire output_13_500, output_13_5, output_12_500;
mixer gate_output_12_500(.a(output_13_500), .b(output_13_5), .y(output_12_500));
wire output_14_500, output_14_5, output_13_500;
mixer gate_output_13_500(.a(output_14_500), .b(output_14_5), .y(output_13_500));
wire output_15_500, output_15_5, output_14_500;
mixer gate_output_14_500(.a(output_15_500), .b(output_15_5), .y(output_14_500));
wire output_16_500, output_16_5, output_15_500;
mixer gate_output_15_500(.a(output_16_500), .b(output_16_5), .y(output_15_500));
wire output_1_501, output_1_6, output_0_501;
mixer gate_output_0_501(.a(output_1_501), .b(output_1_6), .y(output_0_501));
wire output_2_501, output_2_6, output_1_501;
mixer gate_output_1_501(.a(output_2_501), .b(output_2_6), .y(output_1_501));
wire output_3_501, output_3_6, output_2_501;
mixer gate_output_2_501(.a(output_3_501), .b(output_3_6), .y(output_2_501));
wire output_4_501, output_4_6, output_3_501;
mixer gate_output_3_501(.a(output_4_501), .b(output_4_6), .y(output_3_501));
wire output_5_501, output_5_6, output_4_501;
mixer gate_output_4_501(.a(output_5_501), .b(output_5_6), .y(output_4_501));
wire output_6_501, output_6_6, output_5_501;
mixer gate_output_5_501(.a(output_6_501), .b(output_6_6), .y(output_5_501));
wire output_7_501, output_7_6, output_6_501;
mixer gate_output_6_501(.a(output_7_501), .b(output_7_6), .y(output_6_501));
wire output_8_501, output_8_6, output_7_501;
mixer gate_output_7_501(.a(output_8_501), .b(output_8_6), .y(output_7_501));
wire output_9_501, output_9_6, output_8_501;
mixer gate_output_8_501(.a(output_9_501), .b(output_9_6), .y(output_8_501));
wire output_10_501, output_10_6, output_9_501;
mixer gate_output_9_501(.a(output_10_501), .b(output_10_6), .y(output_9_501));
wire output_11_501, output_11_6, output_10_501;
mixer gate_output_10_501(.a(output_11_501), .b(output_11_6), .y(output_10_501));
wire output_12_501, output_12_6, output_11_501;
mixer gate_output_11_501(.a(output_12_501), .b(output_12_6), .y(output_11_501));
wire output_13_501, output_13_6, output_12_501;
mixer gate_output_12_501(.a(output_13_501), .b(output_13_6), .y(output_12_501));
wire output_14_501, output_14_6, output_13_501;
mixer gate_output_13_501(.a(output_14_501), .b(output_14_6), .y(output_13_501));
wire output_15_501, output_15_6, output_14_501;
mixer gate_output_14_501(.a(output_15_501), .b(output_15_6), .y(output_14_501));
wire output_16_501, output_16_6, output_15_501;
mixer gate_output_15_501(.a(output_16_501), .b(output_16_6), .y(output_15_501));
wire output_1_502, output_1_7, output_0_502;
mixer gate_output_0_502(.a(output_1_502), .b(output_1_7), .y(output_0_502));
wire output_2_502, output_2_7, output_1_502;
mixer gate_output_1_502(.a(output_2_502), .b(output_2_7), .y(output_1_502));
wire output_3_502, output_3_7, output_2_502;
mixer gate_output_2_502(.a(output_3_502), .b(output_3_7), .y(output_2_502));
wire output_4_502, output_4_7, output_3_502;
mixer gate_output_3_502(.a(output_4_502), .b(output_4_7), .y(output_3_502));
wire output_5_502, output_5_7, output_4_502;
mixer gate_output_4_502(.a(output_5_502), .b(output_5_7), .y(output_4_502));
wire output_6_502, output_6_7, output_5_502;
mixer gate_output_5_502(.a(output_6_502), .b(output_6_7), .y(output_5_502));
wire output_7_502, output_7_7, output_6_502;
mixer gate_output_6_502(.a(output_7_502), .b(output_7_7), .y(output_6_502));
wire output_8_502, output_8_7, output_7_502;
mixer gate_output_7_502(.a(output_8_502), .b(output_8_7), .y(output_7_502));
wire output_9_502, output_9_7, output_8_502;
mixer gate_output_8_502(.a(output_9_502), .b(output_9_7), .y(output_8_502));
wire output_10_502, output_10_7, output_9_502;
mixer gate_output_9_502(.a(output_10_502), .b(output_10_7), .y(output_9_502));
wire output_11_502, output_11_7, output_10_502;
mixer gate_output_10_502(.a(output_11_502), .b(output_11_7), .y(output_10_502));
wire output_12_502, output_12_7, output_11_502;
mixer gate_output_11_502(.a(output_12_502), .b(output_12_7), .y(output_11_502));
wire output_13_502, output_13_7, output_12_502;
mixer gate_output_12_502(.a(output_13_502), .b(output_13_7), .y(output_12_502));
wire output_14_502, output_14_7, output_13_502;
mixer gate_output_13_502(.a(output_14_502), .b(output_14_7), .y(output_13_502));
wire output_15_502, output_15_7, output_14_502;
mixer gate_output_14_502(.a(output_15_502), .b(output_15_7), .y(output_14_502));
wire output_16_502, output_16_7, output_15_502;
mixer gate_output_15_502(.a(output_16_502), .b(output_16_7), .y(output_15_502));
wire output_1_503, output_1_8, output_0_503;
mixer gate_output_0_503(.a(output_1_503), .b(output_1_8), .y(output_0_503));
wire output_2_503, output_2_8, output_1_503;
mixer gate_output_1_503(.a(output_2_503), .b(output_2_8), .y(output_1_503));
wire output_3_503, output_3_8, output_2_503;
mixer gate_output_2_503(.a(output_3_503), .b(output_3_8), .y(output_2_503));
wire output_4_503, output_4_8, output_3_503;
mixer gate_output_3_503(.a(output_4_503), .b(output_4_8), .y(output_3_503));
wire output_5_503, output_5_8, output_4_503;
mixer gate_output_4_503(.a(output_5_503), .b(output_5_8), .y(output_4_503));
wire output_6_503, output_6_8, output_5_503;
mixer gate_output_5_503(.a(output_6_503), .b(output_6_8), .y(output_5_503));
wire output_7_503, output_7_8, output_6_503;
mixer gate_output_6_503(.a(output_7_503), .b(output_7_8), .y(output_6_503));
wire output_8_503, output_8_8, output_7_503;
mixer gate_output_7_503(.a(output_8_503), .b(output_8_8), .y(output_7_503));
wire output_9_503, output_9_8, output_8_503;
mixer gate_output_8_503(.a(output_9_503), .b(output_9_8), .y(output_8_503));
wire output_10_503, output_10_8, output_9_503;
mixer gate_output_9_503(.a(output_10_503), .b(output_10_8), .y(output_9_503));
wire output_11_503, output_11_8, output_10_503;
mixer gate_output_10_503(.a(output_11_503), .b(output_11_8), .y(output_10_503));
wire output_12_503, output_12_8, output_11_503;
mixer gate_output_11_503(.a(output_12_503), .b(output_12_8), .y(output_11_503));
wire output_13_503, output_13_8, output_12_503;
mixer gate_output_12_503(.a(output_13_503), .b(output_13_8), .y(output_12_503));
wire output_14_503, output_14_8, output_13_503;
mixer gate_output_13_503(.a(output_14_503), .b(output_14_8), .y(output_13_503));
wire output_15_503, output_15_8, output_14_503;
mixer gate_output_14_503(.a(output_15_503), .b(output_15_8), .y(output_14_503));
wire output_16_503, output_16_8, output_15_503;
mixer gate_output_15_503(.a(output_16_503), .b(output_16_8), .y(output_15_503));
wire output_1_504, output_1_9, output_0_504;
mixer gate_output_0_504(.a(output_1_504), .b(output_1_9), .y(output_0_504));
wire output_2_504, output_2_9, output_1_504;
mixer gate_output_1_504(.a(output_2_504), .b(output_2_9), .y(output_1_504));
wire output_3_504, output_3_9, output_2_504;
mixer gate_output_2_504(.a(output_3_504), .b(output_3_9), .y(output_2_504));
wire output_4_504, output_4_9, output_3_504;
mixer gate_output_3_504(.a(output_4_504), .b(output_4_9), .y(output_3_504));
wire output_5_504, output_5_9, output_4_504;
mixer gate_output_4_504(.a(output_5_504), .b(output_5_9), .y(output_4_504));
wire output_6_504, output_6_9, output_5_504;
mixer gate_output_5_504(.a(output_6_504), .b(output_6_9), .y(output_5_504));
wire output_7_504, output_7_9, output_6_504;
mixer gate_output_6_504(.a(output_7_504), .b(output_7_9), .y(output_6_504));
wire output_8_504, output_8_9, output_7_504;
mixer gate_output_7_504(.a(output_8_504), .b(output_8_9), .y(output_7_504));
wire output_9_504, output_9_9, output_8_504;
mixer gate_output_8_504(.a(output_9_504), .b(output_9_9), .y(output_8_504));
wire output_10_504, output_10_9, output_9_504;
mixer gate_output_9_504(.a(output_10_504), .b(output_10_9), .y(output_9_504));
wire output_11_504, output_11_9, output_10_504;
mixer gate_output_10_504(.a(output_11_504), .b(output_11_9), .y(output_10_504));
wire output_12_504, output_12_9, output_11_504;
mixer gate_output_11_504(.a(output_12_504), .b(output_12_9), .y(output_11_504));
wire output_13_504, output_13_9, output_12_504;
mixer gate_output_12_504(.a(output_13_504), .b(output_13_9), .y(output_12_504));
wire output_14_504, output_14_9, output_13_504;
mixer gate_output_13_504(.a(output_14_504), .b(output_14_9), .y(output_13_504));
wire output_15_504, output_15_9, output_14_504;
mixer gate_output_14_504(.a(output_15_504), .b(output_15_9), .y(output_14_504));
wire output_16_504, output_16_9, output_15_504;
mixer gate_output_15_504(.a(output_16_504), .b(output_16_9), .y(output_15_504));
wire output_1_505, output_1_10, output_0_505;
mixer gate_output_0_505(.a(output_1_505), .b(output_1_10), .y(output_0_505));
wire output_2_505, output_2_10, output_1_505;
mixer gate_output_1_505(.a(output_2_505), .b(output_2_10), .y(output_1_505));
wire output_3_505, output_3_10, output_2_505;
mixer gate_output_2_505(.a(output_3_505), .b(output_3_10), .y(output_2_505));
wire output_4_505, output_4_10, output_3_505;
mixer gate_output_3_505(.a(output_4_505), .b(output_4_10), .y(output_3_505));
wire output_5_505, output_5_10, output_4_505;
mixer gate_output_4_505(.a(output_5_505), .b(output_5_10), .y(output_4_505));
wire output_6_505, output_6_10, output_5_505;
mixer gate_output_5_505(.a(output_6_505), .b(output_6_10), .y(output_5_505));
wire output_7_505, output_7_10, output_6_505;
mixer gate_output_6_505(.a(output_7_505), .b(output_7_10), .y(output_6_505));
wire output_8_505, output_8_10, output_7_505;
mixer gate_output_7_505(.a(output_8_505), .b(output_8_10), .y(output_7_505));
wire output_9_505, output_9_10, output_8_505;
mixer gate_output_8_505(.a(output_9_505), .b(output_9_10), .y(output_8_505));
wire output_10_505, output_10_10, output_9_505;
mixer gate_output_9_505(.a(output_10_505), .b(output_10_10), .y(output_9_505));
wire output_11_505, output_11_10, output_10_505;
mixer gate_output_10_505(.a(output_11_505), .b(output_11_10), .y(output_10_505));
wire output_12_505, output_12_10, output_11_505;
mixer gate_output_11_505(.a(output_12_505), .b(output_12_10), .y(output_11_505));
wire output_13_505, output_13_10, output_12_505;
mixer gate_output_12_505(.a(output_13_505), .b(output_13_10), .y(output_12_505));
wire output_14_505, output_14_10, output_13_505;
mixer gate_output_13_505(.a(output_14_505), .b(output_14_10), .y(output_13_505));
wire output_15_505, output_15_10, output_14_505;
mixer gate_output_14_505(.a(output_15_505), .b(output_15_10), .y(output_14_505));
wire output_16_505, output_16_10, output_15_505;
mixer gate_output_15_505(.a(output_16_505), .b(output_16_10), .y(output_15_505));
wire output_1_506, output_1_11, output_0_506;
mixer gate_output_0_506(.a(output_1_506), .b(output_1_11), .y(output_0_506));
wire output_2_506, output_2_11, output_1_506;
mixer gate_output_1_506(.a(output_2_506), .b(output_2_11), .y(output_1_506));
wire output_3_506, output_3_11, output_2_506;
mixer gate_output_2_506(.a(output_3_506), .b(output_3_11), .y(output_2_506));
wire output_4_506, output_4_11, output_3_506;
mixer gate_output_3_506(.a(output_4_506), .b(output_4_11), .y(output_3_506));
wire output_5_506, output_5_11, output_4_506;
mixer gate_output_4_506(.a(output_5_506), .b(output_5_11), .y(output_4_506));
wire output_6_506, output_6_11, output_5_506;
mixer gate_output_5_506(.a(output_6_506), .b(output_6_11), .y(output_5_506));
wire output_7_506, output_7_11, output_6_506;
mixer gate_output_6_506(.a(output_7_506), .b(output_7_11), .y(output_6_506));
wire output_8_506, output_8_11, output_7_506;
mixer gate_output_7_506(.a(output_8_506), .b(output_8_11), .y(output_7_506));
wire output_9_506, output_9_11, output_8_506;
mixer gate_output_8_506(.a(output_9_506), .b(output_9_11), .y(output_8_506));
wire output_10_506, output_10_11, output_9_506;
mixer gate_output_9_506(.a(output_10_506), .b(output_10_11), .y(output_9_506));
wire output_11_506, output_11_11, output_10_506;
mixer gate_output_10_506(.a(output_11_506), .b(output_11_11), .y(output_10_506));
wire output_12_506, output_12_11, output_11_506;
mixer gate_output_11_506(.a(output_12_506), .b(output_12_11), .y(output_11_506));
wire output_13_506, output_13_11, output_12_506;
mixer gate_output_12_506(.a(output_13_506), .b(output_13_11), .y(output_12_506));
wire output_14_506, output_14_11, output_13_506;
mixer gate_output_13_506(.a(output_14_506), .b(output_14_11), .y(output_13_506));
wire output_15_506, output_15_11, output_14_506;
mixer gate_output_14_506(.a(output_15_506), .b(output_15_11), .y(output_14_506));
wire output_16_506, output_16_11, output_15_506;
mixer gate_output_15_506(.a(output_16_506), .b(output_16_11), .y(output_15_506));
wire output_1_507, output_1_12, output_0_507;
mixer gate_output_0_507(.a(output_1_507), .b(output_1_12), .y(output_0_507));
wire output_2_507, output_2_12, output_1_507;
mixer gate_output_1_507(.a(output_2_507), .b(output_2_12), .y(output_1_507));
wire output_3_507, output_3_12, output_2_507;
mixer gate_output_2_507(.a(output_3_507), .b(output_3_12), .y(output_2_507));
wire output_4_507, output_4_12, output_3_507;
mixer gate_output_3_507(.a(output_4_507), .b(output_4_12), .y(output_3_507));
wire output_5_507, output_5_12, output_4_507;
mixer gate_output_4_507(.a(output_5_507), .b(output_5_12), .y(output_4_507));
wire output_6_507, output_6_12, output_5_507;
mixer gate_output_5_507(.a(output_6_507), .b(output_6_12), .y(output_5_507));
wire output_7_507, output_7_12, output_6_507;
mixer gate_output_6_507(.a(output_7_507), .b(output_7_12), .y(output_6_507));
wire output_8_507, output_8_12, output_7_507;
mixer gate_output_7_507(.a(output_8_507), .b(output_8_12), .y(output_7_507));
wire output_9_507, output_9_12, output_8_507;
mixer gate_output_8_507(.a(output_9_507), .b(output_9_12), .y(output_8_507));
wire output_10_507, output_10_12, output_9_507;
mixer gate_output_9_507(.a(output_10_507), .b(output_10_12), .y(output_9_507));
wire output_11_507, output_11_12, output_10_507;
mixer gate_output_10_507(.a(output_11_507), .b(output_11_12), .y(output_10_507));
wire output_12_507, output_12_12, output_11_507;
mixer gate_output_11_507(.a(output_12_507), .b(output_12_12), .y(output_11_507));
wire output_13_507, output_13_12, output_12_507;
mixer gate_output_12_507(.a(output_13_507), .b(output_13_12), .y(output_12_507));
wire output_14_507, output_14_12, output_13_507;
mixer gate_output_13_507(.a(output_14_507), .b(output_14_12), .y(output_13_507));
wire output_15_507, output_15_12, output_14_507;
mixer gate_output_14_507(.a(output_15_507), .b(output_15_12), .y(output_14_507));
wire output_16_507, output_16_12, output_15_507;
mixer gate_output_15_507(.a(output_16_507), .b(output_16_12), .y(output_15_507));
wire output_1_508, output_1_13, output_0_508;
mixer gate_output_0_508(.a(output_1_508), .b(output_1_13), .y(output_0_508));
wire output_2_508, output_2_13, output_1_508;
mixer gate_output_1_508(.a(output_2_508), .b(output_2_13), .y(output_1_508));
wire output_3_508, output_3_13, output_2_508;
mixer gate_output_2_508(.a(output_3_508), .b(output_3_13), .y(output_2_508));
wire output_4_508, output_4_13, output_3_508;
mixer gate_output_3_508(.a(output_4_508), .b(output_4_13), .y(output_3_508));
wire output_5_508, output_5_13, output_4_508;
mixer gate_output_4_508(.a(output_5_508), .b(output_5_13), .y(output_4_508));
wire output_6_508, output_6_13, output_5_508;
mixer gate_output_5_508(.a(output_6_508), .b(output_6_13), .y(output_5_508));
wire output_7_508, output_7_13, output_6_508;
mixer gate_output_6_508(.a(output_7_508), .b(output_7_13), .y(output_6_508));
wire output_8_508, output_8_13, output_7_508;
mixer gate_output_7_508(.a(output_8_508), .b(output_8_13), .y(output_7_508));
wire output_9_508, output_9_13, output_8_508;
mixer gate_output_8_508(.a(output_9_508), .b(output_9_13), .y(output_8_508));
wire output_10_508, output_10_13, output_9_508;
mixer gate_output_9_508(.a(output_10_508), .b(output_10_13), .y(output_9_508));
wire output_11_508, output_11_13, output_10_508;
mixer gate_output_10_508(.a(output_11_508), .b(output_11_13), .y(output_10_508));
wire output_12_508, output_12_13, output_11_508;
mixer gate_output_11_508(.a(output_12_508), .b(output_12_13), .y(output_11_508));
wire output_13_508, output_13_13, output_12_508;
mixer gate_output_12_508(.a(output_13_508), .b(output_13_13), .y(output_12_508));
wire output_14_508, output_14_13, output_13_508;
mixer gate_output_13_508(.a(output_14_508), .b(output_14_13), .y(output_13_508));
wire output_15_508, output_15_13, output_14_508;
mixer gate_output_14_508(.a(output_15_508), .b(output_15_13), .y(output_14_508));
wire output_16_508, output_16_13, output_15_508;
mixer gate_output_15_508(.a(output_16_508), .b(output_16_13), .y(output_15_508));
wire output_1_509, output_1_14, output_0_509;
mixer gate_output_0_509(.a(output_1_509), .b(output_1_14), .y(output_0_509));
wire output_2_509, output_2_14, output_1_509;
mixer gate_output_1_509(.a(output_2_509), .b(output_2_14), .y(output_1_509));
wire output_3_509, output_3_14, output_2_509;
mixer gate_output_2_509(.a(output_3_509), .b(output_3_14), .y(output_2_509));
wire output_4_509, output_4_14, output_3_509;
mixer gate_output_3_509(.a(output_4_509), .b(output_4_14), .y(output_3_509));
wire output_5_509, output_5_14, output_4_509;
mixer gate_output_4_509(.a(output_5_509), .b(output_5_14), .y(output_4_509));
wire output_6_509, output_6_14, output_5_509;
mixer gate_output_5_509(.a(output_6_509), .b(output_6_14), .y(output_5_509));
wire output_7_509, output_7_14, output_6_509;
mixer gate_output_6_509(.a(output_7_509), .b(output_7_14), .y(output_6_509));
wire output_8_509, output_8_14, output_7_509;
mixer gate_output_7_509(.a(output_8_509), .b(output_8_14), .y(output_7_509));
wire output_9_509, output_9_14, output_8_509;
mixer gate_output_8_509(.a(output_9_509), .b(output_9_14), .y(output_8_509));
wire output_10_509, output_10_14, output_9_509;
mixer gate_output_9_509(.a(output_10_509), .b(output_10_14), .y(output_9_509));
wire output_11_509, output_11_14, output_10_509;
mixer gate_output_10_509(.a(output_11_509), .b(output_11_14), .y(output_10_509));
wire output_12_509, output_12_14, output_11_509;
mixer gate_output_11_509(.a(output_12_509), .b(output_12_14), .y(output_11_509));
wire output_13_509, output_13_14, output_12_509;
mixer gate_output_12_509(.a(output_13_509), .b(output_13_14), .y(output_12_509));
wire output_14_509, output_14_14, output_13_509;
mixer gate_output_13_509(.a(output_14_509), .b(output_14_14), .y(output_13_509));
wire output_15_509, output_15_14, output_14_509;
mixer gate_output_14_509(.a(output_15_509), .b(output_15_14), .y(output_14_509));
wire output_16_509, output_16_14, output_15_509;
mixer gate_output_15_509(.a(output_16_509), .b(output_16_14), .y(output_15_509));
wire output_1_510, output_1_15, output_0_510;
mixer gate_output_0_510(.a(output_1_510), .b(output_1_15), .y(output_0_510));
wire output_2_510, output_2_15, output_1_510;
mixer gate_output_1_510(.a(output_2_510), .b(output_2_15), .y(output_1_510));
wire output_3_510, output_3_15, output_2_510;
mixer gate_output_2_510(.a(output_3_510), .b(output_3_15), .y(output_2_510));
wire output_4_510, output_4_15, output_3_510;
mixer gate_output_3_510(.a(output_4_510), .b(output_4_15), .y(output_3_510));
wire output_5_510, output_5_15, output_4_510;
mixer gate_output_4_510(.a(output_5_510), .b(output_5_15), .y(output_4_510));
wire output_6_510, output_6_15, output_5_510;
mixer gate_output_5_510(.a(output_6_510), .b(output_6_15), .y(output_5_510));
wire output_7_510, output_7_15, output_6_510;
mixer gate_output_6_510(.a(output_7_510), .b(output_7_15), .y(output_6_510));
wire output_8_510, output_8_15, output_7_510;
mixer gate_output_7_510(.a(output_8_510), .b(output_8_15), .y(output_7_510));
wire output_9_510, output_9_15, output_8_510;
mixer gate_output_8_510(.a(output_9_510), .b(output_9_15), .y(output_8_510));
wire output_10_510, output_10_15, output_9_510;
mixer gate_output_9_510(.a(output_10_510), .b(output_10_15), .y(output_9_510));
wire output_11_510, output_11_15, output_10_510;
mixer gate_output_10_510(.a(output_11_510), .b(output_11_15), .y(output_10_510));
wire output_12_510, output_12_15, output_11_510;
mixer gate_output_11_510(.a(output_12_510), .b(output_12_15), .y(output_11_510));
wire output_13_510, output_13_15, output_12_510;
mixer gate_output_12_510(.a(output_13_510), .b(output_13_15), .y(output_12_510));
wire output_14_510, output_14_15, output_13_510;
mixer gate_output_13_510(.a(output_14_510), .b(output_14_15), .y(output_13_510));
wire output_15_510, output_15_15, output_14_510;
mixer gate_output_14_510(.a(output_15_510), .b(output_15_15), .y(output_14_510));
wire output_16_510, output_16_15, output_15_510;
mixer gate_output_15_510(.a(output_16_510), .b(output_16_15), .y(output_15_510));
wire output_1_511, output_1_0, output_0_511;
mixer gate_output_0_511(.a(output_1_511), .b(output_1_0), .y(output_0_511));
wire output_2_511, output_2_0, output_1_511;
mixer gate_output_1_511(.a(output_2_511), .b(output_2_0), .y(output_1_511));
wire output_3_511, output_3_0, output_2_511;
mixer gate_output_2_511(.a(output_3_511), .b(output_3_0), .y(output_2_511));
wire output_4_511, output_4_0, output_3_511;
mixer gate_output_3_511(.a(output_4_511), .b(output_4_0), .y(output_3_511));
wire output_5_511, output_5_0, output_4_511;
mixer gate_output_4_511(.a(output_5_511), .b(output_5_0), .y(output_4_511));
wire output_6_511, output_6_0, output_5_511;
mixer gate_output_5_511(.a(output_6_511), .b(output_6_0), .y(output_5_511));
wire output_7_511, output_7_0, output_6_511;
mixer gate_output_6_511(.a(output_7_511), .b(output_7_0), .y(output_6_511));
wire output_8_511, output_8_0, output_7_511;
mixer gate_output_7_511(.a(output_8_511), .b(output_8_0), .y(output_7_511));
wire output_9_511, output_9_0, output_8_511;
mixer gate_output_8_511(.a(output_9_511), .b(output_9_0), .y(output_8_511));
wire output_10_511, output_10_0, output_9_511;
mixer gate_output_9_511(.a(output_10_511), .b(output_10_0), .y(output_9_511));
wire output_11_511, output_11_0, output_10_511;
mixer gate_output_10_511(.a(output_11_511), .b(output_11_0), .y(output_10_511));
wire output_12_511, output_12_0, output_11_511;
mixer gate_output_11_511(.a(output_12_511), .b(output_12_0), .y(output_11_511));
wire output_13_511, output_13_0, output_12_511;
mixer gate_output_12_511(.a(output_13_511), .b(output_13_0), .y(output_12_511));
wire output_14_511, output_14_0, output_13_511;
mixer gate_output_13_511(.a(output_14_511), .b(output_14_0), .y(output_13_511));
wire output_15_511, output_15_0, output_14_511;
mixer gate_output_14_511(.a(output_15_511), .b(output_15_0), .y(output_14_511));
wire output_16_511, output_16_0, output_15_511;
mixer gate_output_15_511(.a(output_16_511), .b(output_16_0), .y(output_15_511));
wire output_1_512, output_1_1, output_0_512;
mixer gate_output_0_512(.a(output_1_512), .b(output_1_1), .y(output_0_512));
wire output_2_512, output_2_1, output_1_512;
mixer gate_output_1_512(.a(output_2_512), .b(output_2_1), .y(output_1_512));
wire output_3_512, output_3_1, output_2_512;
mixer gate_output_2_512(.a(output_3_512), .b(output_3_1), .y(output_2_512));
wire output_4_512, output_4_1, output_3_512;
mixer gate_output_3_512(.a(output_4_512), .b(output_4_1), .y(output_3_512));
wire output_5_512, output_5_1, output_4_512;
mixer gate_output_4_512(.a(output_5_512), .b(output_5_1), .y(output_4_512));
wire output_6_512, output_6_1, output_5_512;
mixer gate_output_5_512(.a(output_6_512), .b(output_6_1), .y(output_5_512));
wire output_7_512, output_7_1, output_6_512;
mixer gate_output_6_512(.a(output_7_512), .b(output_7_1), .y(output_6_512));
wire output_8_512, output_8_1, output_7_512;
mixer gate_output_7_512(.a(output_8_512), .b(output_8_1), .y(output_7_512));
wire output_9_512, output_9_1, output_8_512;
mixer gate_output_8_512(.a(output_9_512), .b(output_9_1), .y(output_8_512));
wire output_10_512, output_10_1, output_9_512;
mixer gate_output_9_512(.a(output_10_512), .b(output_10_1), .y(output_9_512));
wire output_11_512, output_11_1, output_10_512;
mixer gate_output_10_512(.a(output_11_512), .b(output_11_1), .y(output_10_512));
wire output_12_512, output_12_1, output_11_512;
mixer gate_output_11_512(.a(output_12_512), .b(output_12_1), .y(output_11_512));
wire output_13_512, output_13_1, output_12_512;
mixer gate_output_12_512(.a(output_13_512), .b(output_13_1), .y(output_12_512));
wire output_14_512, output_14_1, output_13_512;
mixer gate_output_13_512(.a(output_14_512), .b(output_14_1), .y(output_13_512));
wire output_15_512, output_15_1, output_14_512;
mixer gate_output_14_512(.a(output_15_512), .b(output_15_1), .y(output_14_512));
wire output_16_512, output_16_1, output_15_512;
mixer gate_output_15_512(.a(output_16_512), .b(output_16_1), .y(output_15_512));
wire output_1_513, output_1_2, output_0_513;
mixer gate_output_0_513(.a(output_1_513), .b(output_1_2), .y(output_0_513));
wire output_2_513, output_2_2, output_1_513;
mixer gate_output_1_513(.a(output_2_513), .b(output_2_2), .y(output_1_513));
wire output_3_513, output_3_2, output_2_513;
mixer gate_output_2_513(.a(output_3_513), .b(output_3_2), .y(output_2_513));
wire output_4_513, output_4_2, output_3_513;
mixer gate_output_3_513(.a(output_4_513), .b(output_4_2), .y(output_3_513));
wire output_5_513, output_5_2, output_4_513;
mixer gate_output_4_513(.a(output_5_513), .b(output_5_2), .y(output_4_513));
wire output_6_513, output_6_2, output_5_513;
mixer gate_output_5_513(.a(output_6_513), .b(output_6_2), .y(output_5_513));
wire output_7_513, output_7_2, output_6_513;
mixer gate_output_6_513(.a(output_7_513), .b(output_7_2), .y(output_6_513));
wire output_8_513, output_8_2, output_7_513;
mixer gate_output_7_513(.a(output_8_513), .b(output_8_2), .y(output_7_513));
wire output_9_513, output_9_2, output_8_513;
mixer gate_output_8_513(.a(output_9_513), .b(output_9_2), .y(output_8_513));
wire output_10_513, output_10_2, output_9_513;
mixer gate_output_9_513(.a(output_10_513), .b(output_10_2), .y(output_9_513));
wire output_11_513, output_11_2, output_10_513;
mixer gate_output_10_513(.a(output_11_513), .b(output_11_2), .y(output_10_513));
wire output_12_513, output_12_2, output_11_513;
mixer gate_output_11_513(.a(output_12_513), .b(output_12_2), .y(output_11_513));
wire output_13_513, output_13_2, output_12_513;
mixer gate_output_12_513(.a(output_13_513), .b(output_13_2), .y(output_12_513));
wire output_14_513, output_14_2, output_13_513;
mixer gate_output_13_513(.a(output_14_513), .b(output_14_2), .y(output_13_513));
wire output_15_513, output_15_2, output_14_513;
mixer gate_output_14_513(.a(output_15_513), .b(output_15_2), .y(output_14_513));
wire output_16_513, output_16_2, output_15_513;
mixer gate_output_15_513(.a(output_16_513), .b(output_16_2), .y(output_15_513));
wire output_1_514, output_1_3, output_0_514;
mixer gate_output_0_514(.a(output_1_514), .b(output_1_3), .y(output_0_514));
wire output_2_514, output_2_3, output_1_514;
mixer gate_output_1_514(.a(output_2_514), .b(output_2_3), .y(output_1_514));
wire output_3_514, output_3_3, output_2_514;
mixer gate_output_2_514(.a(output_3_514), .b(output_3_3), .y(output_2_514));
wire output_4_514, output_4_3, output_3_514;
mixer gate_output_3_514(.a(output_4_514), .b(output_4_3), .y(output_3_514));
wire output_5_514, output_5_3, output_4_514;
mixer gate_output_4_514(.a(output_5_514), .b(output_5_3), .y(output_4_514));
wire output_6_514, output_6_3, output_5_514;
mixer gate_output_5_514(.a(output_6_514), .b(output_6_3), .y(output_5_514));
wire output_7_514, output_7_3, output_6_514;
mixer gate_output_6_514(.a(output_7_514), .b(output_7_3), .y(output_6_514));
wire output_8_514, output_8_3, output_7_514;
mixer gate_output_7_514(.a(output_8_514), .b(output_8_3), .y(output_7_514));
wire output_9_514, output_9_3, output_8_514;
mixer gate_output_8_514(.a(output_9_514), .b(output_9_3), .y(output_8_514));
wire output_10_514, output_10_3, output_9_514;
mixer gate_output_9_514(.a(output_10_514), .b(output_10_3), .y(output_9_514));
wire output_11_514, output_11_3, output_10_514;
mixer gate_output_10_514(.a(output_11_514), .b(output_11_3), .y(output_10_514));
wire output_12_514, output_12_3, output_11_514;
mixer gate_output_11_514(.a(output_12_514), .b(output_12_3), .y(output_11_514));
wire output_13_514, output_13_3, output_12_514;
mixer gate_output_12_514(.a(output_13_514), .b(output_13_3), .y(output_12_514));
wire output_14_514, output_14_3, output_13_514;
mixer gate_output_13_514(.a(output_14_514), .b(output_14_3), .y(output_13_514));
wire output_15_514, output_15_3, output_14_514;
mixer gate_output_14_514(.a(output_15_514), .b(output_15_3), .y(output_14_514));
wire output_16_514, output_16_3, output_15_514;
mixer gate_output_15_514(.a(output_16_514), .b(output_16_3), .y(output_15_514));
wire output_1_515, output_1_4, output_0_515;
mixer gate_output_0_515(.a(output_1_515), .b(output_1_4), .y(output_0_515));
wire output_2_515, output_2_4, output_1_515;
mixer gate_output_1_515(.a(output_2_515), .b(output_2_4), .y(output_1_515));
wire output_3_515, output_3_4, output_2_515;
mixer gate_output_2_515(.a(output_3_515), .b(output_3_4), .y(output_2_515));
wire output_4_515, output_4_4, output_3_515;
mixer gate_output_3_515(.a(output_4_515), .b(output_4_4), .y(output_3_515));
wire output_5_515, output_5_4, output_4_515;
mixer gate_output_4_515(.a(output_5_515), .b(output_5_4), .y(output_4_515));
wire output_6_515, output_6_4, output_5_515;
mixer gate_output_5_515(.a(output_6_515), .b(output_6_4), .y(output_5_515));
wire output_7_515, output_7_4, output_6_515;
mixer gate_output_6_515(.a(output_7_515), .b(output_7_4), .y(output_6_515));
wire output_8_515, output_8_4, output_7_515;
mixer gate_output_7_515(.a(output_8_515), .b(output_8_4), .y(output_7_515));
wire output_9_515, output_9_4, output_8_515;
mixer gate_output_8_515(.a(output_9_515), .b(output_9_4), .y(output_8_515));
wire output_10_515, output_10_4, output_9_515;
mixer gate_output_9_515(.a(output_10_515), .b(output_10_4), .y(output_9_515));
wire output_11_515, output_11_4, output_10_515;
mixer gate_output_10_515(.a(output_11_515), .b(output_11_4), .y(output_10_515));
wire output_12_515, output_12_4, output_11_515;
mixer gate_output_11_515(.a(output_12_515), .b(output_12_4), .y(output_11_515));
wire output_13_515, output_13_4, output_12_515;
mixer gate_output_12_515(.a(output_13_515), .b(output_13_4), .y(output_12_515));
wire output_14_515, output_14_4, output_13_515;
mixer gate_output_13_515(.a(output_14_515), .b(output_14_4), .y(output_13_515));
wire output_15_515, output_15_4, output_14_515;
mixer gate_output_14_515(.a(output_15_515), .b(output_15_4), .y(output_14_515));
wire output_16_515, output_16_4, output_15_515;
mixer gate_output_15_515(.a(output_16_515), .b(output_16_4), .y(output_15_515));
wire output_1_516, output_1_5, output_0_516;
mixer gate_output_0_516(.a(output_1_516), .b(output_1_5), .y(output_0_516));
wire output_2_516, output_2_5, output_1_516;
mixer gate_output_1_516(.a(output_2_516), .b(output_2_5), .y(output_1_516));
wire output_3_516, output_3_5, output_2_516;
mixer gate_output_2_516(.a(output_3_516), .b(output_3_5), .y(output_2_516));
wire output_4_516, output_4_5, output_3_516;
mixer gate_output_3_516(.a(output_4_516), .b(output_4_5), .y(output_3_516));
wire output_5_516, output_5_5, output_4_516;
mixer gate_output_4_516(.a(output_5_516), .b(output_5_5), .y(output_4_516));
wire output_6_516, output_6_5, output_5_516;
mixer gate_output_5_516(.a(output_6_516), .b(output_6_5), .y(output_5_516));
wire output_7_516, output_7_5, output_6_516;
mixer gate_output_6_516(.a(output_7_516), .b(output_7_5), .y(output_6_516));
wire output_8_516, output_8_5, output_7_516;
mixer gate_output_7_516(.a(output_8_516), .b(output_8_5), .y(output_7_516));
wire output_9_516, output_9_5, output_8_516;
mixer gate_output_8_516(.a(output_9_516), .b(output_9_5), .y(output_8_516));
wire output_10_516, output_10_5, output_9_516;
mixer gate_output_9_516(.a(output_10_516), .b(output_10_5), .y(output_9_516));
wire output_11_516, output_11_5, output_10_516;
mixer gate_output_10_516(.a(output_11_516), .b(output_11_5), .y(output_10_516));
wire output_12_516, output_12_5, output_11_516;
mixer gate_output_11_516(.a(output_12_516), .b(output_12_5), .y(output_11_516));
wire output_13_516, output_13_5, output_12_516;
mixer gate_output_12_516(.a(output_13_516), .b(output_13_5), .y(output_12_516));
wire output_14_516, output_14_5, output_13_516;
mixer gate_output_13_516(.a(output_14_516), .b(output_14_5), .y(output_13_516));
wire output_15_516, output_15_5, output_14_516;
mixer gate_output_14_516(.a(output_15_516), .b(output_15_5), .y(output_14_516));
wire output_16_516, output_16_5, output_15_516;
mixer gate_output_15_516(.a(output_16_516), .b(output_16_5), .y(output_15_516));
wire output_1_517, output_1_6, output_0_517;
mixer gate_output_0_517(.a(output_1_517), .b(output_1_6), .y(output_0_517));
wire output_2_517, output_2_6, output_1_517;
mixer gate_output_1_517(.a(output_2_517), .b(output_2_6), .y(output_1_517));
wire output_3_517, output_3_6, output_2_517;
mixer gate_output_2_517(.a(output_3_517), .b(output_3_6), .y(output_2_517));
wire output_4_517, output_4_6, output_3_517;
mixer gate_output_3_517(.a(output_4_517), .b(output_4_6), .y(output_3_517));
wire output_5_517, output_5_6, output_4_517;
mixer gate_output_4_517(.a(output_5_517), .b(output_5_6), .y(output_4_517));
wire output_6_517, output_6_6, output_5_517;
mixer gate_output_5_517(.a(output_6_517), .b(output_6_6), .y(output_5_517));
wire output_7_517, output_7_6, output_6_517;
mixer gate_output_6_517(.a(output_7_517), .b(output_7_6), .y(output_6_517));
wire output_8_517, output_8_6, output_7_517;
mixer gate_output_7_517(.a(output_8_517), .b(output_8_6), .y(output_7_517));
wire output_9_517, output_9_6, output_8_517;
mixer gate_output_8_517(.a(output_9_517), .b(output_9_6), .y(output_8_517));
wire output_10_517, output_10_6, output_9_517;
mixer gate_output_9_517(.a(output_10_517), .b(output_10_6), .y(output_9_517));
wire output_11_517, output_11_6, output_10_517;
mixer gate_output_10_517(.a(output_11_517), .b(output_11_6), .y(output_10_517));
wire output_12_517, output_12_6, output_11_517;
mixer gate_output_11_517(.a(output_12_517), .b(output_12_6), .y(output_11_517));
wire output_13_517, output_13_6, output_12_517;
mixer gate_output_12_517(.a(output_13_517), .b(output_13_6), .y(output_12_517));
wire output_14_517, output_14_6, output_13_517;
mixer gate_output_13_517(.a(output_14_517), .b(output_14_6), .y(output_13_517));
wire output_15_517, output_15_6, output_14_517;
mixer gate_output_14_517(.a(output_15_517), .b(output_15_6), .y(output_14_517));
wire output_16_517, output_16_6, output_15_517;
mixer gate_output_15_517(.a(output_16_517), .b(output_16_6), .y(output_15_517));
wire output_1_518, output_1_7, output_0_518;
mixer gate_output_0_518(.a(output_1_518), .b(output_1_7), .y(output_0_518));
wire output_2_518, output_2_7, output_1_518;
mixer gate_output_1_518(.a(output_2_518), .b(output_2_7), .y(output_1_518));
wire output_3_518, output_3_7, output_2_518;
mixer gate_output_2_518(.a(output_3_518), .b(output_3_7), .y(output_2_518));
wire output_4_518, output_4_7, output_3_518;
mixer gate_output_3_518(.a(output_4_518), .b(output_4_7), .y(output_3_518));
wire output_5_518, output_5_7, output_4_518;
mixer gate_output_4_518(.a(output_5_518), .b(output_5_7), .y(output_4_518));
wire output_6_518, output_6_7, output_5_518;
mixer gate_output_5_518(.a(output_6_518), .b(output_6_7), .y(output_5_518));
wire output_7_518, output_7_7, output_6_518;
mixer gate_output_6_518(.a(output_7_518), .b(output_7_7), .y(output_6_518));
wire output_8_518, output_8_7, output_7_518;
mixer gate_output_7_518(.a(output_8_518), .b(output_8_7), .y(output_7_518));
wire output_9_518, output_9_7, output_8_518;
mixer gate_output_8_518(.a(output_9_518), .b(output_9_7), .y(output_8_518));
wire output_10_518, output_10_7, output_9_518;
mixer gate_output_9_518(.a(output_10_518), .b(output_10_7), .y(output_9_518));
wire output_11_518, output_11_7, output_10_518;
mixer gate_output_10_518(.a(output_11_518), .b(output_11_7), .y(output_10_518));
wire output_12_518, output_12_7, output_11_518;
mixer gate_output_11_518(.a(output_12_518), .b(output_12_7), .y(output_11_518));
wire output_13_518, output_13_7, output_12_518;
mixer gate_output_12_518(.a(output_13_518), .b(output_13_7), .y(output_12_518));
wire output_14_518, output_14_7, output_13_518;
mixer gate_output_13_518(.a(output_14_518), .b(output_14_7), .y(output_13_518));
wire output_15_518, output_15_7, output_14_518;
mixer gate_output_14_518(.a(output_15_518), .b(output_15_7), .y(output_14_518));
wire output_16_518, output_16_7, output_15_518;
mixer gate_output_15_518(.a(output_16_518), .b(output_16_7), .y(output_15_518));
wire output_1_519, output_1_8, output_0_519;
mixer gate_output_0_519(.a(output_1_519), .b(output_1_8), .y(output_0_519));
wire output_2_519, output_2_8, output_1_519;
mixer gate_output_1_519(.a(output_2_519), .b(output_2_8), .y(output_1_519));
wire output_3_519, output_3_8, output_2_519;
mixer gate_output_2_519(.a(output_3_519), .b(output_3_8), .y(output_2_519));
wire output_4_519, output_4_8, output_3_519;
mixer gate_output_3_519(.a(output_4_519), .b(output_4_8), .y(output_3_519));
wire output_5_519, output_5_8, output_4_519;
mixer gate_output_4_519(.a(output_5_519), .b(output_5_8), .y(output_4_519));
wire output_6_519, output_6_8, output_5_519;
mixer gate_output_5_519(.a(output_6_519), .b(output_6_8), .y(output_5_519));
wire output_7_519, output_7_8, output_6_519;
mixer gate_output_6_519(.a(output_7_519), .b(output_7_8), .y(output_6_519));
wire output_8_519, output_8_8, output_7_519;
mixer gate_output_7_519(.a(output_8_519), .b(output_8_8), .y(output_7_519));
wire output_9_519, output_9_8, output_8_519;
mixer gate_output_8_519(.a(output_9_519), .b(output_9_8), .y(output_8_519));
wire output_10_519, output_10_8, output_9_519;
mixer gate_output_9_519(.a(output_10_519), .b(output_10_8), .y(output_9_519));
wire output_11_519, output_11_8, output_10_519;
mixer gate_output_10_519(.a(output_11_519), .b(output_11_8), .y(output_10_519));
wire output_12_519, output_12_8, output_11_519;
mixer gate_output_11_519(.a(output_12_519), .b(output_12_8), .y(output_11_519));
wire output_13_519, output_13_8, output_12_519;
mixer gate_output_12_519(.a(output_13_519), .b(output_13_8), .y(output_12_519));
wire output_14_519, output_14_8, output_13_519;
mixer gate_output_13_519(.a(output_14_519), .b(output_14_8), .y(output_13_519));
wire output_15_519, output_15_8, output_14_519;
mixer gate_output_14_519(.a(output_15_519), .b(output_15_8), .y(output_14_519));
wire output_16_519, output_16_8, output_15_519;
mixer gate_output_15_519(.a(output_16_519), .b(output_16_8), .y(output_15_519));
wire output_1_520, output_1_9, output_0_520;
mixer gate_output_0_520(.a(output_1_520), .b(output_1_9), .y(output_0_520));
wire output_2_520, output_2_9, output_1_520;
mixer gate_output_1_520(.a(output_2_520), .b(output_2_9), .y(output_1_520));
wire output_3_520, output_3_9, output_2_520;
mixer gate_output_2_520(.a(output_3_520), .b(output_3_9), .y(output_2_520));
wire output_4_520, output_4_9, output_3_520;
mixer gate_output_3_520(.a(output_4_520), .b(output_4_9), .y(output_3_520));
wire output_5_520, output_5_9, output_4_520;
mixer gate_output_4_520(.a(output_5_520), .b(output_5_9), .y(output_4_520));
wire output_6_520, output_6_9, output_5_520;
mixer gate_output_5_520(.a(output_6_520), .b(output_6_9), .y(output_5_520));
wire output_7_520, output_7_9, output_6_520;
mixer gate_output_6_520(.a(output_7_520), .b(output_7_9), .y(output_6_520));
wire output_8_520, output_8_9, output_7_520;
mixer gate_output_7_520(.a(output_8_520), .b(output_8_9), .y(output_7_520));
wire output_9_520, output_9_9, output_8_520;
mixer gate_output_8_520(.a(output_9_520), .b(output_9_9), .y(output_8_520));
wire output_10_520, output_10_9, output_9_520;
mixer gate_output_9_520(.a(output_10_520), .b(output_10_9), .y(output_9_520));
wire output_11_520, output_11_9, output_10_520;
mixer gate_output_10_520(.a(output_11_520), .b(output_11_9), .y(output_10_520));
wire output_12_520, output_12_9, output_11_520;
mixer gate_output_11_520(.a(output_12_520), .b(output_12_9), .y(output_11_520));
wire output_13_520, output_13_9, output_12_520;
mixer gate_output_12_520(.a(output_13_520), .b(output_13_9), .y(output_12_520));
wire output_14_520, output_14_9, output_13_520;
mixer gate_output_13_520(.a(output_14_520), .b(output_14_9), .y(output_13_520));
wire output_15_520, output_15_9, output_14_520;
mixer gate_output_14_520(.a(output_15_520), .b(output_15_9), .y(output_14_520));
wire output_16_520, output_16_9, output_15_520;
mixer gate_output_15_520(.a(output_16_520), .b(output_16_9), .y(output_15_520));
wire output_1_521, output_1_10, output_0_521;
mixer gate_output_0_521(.a(output_1_521), .b(output_1_10), .y(output_0_521));
wire output_2_521, output_2_10, output_1_521;
mixer gate_output_1_521(.a(output_2_521), .b(output_2_10), .y(output_1_521));
wire output_3_521, output_3_10, output_2_521;
mixer gate_output_2_521(.a(output_3_521), .b(output_3_10), .y(output_2_521));
wire output_4_521, output_4_10, output_3_521;
mixer gate_output_3_521(.a(output_4_521), .b(output_4_10), .y(output_3_521));
wire output_5_521, output_5_10, output_4_521;
mixer gate_output_4_521(.a(output_5_521), .b(output_5_10), .y(output_4_521));
wire output_6_521, output_6_10, output_5_521;
mixer gate_output_5_521(.a(output_6_521), .b(output_6_10), .y(output_5_521));
wire output_7_521, output_7_10, output_6_521;
mixer gate_output_6_521(.a(output_7_521), .b(output_7_10), .y(output_6_521));
wire output_8_521, output_8_10, output_7_521;
mixer gate_output_7_521(.a(output_8_521), .b(output_8_10), .y(output_7_521));
wire output_9_521, output_9_10, output_8_521;
mixer gate_output_8_521(.a(output_9_521), .b(output_9_10), .y(output_8_521));
wire output_10_521, output_10_10, output_9_521;
mixer gate_output_9_521(.a(output_10_521), .b(output_10_10), .y(output_9_521));
wire output_11_521, output_11_10, output_10_521;
mixer gate_output_10_521(.a(output_11_521), .b(output_11_10), .y(output_10_521));
wire output_12_521, output_12_10, output_11_521;
mixer gate_output_11_521(.a(output_12_521), .b(output_12_10), .y(output_11_521));
wire output_13_521, output_13_10, output_12_521;
mixer gate_output_12_521(.a(output_13_521), .b(output_13_10), .y(output_12_521));
wire output_14_521, output_14_10, output_13_521;
mixer gate_output_13_521(.a(output_14_521), .b(output_14_10), .y(output_13_521));
wire output_15_521, output_15_10, output_14_521;
mixer gate_output_14_521(.a(output_15_521), .b(output_15_10), .y(output_14_521));
wire output_16_521, output_16_10, output_15_521;
mixer gate_output_15_521(.a(output_16_521), .b(output_16_10), .y(output_15_521));
wire output_1_522, output_1_11, output_0_522;
mixer gate_output_0_522(.a(output_1_522), .b(output_1_11), .y(output_0_522));
wire output_2_522, output_2_11, output_1_522;
mixer gate_output_1_522(.a(output_2_522), .b(output_2_11), .y(output_1_522));
wire output_3_522, output_3_11, output_2_522;
mixer gate_output_2_522(.a(output_3_522), .b(output_3_11), .y(output_2_522));
wire output_4_522, output_4_11, output_3_522;
mixer gate_output_3_522(.a(output_4_522), .b(output_4_11), .y(output_3_522));
wire output_5_522, output_5_11, output_4_522;
mixer gate_output_4_522(.a(output_5_522), .b(output_5_11), .y(output_4_522));
wire output_6_522, output_6_11, output_5_522;
mixer gate_output_5_522(.a(output_6_522), .b(output_6_11), .y(output_5_522));
wire output_7_522, output_7_11, output_6_522;
mixer gate_output_6_522(.a(output_7_522), .b(output_7_11), .y(output_6_522));
wire output_8_522, output_8_11, output_7_522;
mixer gate_output_7_522(.a(output_8_522), .b(output_8_11), .y(output_7_522));
wire output_9_522, output_9_11, output_8_522;
mixer gate_output_8_522(.a(output_9_522), .b(output_9_11), .y(output_8_522));
wire output_10_522, output_10_11, output_9_522;
mixer gate_output_9_522(.a(output_10_522), .b(output_10_11), .y(output_9_522));
wire output_11_522, output_11_11, output_10_522;
mixer gate_output_10_522(.a(output_11_522), .b(output_11_11), .y(output_10_522));
wire output_12_522, output_12_11, output_11_522;
mixer gate_output_11_522(.a(output_12_522), .b(output_12_11), .y(output_11_522));
wire output_13_522, output_13_11, output_12_522;
mixer gate_output_12_522(.a(output_13_522), .b(output_13_11), .y(output_12_522));
wire output_14_522, output_14_11, output_13_522;
mixer gate_output_13_522(.a(output_14_522), .b(output_14_11), .y(output_13_522));
wire output_15_522, output_15_11, output_14_522;
mixer gate_output_14_522(.a(output_15_522), .b(output_15_11), .y(output_14_522));
wire output_16_522, output_16_11, output_15_522;
mixer gate_output_15_522(.a(output_16_522), .b(output_16_11), .y(output_15_522));
wire output_1_523, output_1_12, output_0_523;
mixer gate_output_0_523(.a(output_1_523), .b(output_1_12), .y(output_0_523));
wire output_2_523, output_2_12, output_1_523;
mixer gate_output_1_523(.a(output_2_523), .b(output_2_12), .y(output_1_523));
wire output_3_523, output_3_12, output_2_523;
mixer gate_output_2_523(.a(output_3_523), .b(output_3_12), .y(output_2_523));
wire output_4_523, output_4_12, output_3_523;
mixer gate_output_3_523(.a(output_4_523), .b(output_4_12), .y(output_3_523));
wire output_5_523, output_5_12, output_4_523;
mixer gate_output_4_523(.a(output_5_523), .b(output_5_12), .y(output_4_523));
wire output_6_523, output_6_12, output_5_523;
mixer gate_output_5_523(.a(output_6_523), .b(output_6_12), .y(output_5_523));
wire output_7_523, output_7_12, output_6_523;
mixer gate_output_6_523(.a(output_7_523), .b(output_7_12), .y(output_6_523));
wire output_8_523, output_8_12, output_7_523;
mixer gate_output_7_523(.a(output_8_523), .b(output_8_12), .y(output_7_523));
wire output_9_523, output_9_12, output_8_523;
mixer gate_output_8_523(.a(output_9_523), .b(output_9_12), .y(output_8_523));
wire output_10_523, output_10_12, output_9_523;
mixer gate_output_9_523(.a(output_10_523), .b(output_10_12), .y(output_9_523));
wire output_11_523, output_11_12, output_10_523;
mixer gate_output_10_523(.a(output_11_523), .b(output_11_12), .y(output_10_523));
wire output_12_523, output_12_12, output_11_523;
mixer gate_output_11_523(.a(output_12_523), .b(output_12_12), .y(output_11_523));
wire output_13_523, output_13_12, output_12_523;
mixer gate_output_12_523(.a(output_13_523), .b(output_13_12), .y(output_12_523));
wire output_14_523, output_14_12, output_13_523;
mixer gate_output_13_523(.a(output_14_523), .b(output_14_12), .y(output_13_523));
wire output_15_523, output_15_12, output_14_523;
mixer gate_output_14_523(.a(output_15_523), .b(output_15_12), .y(output_14_523));
wire output_16_523, output_16_12, output_15_523;
mixer gate_output_15_523(.a(output_16_523), .b(output_16_12), .y(output_15_523));
wire output_1_524, output_1_13, output_0_524;
mixer gate_output_0_524(.a(output_1_524), .b(output_1_13), .y(output_0_524));
wire output_2_524, output_2_13, output_1_524;
mixer gate_output_1_524(.a(output_2_524), .b(output_2_13), .y(output_1_524));
wire output_3_524, output_3_13, output_2_524;
mixer gate_output_2_524(.a(output_3_524), .b(output_3_13), .y(output_2_524));
wire output_4_524, output_4_13, output_3_524;
mixer gate_output_3_524(.a(output_4_524), .b(output_4_13), .y(output_3_524));
wire output_5_524, output_5_13, output_4_524;
mixer gate_output_4_524(.a(output_5_524), .b(output_5_13), .y(output_4_524));
wire output_6_524, output_6_13, output_5_524;
mixer gate_output_5_524(.a(output_6_524), .b(output_6_13), .y(output_5_524));
wire output_7_524, output_7_13, output_6_524;
mixer gate_output_6_524(.a(output_7_524), .b(output_7_13), .y(output_6_524));
wire output_8_524, output_8_13, output_7_524;
mixer gate_output_7_524(.a(output_8_524), .b(output_8_13), .y(output_7_524));
wire output_9_524, output_9_13, output_8_524;
mixer gate_output_8_524(.a(output_9_524), .b(output_9_13), .y(output_8_524));
wire output_10_524, output_10_13, output_9_524;
mixer gate_output_9_524(.a(output_10_524), .b(output_10_13), .y(output_9_524));
wire output_11_524, output_11_13, output_10_524;
mixer gate_output_10_524(.a(output_11_524), .b(output_11_13), .y(output_10_524));
wire output_12_524, output_12_13, output_11_524;
mixer gate_output_11_524(.a(output_12_524), .b(output_12_13), .y(output_11_524));
wire output_13_524, output_13_13, output_12_524;
mixer gate_output_12_524(.a(output_13_524), .b(output_13_13), .y(output_12_524));
wire output_14_524, output_14_13, output_13_524;
mixer gate_output_13_524(.a(output_14_524), .b(output_14_13), .y(output_13_524));
wire output_15_524, output_15_13, output_14_524;
mixer gate_output_14_524(.a(output_15_524), .b(output_15_13), .y(output_14_524));
wire output_16_524, output_16_13, output_15_524;
mixer gate_output_15_524(.a(output_16_524), .b(output_16_13), .y(output_15_524));
wire output_1_525, output_1_14, output_0_525;
mixer gate_output_0_525(.a(output_1_525), .b(output_1_14), .y(output_0_525));
wire output_2_525, output_2_14, output_1_525;
mixer gate_output_1_525(.a(output_2_525), .b(output_2_14), .y(output_1_525));
wire output_3_525, output_3_14, output_2_525;
mixer gate_output_2_525(.a(output_3_525), .b(output_3_14), .y(output_2_525));
wire output_4_525, output_4_14, output_3_525;
mixer gate_output_3_525(.a(output_4_525), .b(output_4_14), .y(output_3_525));
wire output_5_525, output_5_14, output_4_525;
mixer gate_output_4_525(.a(output_5_525), .b(output_5_14), .y(output_4_525));
wire output_6_525, output_6_14, output_5_525;
mixer gate_output_5_525(.a(output_6_525), .b(output_6_14), .y(output_5_525));
wire output_7_525, output_7_14, output_6_525;
mixer gate_output_6_525(.a(output_7_525), .b(output_7_14), .y(output_6_525));
wire output_8_525, output_8_14, output_7_525;
mixer gate_output_7_525(.a(output_8_525), .b(output_8_14), .y(output_7_525));
wire output_9_525, output_9_14, output_8_525;
mixer gate_output_8_525(.a(output_9_525), .b(output_9_14), .y(output_8_525));
wire output_10_525, output_10_14, output_9_525;
mixer gate_output_9_525(.a(output_10_525), .b(output_10_14), .y(output_9_525));
wire output_11_525, output_11_14, output_10_525;
mixer gate_output_10_525(.a(output_11_525), .b(output_11_14), .y(output_10_525));
wire output_12_525, output_12_14, output_11_525;
mixer gate_output_11_525(.a(output_12_525), .b(output_12_14), .y(output_11_525));
wire output_13_525, output_13_14, output_12_525;
mixer gate_output_12_525(.a(output_13_525), .b(output_13_14), .y(output_12_525));
wire output_14_525, output_14_14, output_13_525;
mixer gate_output_13_525(.a(output_14_525), .b(output_14_14), .y(output_13_525));
wire output_15_525, output_15_14, output_14_525;
mixer gate_output_14_525(.a(output_15_525), .b(output_15_14), .y(output_14_525));
wire output_16_525, output_16_14, output_15_525;
mixer gate_output_15_525(.a(output_16_525), .b(output_16_14), .y(output_15_525));
wire output_1_526, output_1_15, output_0_526;
mixer gate_output_0_526(.a(output_1_526), .b(output_1_15), .y(output_0_526));
wire output_2_526, output_2_15, output_1_526;
mixer gate_output_1_526(.a(output_2_526), .b(output_2_15), .y(output_1_526));
wire output_3_526, output_3_15, output_2_526;
mixer gate_output_2_526(.a(output_3_526), .b(output_3_15), .y(output_2_526));
wire output_4_526, output_4_15, output_3_526;
mixer gate_output_3_526(.a(output_4_526), .b(output_4_15), .y(output_3_526));
wire output_5_526, output_5_15, output_4_526;
mixer gate_output_4_526(.a(output_5_526), .b(output_5_15), .y(output_4_526));
wire output_6_526, output_6_15, output_5_526;
mixer gate_output_5_526(.a(output_6_526), .b(output_6_15), .y(output_5_526));
wire output_7_526, output_7_15, output_6_526;
mixer gate_output_6_526(.a(output_7_526), .b(output_7_15), .y(output_6_526));
wire output_8_526, output_8_15, output_7_526;
mixer gate_output_7_526(.a(output_8_526), .b(output_8_15), .y(output_7_526));
wire output_9_526, output_9_15, output_8_526;
mixer gate_output_8_526(.a(output_9_526), .b(output_9_15), .y(output_8_526));
wire output_10_526, output_10_15, output_9_526;
mixer gate_output_9_526(.a(output_10_526), .b(output_10_15), .y(output_9_526));
wire output_11_526, output_11_15, output_10_526;
mixer gate_output_10_526(.a(output_11_526), .b(output_11_15), .y(output_10_526));
wire output_12_526, output_12_15, output_11_526;
mixer gate_output_11_526(.a(output_12_526), .b(output_12_15), .y(output_11_526));
wire output_13_526, output_13_15, output_12_526;
mixer gate_output_12_526(.a(output_13_526), .b(output_13_15), .y(output_12_526));
wire output_14_526, output_14_15, output_13_526;
mixer gate_output_13_526(.a(output_14_526), .b(output_14_15), .y(output_13_526));
wire output_15_526, output_15_15, output_14_526;
mixer gate_output_14_526(.a(output_15_526), .b(output_15_15), .y(output_14_526));
wire output_16_526, output_16_15, output_15_526;
mixer gate_output_15_526(.a(output_16_526), .b(output_16_15), .y(output_15_526));
wire output_1_527, output_1_0, output_0_527;
mixer gate_output_0_527(.a(output_1_527), .b(output_1_0), .y(output_0_527));
wire output_2_527, output_2_0, output_1_527;
mixer gate_output_1_527(.a(output_2_527), .b(output_2_0), .y(output_1_527));
wire output_3_527, output_3_0, output_2_527;
mixer gate_output_2_527(.a(output_3_527), .b(output_3_0), .y(output_2_527));
wire output_4_527, output_4_0, output_3_527;
mixer gate_output_3_527(.a(output_4_527), .b(output_4_0), .y(output_3_527));
wire output_5_527, output_5_0, output_4_527;
mixer gate_output_4_527(.a(output_5_527), .b(output_5_0), .y(output_4_527));
wire output_6_527, output_6_0, output_5_527;
mixer gate_output_5_527(.a(output_6_527), .b(output_6_0), .y(output_5_527));
wire output_7_527, output_7_0, output_6_527;
mixer gate_output_6_527(.a(output_7_527), .b(output_7_0), .y(output_6_527));
wire output_8_527, output_8_0, output_7_527;
mixer gate_output_7_527(.a(output_8_527), .b(output_8_0), .y(output_7_527));
wire output_9_527, output_9_0, output_8_527;
mixer gate_output_8_527(.a(output_9_527), .b(output_9_0), .y(output_8_527));
wire output_10_527, output_10_0, output_9_527;
mixer gate_output_9_527(.a(output_10_527), .b(output_10_0), .y(output_9_527));
wire output_11_527, output_11_0, output_10_527;
mixer gate_output_10_527(.a(output_11_527), .b(output_11_0), .y(output_10_527));
wire output_12_527, output_12_0, output_11_527;
mixer gate_output_11_527(.a(output_12_527), .b(output_12_0), .y(output_11_527));
wire output_13_527, output_13_0, output_12_527;
mixer gate_output_12_527(.a(output_13_527), .b(output_13_0), .y(output_12_527));
wire output_14_527, output_14_0, output_13_527;
mixer gate_output_13_527(.a(output_14_527), .b(output_14_0), .y(output_13_527));
wire output_15_527, output_15_0, output_14_527;
mixer gate_output_14_527(.a(output_15_527), .b(output_15_0), .y(output_14_527));
wire output_16_527, output_16_0, output_15_527;
mixer gate_output_15_527(.a(output_16_527), .b(output_16_0), .y(output_15_527));
wire output_1_528, output_1_1, output_0_528;
mixer gate_output_0_528(.a(output_1_528), .b(output_1_1), .y(output_0_528));
wire output_2_528, output_2_1, output_1_528;
mixer gate_output_1_528(.a(output_2_528), .b(output_2_1), .y(output_1_528));
wire output_3_528, output_3_1, output_2_528;
mixer gate_output_2_528(.a(output_3_528), .b(output_3_1), .y(output_2_528));
wire output_4_528, output_4_1, output_3_528;
mixer gate_output_3_528(.a(output_4_528), .b(output_4_1), .y(output_3_528));
wire output_5_528, output_5_1, output_4_528;
mixer gate_output_4_528(.a(output_5_528), .b(output_5_1), .y(output_4_528));
wire output_6_528, output_6_1, output_5_528;
mixer gate_output_5_528(.a(output_6_528), .b(output_6_1), .y(output_5_528));
wire output_7_528, output_7_1, output_6_528;
mixer gate_output_6_528(.a(output_7_528), .b(output_7_1), .y(output_6_528));
wire output_8_528, output_8_1, output_7_528;
mixer gate_output_7_528(.a(output_8_528), .b(output_8_1), .y(output_7_528));
wire output_9_528, output_9_1, output_8_528;
mixer gate_output_8_528(.a(output_9_528), .b(output_9_1), .y(output_8_528));
wire output_10_528, output_10_1, output_9_528;
mixer gate_output_9_528(.a(output_10_528), .b(output_10_1), .y(output_9_528));
wire output_11_528, output_11_1, output_10_528;
mixer gate_output_10_528(.a(output_11_528), .b(output_11_1), .y(output_10_528));
wire output_12_528, output_12_1, output_11_528;
mixer gate_output_11_528(.a(output_12_528), .b(output_12_1), .y(output_11_528));
wire output_13_528, output_13_1, output_12_528;
mixer gate_output_12_528(.a(output_13_528), .b(output_13_1), .y(output_12_528));
wire output_14_528, output_14_1, output_13_528;
mixer gate_output_13_528(.a(output_14_528), .b(output_14_1), .y(output_13_528));
wire output_15_528, output_15_1, output_14_528;
mixer gate_output_14_528(.a(output_15_528), .b(output_15_1), .y(output_14_528));
wire output_16_528, output_16_1, output_15_528;
mixer gate_output_15_528(.a(output_16_528), .b(output_16_1), .y(output_15_528));
wire output_1_529, output_1_2, output_0_529;
mixer gate_output_0_529(.a(output_1_529), .b(output_1_2), .y(output_0_529));
wire output_2_529, output_2_2, output_1_529;
mixer gate_output_1_529(.a(output_2_529), .b(output_2_2), .y(output_1_529));
wire output_3_529, output_3_2, output_2_529;
mixer gate_output_2_529(.a(output_3_529), .b(output_3_2), .y(output_2_529));
wire output_4_529, output_4_2, output_3_529;
mixer gate_output_3_529(.a(output_4_529), .b(output_4_2), .y(output_3_529));
wire output_5_529, output_5_2, output_4_529;
mixer gate_output_4_529(.a(output_5_529), .b(output_5_2), .y(output_4_529));
wire output_6_529, output_6_2, output_5_529;
mixer gate_output_5_529(.a(output_6_529), .b(output_6_2), .y(output_5_529));
wire output_7_529, output_7_2, output_6_529;
mixer gate_output_6_529(.a(output_7_529), .b(output_7_2), .y(output_6_529));
wire output_8_529, output_8_2, output_7_529;
mixer gate_output_7_529(.a(output_8_529), .b(output_8_2), .y(output_7_529));
wire output_9_529, output_9_2, output_8_529;
mixer gate_output_8_529(.a(output_9_529), .b(output_9_2), .y(output_8_529));
wire output_10_529, output_10_2, output_9_529;
mixer gate_output_9_529(.a(output_10_529), .b(output_10_2), .y(output_9_529));
wire output_11_529, output_11_2, output_10_529;
mixer gate_output_10_529(.a(output_11_529), .b(output_11_2), .y(output_10_529));
wire output_12_529, output_12_2, output_11_529;
mixer gate_output_11_529(.a(output_12_529), .b(output_12_2), .y(output_11_529));
wire output_13_529, output_13_2, output_12_529;
mixer gate_output_12_529(.a(output_13_529), .b(output_13_2), .y(output_12_529));
wire output_14_529, output_14_2, output_13_529;
mixer gate_output_13_529(.a(output_14_529), .b(output_14_2), .y(output_13_529));
wire output_15_529, output_15_2, output_14_529;
mixer gate_output_14_529(.a(output_15_529), .b(output_15_2), .y(output_14_529));
wire output_16_529, output_16_2, output_15_529;
mixer gate_output_15_529(.a(output_16_529), .b(output_16_2), .y(output_15_529));
wire output_1_530, output_1_3, output_0_530;
mixer gate_output_0_530(.a(output_1_530), .b(output_1_3), .y(output_0_530));
wire output_2_530, output_2_3, output_1_530;
mixer gate_output_1_530(.a(output_2_530), .b(output_2_3), .y(output_1_530));
wire output_3_530, output_3_3, output_2_530;
mixer gate_output_2_530(.a(output_3_530), .b(output_3_3), .y(output_2_530));
wire output_4_530, output_4_3, output_3_530;
mixer gate_output_3_530(.a(output_4_530), .b(output_4_3), .y(output_3_530));
wire output_5_530, output_5_3, output_4_530;
mixer gate_output_4_530(.a(output_5_530), .b(output_5_3), .y(output_4_530));
wire output_6_530, output_6_3, output_5_530;
mixer gate_output_5_530(.a(output_6_530), .b(output_6_3), .y(output_5_530));
wire output_7_530, output_7_3, output_6_530;
mixer gate_output_6_530(.a(output_7_530), .b(output_7_3), .y(output_6_530));
wire output_8_530, output_8_3, output_7_530;
mixer gate_output_7_530(.a(output_8_530), .b(output_8_3), .y(output_7_530));
wire output_9_530, output_9_3, output_8_530;
mixer gate_output_8_530(.a(output_9_530), .b(output_9_3), .y(output_8_530));
wire output_10_530, output_10_3, output_9_530;
mixer gate_output_9_530(.a(output_10_530), .b(output_10_3), .y(output_9_530));
wire output_11_530, output_11_3, output_10_530;
mixer gate_output_10_530(.a(output_11_530), .b(output_11_3), .y(output_10_530));
wire output_12_530, output_12_3, output_11_530;
mixer gate_output_11_530(.a(output_12_530), .b(output_12_3), .y(output_11_530));
wire output_13_530, output_13_3, output_12_530;
mixer gate_output_12_530(.a(output_13_530), .b(output_13_3), .y(output_12_530));
wire output_14_530, output_14_3, output_13_530;
mixer gate_output_13_530(.a(output_14_530), .b(output_14_3), .y(output_13_530));
wire output_15_530, output_15_3, output_14_530;
mixer gate_output_14_530(.a(output_15_530), .b(output_15_3), .y(output_14_530));
wire output_16_530, output_16_3, output_15_530;
mixer gate_output_15_530(.a(output_16_530), .b(output_16_3), .y(output_15_530));
wire output_1_531, output_1_4, output_0_531;
mixer gate_output_0_531(.a(output_1_531), .b(output_1_4), .y(output_0_531));
wire output_2_531, output_2_4, output_1_531;
mixer gate_output_1_531(.a(output_2_531), .b(output_2_4), .y(output_1_531));
wire output_3_531, output_3_4, output_2_531;
mixer gate_output_2_531(.a(output_3_531), .b(output_3_4), .y(output_2_531));
wire output_4_531, output_4_4, output_3_531;
mixer gate_output_3_531(.a(output_4_531), .b(output_4_4), .y(output_3_531));
wire output_5_531, output_5_4, output_4_531;
mixer gate_output_4_531(.a(output_5_531), .b(output_5_4), .y(output_4_531));
wire output_6_531, output_6_4, output_5_531;
mixer gate_output_5_531(.a(output_6_531), .b(output_6_4), .y(output_5_531));
wire output_7_531, output_7_4, output_6_531;
mixer gate_output_6_531(.a(output_7_531), .b(output_7_4), .y(output_6_531));
wire output_8_531, output_8_4, output_7_531;
mixer gate_output_7_531(.a(output_8_531), .b(output_8_4), .y(output_7_531));
wire output_9_531, output_9_4, output_8_531;
mixer gate_output_8_531(.a(output_9_531), .b(output_9_4), .y(output_8_531));
wire output_10_531, output_10_4, output_9_531;
mixer gate_output_9_531(.a(output_10_531), .b(output_10_4), .y(output_9_531));
wire output_11_531, output_11_4, output_10_531;
mixer gate_output_10_531(.a(output_11_531), .b(output_11_4), .y(output_10_531));
wire output_12_531, output_12_4, output_11_531;
mixer gate_output_11_531(.a(output_12_531), .b(output_12_4), .y(output_11_531));
wire output_13_531, output_13_4, output_12_531;
mixer gate_output_12_531(.a(output_13_531), .b(output_13_4), .y(output_12_531));
wire output_14_531, output_14_4, output_13_531;
mixer gate_output_13_531(.a(output_14_531), .b(output_14_4), .y(output_13_531));
wire output_15_531, output_15_4, output_14_531;
mixer gate_output_14_531(.a(output_15_531), .b(output_15_4), .y(output_14_531));
wire output_16_531, output_16_4, output_15_531;
mixer gate_output_15_531(.a(output_16_531), .b(output_16_4), .y(output_15_531));
wire output_1_532, output_1_5, output_0_532;
mixer gate_output_0_532(.a(output_1_532), .b(output_1_5), .y(output_0_532));
wire output_2_532, output_2_5, output_1_532;
mixer gate_output_1_532(.a(output_2_532), .b(output_2_5), .y(output_1_532));
wire output_3_532, output_3_5, output_2_532;
mixer gate_output_2_532(.a(output_3_532), .b(output_3_5), .y(output_2_532));
wire output_4_532, output_4_5, output_3_532;
mixer gate_output_3_532(.a(output_4_532), .b(output_4_5), .y(output_3_532));
wire output_5_532, output_5_5, output_4_532;
mixer gate_output_4_532(.a(output_5_532), .b(output_5_5), .y(output_4_532));
wire output_6_532, output_6_5, output_5_532;
mixer gate_output_5_532(.a(output_6_532), .b(output_6_5), .y(output_5_532));
wire output_7_532, output_7_5, output_6_532;
mixer gate_output_6_532(.a(output_7_532), .b(output_7_5), .y(output_6_532));
wire output_8_532, output_8_5, output_7_532;
mixer gate_output_7_532(.a(output_8_532), .b(output_8_5), .y(output_7_532));
wire output_9_532, output_9_5, output_8_532;
mixer gate_output_8_532(.a(output_9_532), .b(output_9_5), .y(output_8_532));
wire output_10_532, output_10_5, output_9_532;
mixer gate_output_9_532(.a(output_10_532), .b(output_10_5), .y(output_9_532));
wire output_11_532, output_11_5, output_10_532;
mixer gate_output_10_532(.a(output_11_532), .b(output_11_5), .y(output_10_532));
wire output_12_532, output_12_5, output_11_532;
mixer gate_output_11_532(.a(output_12_532), .b(output_12_5), .y(output_11_532));
wire output_13_532, output_13_5, output_12_532;
mixer gate_output_12_532(.a(output_13_532), .b(output_13_5), .y(output_12_532));
wire output_14_532, output_14_5, output_13_532;
mixer gate_output_13_532(.a(output_14_532), .b(output_14_5), .y(output_13_532));
wire output_15_532, output_15_5, output_14_532;
mixer gate_output_14_532(.a(output_15_532), .b(output_15_5), .y(output_14_532));
wire output_16_532, output_16_5, output_15_532;
mixer gate_output_15_532(.a(output_16_532), .b(output_16_5), .y(output_15_532));
wire output_1_533, output_1_6, output_0_533;
mixer gate_output_0_533(.a(output_1_533), .b(output_1_6), .y(output_0_533));
wire output_2_533, output_2_6, output_1_533;
mixer gate_output_1_533(.a(output_2_533), .b(output_2_6), .y(output_1_533));
wire output_3_533, output_3_6, output_2_533;
mixer gate_output_2_533(.a(output_3_533), .b(output_3_6), .y(output_2_533));
wire output_4_533, output_4_6, output_3_533;
mixer gate_output_3_533(.a(output_4_533), .b(output_4_6), .y(output_3_533));
wire output_5_533, output_5_6, output_4_533;
mixer gate_output_4_533(.a(output_5_533), .b(output_5_6), .y(output_4_533));
wire output_6_533, output_6_6, output_5_533;
mixer gate_output_5_533(.a(output_6_533), .b(output_6_6), .y(output_5_533));
wire output_7_533, output_7_6, output_6_533;
mixer gate_output_6_533(.a(output_7_533), .b(output_7_6), .y(output_6_533));
wire output_8_533, output_8_6, output_7_533;
mixer gate_output_7_533(.a(output_8_533), .b(output_8_6), .y(output_7_533));
wire output_9_533, output_9_6, output_8_533;
mixer gate_output_8_533(.a(output_9_533), .b(output_9_6), .y(output_8_533));
wire output_10_533, output_10_6, output_9_533;
mixer gate_output_9_533(.a(output_10_533), .b(output_10_6), .y(output_9_533));
wire output_11_533, output_11_6, output_10_533;
mixer gate_output_10_533(.a(output_11_533), .b(output_11_6), .y(output_10_533));
wire output_12_533, output_12_6, output_11_533;
mixer gate_output_11_533(.a(output_12_533), .b(output_12_6), .y(output_11_533));
wire output_13_533, output_13_6, output_12_533;
mixer gate_output_12_533(.a(output_13_533), .b(output_13_6), .y(output_12_533));
wire output_14_533, output_14_6, output_13_533;
mixer gate_output_13_533(.a(output_14_533), .b(output_14_6), .y(output_13_533));
wire output_15_533, output_15_6, output_14_533;
mixer gate_output_14_533(.a(output_15_533), .b(output_15_6), .y(output_14_533));
wire output_16_533, output_16_6, output_15_533;
mixer gate_output_15_533(.a(output_16_533), .b(output_16_6), .y(output_15_533));
wire output_1_534, output_1_7, output_0_534;
mixer gate_output_0_534(.a(output_1_534), .b(output_1_7), .y(output_0_534));
wire output_2_534, output_2_7, output_1_534;
mixer gate_output_1_534(.a(output_2_534), .b(output_2_7), .y(output_1_534));
wire output_3_534, output_3_7, output_2_534;
mixer gate_output_2_534(.a(output_3_534), .b(output_3_7), .y(output_2_534));
wire output_4_534, output_4_7, output_3_534;
mixer gate_output_3_534(.a(output_4_534), .b(output_4_7), .y(output_3_534));
wire output_5_534, output_5_7, output_4_534;
mixer gate_output_4_534(.a(output_5_534), .b(output_5_7), .y(output_4_534));
wire output_6_534, output_6_7, output_5_534;
mixer gate_output_5_534(.a(output_6_534), .b(output_6_7), .y(output_5_534));
wire output_7_534, output_7_7, output_6_534;
mixer gate_output_6_534(.a(output_7_534), .b(output_7_7), .y(output_6_534));
wire output_8_534, output_8_7, output_7_534;
mixer gate_output_7_534(.a(output_8_534), .b(output_8_7), .y(output_7_534));
wire output_9_534, output_9_7, output_8_534;
mixer gate_output_8_534(.a(output_9_534), .b(output_9_7), .y(output_8_534));
wire output_10_534, output_10_7, output_9_534;
mixer gate_output_9_534(.a(output_10_534), .b(output_10_7), .y(output_9_534));
wire output_11_534, output_11_7, output_10_534;
mixer gate_output_10_534(.a(output_11_534), .b(output_11_7), .y(output_10_534));
wire output_12_534, output_12_7, output_11_534;
mixer gate_output_11_534(.a(output_12_534), .b(output_12_7), .y(output_11_534));
wire output_13_534, output_13_7, output_12_534;
mixer gate_output_12_534(.a(output_13_534), .b(output_13_7), .y(output_12_534));
wire output_14_534, output_14_7, output_13_534;
mixer gate_output_13_534(.a(output_14_534), .b(output_14_7), .y(output_13_534));
wire output_15_534, output_15_7, output_14_534;
mixer gate_output_14_534(.a(output_15_534), .b(output_15_7), .y(output_14_534));
wire output_16_534, output_16_7, output_15_534;
mixer gate_output_15_534(.a(output_16_534), .b(output_16_7), .y(output_15_534));
wire output_1_535, output_1_8, output_0_535;
mixer gate_output_0_535(.a(output_1_535), .b(output_1_8), .y(output_0_535));
wire output_2_535, output_2_8, output_1_535;
mixer gate_output_1_535(.a(output_2_535), .b(output_2_8), .y(output_1_535));
wire output_3_535, output_3_8, output_2_535;
mixer gate_output_2_535(.a(output_3_535), .b(output_3_8), .y(output_2_535));
wire output_4_535, output_4_8, output_3_535;
mixer gate_output_3_535(.a(output_4_535), .b(output_4_8), .y(output_3_535));
wire output_5_535, output_5_8, output_4_535;
mixer gate_output_4_535(.a(output_5_535), .b(output_5_8), .y(output_4_535));
wire output_6_535, output_6_8, output_5_535;
mixer gate_output_5_535(.a(output_6_535), .b(output_6_8), .y(output_5_535));
wire output_7_535, output_7_8, output_6_535;
mixer gate_output_6_535(.a(output_7_535), .b(output_7_8), .y(output_6_535));
wire output_8_535, output_8_8, output_7_535;
mixer gate_output_7_535(.a(output_8_535), .b(output_8_8), .y(output_7_535));
wire output_9_535, output_9_8, output_8_535;
mixer gate_output_8_535(.a(output_9_535), .b(output_9_8), .y(output_8_535));
wire output_10_535, output_10_8, output_9_535;
mixer gate_output_9_535(.a(output_10_535), .b(output_10_8), .y(output_9_535));
wire output_11_535, output_11_8, output_10_535;
mixer gate_output_10_535(.a(output_11_535), .b(output_11_8), .y(output_10_535));
wire output_12_535, output_12_8, output_11_535;
mixer gate_output_11_535(.a(output_12_535), .b(output_12_8), .y(output_11_535));
wire output_13_535, output_13_8, output_12_535;
mixer gate_output_12_535(.a(output_13_535), .b(output_13_8), .y(output_12_535));
wire output_14_535, output_14_8, output_13_535;
mixer gate_output_13_535(.a(output_14_535), .b(output_14_8), .y(output_13_535));
wire output_15_535, output_15_8, output_14_535;
mixer gate_output_14_535(.a(output_15_535), .b(output_15_8), .y(output_14_535));
wire output_16_535, output_16_8, output_15_535;
mixer gate_output_15_535(.a(output_16_535), .b(output_16_8), .y(output_15_535));
wire output_1_536, output_1_9, output_0_536;
mixer gate_output_0_536(.a(output_1_536), .b(output_1_9), .y(output_0_536));
wire output_2_536, output_2_9, output_1_536;
mixer gate_output_1_536(.a(output_2_536), .b(output_2_9), .y(output_1_536));
wire output_3_536, output_3_9, output_2_536;
mixer gate_output_2_536(.a(output_3_536), .b(output_3_9), .y(output_2_536));
wire output_4_536, output_4_9, output_3_536;
mixer gate_output_3_536(.a(output_4_536), .b(output_4_9), .y(output_3_536));
wire output_5_536, output_5_9, output_4_536;
mixer gate_output_4_536(.a(output_5_536), .b(output_5_9), .y(output_4_536));
wire output_6_536, output_6_9, output_5_536;
mixer gate_output_5_536(.a(output_6_536), .b(output_6_9), .y(output_5_536));
wire output_7_536, output_7_9, output_6_536;
mixer gate_output_6_536(.a(output_7_536), .b(output_7_9), .y(output_6_536));
wire output_8_536, output_8_9, output_7_536;
mixer gate_output_7_536(.a(output_8_536), .b(output_8_9), .y(output_7_536));
wire output_9_536, output_9_9, output_8_536;
mixer gate_output_8_536(.a(output_9_536), .b(output_9_9), .y(output_8_536));
wire output_10_536, output_10_9, output_9_536;
mixer gate_output_9_536(.a(output_10_536), .b(output_10_9), .y(output_9_536));
wire output_11_536, output_11_9, output_10_536;
mixer gate_output_10_536(.a(output_11_536), .b(output_11_9), .y(output_10_536));
wire output_12_536, output_12_9, output_11_536;
mixer gate_output_11_536(.a(output_12_536), .b(output_12_9), .y(output_11_536));
wire output_13_536, output_13_9, output_12_536;
mixer gate_output_12_536(.a(output_13_536), .b(output_13_9), .y(output_12_536));
wire output_14_536, output_14_9, output_13_536;
mixer gate_output_13_536(.a(output_14_536), .b(output_14_9), .y(output_13_536));
wire output_15_536, output_15_9, output_14_536;
mixer gate_output_14_536(.a(output_15_536), .b(output_15_9), .y(output_14_536));
wire output_16_536, output_16_9, output_15_536;
mixer gate_output_15_536(.a(output_16_536), .b(output_16_9), .y(output_15_536));
wire output_1_537, output_1_10, output_0_537;
mixer gate_output_0_537(.a(output_1_537), .b(output_1_10), .y(output_0_537));
wire output_2_537, output_2_10, output_1_537;
mixer gate_output_1_537(.a(output_2_537), .b(output_2_10), .y(output_1_537));
wire output_3_537, output_3_10, output_2_537;
mixer gate_output_2_537(.a(output_3_537), .b(output_3_10), .y(output_2_537));
wire output_4_537, output_4_10, output_3_537;
mixer gate_output_3_537(.a(output_4_537), .b(output_4_10), .y(output_3_537));
wire output_5_537, output_5_10, output_4_537;
mixer gate_output_4_537(.a(output_5_537), .b(output_5_10), .y(output_4_537));
wire output_6_537, output_6_10, output_5_537;
mixer gate_output_5_537(.a(output_6_537), .b(output_6_10), .y(output_5_537));
wire output_7_537, output_7_10, output_6_537;
mixer gate_output_6_537(.a(output_7_537), .b(output_7_10), .y(output_6_537));
wire output_8_537, output_8_10, output_7_537;
mixer gate_output_7_537(.a(output_8_537), .b(output_8_10), .y(output_7_537));
wire output_9_537, output_9_10, output_8_537;
mixer gate_output_8_537(.a(output_9_537), .b(output_9_10), .y(output_8_537));
wire output_10_537, output_10_10, output_9_537;
mixer gate_output_9_537(.a(output_10_537), .b(output_10_10), .y(output_9_537));
wire output_11_537, output_11_10, output_10_537;
mixer gate_output_10_537(.a(output_11_537), .b(output_11_10), .y(output_10_537));
wire output_12_537, output_12_10, output_11_537;
mixer gate_output_11_537(.a(output_12_537), .b(output_12_10), .y(output_11_537));
wire output_13_537, output_13_10, output_12_537;
mixer gate_output_12_537(.a(output_13_537), .b(output_13_10), .y(output_12_537));
wire output_14_537, output_14_10, output_13_537;
mixer gate_output_13_537(.a(output_14_537), .b(output_14_10), .y(output_13_537));
wire output_15_537, output_15_10, output_14_537;
mixer gate_output_14_537(.a(output_15_537), .b(output_15_10), .y(output_14_537));
wire output_16_537, output_16_10, output_15_537;
mixer gate_output_15_537(.a(output_16_537), .b(output_16_10), .y(output_15_537));
wire output_1_538, output_1_11, output_0_538;
mixer gate_output_0_538(.a(output_1_538), .b(output_1_11), .y(output_0_538));
wire output_2_538, output_2_11, output_1_538;
mixer gate_output_1_538(.a(output_2_538), .b(output_2_11), .y(output_1_538));
wire output_3_538, output_3_11, output_2_538;
mixer gate_output_2_538(.a(output_3_538), .b(output_3_11), .y(output_2_538));
wire output_4_538, output_4_11, output_3_538;
mixer gate_output_3_538(.a(output_4_538), .b(output_4_11), .y(output_3_538));
wire output_5_538, output_5_11, output_4_538;
mixer gate_output_4_538(.a(output_5_538), .b(output_5_11), .y(output_4_538));
wire output_6_538, output_6_11, output_5_538;
mixer gate_output_5_538(.a(output_6_538), .b(output_6_11), .y(output_5_538));
wire output_7_538, output_7_11, output_6_538;
mixer gate_output_6_538(.a(output_7_538), .b(output_7_11), .y(output_6_538));
wire output_8_538, output_8_11, output_7_538;
mixer gate_output_7_538(.a(output_8_538), .b(output_8_11), .y(output_7_538));
wire output_9_538, output_9_11, output_8_538;
mixer gate_output_8_538(.a(output_9_538), .b(output_9_11), .y(output_8_538));
wire output_10_538, output_10_11, output_9_538;
mixer gate_output_9_538(.a(output_10_538), .b(output_10_11), .y(output_9_538));
wire output_11_538, output_11_11, output_10_538;
mixer gate_output_10_538(.a(output_11_538), .b(output_11_11), .y(output_10_538));
wire output_12_538, output_12_11, output_11_538;
mixer gate_output_11_538(.a(output_12_538), .b(output_12_11), .y(output_11_538));
wire output_13_538, output_13_11, output_12_538;
mixer gate_output_12_538(.a(output_13_538), .b(output_13_11), .y(output_12_538));
wire output_14_538, output_14_11, output_13_538;
mixer gate_output_13_538(.a(output_14_538), .b(output_14_11), .y(output_13_538));
wire output_15_538, output_15_11, output_14_538;
mixer gate_output_14_538(.a(output_15_538), .b(output_15_11), .y(output_14_538));
wire output_16_538, output_16_11, output_15_538;
mixer gate_output_15_538(.a(output_16_538), .b(output_16_11), .y(output_15_538));
wire output_1_539, output_1_12, output_0_539;
mixer gate_output_0_539(.a(output_1_539), .b(output_1_12), .y(output_0_539));
wire output_2_539, output_2_12, output_1_539;
mixer gate_output_1_539(.a(output_2_539), .b(output_2_12), .y(output_1_539));
wire output_3_539, output_3_12, output_2_539;
mixer gate_output_2_539(.a(output_3_539), .b(output_3_12), .y(output_2_539));
wire output_4_539, output_4_12, output_3_539;
mixer gate_output_3_539(.a(output_4_539), .b(output_4_12), .y(output_3_539));
wire output_5_539, output_5_12, output_4_539;
mixer gate_output_4_539(.a(output_5_539), .b(output_5_12), .y(output_4_539));
wire output_6_539, output_6_12, output_5_539;
mixer gate_output_5_539(.a(output_6_539), .b(output_6_12), .y(output_5_539));
wire output_7_539, output_7_12, output_6_539;
mixer gate_output_6_539(.a(output_7_539), .b(output_7_12), .y(output_6_539));
wire output_8_539, output_8_12, output_7_539;
mixer gate_output_7_539(.a(output_8_539), .b(output_8_12), .y(output_7_539));
wire output_9_539, output_9_12, output_8_539;
mixer gate_output_8_539(.a(output_9_539), .b(output_9_12), .y(output_8_539));
wire output_10_539, output_10_12, output_9_539;
mixer gate_output_9_539(.a(output_10_539), .b(output_10_12), .y(output_9_539));
wire output_11_539, output_11_12, output_10_539;
mixer gate_output_10_539(.a(output_11_539), .b(output_11_12), .y(output_10_539));
wire output_12_539, output_12_12, output_11_539;
mixer gate_output_11_539(.a(output_12_539), .b(output_12_12), .y(output_11_539));
wire output_13_539, output_13_12, output_12_539;
mixer gate_output_12_539(.a(output_13_539), .b(output_13_12), .y(output_12_539));
wire output_14_539, output_14_12, output_13_539;
mixer gate_output_13_539(.a(output_14_539), .b(output_14_12), .y(output_13_539));
wire output_15_539, output_15_12, output_14_539;
mixer gate_output_14_539(.a(output_15_539), .b(output_15_12), .y(output_14_539));
wire output_16_539, output_16_12, output_15_539;
mixer gate_output_15_539(.a(output_16_539), .b(output_16_12), .y(output_15_539));
wire output_1_540, output_1_13, output_0_540;
mixer gate_output_0_540(.a(output_1_540), .b(output_1_13), .y(output_0_540));
wire output_2_540, output_2_13, output_1_540;
mixer gate_output_1_540(.a(output_2_540), .b(output_2_13), .y(output_1_540));
wire output_3_540, output_3_13, output_2_540;
mixer gate_output_2_540(.a(output_3_540), .b(output_3_13), .y(output_2_540));
wire output_4_540, output_4_13, output_3_540;
mixer gate_output_3_540(.a(output_4_540), .b(output_4_13), .y(output_3_540));
wire output_5_540, output_5_13, output_4_540;
mixer gate_output_4_540(.a(output_5_540), .b(output_5_13), .y(output_4_540));
wire output_6_540, output_6_13, output_5_540;
mixer gate_output_5_540(.a(output_6_540), .b(output_6_13), .y(output_5_540));
wire output_7_540, output_7_13, output_6_540;
mixer gate_output_6_540(.a(output_7_540), .b(output_7_13), .y(output_6_540));
wire output_8_540, output_8_13, output_7_540;
mixer gate_output_7_540(.a(output_8_540), .b(output_8_13), .y(output_7_540));
wire output_9_540, output_9_13, output_8_540;
mixer gate_output_8_540(.a(output_9_540), .b(output_9_13), .y(output_8_540));
wire output_10_540, output_10_13, output_9_540;
mixer gate_output_9_540(.a(output_10_540), .b(output_10_13), .y(output_9_540));
wire output_11_540, output_11_13, output_10_540;
mixer gate_output_10_540(.a(output_11_540), .b(output_11_13), .y(output_10_540));
wire output_12_540, output_12_13, output_11_540;
mixer gate_output_11_540(.a(output_12_540), .b(output_12_13), .y(output_11_540));
wire output_13_540, output_13_13, output_12_540;
mixer gate_output_12_540(.a(output_13_540), .b(output_13_13), .y(output_12_540));
wire output_14_540, output_14_13, output_13_540;
mixer gate_output_13_540(.a(output_14_540), .b(output_14_13), .y(output_13_540));
wire output_15_540, output_15_13, output_14_540;
mixer gate_output_14_540(.a(output_15_540), .b(output_15_13), .y(output_14_540));
wire output_16_540, output_16_13, output_15_540;
mixer gate_output_15_540(.a(output_16_540), .b(output_16_13), .y(output_15_540));
wire output_1_541, output_1_14, output_0_541;
mixer gate_output_0_541(.a(output_1_541), .b(output_1_14), .y(output_0_541));
wire output_2_541, output_2_14, output_1_541;
mixer gate_output_1_541(.a(output_2_541), .b(output_2_14), .y(output_1_541));
wire output_3_541, output_3_14, output_2_541;
mixer gate_output_2_541(.a(output_3_541), .b(output_3_14), .y(output_2_541));
wire output_4_541, output_4_14, output_3_541;
mixer gate_output_3_541(.a(output_4_541), .b(output_4_14), .y(output_3_541));
wire output_5_541, output_5_14, output_4_541;
mixer gate_output_4_541(.a(output_5_541), .b(output_5_14), .y(output_4_541));
wire output_6_541, output_6_14, output_5_541;
mixer gate_output_5_541(.a(output_6_541), .b(output_6_14), .y(output_5_541));
wire output_7_541, output_7_14, output_6_541;
mixer gate_output_6_541(.a(output_7_541), .b(output_7_14), .y(output_6_541));
wire output_8_541, output_8_14, output_7_541;
mixer gate_output_7_541(.a(output_8_541), .b(output_8_14), .y(output_7_541));
wire output_9_541, output_9_14, output_8_541;
mixer gate_output_8_541(.a(output_9_541), .b(output_9_14), .y(output_8_541));
wire output_10_541, output_10_14, output_9_541;
mixer gate_output_9_541(.a(output_10_541), .b(output_10_14), .y(output_9_541));
wire output_11_541, output_11_14, output_10_541;
mixer gate_output_10_541(.a(output_11_541), .b(output_11_14), .y(output_10_541));
wire output_12_541, output_12_14, output_11_541;
mixer gate_output_11_541(.a(output_12_541), .b(output_12_14), .y(output_11_541));
wire output_13_541, output_13_14, output_12_541;
mixer gate_output_12_541(.a(output_13_541), .b(output_13_14), .y(output_12_541));
wire output_14_541, output_14_14, output_13_541;
mixer gate_output_13_541(.a(output_14_541), .b(output_14_14), .y(output_13_541));
wire output_15_541, output_15_14, output_14_541;
mixer gate_output_14_541(.a(output_15_541), .b(output_15_14), .y(output_14_541));
wire output_16_541, output_16_14, output_15_541;
mixer gate_output_15_541(.a(output_16_541), .b(output_16_14), .y(output_15_541));
wire output_1_542, output_1_15, output_0_542;
mixer gate_output_0_542(.a(output_1_542), .b(output_1_15), .y(output_0_542));
wire output_2_542, output_2_15, output_1_542;
mixer gate_output_1_542(.a(output_2_542), .b(output_2_15), .y(output_1_542));
wire output_3_542, output_3_15, output_2_542;
mixer gate_output_2_542(.a(output_3_542), .b(output_3_15), .y(output_2_542));
wire output_4_542, output_4_15, output_3_542;
mixer gate_output_3_542(.a(output_4_542), .b(output_4_15), .y(output_3_542));
wire output_5_542, output_5_15, output_4_542;
mixer gate_output_4_542(.a(output_5_542), .b(output_5_15), .y(output_4_542));
wire output_6_542, output_6_15, output_5_542;
mixer gate_output_5_542(.a(output_6_542), .b(output_6_15), .y(output_5_542));
wire output_7_542, output_7_15, output_6_542;
mixer gate_output_6_542(.a(output_7_542), .b(output_7_15), .y(output_6_542));
wire output_8_542, output_8_15, output_7_542;
mixer gate_output_7_542(.a(output_8_542), .b(output_8_15), .y(output_7_542));
wire output_9_542, output_9_15, output_8_542;
mixer gate_output_8_542(.a(output_9_542), .b(output_9_15), .y(output_8_542));
wire output_10_542, output_10_15, output_9_542;
mixer gate_output_9_542(.a(output_10_542), .b(output_10_15), .y(output_9_542));
wire output_11_542, output_11_15, output_10_542;
mixer gate_output_10_542(.a(output_11_542), .b(output_11_15), .y(output_10_542));
wire output_12_542, output_12_15, output_11_542;
mixer gate_output_11_542(.a(output_12_542), .b(output_12_15), .y(output_11_542));
wire output_13_542, output_13_15, output_12_542;
mixer gate_output_12_542(.a(output_13_542), .b(output_13_15), .y(output_12_542));
wire output_14_542, output_14_15, output_13_542;
mixer gate_output_13_542(.a(output_14_542), .b(output_14_15), .y(output_13_542));
wire output_15_542, output_15_15, output_14_542;
mixer gate_output_14_542(.a(output_15_542), .b(output_15_15), .y(output_14_542));
wire output_16_542, output_16_15, output_15_542;
mixer gate_output_15_542(.a(output_16_542), .b(output_16_15), .y(output_15_542));
wire output_1_543, output_1_0, output_0_543;
mixer gate_output_0_543(.a(output_1_543), .b(output_1_0), .y(output_0_543));
wire output_2_543, output_2_0, output_1_543;
mixer gate_output_1_543(.a(output_2_543), .b(output_2_0), .y(output_1_543));
wire output_3_543, output_3_0, output_2_543;
mixer gate_output_2_543(.a(output_3_543), .b(output_3_0), .y(output_2_543));
wire output_4_543, output_4_0, output_3_543;
mixer gate_output_3_543(.a(output_4_543), .b(output_4_0), .y(output_3_543));
wire output_5_543, output_5_0, output_4_543;
mixer gate_output_4_543(.a(output_5_543), .b(output_5_0), .y(output_4_543));
wire output_6_543, output_6_0, output_5_543;
mixer gate_output_5_543(.a(output_6_543), .b(output_6_0), .y(output_5_543));
wire output_7_543, output_7_0, output_6_543;
mixer gate_output_6_543(.a(output_7_543), .b(output_7_0), .y(output_6_543));
wire output_8_543, output_8_0, output_7_543;
mixer gate_output_7_543(.a(output_8_543), .b(output_8_0), .y(output_7_543));
wire output_9_543, output_9_0, output_8_543;
mixer gate_output_8_543(.a(output_9_543), .b(output_9_0), .y(output_8_543));
wire output_10_543, output_10_0, output_9_543;
mixer gate_output_9_543(.a(output_10_543), .b(output_10_0), .y(output_9_543));
wire output_11_543, output_11_0, output_10_543;
mixer gate_output_10_543(.a(output_11_543), .b(output_11_0), .y(output_10_543));
wire output_12_543, output_12_0, output_11_543;
mixer gate_output_11_543(.a(output_12_543), .b(output_12_0), .y(output_11_543));
wire output_13_543, output_13_0, output_12_543;
mixer gate_output_12_543(.a(output_13_543), .b(output_13_0), .y(output_12_543));
wire output_14_543, output_14_0, output_13_543;
mixer gate_output_13_543(.a(output_14_543), .b(output_14_0), .y(output_13_543));
wire output_15_543, output_15_0, output_14_543;
mixer gate_output_14_543(.a(output_15_543), .b(output_15_0), .y(output_14_543));
wire output_16_543, output_16_0, output_15_543;
mixer gate_output_15_543(.a(output_16_543), .b(output_16_0), .y(output_15_543));
wire output_1_544, output_1_1, output_0_544;
mixer gate_output_0_544(.a(output_1_544), .b(output_1_1), .y(output_0_544));
wire output_2_544, output_2_1, output_1_544;
mixer gate_output_1_544(.a(output_2_544), .b(output_2_1), .y(output_1_544));
wire output_3_544, output_3_1, output_2_544;
mixer gate_output_2_544(.a(output_3_544), .b(output_3_1), .y(output_2_544));
wire output_4_544, output_4_1, output_3_544;
mixer gate_output_3_544(.a(output_4_544), .b(output_4_1), .y(output_3_544));
wire output_5_544, output_5_1, output_4_544;
mixer gate_output_4_544(.a(output_5_544), .b(output_5_1), .y(output_4_544));
wire output_6_544, output_6_1, output_5_544;
mixer gate_output_5_544(.a(output_6_544), .b(output_6_1), .y(output_5_544));
wire output_7_544, output_7_1, output_6_544;
mixer gate_output_6_544(.a(output_7_544), .b(output_7_1), .y(output_6_544));
wire output_8_544, output_8_1, output_7_544;
mixer gate_output_7_544(.a(output_8_544), .b(output_8_1), .y(output_7_544));
wire output_9_544, output_9_1, output_8_544;
mixer gate_output_8_544(.a(output_9_544), .b(output_9_1), .y(output_8_544));
wire output_10_544, output_10_1, output_9_544;
mixer gate_output_9_544(.a(output_10_544), .b(output_10_1), .y(output_9_544));
wire output_11_544, output_11_1, output_10_544;
mixer gate_output_10_544(.a(output_11_544), .b(output_11_1), .y(output_10_544));
wire output_12_544, output_12_1, output_11_544;
mixer gate_output_11_544(.a(output_12_544), .b(output_12_1), .y(output_11_544));
wire output_13_544, output_13_1, output_12_544;
mixer gate_output_12_544(.a(output_13_544), .b(output_13_1), .y(output_12_544));
wire output_14_544, output_14_1, output_13_544;
mixer gate_output_13_544(.a(output_14_544), .b(output_14_1), .y(output_13_544));
wire output_15_544, output_15_1, output_14_544;
mixer gate_output_14_544(.a(output_15_544), .b(output_15_1), .y(output_14_544));
wire output_16_544, output_16_1, output_15_544;
mixer gate_output_15_544(.a(output_16_544), .b(output_16_1), .y(output_15_544));
wire output_1_545, output_1_2, output_0_545;
mixer gate_output_0_545(.a(output_1_545), .b(output_1_2), .y(output_0_545));
wire output_2_545, output_2_2, output_1_545;
mixer gate_output_1_545(.a(output_2_545), .b(output_2_2), .y(output_1_545));
wire output_3_545, output_3_2, output_2_545;
mixer gate_output_2_545(.a(output_3_545), .b(output_3_2), .y(output_2_545));
wire output_4_545, output_4_2, output_3_545;
mixer gate_output_3_545(.a(output_4_545), .b(output_4_2), .y(output_3_545));
wire output_5_545, output_5_2, output_4_545;
mixer gate_output_4_545(.a(output_5_545), .b(output_5_2), .y(output_4_545));
wire output_6_545, output_6_2, output_5_545;
mixer gate_output_5_545(.a(output_6_545), .b(output_6_2), .y(output_5_545));
wire output_7_545, output_7_2, output_6_545;
mixer gate_output_6_545(.a(output_7_545), .b(output_7_2), .y(output_6_545));
wire output_8_545, output_8_2, output_7_545;
mixer gate_output_7_545(.a(output_8_545), .b(output_8_2), .y(output_7_545));
wire output_9_545, output_9_2, output_8_545;
mixer gate_output_8_545(.a(output_9_545), .b(output_9_2), .y(output_8_545));
wire output_10_545, output_10_2, output_9_545;
mixer gate_output_9_545(.a(output_10_545), .b(output_10_2), .y(output_9_545));
wire output_11_545, output_11_2, output_10_545;
mixer gate_output_10_545(.a(output_11_545), .b(output_11_2), .y(output_10_545));
wire output_12_545, output_12_2, output_11_545;
mixer gate_output_11_545(.a(output_12_545), .b(output_12_2), .y(output_11_545));
wire output_13_545, output_13_2, output_12_545;
mixer gate_output_12_545(.a(output_13_545), .b(output_13_2), .y(output_12_545));
wire output_14_545, output_14_2, output_13_545;
mixer gate_output_13_545(.a(output_14_545), .b(output_14_2), .y(output_13_545));
wire output_15_545, output_15_2, output_14_545;
mixer gate_output_14_545(.a(output_15_545), .b(output_15_2), .y(output_14_545));
wire output_16_545, output_16_2, output_15_545;
mixer gate_output_15_545(.a(output_16_545), .b(output_16_2), .y(output_15_545));
wire output_1_546, output_1_3, output_0_546;
mixer gate_output_0_546(.a(output_1_546), .b(output_1_3), .y(output_0_546));
wire output_2_546, output_2_3, output_1_546;
mixer gate_output_1_546(.a(output_2_546), .b(output_2_3), .y(output_1_546));
wire output_3_546, output_3_3, output_2_546;
mixer gate_output_2_546(.a(output_3_546), .b(output_3_3), .y(output_2_546));
wire output_4_546, output_4_3, output_3_546;
mixer gate_output_3_546(.a(output_4_546), .b(output_4_3), .y(output_3_546));
wire output_5_546, output_5_3, output_4_546;
mixer gate_output_4_546(.a(output_5_546), .b(output_5_3), .y(output_4_546));
wire output_6_546, output_6_3, output_5_546;
mixer gate_output_5_546(.a(output_6_546), .b(output_6_3), .y(output_5_546));
wire output_7_546, output_7_3, output_6_546;
mixer gate_output_6_546(.a(output_7_546), .b(output_7_3), .y(output_6_546));
wire output_8_546, output_8_3, output_7_546;
mixer gate_output_7_546(.a(output_8_546), .b(output_8_3), .y(output_7_546));
wire output_9_546, output_9_3, output_8_546;
mixer gate_output_8_546(.a(output_9_546), .b(output_9_3), .y(output_8_546));
wire output_10_546, output_10_3, output_9_546;
mixer gate_output_9_546(.a(output_10_546), .b(output_10_3), .y(output_9_546));
wire output_11_546, output_11_3, output_10_546;
mixer gate_output_10_546(.a(output_11_546), .b(output_11_3), .y(output_10_546));
wire output_12_546, output_12_3, output_11_546;
mixer gate_output_11_546(.a(output_12_546), .b(output_12_3), .y(output_11_546));
wire output_13_546, output_13_3, output_12_546;
mixer gate_output_12_546(.a(output_13_546), .b(output_13_3), .y(output_12_546));
wire output_14_546, output_14_3, output_13_546;
mixer gate_output_13_546(.a(output_14_546), .b(output_14_3), .y(output_13_546));
wire output_15_546, output_15_3, output_14_546;
mixer gate_output_14_546(.a(output_15_546), .b(output_15_3), .y(output_14_546));
wire output_16_546, output_16_3, output_15_546;
mixer gate_output_15_546(.a(output_16_546), .b(output_16_3), .y(output_15_546));
wire output_1_547, output_1_4, output_0_547;
mixer gate_output_0_547(.a(output_1_547), .b(output_1_4), .y(output_0_547));
wire output_2_547, output_2_4, output_1_547;
mixer gate_output_1_547(.a(output_2_547), .b(output_2_4), .y(output_1_547));
wire output_3_547, output_3_4, output_2_547;
mixer gate_output_2_547(.a(output_3_547), .b(output_3_4), .y(output_2_547));
wire output_4_547, output_4_4, output_3_547;
mixer gate_output_3_547(.a(output_4_547), .b(output_4_4), .y(output_3_547));
wire output_5_547, output_5_4, output_4_547;
mixer gate_output_4_547(.a(output_5_547), .b(output_5_4), .y(output_4_547));
wire output_6_547, output_6_4, output_5_547;
mixer gate_output_5_547(.a(output_6_547), .b(output_6_4), .y(output_5_547));
wire output_7_547, output_7_4, output_6_547;
mixer gate_output_6_547(.a(output_7_547), .b(output_7_4), .y(output_6_547));
wire output_8_547, output_8_4, output_7_547;
mixer gate_output_7_547(.a(output_8_547), .b(output_8_4), .y(output_7_547));
wire output_9_547, output_9_4, output_8_547;
mixer gate_output_8_547(.a(output_9_547), .b(output_9_4), .y(output_8_547));
wire output_10_547, output_10_4, output_9_547;
mixer gate_output_9_547(.a(output_10_547), .b(output_10_4), .y(output_9_547));
wire output_11_547, output_11_4, output_10_547;
mixer gate_output_10_547(.a(output_11_547), .b(output_11_4), .y(output_10_547));
wire output_12_547, output_12_4, output_11_547;
mixer gate_output_11_547(.a(output_12_547), .b(output_12_4), .y(output_11_547));
wire output_13_547, output_13_4, output_12_547;
mixer gate_output_12_547(.a(output_13_547), .b(output_13_4), .y(output_12_547));
wire output_14_547, output_14_4, output_13_547;
mixer gate_output_13_547(.a(output_14_547), .b(output_14_4), .y(output_13_547));
wire output_15_547, output_15_4, output_14_547;
mixer gate_output_14_547(.a(output_15_547), .b(output_15_4), .y(output_14_547));
wire output_16_547, output_16_4, output_15_547;
mixer gate_output_15_547(.a(output_16_547), .b(output_16_4), .y(output_15_547));
wire output_1_548, output_1_5, output_0_548;
mixer gate_output_0_548(.a(output_1_548), .b(output_1_5), .y(output_0_548));
wire output_2_548, output_2_5, output_1_548;
mixer gate_output_1_548(.a(output_2_548), .b(output_2_5), .y(output_1_548));
wire output_3_548, output_3_5, output_2_548;
mixer gate_output_2_548(.a(output_3_548), .b(output_3_5), .y(output_2_548));
wire output_4_548, output_4_5, output_3_548;
mixer gate_output_3_548(.a(output_4_548), .b(output_4_5), .y(output_3_548));
wire output_5_548, output_5_5, output_4_548;
mixer gate_output_4_548(.a(output_5_548), .b(output_5_5), .y(output_4_548));
wire output_6_548, output_6_5, output_5_548;
mixer gate_output_5_548(.a(output_6_548), .b(output_6_5), .y(output_5_548));
wire output_7_548, output_7_5, output_6_548;
mixer gate_output_6_548(.a(output_7_548), .b(output_7_5), .y(output_6_548));
wire output_8_548, output_8_5, output_7_548;
mixer gate_output_7_548(.a(output_8_548), .b(output_8_5), .y(output_7_548));
wire output_9_548, output_9_5, output_8_548;
mixer gate_output_8_548(.a(output_9_548), .b(output_9_5), .y(output_8_548));
wire output_10_548, output_10_5, output_9_548;
mixer gate_output_9_548(.a(output_10_548), .b(output_10_5), .y(output_9_548));
wire output_11_548, output_11_5, output_10_548;
mixer gate_output_10_548(.a(output_11_548), .b(output_11_5), .y(output_10_548));
wire output_12_548, output_12_5, output_11_548;
mixer gate_output_11_548(.a(output_12_548), .b(output_12_5), .y(output_11_548));
wire output_13_548, output_13_5, output_12_548;
mixer gate_output_12_548(.a(output_13_548), .b(output_13_5), .y(output_12_548));
wire output_14_548, output_14_5, output_13_548;
mixer gate_output_13_548(.a(output_14_548), .b(output_14_5), .y(output_13_548));
wire output_15_548, output_15_5, output_14_548;
mixer gate_output_14_548(.a(output_15_548), .b(output_15_5), .y(output_14_548));
wire output_16_548, output_16_5, output_15_548;
mixer gate_output_15_548(.a(output_16_548), .b(output_16_5), .y(output_15_548));
wire output_1_549, output_1_6, output_0_549;
mixer gate_output_0_549(.a(output_1_549), .b(output_1_6), .y(output_0_549));
wire output_2_549, output_2_6, output_1_549;
mixer gate_output_1_549(.a(output_2_549), .b(output_2_6), .y(output_1_549));
wire output_3_549, output_3_6, output_2_549;
mixer gate_output_2_549(.a(output_3_549), .b(output_3_6), .y(output_2_549));
wire output_4_549, output_4_6, output_3_549;
mixer gate_output_3_549(.a(output_4_549), .b(output_4_6), .y(output_3_549));
wire output_5_549, output_5_6, output_4_549;
mixer gate_output_4_549(.a(output_5_549), .b(output_5_6), .y(output_4_549));
wire output_6_549, output_6_6, output_5_549;
mixer gate_output_5_549(.a(output_6_549), .b(output_6_6), .y(output_5_549));
wire output_7_549, output_7_6, output_6_549;
mixer gate_output_6_549(.a(output_7_549), .b(output_7_6), .y(output_6_549));
wire output_8_549, output_8_6, output_7_549;
mixer gate_output_7_549(.a(output_8_549), .b(output_8_6), .y(output_7_549));
wire output_9_549, output_9_6, output_8_549;
mixer gate_output_8_549(.a(output_9_549), .b(output_9_6), .y(output_8_549));
wire output_10_549, output_10_6, output_9_549;
mixer gate_output_9_549(.a(output_10_549), .b(output_10_6), .y(output_9_549));
wire output_11_549, output_11_6, output_10_549;
mixer gate_output_10_549(.a(output_11_549), .b(output_11_6), .y(output_10_549));
wire output_12_549, output_12_6, output_11_549;
mixer gate_output_11_549(.a(output_12_549), .b(output_12_6), .y(output_11_549));
wire output_13_549, output_13_6, output_12_549;
mixer gate_output_12_549(.a(output_13_549), .b(output_13_6), .y(output_12_549));
wire output_14_549, output_14_6, output_13_549;
mixer gate_output_13_549(.a(output_14_549), .b(output_14_6), .y(output_13_549));
wire output_15_549, output_15_6, output_14_549;
mixer gate_output_14_549(.a(output_15_549), .b(output_15_6), .y(output_14_549));
wire output_16_549, output_16_6, output_15_549;
mixer gate_output_15_549(.a(output_16_549), .b(output_16_6), .y(output_15_549));
wire output_1_550, output_1_7, output_0_550;
mixer gate_output_0_550(.a(output_1_550), .b(output_1_7), .y(output_0_550));
wire output_2_550, output_2_7, output_1_550;
mixer gate_output_1_550(.a(output_2_550), .b(output_2_7), .y(output_1_550));
wire output_3_550, output_3_7, output_2_550;
mixer gate_output_2_550(.a(output_3_550), .b(output_3_7), .y(output_2_550));
wire output_4_550, output_4_7, output_3_550;
mixer gate_output_3_550(.a(output_4_550), .b(output_4_7), .y(output_3_550));
wire output_5_550, output_5_7, output_4_550;
mixer gate_output_4_550(.a(output_5_550), .b(output_5_7), .y(output_4_550));
wire output_6_550, output_6_7, output_5_550;
mixer gate_output_5_550(.a(output_6_550), .b(output_6_7), .y(output_5_550));
wire output_7_550, output_7_7, output_6_550;
mixer gate_output_6_550(.a(output_7_550), .b(output_7_7), .y(output_6_550));
wire output_8_550, output_8_7, output_7_550;
mixer gate_output_7_550(.a(output_8_550), .b(output_8_7), .y(output_7_550));
wire output_9_550, output_9_7, output_8_550;
mixer gate_output_8_550(.a(output_9_550), .b(output_9_7), .y(output_8_550));
wire output_10_550, output_10_7, output_9_550;
mixer gate_output_9_550(.a(output_10_550), .b(output_10_7), .y(output_9_550));
wire output_11_550, output_11_7, output_10_550;
mixer gate_output_10_550(.a(output_11_550), .b(output_11_7), .y(output_10_550));
wire output_12_550, output_12_7, output_11_550;
mixer gate_output_11_550(.a(output_12_550), .b(output_12_7), .y(output_11_550));
wire output_13_550, output_13_7, output_12_550;
mixer gate_output_12_550(.a(output_13_550), .b(output_13_7), .y(output_12_550));
wire output_14_550, output_14_7, output_13_550;
mixer gate_output_13_550(.a(output_14_550), .b(output_14_7), .y(output_13_550));
wire output_15_550, output_15_7, output_14_550;
mixer gate_output_14_550(.a(output_15_550), .b(output_15_7), .y(output_14_550));
wire output_16_550, output_16_7, output_15_550;
mixer gate_output_15_550(.a(output_16_550), .b(output_16_7), .y(output_15_550));
wire output_1_551, output_1_8, output_0_551;
mixer gate_output_0_551(.a(output_1_551), .b(output_1_8), .y(output_0_551));
wire output_2_551, output_2_8, output_1_551;
mixer gate_output_1_551(.a(output_2_551), .b(output_2_8), .y(output_1_551));
wire output_3_551, output_3_8, output_2_551;
mixer gate_output_2_551(.a(output_3_551), .b(output_3_8), .y(output_2_551));
wire output_4_551, output_4_8, output_3_551;
mixer gate_output_3_551(.a(output_4_551), .b(output_4_8), .y(output_3_551));
wire output_5_551, output_5_8, output_4_551;
mixer gate_output_4_551(.a(output_5_551), .b(output_5_8), .y(output_4_551));
wire output_6_551, output_6_8, output_5_551;
mixer gate_output_5_551(.a(output_6_551), .b(output_6_8), .y(output_5_551));
wire output_7_551, output_7_8, output_6_551;
mixer gate_output_6_551(.a(output_7_551), .b(output_7_8), .y(output_6_551));
wire output_8_551, output_8_8, output_7_551;
mixer gate_output_7_551(.a(output_8_551), .b(output_8_8), .y(output_7_551));
wire output_9_551, output_9_8, output_8_551;
mixer gate_output_8_551(.a(output_9_551), .b(output_9_8), .y(output_8_551));
wire output_10_551, output_10_8, output_9_551;
mixer gate_output_9_551(.a(output_10_551), .b(output_10_8), .y(output_9_551));
wire output_11_551, output_11_8, output_10_551;
mixer gate_output_10_551(.a(output_11_551), .b(output_11_8), .y(output_10_551));
wire output_12_551, output_12_8, output_11_551;
mixer gate_output_11_551(.a(output_12_551), .b(output_12_8), .y(output_11_551));
wire output_13_551, output_13_8, output_12_551;
mixer gate_output_12_551(.a(output_13_551), .b(output_13_8), .y(output_12_551));
wire output_14_551, output_14_8, output_13_551;
mixer gate_output_13_551(.a(output_14_551), .b(output_14_8), .y(output_13_551));
wire output_15_551, output_15_8, output_14_551;
mixer gate_output_14_551(.a(output_15_551), .b(output_15_8), .y(output_14_551));
wire output_16_551, output_16_8, output_15_551;
mixer gate_output_15_551(.a(output_16_551), .b(output_16_8), .y(output_15_551));
wire output_1_552, output_1_9, output_0_552;
mixer gate_output_0_552(.a(output_1_552), .b(output_1_9), .y(output_0_552));
wire output_2_552, output_2_9, output_1_552;
mixer gate_output_1_552(.a(output_2_552), .b(output_2_9), .y(output_1_552));
wire output_3_552, output_3_9, output_2_552;
mixer gate_output_2_552(.a(output_3_552), .b(output_3_9), .y(output_2_552));
wire output_4_552, output_4_9, output_3_552;
mixer gate_output_3_552(.a(output_4_552), .b(output_4_9), .y(output_3_552));
wire output_5_552, output_5_9, output_4_552;
mixer gate_output_4_552(.a(output_5_552), .b(output_5_9), .y(output_4_552));
wire output_6_552, output_6_9, output_5_552;
mixer gate_output_5_552(.a(output_6_552), .b(output_6_9), .y(output_5_552));
wire output_7_552, output_7_9, output_6_552;
mixer gate_output_6_552(.a(output_7_552), .b(output_7_9), .y(output_6_552));
wire output_8_552, output_8_9, output_7_552;
mixer gate_output_7_552(.a(output_8_552), .b(output_8_9), .y(output_7_552));
wire output_9_552, output_9_9, output_8_552;
mixer gate_output_8_552(.a(output_9_552), .b(output_9_9), .y(output_8_552));
wire output_10_552, output_10_9, output_9_552;
mixer gate_output_9_552(.a(output_10_552), .b(output_10_9), .y(output_9_552));
wire output_11_552, output_11_9, output_10_552;
mixer gate_output_10_552(.a(output_11_552), .b(output_11_9), .y(output_10_552));
wire output_12_552, output_12_9, output_11_552;
mixer gate_output_11_552(.a(output_12_552), .b(output_12_9), .y(output_11_552));
wire output_13_552, output_13_9, output_12_552;
mixer gate_output_12_552(.a(output_13_552), .b(output_13_9), .y(output_12_552));
wire output_14_552, output_14_9, output_13_552;
mixer gate_output_13_552(.a(output_14_552), .b(output_14_9), .y(output_13_552));
wire output_15_552, output_15_9, output_14_552;
mixer gate_output_14_552(.a(output_15_552), .b(output_15_9), .y(output_14_552));
wire output_16_552, output_16_9, output_15_552;
mixer gate_output_15_552(.a(output_16_552), .b(output_16_9), .y(output_15_552));
wire output_1_553, output_1_10, output_0_553;
mixer gate_output_0_553(.a(output_1_553), .b(output_1_10), .y(output_0_553));
wire output_2_553, output_2_10, output_1_553;
mixer gate_output_1_553(.a(output_2_553), .b(output_2_10), .y(output_1_553));
wire output_3_553, output_3_10, output_2_553;
mixer gate_output_2_553(.a(output_3_553), .b(output_3_10), .y(output_2_553));
wire output_4_553, output_4_10, output_3_553;
mixer gate_output_3_553(.a(output_4_553), .b(output_4_10), .y(output_3_553));
wire output_5_553, output_5_10, output_4_553;
mixer gate_output_4_553(.a(output_5_553), .b(output_5_10), .y(output_4_553));
wire output_6_553, output_6_10, output_5_553;
mixer gate_output_5_553(.a(output_6_553), .b(output_6_10), .y(output_5_553));
wire output_7_553, output_7_10, output_6_553;
mixer gate_output_6_553(.a(output_7_553), .b(output_7_10), .y(output_6_553));
wire output_8_553, output_8_10, output_7_553;
mixer gate_output_7_553(.a(output_8_553), .b(output_8_10), .y(output_7_553));
wire output_9_553, output_9_10, output_8_553;
mixer gate_output_8_553(.a(output_9_553), .b(output_9_10), .y(output_8_553));
wire output_10_553, output_10_10, output_9_553;
mixer gate_output_9_553(.a(output_10_553), .b(output_10_10), .y(output_9_553));
wire output_11_553, output_11_10, output_10_553;
mixer gate_output_10_553(.a(output_11_553), .b(output_11_10), .y(output_10_553));
wire output_12_553, output_12_10, output_11_553;
mixer gate_output_11_553(.a(output_12_553), .b(output_12_10), .y(output_11_553));
wire output_13_553, output_13_10, output_12_553;
mixer gate_output_12_553(.a(output_13_553), .b(output_13_10), .y(output_12_553));
wire output_14_553, output_14_10, output_13_553;
mixer gate_output_13_553(.a(output_14_553), .b(output_14_10), .y(output_13_553));
wire output_15_553, output_15_10, output_14_553;
mixer gate_output_14_553(.a(output_15_553), .b(output_15_10), .y(output_14_553));
wire output_16_553, output_16_10, output_15_553;
mixer gate_output_15_553(.a(output_16_553), .b(output_16_10), .y(output_15_553));
wire output_1_554, output_1_11, output_0_554;
mixer gate_output_0_554(.a(output_1_554), .b(output_1_11), .y(output_0_554));
wire output_2_554, output_2_11, output_1_554;
mixer gate_output_1_554(.a(output_2_554), .b(output_2_11), .y(output_1_554));
wire output_3_554, output_3_11, output_2_554;
mixer gate_output_2_554(.a(output_3_554), .b(output_3_11), .y(output_2_554));
wire output_4_554, output_4_11, output_3_554;
mixer gate_output_3_554(.a(output_4_554), .b(output_4_11), .y(output_3_554));
wire output_5_554, output_5_11, output_4_554;
mixer gate_output_4_554(.a(output_5_554), .b(output_5_11), .y(output_4_554));
wire output_6_554, output_6_11, output_5_554;
mixer gate_output_5_554(.a(output_6_554), .b(output_6_11), .y(output_5_554));
wire output_7_554, output_7_11, output_6_554;
mixer gate_output_6_554(.a(output_7_554), .b(output_7_11), .y(output_6_554));
wire output_8_554, output_8_11, output_7_554;
mixer gate_output_7_554(.a(output_8_554), .b(output_8_11), .y(output_7_554));
wire output_9_554, output_9_11, output_8_554;
mixer gate_output_8_554(.a(output_9_554), .b(output_9_11), .y(output_8_554));
wire output_10_554, output_10_11, output_9_554;
mixer gate_output_9_554(.a(output_10_554), .b(output_10_11), .y(output_9_554));
wire output_11_554, output_11_11, output_10_554;
mixer gate_output_10_554(.a(output_11_554), .b(output_11_11), .y(output_10_554));
wire output_12_554, output_12_11, output_11_554;
mixer gate_output_11_554(.a(output_12_554), .b(output_12_11), .y(output_11_554));
wire output_13_554, output_13_11, output_12_554;
mixer gate_output_12_554(.a(output_13_554), .b(output_13_11), .y(output_12_554));
wire output_14_554, output_14_11, output_13_554;
mixer gate_output_13_554(.a(output_14_554), .b(output_14_11), .y(output_13_554));
wire output_15_554, output_15_11, output_14_554;
mixer gate_output_14_554(.a(output_15_554), .b(output_15_11), .y(output_14_554));
wire output_16_554, output_16_11, output_15_554;
mixer gate_output_15_554(.a(output_16_554), .b(output_16_11), .y(output_15_554));
wire output_1_555, output_1_12, output_0_555;
mixer gate_output_0_555(.a(output_1_555), .b(output_1_12), .y(output_0_555));
wire output_2_555, output_2_12, output_1_555;
mixer gate_output_1_555(.a(output_2_555), .b(output_2_12), .y(output_1_555));
wire output_3_555, output_3_12, output_2_555;
mixer gate_output_2_555(.a(output_3_555), .b(output_3_12), .y(output_2_555));
wire output_4_555, output_4_12, output_3_555;
mixer gate_output_3_555(.a(output_4_555), .b(output_4_12), .y(output_3_555));
wire output_5_555, output_5_12, output_4_555;
mixer gate_output_4_555(.a(output_5_555), .b(output_5_12), .y(output_4_555));
wire output_6_555, output_6_12, output_5_555;
mixer gate_output_5_555(.a(output_6_555), .b(output_6_12), .y(output_5_555));
wire output_7_555, output_7_12, output_6_555;
mixer gate_output_6_555(.a(output_7_555), .b(output_7_12), .y(output_6_555));
wire output_8_555, output_8_12, output_7_555;
mixer gate_output_7_555(.a(output_8_555), .b(output_8_12), .y(output_7_555));
wire output_9_555, output_9_12, output_8_555;
mixer gate_output_8_555(.a(output_9_555), .b(output_9_12), .y(output_8_555));
wire output_10_555, output_10_12, output_9_555;
mixer gate_output_9_555(.a(output_10_555), .b(output_10_12), .y(output_9_555));
wire output_11_555, output_11_12, output_10_555;
mixer gate_output_10_555(.a(output_11_555), .b(output_11_12), .y(output_10_555));
wire output_12_555, output_12_12, output_11_555;
mixer gate_output_11_555(.a(output_12_555), .b(output_12_12), .y(output_11_555));
wire output_13_555, output_13_12, output_12_555;
mixer gate_output_12_555(.a(output_13_555), .b(output_13_12), .y(output_12_555));
wire output_14_555, output_14_12, output_13_555;
mixer gate_output_13_555(.a(output_14_555), .b(output_14_12), .y(output_13_555));
wire output_15_555, output_15_12, output_14_555;
mixer gate_output_14_555(.a(output_15_555), .b(output_15_12), .y(output_14_555));
wire output_16_555, output_16_12, output_15_555;
mixer gate_output_15_555(.a(output_16_555), .b(output_16_12), .y(output_15_555));
wire output_1_556, output_1_13, output_0_556;
mixer gate_output_0_556(.a(output_1_556), .b(output_1_13), .y(output_0_556));
wire output_2_556, output_2_13, output_1_556;
mixer gate_output_1_556(.a(output_2_556), .b(output_2_13), .y(output_1_556));
wire output_3_556, output_3_13, output_2_556;
mixer gate_output_2_556(.a(output_3_556), .b(output_3_13), .y(output_2_556));
wire output_4_556, output_4_13, output_3_556;
mixer gate_output_3_556(.a(output_4_556), .b(output_4_13), .y(output_3_556));
wire output_5_556, output_5_13, output_4_556;
mixer gate_output_4_556(.a(output_5_556), .b(output_5_13), .y(output_4_556));
wire output_6_556, output_6_13, output_5_556;
mixer gate_output_5_556(.a(output_6_556), .b(output_6_13), .y(output_5_556));
wire output_7_556, output_7_13, output_6_556;
mixer gate_output_6_556(.a(output_7_556), .b(output_7_13), .y(output_6_556));
wire output_8_556, output_8_13, output_7_556;
mixer gate_output_7_556(.a(output_8_556), .b(output_8_13), .y(output_7_556));
wire output_9_556, output_9_13, output_8_556;
mixer gate_output_8_556(.a(output_9_556), .b(output_9_13), .y(output_8_556));
wire output_10_556, output_10_13, output_9_556;
mixer gate_output_9_556(.a(output_10_556), .b(output_10_13), .y(output_9_556));
wire output_11_556, output_11_13, output_10_556;
mixer gate_output_10_556(.a(output_11_556), .b(output_11_13), .y(output_10_556));
wire output_12_556, output_12_13, output_11_556;
mixer gate_output_11_556(.a(output_12_556), .b(output_12_13), .y(output_11_556));
wire output_13_556, output_13_13, output_12_556;
mixer gate_output_12_556(.a(output_13_556), .b(output_13_13), .y(output_12_556));
wire output_14_556, output_14_13, output_13_556;
mixer gate_output_13_556(.a(output_14_556), .b(output_14_13), .y(output_13_556));
wire output_15_556, output_15_13, output_14_556;
mixer gate_output_14_556(.a(output_15_556), .b(output_15_13), .y(output_14_556));
wire output_16_556, output_16_13, output_15_556;
mixer gate_output_15_556(.a(output_16_556), .b(output_16_13), .y(output_15_556));
wire output_1_557, output_1_14, output_0_557;
mixer gate_output_0_557(.a(output_1_557), .b(output_1_14), .y(output_0_557));
wire output_2_557, output_2_14, output_1_557;
mixer gate_output_1_557(.a(output_2_557), .b(output_2_14), .y(output_1_557));
wire output_3_557, output_3_14, output_2_557;
mixer gate_output_2_557(.a(output_3_557), .b(output_3_14), .y(output_2_557));
wire output_4_557, output_4_14, output_3_557;
mixer gate_output_3_557(.a(output_4_557), .b(output_4_14), .y(output_3_557));
wire output_5_557, output_5_14, output_4_557;
mixer gate_output_4_557(.a(output_5_557), .b(output_5_14), .y(output_4_557));
wire output_6_557, output_6_14, output_5_557;
mixer gate_output_5_557(.a(output_6_557), .b(output_6_14), .y(output_5_557));
wire output_7_557, output_7_14, output_6_557;
mixer gate_output_6_557(.a(output_7_557), .b(output_7_14), .y(output_6_557));
wire output_8_557, output_8_14, output_7_557;
mixer gate_output_7_557(.a(output_8_557), .b(output_8_14), .y(output_7_557));
wire output_9_557, output_9_14, output_8_557;
mixer gate_output_8_557(.a(output_9_557), .b(output_9_14), .y(output_8_557));
wire output_10_557, output_10_14, output_9_557;
mixer gate_output_9_557(.a(output_10_557), .b(output_10_14), .y(output_9_557));
wire output_11_557, output_11_14, output_10_557;
mixer gate_output_10_557(.a(output_11_557), .b(output_11_14), .y(output_10_557));
wire output_12_557, output_12_14, output_11_557;
mixer gate_output_11_557(.a(output_12_557), .b(output_12_14), .y(output_11_557));
wire output_13_557, output_13_14, output_12_557;
mixer gate_output_12_557(.a(output_13_557), .b(output_13_14), .y(output_12_557));
wire output_14_557, output_14_14, output_13_557;
mixer gate_output_13_557(.a(output_14_557), .b(output_14_14), .y(output_13_557));
wire output_15_557, output_15_14, output_14_557;
mixer gate_output_14_557(.a(output_15_557), .b(output_15_14), .y(output_14_557));
wire output_16_557, output_16_14, output_15_557;
mixer gate_output_15_557(.a(output_16_557), .b(output_16_14), .y(output_15_557));
wire output_1_558, output_1_15, output_0_558;
mixer gate_output_0_558(.a(output_1_558), .b(output_1_15), .y(output_0_558));
wire output_2_558, output_2_15, output_1_558;
mixer gate_output_1_558(.a(output_2_558), .b(output_2_15), .y(output_1_558));
wire output_3_558, output_3_15, output_2_558;
mixer gate_output_2_558(.a(output_3_558), .b(output_3_15), .y(output_2_558));
wire output_4_558, output_4_15, output_3_558;
mixer gate_output_3_558(.a(output_4_558), .b(output_4_15), .y(output_3_558));
wire output_5_558, output_5_15, output_4_558;
mixer gate_output_4_558(.a(output_5_558), .b(output_5_15), .y(output_4_558));
wire output_6_558, output_6_15, output_5_558;
mixer gate_output_5_558(.a(output_6_558), .b(output_6_15), .y(output_5_558));
wire output_7_558, output_7_15, output_6_558;
mixer gate_output_6_558(.a(output_7_558), .b(output_7_15), .y(output_6_558));
wire output_8_558, output_8_15, output_7_558;
mixer gate_output_7_558(.a(output_8_558), .b(output_8_15), .y(output_7_558));
wire output_9_558, output_9_15, output_8_558;
mixer gate_output_8_558(.a(output_9_558), .b(output_9_15), .y(output_8_558));
wire output_10_558, output_10_15, output_9_558;
mixer gate_output_9_558(.a(output_10_558), .b(output_10_15), .y(output_9_558));
wire output_11_558, output_11_15, output_10_558;
mixer gate_output_10_558(.a(output_11_558), .b(output_11_15), .y(output_10_558));
wire output_12_558, output_12_15, output_11_558;
mixer gate_output_11_558(.a(output_12_558), .b(output_12_15), .y(output_11_558));
wire output_13_558, output_13_15, output_12_558;
mixer gate_output_12_558(.a(output_13_558), .b(output_13_15), .y(output_12_558));
wire output_14_558, output_14_15, output_13_558;
mixer gate_output_13_558(.a(output_14_558), .b(output_14_15), .y(output_13_558));
wire output_15_558, output_15_15, output_14_558;
mixer gate_output_14_558(.a(output_15_558), .b(output_15_15), .y(output_14_558));
wire output_16_558, output_16_15, output_15_558;
mixer gate_output_15_558(.a(output_16_558), .b(output_16_15), .y(output_15_558));
wire output_1_559, output_1_0, output_0_559;
mixer gate_output_0_559(.a(output_1_559), .b(output_1_0), .y(output_0_559));
wire output_2_559, output_2_0, output_1_559;
mixer gate_output_1_559(.a(output_2_559), .b(output_2_0), .y(output_1_559));
wire output_3_559, output_3_0, output_2_559;
mixer gate_output_2_559(.a(output_3_559), .b(output_3_0), .y(output_2_559));
wire output_4_559, output_4_0, output_3_559;
mixer gate_output_3_559(.a(output_4_559), .b(output_4_0), .y(output_3_559));
wire output_5_559, output_5_0, output_4_559;
mixer gate_output_4_559(.a(output_5_559), .b(output_5_0), .y(output_4_559));
wire output_6_559, output_6_0, output_5_559;
mixer gate_output_5_559(.a(output_6_559), .b(output_6_0), .y(output_5_559));
wire output_7_559, output_7_0, output_6_559;
mixer gate_output_6_559(.a(output_7_559), .b(output_7_0), .y(output_6_559));
wire output_8_559, output_8_0, output_7_559;
mixer gate_output_7_559(.a(output_8_559), .b(output_8_0), .y(output_7_559));
wire output_9_559, output_9_0, output_8_559;
mixer gate_output_8_559(.a(output_9_559), .b(output_9_0), .y(output_8_559));
wire output_10_559, output_10_0, output_9_559;
mixer gate_output_9_559(.a(output_10_559), .b(output_10_0), .y(output_9_559));
wire output_11_559, output_11_0, output_10_559;
mixer gate_output_10_559(.a(output_11_559), .b(output_11_0), .y(output_10_559));
wire output_12_559, output_12_0, output_11_559;
mixer gate_output_11_559(.a(output_12_559), .b(output_12_0), .y(output_11_559));
wire output_13_559, output_13_0, output_12_559;
mixer gate_output_12_559(.a(output_13_559), .b(output_13_0), .y(output_12_559));
wire output_14_559, output_14_0, output_13_559;
mixer gate_output_13_559(.a(output_14_559), .b(output_14_0), .y(output_13_559));
wire output_15_559, output_15_0, output_14_559;
mixer gate_output_14_559(.a(output_15_559), .b(output_15_0), .y(output_14_559));
wire output_16_559, output_16_0, output_15_559;
mixer gate_output_15_559(.a(output_16_559), .b(output_16_0), .y(output_15_559));
wire output_1_560, output_1_1, output_0_560;
mixer gate_output_0_560(.a(output_1_560), .b(output_1_1), .y(output_0_560));
wire output_2_560, output_2_1, output_1_560;
mixer gate_output_1_560(.a(output_2_560), .b(output_2_1), .y(output_1_560));
wire output_3_560, output_3_1, output_2_560;
mixer gate_output_2_560(.a(output_3_560), .b(output_3_1), .y(output_2_560));
wire output_4_560, output_4_1, output_3_560;
mixer gate_output_3_560(.a(output_4_560), .b(output_4_1), .y(output_3_560));
wire output_5_560, output_5_1, output_4_560;
mixer gate_output_4_560(.a(output_5_560), .b(output_5_1), .y(output_4_560));
wire output_6_560, output_6_1, output_5_560;
mixer gate_output_5_560(.a(output_6_560), .b(output_6_1), .y(output_5_560));
wire output_7_560, output_7_1, output_6_560;
mixer gate_output_6_560(.a(output_7_560), .b(output_7_1), .y(output_6_560));
wire output_8_560, output_8_1, output_7_560;
mixer gate_output_7_560(.a(output_8_560), .b(output_8_1), .y(output_7_560));
wire output_9_560, output_9_1, output_8_560;
mixer gate_output_8_560(.a(output_9_560), .b(output_9_1), .y(output_8_560));
wire output_10_560, output_10_1, output_9_560;
mixer gate_output_9_560(.a(output_10_560), .b(output_10_1), .y(output_9_560));
wire output_11_560, output_11_1, output_10_560;
mixer gate_output_10_560(.a(output_11_560), .b(output_11_1), .y(output_10_560));
wire output_12_560, output_12_1, output_11_560;
mixer gate_output_11_560(.a(output_12_560), .b(output_12_1), .y(output_11_560));
wire output_13_560, output_13_1, output_12_560;
mixer gate_output_12_560(.a(output_13_560), .b(output_13_1), .y(output_12_560));
wire output_14_560, output_14_1, output_13_560;
mixer gate_output_13_560(.a(output_14_560), .b(output_14_1), .y(output_13_560));
wire output_15_560, output_15_1, output_14_560;
mixer gate_output_14_560(.a(output_15_560), .b(output_15_1), .y(output_14_560));
wire output_16_560, output_16_1, output_15_560;
mixer gate_output_15_560(.a(output_16_560), .b(output_16_1), .y(output_15_560));
wire output_1_561, output_1_2, output_0_561;
mixer gate_output_0_561(.a(output_1_561), .b(output_1_2), .y(output_0_561));
wire output_2_561, output_2_2, output_1_561;
mixer gate_output_1_561(.a(output_2_561), .b(output_2_2), .y(output_1_561));
wire output_3_561, output_3_2, output_2_561;
mixer gate_output_2_561(.a(output_3_561), .b(output_3_2), .y(output_2_561));
wire output_4_561, output_4_2, output_3_561;
mixer gate_output_3_561(.a(output_4_561), .b(output_4_2), .y(output_3_561));
wire output_5_561, output_5_2, output_4_561;
mixer gate_output_4_561(.a(output_5_561), .b(output_5_2), .y(output_4_561));
wire output_6_561, output_6_2, output_5_561;
mixer gate_output_5_561(.a(output_6_561), .b(output_6_2), .y(output_5_561));
wire output_7_561, output_7_2, output_6_561;
mixer gate_output_6_561(.a(output_7_561), .b(output_7_2), .y(output_6_561));
wire output_8_561, output_8_2, output_7_561;
mixer gate_output_7_561(.a(output_8_561), .b(output_8_2), .y(output_7_561));
wire output_9_561, output_9_2, output_8_561;
mixer gate_output_8_561(.a(output_9_561), .b(output_9_2), .y(output_8_561));
wire output_10_561, output_10_2, output_9_561;
mixer gate_output_9_561(.a(output_10_561), .b(output_10_2), .y(output_9_561));
wire output_11_561, output_11_2, output_10_561;
mixer gate_output_10_561(.a(output_11_561), .b(output_11_2), .y(output_10_561));
wire output_12_561, output_12_2, output_11_561;
mixer gate_output_11_561(.a(output_12_561), .b(output_12_2), .y(output_11_561));
wire output_13_561, output_13_2, output_12_561;
mixer gate_output_12_561(.a(output_13_561), .b(output_13_2), .y(output_12_561));
wire output_14_561, output_14_2, output_13_561;
mixer gate_output_13_561(.a(output_14_561), .b(output_14_2), .y(output_13_561));
wire output_15_561, output_15_2, output_14_561;
mixer gate_output_14_561(.a(output_15_561), .b(output_15_2), .y(output_14_561));
wire output_16_561, output_16_2, output_15_561;
mixer gate_output_15_561(.a(output_16_561), .b(output_16_2), .y(output_15_561));
wire output_1_562, output_1_3, output_0_562;
mixer gate_output_0_562(.a(output_1_562), .b(output_1_3), .y(output_0_562));
wire output_2_562, output_2_3, output_1_562;
mixer gate_output_1_562(.a(output_2_562), .b(output_2_3), .y(output_1_562));
wire output_3_562, output_3_3, output_2_562;
mixer gate_output_2_562(.a(output_3_562), .b(output_3_3), .y(output_2_562));
wire output_4_562, output_4_3, output_3_562;
mixer gate_output_3_562(.a(output_4_562), .b(output_4_3), .y(output_3_562));
wire output_5_562, output_5_3, output_4_562;
mixer gate_output_4_562(.a(output_5_562), .b(output_5_3), .y(output_4_562));
wire output_6_562, output_6_3, output_5_562;
mixer gate_output_5_562(.a(output_6_562), .b(output_6_3), .y(output_5_562));
wire output_7_562, output_7_3, output_6_562;
mixer gate_output_6_562(.a(output_7_562), .b(output_7_3), .y(output_6_562));
wire output_8_562, output_8_3, output_7_562;
mixer gate_output_7_562(.a(output_8_562), .b(output_8_3), .y(output_7_562));
wire output_9_562, output_9_3, output_8_562;
mixer gate_output_8_562(.a(output_9_562), .b(output_9_3), .y(output_8_562));
wire output_10_562, output_10_3, output_9_562;
mixer gate_output_9_562(.a(output_10_562), .b(output_10_3), .y(output_9_562));
wire output_11_562, output_11_3, output_10_562;
mixer gate_output_10_562(.a(output_11_562), .b(output_11_3), .y(output_10_562));
wire output_12_562, output_12_3, output_11_562;
mixer gate_output_11_562(.a(output_12_562), .b(output_12_3), .y(output_11_562));
wire output_13_562, output_13_3, output_12_562;
mixer gate_output_12_562(.a(output_13_562), .b(output_13_3), .y(output_12_562));
wire output_14_562, output_14_3, output_13_562;
mixer gate_output_13_562(.a(output_14_562), .b(output_14_3), .y(output_13_562));
wire output_15_562, output_15_3, output_14_562;
mixer gate_output_14_562(.a(output_15_562), .b(output_15_3), .y(output_14_562));
wire output_16_562, output_16_3, output_15_562;
mixer gate_output_15_562(.a(output_16_562), .b(output_16_3), .y(output_15_562));
wire output_1_563, output_1_4, output_0_563;
mixer gate_output_0_563(.a(output_1_563), .b(output_1_4), .y(output_0_563));
wire output_2_563, output_2_4, output_1_563;
mixer gate_output_1_563(.a(output_2_563), .b(output_2_4), .y(output_1_563));
wire output_3_563, output_3_4, output_2_563;
mixer gate_output_2_563(.a(output_3_563), .b(output_3_4), .y(output_2_563));
wire output_4_563, output_4_4, output_3_563;
mixer gate_output_3_563(.a(output_4_563), .b(output_4_4), .y(output_3_563));
wire output_5_563, output_5_4, output_4_563;
mixer gate_output_4_563(.a(output_5_563), .b(output_5_4), .y(output_4_563));
wire output_6_563, output_6_4, output_5_563;
mixer gate_output_5_563(.a(output_6_563), .b(output_6_4), .y(output_5_563));
wire output_7_563, output_7_4, output_6_563;
mixer gate_output_6_563(.a(output_7_563), .b(output_7_4), .y(output_6_563));
wire output_8_563, output_8_4, output_7_563;
mixer gate_output_7_563(.a(output_8_563), .b(output_8_4), .y(output_7_563));
wire output_9_563, output_9_4, output_8_563;
mixer gate_output_8_563(.a(output_9_563), .b(output_9_4), .y(output_8_563));
wire output_10_563, output_10_4, output_9_563;
mixer gate_output_9_563(.a(output_10_563), .b(output_10_4), .y(output_9_563));
wire output_11_563, output_11_4, output_10_563;
mixer gate_output_10_563(.a(output_11_563), .b(output_11_4), .y(output_10_563));
wire output_12_563, output_12_4, output_11_563;
mixer gate_output_11_563(.a(output_12_563), .b(output_12_4), .y(output_11_563));
wire output_13_563, output_13_4, output_12_563;
mixer gate_output_12_563(.a(output_13_563), .b(output_13_4), .y(output_12_563));
wire output_14_563, output_14_4, output_13_563;
mixer gate_output_13_563(.a(output_14_563), .b(output_14_4), .y(output_13_563));
wire output_15_563, output_15_4, output_14_563;
mixer gate_output_14_563(.a(output_15_563), .b(output_15_4), .y(output_14_563));
wire output_16_563, output_16_4, output_15_563;
mixer gate_output_15_563(.a(output_16_563), .b(output_16_4), .y(output_15_563));
wire output_1_564, output_1_5, output_0_564;
mixer gate_output_0_564(.a(output_1_564), .b(output_1_5), .y(output_0_564));
wire output_2_564, output_2_5, output_1_564;
mixer gate_output_1_564(.a(output_2_564), .b(output_2_5), .y(output_1_564));
wire output_3_564, output_3_5, output_2_564;
mixer gate_output_2_564(.a(output_3_564), .b(output_3_5), .y(output_2_564));
wire output_4_564, output_4_5, output_3_564;
mixer gate_output_3_564(.a(output_4_564), .b(output_4_5), .y(output_3_564));
wire output_5_564, output_5_5, output_4_564;
mixer gate_output_4_564(.a(output_5_564), .b(output_5_5), .y(output_4_564));
wire output_6_564, output_6_5, output_5_564;
mixer gate_output_5_564(.a(output_6_564), .b(output_6_5), .y(output_5_564));
wire output_7_564, output_7_5, output_6_564;
mixer gate_output_6_564(.a(output_7_564), .b(output_7_5), .y(output_6_564));
wire output_8_564, output_8_5, output_7_564;
mixer gate_output_7_564(.a(output_8_564), .b(output_8_5), .y(output_7_564));
wire output_9_564, output_9_5, output_8_564;
mixer gate_output_8_564(.a(output_9_564), .b(output_9_5), .y(output_8_564));
wire output_10_564, output_10_5, output_9_564;
mixer gate_output_9_564(.a(output_10_564), .b(output_10_5), .y(output_9_564));
wire output_11_564, output_11_5, output_10_564;
mixer gate_output_10_564(.a(output_11_564), .b(output_11_5), .y(output_10_564));
wire output_12_564, output_12_5, output_11_564;
mixer gate_output_11_564(.a(output_12_564), .b(output_12_5), .y(output_11_564));
wire output_13_564, output_13_5, output_12_564;
mixer gate_output_12_564(.a(output_13_564), .b(output_13_5), .y(output_12_564));
wire output_14_564, output_14_5, output_13_564;
mixer gate_output_13_564(.a(output_14_564), .b(output_14_5), .y(output_13_564));
wire output_15_564, output_15_5, output_14_564;
mixer gate_output_14_564(.a(output_15_564), .b(output_15_5), .y(output_14_564));
wire output_16_564, output_16_5, output_15_564;
mixer gate_output_15_564(.a(output_16_564), .b(output_16_5), .y(output_15_564));
wire output_1_565, output_1_6, output_0_565;
mixer gate_output_0_565(.a(output_1_565), .b(output_1_6), .y(output_0_565));
wire output_2_565, output_2_6, output_1_565;
mixer gate_output_1_565(.a(output_2_565), .b(output_2_6), .y(output_1_565));
wire output_3_565, output_3_6, output_2_565;
mixer gate_output_2_565(.a(output_3_565), .b(output_3_6), .y(output_2_565));
wire output_4_565, output_4_6, output_3_565;
mixer gate_output_3_565(.a(output_4_565), .b(output_4_6), .y(output_3_565));
wire output_5_565, output_5_6, output_4_565;
mixer gate_output_4_565(.a(output_5_565), .b(output_5_6), .y(output_4_565));
wire output_6_565, output_6_6, output_5_565;
mixer gate_output_5_565(.a(output_6_565), .b(output_6_6), .y(output_5_565));
wire output_7_565, output_7_6, output_6_565;
mixer gate_output_6_565(.a(output_7_565), .b(output_7_6), .y(output_6_565));
wire output_8_565, output_8_6, output_7_565;
mixer gate_output_7_565(.a(output_8_565), .b(output_8_6), .y(output_7_565));
wire output_9_565, output_9_6, output_8_565;
mixer gate_output_8_565(.a(output_9_565), .b(output_9_6), .y(output_8_565));
wire output_10_565, output_10_6, output_9_565;
mixer gate_output_9_565(.a(output_10_565), .b(output_10_6), .y(output_9_565));
wire output_11_565, output_11_6, output_10_565;
mixer gate_output_10_565(.a(output_11_565), .b(output_11_6), .y(output_10_565));
wire output_12_565, output_12_6, output_11_565;
mixer gate_output_11_565(.a(output_12_565), .b(output_12_6), .y(output_11_565));
wire output_13_565, output_13_6, output_12_565;
mixer gate_output_12_565(.a(output_13_565), .b(output_13_6), .y(output_12_565));
wire output_14_565, output_14_6, output_13_565;
mixer gate_output_13_565(.a(output_14_565), .b(output_14_6), .y(output_13_565));
wire output_15_565, output_15_6, output_14_565;
mixer gate_output_14_565(.a(output_15_565), .b(output_15_6), .y(output_14_565));
wire output_16_565, output_16_6, output_15_565;
mixer gate_output_15_565(.a(output_16_565), .b(output_16_6), .y(output_15_565));
wire output_1_566, output_1_7, output_0_566;
mixer gate_output_0_566(.a(output_1_566), .b(output_1_7), .y(output_0_566));
wire output_2_566, output_2_7, output_1_566;
mixer gate_output_1_566(.a(output_2_566), .b(output_2_7), .y(output_1_566));
wire output_3_566, output_3_7, output_2_566;
mixer gate_output_2_566(.a(output_3_566), .b(output_3_7), .y(output_2_566));
wire output_4_566, output_4_7, output_3_566;
mixer gate_output_3_566(.a(output_4_566), .b(output_4_7), .y(output_3_566));
wire output_5_566, output_5_7, output_4_566;
mixer gate_output_4_566(.a(output_5_566), .b(output_5_7), .y(output_4_566));
wire output_6_566, output_6_7, output_5_566;
mixer gate_output_5_566(.a(output_6_566), .b(output_6_7), .y(output_5_566));
wire output_7_566, output_7_7, output_6_566;
mixer gate_output_6_566(.a(output_7_566), .b(output_7_7), .y(output_6_566));
wire output_8_566, output_8_7, output_7_566;
mixer gate_output_7_566(.a(output_8_566), .b(output_8_7), .y(output_7_566));
wire output_9_566, output_9_7, output_8_566;
mixer gate_output_8_566(.a(output_9_566), .b(output_9_7), .y(output_8_566));
wire output_10_566, output_10_7, output_9_566;
mixer gate_output_9_566(.a(output_10_566), .b(output_10_7), .y(output_9_566));
wire output_11_566, output_11_7, output_10_566;
mixer gate_output_10_566(.a(output_11_566), .b(output_11_7), .y(output_10_566));
wire output_12_566, output_12_7, output_11_566;
mixer gate_output_11_566(.a(output_12_566), .b(output_12_7), .y(output_11_566));
wire output_13_566, output_13_7, output_12_566;
mixer gate_output_12_566(.a(output_13_566), .b(output_13_7), .y(output_12_566));
wire output_14_566, output_14_7, output_13_566;
mixer gate_output_13_566(.a(output_14_566), .b(output_14_7), .y(output_13_566));
wire output_15_566, output_15_7, output_14_566;
mixer gate_output_14_566(.a(output_15_566), .b(output_15_7), .y(output_14_566));
wire output_16_566, output_16_7, output_15_566;
mixer gate_output_15_566(.a(output_16_566), .b(output_16_7), .y(output_15_566));
wire output_1_567, output_1_8, output_0_567;
mixer gate_output_0_567(.a(output_1_567), .b(output_1_8), .y(output_0_567));
wire output_2_567, output_2_8, output_1_567;
mixer gate_output_1_567(.a(output_2_567), .b(output_2_8), .y(output_1_567));
wire output_3_567, output_3_8, output_2_567;
mixer gate_output_2_567(.a(output_3_567), .b(output_3_8), .y(output_2_567));
wire output_4_567, output_4_8, output_3_567;
mixer gate_output_3_567(.a(output_4_567), .b(output_4_8), .y(output_3_567));
wire output_5_567, output_5_8, output_4_567;
mixer gate_output_4_567(.a(output_5_567), .b(output_5_8), .y(output_4_567));
wire output_6_567, output_6_8, output_5_567;
mixer gate_output_5_567(.a(output_6_567), .b(output_6_8), .y(output_5_567));
wire output_7_567, output_7_8, output_6_567;
mixer gate_output_6_567(.a(output_7_567), .b(output_7_8), .y(output_6_567));
wire output_8_567, output_8_8, output_7_567;
mixer gate_output_7_567(.a(output_8_567), .b(output_8_8), .y(output_7_567));
wire output_9_567, output_9_8, output_8_567;
mixer gate_output_8_567(.a(output_9_567), .b(output_9_8), .y(output_8_567));
wire output_10_567, output_10_8, output_9_567;
mixer gate_output_9_567(.a(output_10_567), .b(output_10_8), .y(output_9_567));
wire output_11_567, output_11_8, output_10_567;
mixer gate_output_10_567(.a(output_11_567), .b(output_11_8), .y(output_10_567));
wire output_12_567, output_12_8, output_11_567;
mixer gate_output_11_567(.a(output_12_567), .b(output_12_8), .y(output_11_567));
wire output_13_567, output_13_8, output_12_567;
mixer gate_output_12_567(.a(output_13_567), .b(output_13_8), .y(output_12_567));
wire output_14_567, output_14_8, output_13_567;
mixer gate_output_13_567(.a(output_14_567), .b(output_14_8), .y(output_13_567));
wire output_15_567, output_15_8, output_14_567;
mixer gate_output_14_567(.a(output_15_567), .b(output_15_8), .y(output_14_567));
wire output_16_567, output_16_8, output_15_567;
mixer gate_output_15_567(.a(output_16_567), .b(output_16_8), .y(output_15_567));
wire output_1_568, output_1_9, output_0_568;
mixer gate_output_0_568(.a(output_1_568), .b(output_1_9), .y(output_0_568));
wire output_2_568, output_2_9, output_1_568;
mixer gate_output_1_568(.a(output_2_568), .b(output_2_9), .y(output_1_568));
wire output_3_568, output_3_9, output_2_568;
mixer gate_output_2_568(.a(output_3_568), .b(output_3_9), .y(output_2_568));
wire output_4_568, output_4_9, output_3_568;
mixer gate_output_3_568(.a(output_4_568), .b(output_4_9), .y(output_3_568));
wire output_5_568, output_5_9, output_4_568;
mixer gate_output_4_568(.a(output_5_568), .b(output_5_9), .y(output_4_568));
wire output_6_568, output_6_9, output_5_568;
mixer gate_output_5_568(.a(output_6_568), .b(output_6_9), .y(output_5_568));
wire output_7_568, output_7_9, output_6_568;
mixer gate_output_6_568(.a(output_7_568), .b(output_7_9), .y(output_6_568));
wire output_8_568, output_8_9, output_7_568;
mixer gate_output_7_568(.a(output_8_568), .b(output_8_9), .y(output_7_568));
wire output_9_568, output_9_9, output_8_568;
mixer gate_output_8_568(.a(output_9_568), .b(output_9_9), .y(output_8_568));
wire output_10_568, output_10_9, output_9_568;
mixer gate_output_9_568(.a(output_10_568), .b(output_10_9), .y(output_9_568));
wire output_11_568, output_11_9, output_10_568;
mixer gate_output_10_568(.a(output_11_568), .b(output_11_9), .y(output_10_568));
wire output_12_568, output_12_9, output_11_568;
mixer gate_output_11_568(.a(output_12_568), .b(output_12_9), .y(output_11_568));
wire output_13_568, output_13_9, output_12_568;
mixer gate_output_12_568(.a(output_13_568), .b(output_13_9), .y(output_12_568));
wire output_14_568, output_14_9, output_13_568;
mixer gate_output_13_568(.a(output_14_568), .b(output_14_9), .y(output_13_568));
wire output_15_568, output_15_9, output_14_568;
mixer gate_output_14_568(.a(output_15_568), .b(output_15_9), .y(output_14_568));
wire output_16_568, output_16_9, output_15_568;
mixer gate_output_15_568(.a(output_16_568), .b(output_16_9), .y(output_15_568));
wire output_1_569, output_1_10, output_0_569;
mixer gate_output_0_569(.a(output_1_569), .b(output_1_10), .y(output_0_569));
wire output_2_569, output_2_10, output_1_569;
mixer gate_output_1_569(.a(output_2_569), .b(output_2_10), .y(output_1_569));
wire output_3_569, output_3_10, output_2_569;
mixer gate_output_2_569(.a(output_3_569), .b(output_3_10), .y(output_2_569));
wire output_4_569, output_4_10, output_3_569;
mixer gate_output_3_569(.a(output_4_569), .b(output_4_10), .y(output_3_569));
wire output_5_569, output_5_10, output_4_569;
mixer gate_output_4_569(.a(output_5_569), .b(output_5_10), .y(output_4_569));
wire output_6_569, output_6_10, output_5_569;
mixer gate_output_5_569(.a(output_6_569), .b(output_6_10), .y(output_5_569));
wire output_7_569, output_7_10, output_6_569;
mixer gate_output_6_569(.a(output_7_569), .b(output_7_10), .y(output_6_569));
wire output_8_569, output_8_10, output_7_569;
mixer gate_output_7_569(.a(output_8_569), .b(output_8_10), .y(output_7_569));
wire output_9_569, output_9_10, output_8_569;
mixer gate_output_8_569(.a(output_9_569), .b(output_9_10), .y(output_8_569));
wire output_10_569, output_10_10, output_9_569;
mixer gate_output_9_569(.a(output_10_569), .b(output_10_10), .y(output_9_569));
wire output_11_569, output_11_10, output_10_569;
mixer gate_output_10_569(.a(output_11_569), .b(output_11_10), .y(output_10_569));
wire output_12_569, output_12_10, output_11_569;
mixer gate_output_11_569(.a(output_12_569), .b(output_12_10), .y(output_11_569));
wire output_13_569, output_13_10, output_12_569;
mixer gate_output_12_569(.a(output_13_569), .b(output_13_10), .y(output_12_569));
wire output_14_569, output_14_10, output_13_569;
mixer gate_output_13_569(.a(output_14_569), .b(output_14_10), .y(output_13_569));
wire output_15_569, output_15_10, output_14_569;
mixer gate_output_14_569(.a(output_15_569), .b(output_15_10), .y(output_14_569));
wire output_16_569, output_16_10, output_15_569;
mixer gate_output_15_569(.a(output_16_569), .b(output_16_10), .y(output_15_569));
wire output_1_570, output_1_11, output_0_570;
mixer gate_output_0_570(.a(output_1_570), .b(output_1_11), .y(output_0_570));
wire output_2_570, output_2_11, output_1_570;
mixer gate_output_1_570(.a(output_2_570), .b(output_2_11), .y(output_1_570));
wire output_3_570, output_3_11, output_2_570;
mixer gate_output_2_570(.a(output_3_570), .b(output_3_11), .y(output_2_570));
wire output_4_570, output_4_11, output_3_570;
mixer gate_output_3_570(.a(output_4_570), .b(output_4_11), .y(output_3_570));
wire output_5_570, output_5_11, output_4_570;
mixer gate_output_4_570(.a(output_5_570), .b(output_5_11), .y(output_4_570));
wire output_6_570, output_6_11, output_5_570;
mixer gate_output_5_570(.a(output_6_570), .b(output_6_11), .y(output_5_570));
wire output_7_570, output_7_11, output_6_570;
mixer gate_output_6_570(.a(output_7_570), .b(output_7_11), .y(output_6_570));
wire output_8_570, output_8_11, output_7_570;
mixer gate_output_7_570(.a(output_8_570), .b(output_8_11), .y(output_7_570));
wire output_9_570, output_9_11, output_8_570;
mixer gate_output_8_570(.a(output_9_570), .b(output_9_11), .y(output_8_570));
wire output_10_570, output_10_11, output_9_570;
mixer gate_output_9_570(.a(output_10_570), .b(output_10_11), .y(output_9_570));
wire output_11_570, output_11_11, output_10_570;
mixer gate_output_10_570(.a(output_11_570), .b(output_11_11), .y(output_10_570));
wire output_12_570, output_12_11, output_11_570;
mixer gate_output_11_570(.a(output_12_570), .b(output_12_11), .y(output_11_570));
wire output_13_570, output_13_11, output_12_570;
mixer gate_output_12_570(.a(output_13_570), .b(output_13_11), .y(output_12_570));
wire output_14_570, output_14_11, output_13_570;
mixer gate_output_13_570(.a(output_14_570), .b(output_14_11), .y(output_13_570));
wire output_15_570, output_15_11, output_14_570;
mixer gate_output_14_570(.a(output_15_570), .b(output_15_11), .y(output_14_570));
wire output_16_570, output_16_11, output_15_570;
mixer gate_output_15_570(.a(output_16_570), .b(output_16_11), .y(output_15_570));
wire output_1_571, output_1_12, output_0_571;
mixer gate_output_0_571(.a(output_1_571), .b(output_1_12), .y(output_0_571));
wire output_2_571, output_2_12, output_1_571;
mixer gate_output_1_571(.a(output_2_571), .b(output_2_12), .y(output_1_571));
wire output_3_571, output_3_12, output_2_571;
mixer gate_output_2_571(.a(output_3_571), .b(output_3_12), .y(output_2_571));
wire output_4_571, output_4_12, output_3_571;
mixer gate_output_3_571(.a(output_4_571), .b(output_4_12), .y(output_3_571));
wire output_5_571, output_5_12, output_4_571;
mixer gate_output_4_571(.a(output_5_571), .b(output_5_12), .y(output_4_571));
wire output_6_571, output_6_12, output_5_571;
mixer gate_output_5_571(.a(output_6_571), .b(output_6_12), .y(output_5_571));
wire output_7_571, output_7_12, output_6_571;
mixer gate_output_6_571(.a(output_7_571), .b(output_7_12), .y(output_6_571));
wire output_8_571, output_8_12, output_7_571;
mixer gate_output_7_571(.a(output_8_571), .b(output_8_12), .y(output_7_571));
wire output_9_571, output_9_12, output_8_571;
mixer gate_output_8_571(.a(output_9_571), .b(output_9_12), .y(output_8_571));
wire output_10_571, output_10_12, output_9_571;
mixer gate_output_9_571(.a(output_10_571), .b(output_10_12), .y(output_9_571));
wire output_11_571, output_11_12, output_10_571;
mixer gate_output_10_571(.a(output_11_571), .b(output_11_12), .y(output_10_571));
wire output_12_571, output_12_12, output_11_571;
mixer gate_output_11_571(.a(output_12_571), .b(output_12_12), .y(output_11_571));
wire output_13_571, output_13_12, output_12_571;
mixer gate_output_12_571(.a(output_13_571), .b(output_13_12), .y(output_12_571));
wire output_14_571, output_14_12, output_13_571;
mixer gate_output_13_571(.a(output_14_571), .b(output_14_12), .y(output_13_571));
wire output_15_571, output_15_12, output_14_571;
mixer gate_output_14_571(.a(output_15_571), .b(output_15_12), .y(output_14_571));
wire output_16_571, output_16_12, output_15_571;
mixer gate_output_15_571(.a(output_16_571), .b(output_16_12), .y(output_15_571));
wire output_1_572, output_1_13, output_0_572;
mixer gate_output_0_572(.a(output_1_572), .b(output_1_13), .y(output_0_572));
wire output_2_572, output_2_13, output_1_572;
mixer gate_output_1_572(.a(output_2_572), .b(output_2_13), .y(output_1_572));
wire output_3_572, output_3_13, output_2_572;
mixer gate_output_2_572(.a(output_3_572), .b(output_3_13), .y(output_2_572));
wire output_4_572, output_4_13, output_3_572;
mixer gate_output_3_572(.a(output_4_572), .b(output_4_13), .y(output_3_572));
wire output_5_572, output_5_13, output_4_572;
mixer gate_output_4_572(.a(output_5_572), .b(output_5_13), .y(output_4_572));
wire output_6_572, output_6_13, output_5_572;
mixer gate_output_5_572(.a(output_6_572), .b(output_6_13), .y(output_5_572));
wire output_7_572, output_7_13, output_6_572;
mixer gate_output_6_572(.a(output_7_572), .b(output_7_13), .y(output_6_572));
wire output_8_572, output_8_13, output_7_572;
mixer gate_output_7_572(.a(output_8_572), .b(output_8_13), .y(output_7_572));
wire output_9_572, output_9_13, output_8_572;
mixer gate_output_8_572(.a(output_9_572), .b(output_9_13), .y(output_8_572));
wire output_10_572, output_10_13, output_9_572;
mixer gate_output_9_572(.a(output_10_572), .b(output_10_13), .y(output_9_572));
wire output_11_572, output_11_13, output_10_572;
mixer gate_output_10_572(.a(output_11_572), .b(output_11_13), .y(output_10_572));
wire output_12_572, output_12_13, output_11_572;
mixer gate_output_11_572(.a(output_12_572), .b(output_12_13), .y(output_11_572));
wire output_13_572, output_13_13, output_12_572;
mixer gate_output_12_572(.a(output_13_572), .b(output_13_13), .y(output_12_572));
wire output_14_572, output_14_13, output_13_572;
mixer gate_output_13_572(.a(output_14_572), .b(output_14_13), .y(output_13_572));
wire output_15_572, output_15_13, output_14_572;
mixer gate_output_14_572(.a(output_15_572), .b(output_15_13), .y(output_14_572));
wire output_16_572, output_16_13, output_15_572;
mixer gate_output_15_572(.a(output_16_572), .b(output_16_13), .y(output_15_572));
wire output_1_573, output_1_14, output_0_573;
mixer gate_output_0_573(.a(output_1_573), .b(output_1_14), .y(output_0_573));
wire output_2_573, output_2_14, output_1_573;
mixer gate_output_1_573(.a(output_2_573), .b(output_2_14), .y(output_1_573));
wire output_3_573, output_3_14, output_2_573;
mixer gate_output_2_573(.a(output_3_573), .b(output_3_14), .y(output_2_573));
wire output_4_573, output_4_14, output_3_573;
mixer gate_output_3_573(.a(output_4_573), .b(output_4_14), .y(output_3_573));
wire output_5_573, output_5_14, output_4_573;
mixer gate_output_4_573(.a(output_5_573), .b(output_5_14), .y(output_4_573));
wire output_6_573, output_6_14, output_5_573;
mixer gate_output_5_573(.a(output_6_573), .b(output_6_14), .y(output_5_573));
wire output_7_573, output_7_14, output_6_573;
mixer gate_output_6_573(.a(output_7_573), .b(output_7_14), .y(output_6_573));
wire output_8_573, output_8_14, output_7_573;
mixer gate_output_7_573(.a(output_8_573), .b(output_8_14), .y(output_7_573));
wire output_9_573, output_9_14, output_8_573;
mixer gate_output_8_573(.a(output_9_573), .b(output_9_14), .y(output_8_573));
wire output_10_573, output_10_14, output_9_573;
mixer gate_output_9_573(.a(output_10_573), .b(output_10_14), .y(output_9_573));
wire output_11_573, output_11_14, output_10_573;
mixer gate_output_10_573(.a(output_11_573), .b(output_11_14), .y(output_10_573));
wire output_12_573, output_12_14, output_11_573;
mixer gate_output_11_573(.a(output_12_573), .b(output_12_14), .y(output_11_573));
wire output_13_573, output_13_14, output_12_573;
mixer gate_output_12_573(.a(output_13_573), .b(output_13_14), .y(output_12_573));
wire output_14_573, output_14_14, output_13_573;
mixer gate_output_13_573(.a(output_14_573), .b(output_14_14), .y(output_13_573));
wire output_15_573, output_15_14, output_14_573;
mixer gate_output_14_573(.a(output_15_573), .b(output_15_14), .y(output_14_573));
wire output_16_573, output_16_14, output_15_573;
mixer gate_output_15_573(.a(output_16_573), .b(output_16_14), .y(output_15_573));
wire output_1_574, output_1_15, output_0_574;
mixer gate_output_0_574(.a(output_1_574), .b(output_1_15), .y(output_0_574));
wire output_2_574, output_2_15, output_1_574;
mixer gate_output_1_574(.a(output_2_574), .b(output_2_15), .y(output_1_574));
wire output_3_574, output_3_15, output_2_574;
mixer gate_output_2_574(.a(output_3_574), .b(output_3_15), .y(output_2_574));
wire output_4_574, output_4_15, output_3_574;
mixer gate_output_3_574(.a(output_4_574), .b(output_4_15), .y(output_3_574));
wire output_5_574, output_5_15, output_4_574;
mixer gate_output_4_574(.a(output_5_574), .b(output_5_15), .y(output_4_574));
wire output_6_574, output_6_15, output_5_574;
mixer gate_output_5_574(.a(output_6_574), .b(output_6_15), .y(output_5_574));
wire output_7_574, output_7_15, output_6_574;
mixer gate_output_6_574(.a(output_7_574), .b(output_7_15), .y(output_6_574));
wire output_8_574, output_8_15, output_7_574;
mixer gate_output_7_574(.a(output_8_574), .b(output_8_15), .y(output_7_574));
wire output_9_574, output_9_15, output_8_574;
mixer gate_output_8_574(.a(output_9_574), .b(output_9_15), .y(output_8_574));
wire output_10_574, output_10_15, output_9_574;
mixer gate_output_9_574(.a(output_10_574), .b(output_10_15), .y(output_9_574));
wire output_11_574, output_11_15, output_10_574;
mixer gate_output_10_574(.a(output_11_574), .b(output_11_15), .y(output_10_574));
wire output_12_574, output_12_15, output_11_574;
mixer gate_output_11_574(.a(output_12_574), .b(output_12_15), .y(output_11_574));
wire output_13_574, output_13_15, output_12_574;
mixer gate_output_12_574(.a(output_13_574), .b(output_13_15), .y(output_12_574));
wire output_14_574, output_14_15, output_13_574;
mixer gate_output_13_574(.a(output_14_574), .b(output_14_15), .y(output_13_574));
wire output_15_574, output_15_15, output_14_574;
mixer gate_output_14_574(.a(output_15_574), .b(output_15_15), .y(output_14_574));
wire output_16_574, output_16_15, output_15_574;
mixer gate_output_15_574(.a(output_16_574), .b(output_16_15), .y(output_15_574));
wire output_1_575, output_1_0, output_0_575;
mixer gate_output_0_575(.a(output_1_575), .b(output_1_0), .y(output_0_575));
wire output_2_575, output_2_0, output_1_575;
mixer gate_output_1_575(.a(output_2_575), .b(output_2_0), .y(output_1_575));
wire output_3_575, output_3_0, output_2_575;
mixer gate_output_2_575(.a(output_3_575), .b(output_3_0), .y(output_2_575));
wire output_4_575, output_4_0, output_3_575;
mixer gate_output_3_575(.a(output_4_575), .b(output_4_0), .y(output_3_575));
wire output_5_575, output_5_0, output_4_575;
mixer gate_output_4_575(.a(output_5_575), .b(output_5_0), .y(output_4_575));
wire output_6_575, output_6_0, output_5_575;
mixer gate_output_5_575(.a(output_6_575), .b(output_6_0), .y(output_5_575));
wire output_7_575, output_7_0, output_6_575;
mixer gate_output_6_575(.a(output_7_575), .b(output_7_0), .y(output_6_575));
wire output_8_575, output_8_0, output_7_575;
mixer gate_output_7_575(.a(output_8_575), .b(output_8_0), .y(output_7_575));
wire output_9_575, output_9_0, output_8_575;
mixer gate_output_8_575(.a(output_9_575), .b(output_9_0), .y(output_8_575));
wire output_10_575, output_10_0, output_9_575;
mixer gate_output_9_575(.a(output_10_575), .b(output_10_0), .y(output_9_575));
wire output_11_575, output_11_0, output_10_575;
mixer gate_output_10_575(.a(output_11_575), .b(output_11_0), .y(output_10_575));
wire output_12_575, output_12_0, output_11_575;
mixer gate_output_11_575(.a(output_12_575), .b(output_12_0), .y(output_11_575));
wire output_13_575, output_13_0, output_12_575;
mixer gate_output_12_575(.a(output_13_575), .b(output_13_0), .y(output_12_575));
wire output_14_575, output_14_0, output_13_575;
mixer gate_output_13_575(.a(output_14_575), .b(output_14_0), .y(output_13_575));
wire output_15_575, output_15_0, output_14_575;
mixer gate_output_14_575(.a(output_15_575), .b(output_15_0), .y(output_14_575));
wire output_16_575, output_16_0, output_15_575;
mixer gate_output_15_575(.a(output_16_575), .b(output_16_0), .y(output_15_575));
wire output_1_576, output_1_1, output_0_576;
mixer gate_output_0_576(.a(output_1_576), .b(output_1_1), .y(output_0_576));
wire output_2_576, output_2_1, output_1_576;
mixer gate_output_1_576(.a(output_2_576), .b(output_2_1), .y(output_1_576));
wire output_3_576, output_3_1, output_2_576;
mixer gate_output_2_576(.a(output_3_576), .b(output_3_1), .y(output_2_576));
wire output_4_576, output_4_1, output_3_576;
mixer gate_output_3_576(.a(output_4_576), .b(output_4_1), .y(output_3_576));
wire output_5_576, output_5_1, output_4_576;
mixer gate_output_4_576(.a(output_5_576), .b(output_5_1), .y(output_4_576));
wire output_6_576, output_6_1, output_5_576;
mixer gate_output_5_576(.a(output_6_576), .b(output_6_1), .y(output_5_576));
wire output_7_576, output_7_1, output_6_576;
mixer gate_output_6_576(.a(output_7_576), .b(output_7_1), .y(output_6_576));
wire output_8_576, output_8_1, output_7_576;
mixer gate_output_7_576(.a(output_8_576), .b(output_8_1), .y(output_7_576));
wire output_9_576, output_9_1, output_8_576;
mixer gate_output_8_576(.a(output_9_576), .b(output_9_1), .y(output_8_576));
wire output_10_576, output_10_1, output_9_576;
mixer gate_output_9_576(.a(output_10_576), .b(output_10_1), .y(output_9_576));
wire output_11_576, output_11_1, output_10_576;
mixer gate_output_10_576(.a(output_11_576), .b(output_11_1), .y(output_10_576));
wire output_12_576, output_12_1, output_11_576;
mixer gate_output_11_576(.a(output_12_576), .b(output_12_1), .y(output_11_576));
wire output_13_576, output_13_1, output_12_576;
mixer gate_output_12_576(.a(output_13_576), .b(output_13_1), .y(output_12_576));
wire output_14_576, output_14_1, output_13_576;
mixer gate_output_13_576(.a(output_14_576), .b(output_14_1), .y(output_13_576));
wire output_15_576, output_15_1, output_14_576;
mixer gate_output_14_576(.a(output_15_576), .b(output_15_1), .y(output_14_576));
wire output_16_576, output_16_1, output_15_576;
mixer gate_output_15_576(.a(output_16_576), .b(output_16_1), .y(output_15_576));
wire output_1_577, output_1_2, output_0_577;
mixer gate_output_0_577(.a(output_1_577), .b(output_1_2), .y(output_0_577));
wire output_2_577, output_2_2, output_1_577;
mixer gate_output_1_577(.a(output_2_577), .b(output_2_2), .y(output_1_577));
wire output_3_577, output_3_2, output_2_577;
mixer gate_output_2_577(.a(output_3_577), .b(output_3_2), .y(output_2_577));
wire output_4_577, output_4_2, output_3_577;
mixer gate_output_3_577(.a(output_4_577), .b(output_4_2), .y(output_3_577));
wire output_5_577, output_5_2, output_4_577;
mixer gate_output_4_577(.a(output_5_577), .b(output_5_2), .y(output_4_577));
wire output_6_577, output_6_2, output_5_577;
mixer gate_output_5_577(.a(output_6_577), .b(output_6_2), .y(output_5_577));
wire output_7_577, output_7_2, output_6_577;
mixer gate_output_6_577(.a(output_7_577), .b(output_7_2), .y(output_6_577));
wire output_8_577, output_8_2, output_7_577;
mixer gate_output_7_577(.a(output_8_577), .b(output_8_2), .y(output_7_577));
wire output_9_577, output_9_2, output_8_577;
mixer gate_output_8_577(.a(output_9_577), .b(output_9_2), .y(output_8_577));
wire output_10_577, output_10_2, output_9_577;
mixer gate_output_9_577(.a(output_10_577), .b(output_10_2), .y(output_9_577));
wire output_11_577, output_11_2, output_10_577;
mixer gate_output_10_577(.a(output_11_577), .b(output_11_2), .y(output_10_577));
wire output_12_577, output_12_2, output_11_577;
mixer gate_output_11_577(.a(output_12_577), .b(output_12_2), .y(output_11_577));
wire output_13_577, output_13_2, output_12_577;
mixer gate_output_12_577(.a(output_13_577), .b(output_13_2), .y(output_12_577));
wire output_14_577, output_14_2, output_13_577;
mixer gate_output_13_577(.a(output_14_577), .b(output_14_2), .y(output_13_577));
wire output_15_577, output_15_2, output_14_577;
mixer gate_output_14_577(.a(output_15_577), .b(output_15_2), .y(output_14_577));
wire output_16_577, output_16_2, output_15_577;
mixer gate_output_15_577(.a(output_16_577), .b(output_16_2), .y(output_15_577));
wire output_1_578, output_1_3, output_0_578;
mixer gate_output_0_578(.a(output_1_578), .b(output_1_3), .y(output_0_578));
wire output_2_578, output_2_3, output_1_578;
mixer gate_output_1_578(.a(output_2_578), .b(output_2_3), .y(output_1_578));
wire output_3_578, output_3_3, output_2_578;
mixer gate_output_2_578(.a(output_3_578), .b(output_3_3), .y(output_2_578));
wire output_4_578, output_4_3, output_3_578;
mixer gate_output_3_578(.a(output_4_578), .b(output_4_3), .y(output_3_578));
wire output_5_578, output_5_3, output_4_578;
mixer gate_output_4_578(.a(output_5_578), .b(output_5_3), .y(output_4_578));
wire output_6_578, output_6_3, output_5_578;
mixer gate_output_5_578(.a(output_6_578), .b(output_6_3), .y(output_5_578));
wire output_7_578, output_7_3, output_6_578;
mixer gate_output_6_578(.a(output_7_578), .b(output_7_3), .y(output_6_578));
wire output_8_578, output_8_3, output_7_578;
mixer gate_output_7_578(.a(output_8_578), .b(output_8_3), .y(output_7_578));
wire output_9_578, output_9_3, output_8_578;
mixer gate_output_8_578(.a(output_9_578), .b(output_9_3), .y(output_8_578));
wire output_10_578, output_10_3, output_9_578;
mixer gate_output_9_578(.a(output_10_578), .b(output_10_3), .y(output_9_578));
wire output_11_578, output_11_3, output_10_578;
mixer gate_output_10_578(.a(output_11_578), .b(output_11_3), .y(output_10_578));
wire output_12_578, output_12_3, output_11_578;
mixer gate_output_11_578(.a(output_12_578), .b(output_12_3), .y(output_11_578));
wire output_13_578, output_13_3, output_12_578;
mixer gate_output_12_578(.a(output_13_578), .b(output_13_3), .y(output_12_578));
wire output_14_578, output_14_3, output_13_578;
mixer gate_output_13_578(.a(output_14_578), .b(output_14_3), .y(output_13_578));
wire output_15_578, output_15_3, output_14_578;
mixer gate_output_14_578(.a(output_15_578), .b(output_15_3), .y(output_14_578));
wire output_16_578, output_16_3, output_15_578;
mixer gate_output_15_578(.a(output_16_578), .b(output_16_3), .y(output_15_578));
wire output_1_579, output_1_4, output_0_579;
mixer gate_output_0_579(.a(output_1_579), .b(output_1_4), .y(output_0_579));
wire output_2_579, output_2_4, output_1_579;
mixer gate_output_1_579(.a(output_2_579), .b(output_2_4), .y(output_1_579));
wire output_3_579, output_3_4, output_2_579;
mixer gate_output_2_579(.a(output_3_579), .b(output_3_4), .y(output_2_579));
wire output_4_579, output_4_4, output_3_579;
mixer gate_output_3_579(.a(output_4_579), .b(output_4_4), .y(output_3_579));
wire output_5_579, output_5_4, output_4_579;
mixer gate_output_4_579(.a(output_5_579), .b(output_5_4), .y(output_4_579));
wire output_6_579, output_6_4, output_5_579;
mixer gate_output_5_579(.a(output_6_579), .b(output_6_4), .y(output_5_579));
wire output_7_579, output_7_4, output_6_579;
mixer gate_output_6_579(.a(output_7_579), .b(output_7_4), .y(output_6_579));
wire output_8_579, output_8_4, output_7_579;
mixer gate_output_7_579(.a(output_8_579), .b(output_8_4), .y(output_7_579));
wire output_9_579, output_9_4, output_8_579;
mixer gate_output_8_579(.a(output_9_579), .b(output_9_4), .y(output_8_579));
wire output_10_579, output_10_4, output_9_579;
mixer gate_output_9_579(.a(output_10_579), .b(output_10_4), .y(output_9_579));
wire output_11_579, output_11_4, output_10_579;
mixer gate_output_10_579(.a(output_11_579), .b(output_11_4), .y(output_10_579));
wire output_12_579, output_12_4, output_11_579;
mixer gate_output_11_579(.a(output_12_579), .b(output_12_4), .y(output_11_579));
wire output_13_579, output_13_4, output_12_579;
mixer gate_output_12_579(.a(output_13_579), .b(output_13_4), .y(output_12_579));
wire output_14_579, output_14_4, output_13_579;
mixer gate_output_13_579(.a(output_14_579), .b(output_14_4), .y(output_13_579));
wire output_15_579, output_15_4, output_14_579;
mixer gate_output_14_579(.a(output_15_579), .b(output_15_4), .y(output_14_579));
wire output_16_579, output_16_4, output_15_579;
mixer gate_output_15_579(.a(output_16_579), .b(output_16_4), .y(output_15_579));
wire output_1_580, output_1_5, output_0_580;
mixer gate_output_0_580(.a(output_1_580), .b(output_1_5), .y(output_0_580));
wire output_2_580, output_2_5, output_1_580;
mixer gate_output_1_580(.a(output_2_580), .b(output_2_5), .y(output_1_580));
wire output_3_580, output_3_5, output_2_580;
mixer gate_output_2_580(.a(output_3_580), .b(output_3_5), .y(output_2_580));
wire output_4_580, output_4_5, output_3_580;
mixer gate_output_3_580(.a(output_4_580), .b(output_4_5), .y(output_3_580));
wire output_5_580, output_5_5, output_4_580;
mixer gate_output_4_580(.a(output_5_580), .b(output_5_5), .y(output_4_580));
wire output_6_580, output_6_5, output_5_580;
mixer gate_output_5_580(.a(output_6_580), .b(output_6_5), .y(output_5_580));
wire output_7_580, output_7_5, output_6_580;
mixer gate_output_6_580(.a(output_7_580), .b(output_7_5), .y(output_6_580));
wire output_8_580, output_8_5, output_7_580;
mixer gate_output_7_580(.a(output_8_580), .b(output_8_5), .y(output_7_580));
wire output_9_580, output_9_5, output_8_580;
mixer gate_output_8_580(.a(output_9_580), .b(output_9_5), .y(output_8_580));
wire output_10_580, output_10_5, output_9_580;
mixer gate_output_9_580(.a(output_10_580), .b(output_10_5), .y(output_9_580));
wire output_11_580, output_11_5, output_10_580;
mixer gate_output_10_580(.a(output_11_580), .b(output_11_5), .y(output_10_580));
wire output_12_580, output_12_5, output_11_580;
mixer gate_output_11_580(.a(output_12_580), .b(output_12_5), .y(output_11_580));
wire output_13_580, output_13_5, output_12_580;
mixer gate_output_12_580(.a(output_13_580), .b(output_13_5), .y(output_12_580));
wire output_14_580, output_14_5, output_13_580;
mixer gate_output_13_580(.a(output_14_580), .b(output_14_5), .y(output_13_580));
wire output_15_580, output_15_5, output_14_580;
mixer gate_output_14_580(.a(output_15_580), .b(output_15_5), .y(output_14_580));
wire output_16_580, output_16_5, output_15_580;
mixer gate_output_15_580(.a(output_16_580), .b(output_16_5), .y(output_15_580));
wire output_1_581, output_1_6, output_0_581;
mixer gate_output_0_581(.a(output_1_581), .b(output_1_6), .y(output_0_581));
wire output_2_581, output_2_6, output_1_581;
mixer gate_output_1_581(.a(output_2_581), .b(output_2_6), .y(output_1_581));
wire output_3_581, output_3_6, output_2_581;
mixer gate_output_2_581(.a(output_3_581), .b(output_3_6), .y(output_2_581));
wire output_4_581, output_4_6, output_3_581;
mixer gate_output_3_581(.a(output_4_581), .b(output_4_6), .y(output_3_581));
wire output_5_581, output_5_6, output_4_581;
mixer gate_output_4_581(.a(output_5_581), .b(output_5_6), .y(output_4_581));
wire output_6_581, output_6_6, output_5_581;
mixer gate_output_5_581(.a(output_6_581), .b(output_6_6), .y(output_5_581));
wire output_7_581, output_7_6, output_6_581;
mixer gate_output_6_581(.a(output_7_581), .b(output_7_6), .y(output_6_581));
wire output_8_581, output_8_6, output_7_581;
mixer gate_output_7_581(.a(output_8_581), .b(output_8_6), .y(output_7_581));
wire output_9_581, output_9_6, output_8_581;
mixer gate_output_8_581(.a(output_9_581), .b(output_9_6), .y(output_8_581));
wire output_10_581, output_10_6, output_9_581;
mixer gate_output_9_581(.a(output_10_581), .b(output_10_6), .y(output_9_581));
wire output_11_581, output_11_6, output_10_581;
mixer gate_output_10_581(.a(output_11_581), .b(output_11_6), .y(output_10_581));
wire output_12_581, output_12_6, output_11_581;
mixer gate_output_11_581(.a(output_12_581), .b(output_12_6), .y(output_11_581));
wire output_13_581, output_13_6, output_12_581;
mixer gate_output_12_581(.a(output_13_581), .b(output_13_6), .y(output_12_581));
wire output_14_581, output_14_6, output_13_581;
mixer gate_output_13_581(.a(output_14_581), .b(output_14_6), .y(output_13_581));
wire output_15_581, output_15_6, output_14_581;
mixer gate_output_14_581(.a(output_15_581), .b(output_15_6), .y(output_14_581));
wire output_16_581, output_16_6, output_15_581;
mixer gate_output_15_581(.a(output_16_581), .b(output_16_6), .y(output_15_581));
wire output_1_582, output_1_7, output_0_582;
mixer gate_output_0_582(.a(output_1_582), .b(output_1_7), .y(output_0_582));
wire output_2_582, output_2_7, output_1_582;
mixer gate_output_1_582(.a(output_2_582), .b(output_2_7), .y(output_1_582));
wire output_3_582, output_3_7, output_2_582;
mixer gate_output_2_582(.a(output_3_582), .b(output_3_7), .y(output_2_582));
wire output_4_582, output_4_7, output_3_582;
mixer gate_output_3_582(.a(output_4_582), .b(output_4_7), .y(output_3_582));
wire output_5_582, output_5_7, output_4_582;
mixer gate_output_4_582(.a(output_5_582), .b(output_5_7), .y(output_4_582));
wire output_6_582, output_6_7, output_5_582;
mixer gate_output_5_582(.a(output_6_582), .b(output_6_7), .y(output_5_582));
wire output_7_582, output_7_7, output_6_582;
mixer gate_output_6_582(.a(output_7_582), .b(output_7_7), .y(output_6_582));
wire output_8_582, output_8_7, output_7_582;
mixer gate_output_7_582(.a(output_8_582), .b(output_8_7), .y(output_7_582));
wire output_9_582, output_9_7, output_8_582;
mixer gate_output_8_582(.a(output_9_582), .b(output_9_7), .y(output_8_582));
wire output_10_582, output_10_7, output_9_582;
mixer gate_output_9_582(.a(output_10_582), .b(output_10_7), .y(output_9_582));
wire output_11_582, output_11_7, output_10_582;
mixer gate_output_10_582(.a(output_11_582), .b(output_11_7), .y(output_10_582));
wire output_12_582, output_12_7, output_11_582;
mixer gate_output_11_582(.a(output_12_582), .b(output_12_7), .y(output_11_582));
wire output_13_582, output_13_7, output_12_582;
mixer gate_output_12_582(.a(output_13_582), .b(output_13_7), .y(output_12_582));
wire output_14_582, output_14_7, output_13_582;
mixer gate_output_13_582(.a(output_14_582), .b(output_14_7), .y(output_13_582));
wire output_15_582, output_15_7, output_14_582;
mixer gate_output_14_582(.a(output_15_582), .b(output_15_7), .y(output_14_582));
wire output_16_582, output_16_7, output_15_582;
mixer gate_output_15_582(.a(output_16_582), .b(output_16_7), .y(output_15_582));
wire output_1_583, output_1_8, output_0_583;
mixer gate_output_0_583(.a(output_1_583), .b(output_1_8), .y(output_0_583));
wire output_2_583, output_2_8, output_1_583;
mixer gate_output_1_583(.a(output_2_583), .b(output_2_8), .y(output_1_583));
wire output_3_583, output_3_8, output_2_583;
mixer gate_output_2_583(.a(output_3_583), .b(output_3_8), .y(output_2_583));
wire output_4_583, output_4_8, output_3_583;
mixer gate_output_3_583(.a(output_4_583), .b(output_4_8), .y(output_3_583));
wire output_5_583, output_5_8, output_4_583;
mixer gate_output_4_583(.a(output_5_583), .b(output_5_8), .y(output_4_583));
wire output_6_583, output_6_8, output_5_583;
mixer gate_output_5_583(.a(output_6_583), .b(output_6_8), .y(output_5_583));
wire output_7_583, output_7_8, output_6_583;
mixer gate_output_6_583(.a(output_7_583), .b(output_7_8), .y(output_6_583));
wire output_8_583, output_8_8, output_7_583;
mixer gate_output_7_583(.a(output_8_583), .b(output_8_8), .y(output_7_583));
wire output_9_583, output_9_8, output_8_583;
mixer gate_output_8_583(.a(output_9_583), .b(output_9_8), .y(output_8_583));
wire output_10_583, output_10_8, output_9_583;
mixer gate_output_9_583(.a(output_10_583), .b(output_10_8), .y(output_9_583));
wire output_11_583, output_11_8, output_10_583;
mixer gate_output_10_583(.a(output_11_583), .b(output_11_8), .y(output_10_583));
wire output_12_583, output_12_8, output_11_583;
mixer gate_output_11_583(.a(output_12_583), .b(output_12_8), .y(output_11_583));
wire output_13_583, output_13_8, output_12_583;
mixer gate_output_12_583(.a(output_13_583), .b(output_13_8), .y(output_12_583));
wire output_14_583, output_14_8, output_13_583;
mixer gate_output_13_583(.a(output_14_583), .b(output_14_8), .y(output_13_583));
wire output_15_583, output_15_8, output_14_583;
mixer gate_output_14_583(.a(output_15_583), .b(output_15_8), .y(output_14_583));
wire output_16_583, output_16_8, output_15_583;
mixer gate_output_15_583(.a(output_16_583), .b(output_16_8), .y(output_15_583));
wire output_1_584, output_1_9, output_0_584;
mixer gate_output_0_584(.a(output_1_584), .b(output_1_9), .y(output_0_584));
wire output_2_584, output_2_9, output_1_584;
mixer gate_output_1_584(.a(output_2_584), .b(output_2_9), .y(output_1_584));
wire output_3_584, output_3_9, output_2_584;
mixer gate_output_2_584(.a(output_3_584), .b(output_3_9), .y(output_2_584));
wire output_4_584, output_4_9, output_3_584;
mixer gate_output_3_584(.a(output_4_584), .b(output_4_9), .y(output_3_584));
wire output_5_584, output_5_9, output_4_584;
mixer gate_output_4_584(.a(output_5_584), .b(output_5_9), .y(output_4_584));
wire output_6_584, output_6_9, output_5_584;
mixer gate_output_5_584(.a(output_6_584), .b(output_6_9), .y(output_5_584));
wire output_7_584, output_7_9, output_6_584;
mixer gate_output_6_584(.a(output_7_584), .b(output_7_9), .y(output_6_584));
wire output_8_584, output_8_9, output_7_584;
mixer gate_output_7_584(.a(output_8_584), .b(output_8_9), .y(output_7_584));
wire output_9_584, output_9_9, output_8_584;
mixer gate_output_8_584(.a(output_9_584), .b(output_9_9), .y(output_8_584));
wire output_10_584, output_10_9, output_9_584;
mixer gate_output_9_584(.a(output_10_584), .b(output_10_9), .y(output_9_584));
wire output_11_584, output_11_9, output_10_584;
mixer gate_output_10_584(.a(output_11_584), .b(output_11_9), .y(output_10_584));
wire output_12_584, output_12_9, output_11_584;
mixer gate_output_11_584(.a(output_12_584), .b(output_12_9), .y(output_11_584));
wire output_13_584, output_13_9, output_12_584;
mixer gate_output_12_584(.a(output_13_584), .b(output_13_9), .y(output_12_584));
wire output_14_584, output_14_9, output_13_584;
mixer gate_output_13_584(.a(output_14_584), .b(output_14_9), .y(output_13_584));
wire output_15_584, output_15_9, output_14_584;
mixer gate_output_14_584(.a(output_15_584), .b(output_15_9), .y(output_14_584));
wire output_16_584, output_16_9, output_15_584;
mixer gate_output_15_584(.a(output_16_584), .b(output_16_9), .y(output_15_584));
wire output_1_585, output_1_10, output_0_585;
mixer gate_output_0_585(.a(output_1_585), .b(output_1_10), .y(output_0_585));
wire output_2_585, output_2_10, output_1_585;
mixer gate_output_1_585(.a(output_2_585), .b(output_2_10), .y(output_1_585));
wire output_3_585, output_3_10, output_2_585;
mixer gate_output_2_585(.a(output_3_585), .b(output_3_10), .y(output_2_585));
wire output_4_585, output_4_10, output_3_585;
mixer gate_output_3_585(.a(output_4_585), .b(output_4_10), .y(output_3_585));
wire output_5_585, output_5_10, output_4_585;
mixer gate_output_4_585(.a(output_5_585), .b(output_5_10), .y(output_4_585));
wire output_6_585, output_6_10, output_5_585;
mixer gate_output_5_585(.a(output_6_585), .b(output_6_10), .y(output_5_585));
wire output_7_585, output_7_10, output_6_585;
mixer gate_output_6_585(.a(output_7_585), .b(output_7_10), .y(output_6_585));
wire output_8_585, output_8_10, output_7_585;
mixer gate_output_7_585(.a(output_8_585), .b(output_8_10), .y(output_7_585));
wire output_9_585, output_9_10, output_8_585;
mixer gate_output_8_585(.a(output_9_585), .b(output_9_10), .y(output_8_585));
wire output_10_585, output_10_10, output_9_585;
mixer gate_output_9_585(.a(output_10_585), .b(output_10_10), .y(output_9_585));
wire output_11_585, output_11_10, output_10_585;
mixer gate_output_10_585(.a(output_11_585), .b(output_11_10), .y(output_10_585));
wire output_12_585, output_12_10, output_11_585;
mixer gate_output_11_585(.a(output_12_585), .b(output_12_10), .y(output_11_585));
wire output_13_585, output_13_10, output_12_585;
mixer gate_output_12_585(.a(output_13_585), .b(output_13_10), .y(output_12_585));
wire output_14_585, output_14_10, output_13_585;
mixer gate_output_13_585(.a(output_14_585), .b(output_14_10), .y(output_13_585));
wire output_15_585, output_15_10, output_14_585;
mixer gate_output_14_585(.a(output_15_585), .b(output_15_10), .y(output_14_585));
wire output_16_585, output_16_10, output_15_585;
mixer gate_output_15_585(.a(output_16_585), .b(output_16_10), .y(output_15_585));
wire output_1_586, output_1_11, output_0_586;
mixer gate_output_0_586(.a(output_1_586), .b(output_1_11), .y(output_0_586));
wire output_2_586, output_2_11, output_1_586;
mixer gate_output_1_586(.a(output_2_586), .b(output_2_11), .y(output_1_586));
wire output_3_586, output_3_11, output_2_586;
mixer gate_output_2_586(.a(output_3_586), .b(output_3_11), .y(output_2_586));
wire output_4_586, output_4_11, output_3_586;
mixer gate_output_3_586(.a(output_4_586), .b(output_4_11), .y(output_3_586));
wire output_5_586, output_5_11, output_4_586;
mixer gate_output_4_586(.a(output_5_586), .b(output_5_11), .y(output_4_586));
wire output_6_586, output_6_11, output_5_586;
mixer gate_output_5_586(.a(output_6_586), .b(output_6_11), .y(output_5_586));
wire output_7_586, output_7_11, output_6_586;
mixer gate_output_6_586(.a(output_7_586), .b(output_7_11), .y(output_6_586));
wire output_8_586, output_8_11, output_7_586;
mixer gate_output_7_586(.a(output_8_586), .b(output_8_11), .y(output_7_586));
wire output_9_586, output_9_11, output_8_586;
mixer gate_output_8_586(.a(output_9_586), .b(output_9_11), .y(output_8_586));
wire output_10_586, output_10_11, output_9_586;
mixer gate_output_9_586(.a(output_10_586), .b(output_10_11), .y(output_9_586));
wire output_11_586, output_11_11, output_10_586;
mixer gate_output_10_586(.a(output_11_586), .b(output_11_11), .y(output_10_586));
wire output_12_586, output_12_11, output_11_586;
mixer gate_output_11_586(.a(output_12_586), .b(output_12_11), .y(output_11_586));
wire output_13_586, output_13_11, output_12_586;
mixer gate_output_12_586(.a(output_13_586), .b(output_13_11), .y(output_12_586));
wire output_14_586, output_14_11, output_13_586;
mixer gate_output_13_586(.a(output_14_586), .b(output_14_11), .y(output_13_586));
wire output_15_586, output_15_11, output_14_586;
mixer gate_output_14_586(.a(output_15_586), .b(output_15_11), .y(output_14_586));
wire output_16_586, output_16_11, output_15_586;
mixer gate_output_15_586(.a(output_16_586), .b(output_16_11), .y(output_15_586));
wire output_1_587, output_1_12, output_0_587;
mixer gate_output_0_587(.a(output_1_587), .b(output_1_12), .y(output_0_587));
wire output_2_587, output_2_12, output_1_587;
mixer gate_output_1_587(.a(output_2_587), .b(output_2_12), .y(output_1_587));
wire output_3_587, output_3_12, output_2_587;
mixer gate_output_2_587(.a(output_3_587), .b(output_3_12), .y(output_2_587));
wire output_4_587, output_4_12, output_3_587;
mixer gate_output_3_587(.a(output_4_587), .b(output_4_12), .y(output_3_587));
wire output_5_587, output_5_12, output_4_587;
mixer gate_output_4_587(.a(output_5_587), .b(output_5_12), .y(output_4_587));
wire output_6_587, output_6_12, output_5_587;
mixer gate_output_5_587(.a(output_6_587), .b(output_6_12), .y(output_5_587));
wire output_7_587, output_7_12, output_6_587;
mixer gate_output_6_587(.a(output_7_587), .b(output_7_12), .y(output_6_587));
wire output_8_587, output_8_12, output_7_587;
mixer gate_output_7_587(.a(output_8_587), .b(output_8_12), .y(output_7_587));
wire output_9_587, output_9_12, output_8_587;
mixer gate_output_8_587(.a(output_9_587), .b(output_9_12), .y(output_8_587));
wire output_10_587, output_10_12, output_9_587;
mixer gate_output_9_587(.a(output_10_587), .b(output_10_12), .y(output_9_587));
wire output_11_587, output_11_12, output_10_587;
mixer gate_output_10_587(.a(output_11_587), .b(output_11_12), .y(output_10_587));
wire output_12_587, output_12_12, output_11_587;
mixer gate_output_11_587(.a(output_12_587), .b(output_12_12), .y(output_11_587));
wire output_13_587, output_13_12, output_12_587;
mixer gate_output_12_587(.a(output_13_587), .b(output_13_12), .y(output_12_587));
wire output_14_587, output_14_12, output_13_587;
mixer gate_output_13_587(.a(output_14_587), .b(output_14_12), .y(output_13_587));
wire output_15_587, output_15_12, output_14_587;
mixer gate_output_14_587(.a(output_15_587), .b(output_15_12), .y(output_14_587));
wire output_16_587, output_16_12, output_15_587;
mixer gate_output_15_587(.a(output_16_587), .b(output_16_12), .y(output_15_587));
wire output_1_588, output_1_13, output_0_588;
mixer gate_output_0_588(.a(output_1_588), .b(output_1_13), .y(output_0_588));
wire output_2_588, output_2_13, output_1_588;
mixer gate_output_1_588(.a(output_2_588), .b(output_2_13), .y(output_1_588));
wire output_3_588, output_3_13, output_2_588;
mixer gate_output_2_588(.a(output_3_588), .b(output_3_13), .y(output_2_588));
wire output_4_588, output_4_13, output_3_588;
mixer gate_output_3_588(.a(output_4_588), .b(output_4_13), .y(output_3_588));
wire output_5_588, output_5_13, output_4_588;
mixer gate_output_4_588(.a(output_5_588), .b(output_5_13), .y(output_4_588));
wire output_6_588, output_6_13, output_5_588;
mixer gate_output_5_588(.a(output_6_588), .b(output_6_13), .y(output_5_588));
wire output_7_588, output_7_13, output_6_588;
mixer gate_output_6_588(.a(output_7_588), .b(output_7_13), .y(output_6_588));
wire output_8_588, output_8_13, output_7_588;
mixer gate_output_7_588(.a(output_8_588), .b(output_8_13), .y(output_7_588));
wire output_9_588, output_9_13, output_8_588;
mixer gate_output_8_588(.a(output_9_588), .b(output_9_13), .y(output_8_588));
wire output_10_588, output_10_13, output_9_588;
mixer gate_output_9_588(.a(output_10_588), .b(output_10_13), .y(output_9_588));
wire output_11_588, output_11_13, output_10_588;
mixer gate_output_10_588(.a(output_11_588), .b(output_11_13), .y(output_10_588));
wire output_12_588, output_12_13, output_11_588;
mixer gate_output_11_588(.a(output_12_588), .b(output_12_13), .y(output_11_588));
wire output_13_588, output_13_13, output_12_588;
mixer gate_output_12_588(.a(output_13_588), .b(output_13_13), .y(output_12_588));
wire output_14_588, output_14_13, output_13_588;
mixer gate_output_13_588(.a(output_14_588), .b(output_14_13), .y(output_13_588));
wire output_15_588, output_15_13, output_14_588;
mixer gate_output_14_588(.a(output_15_588), .b(output_15_13), .y(output_14_588));
wire output_16_588, output_16_13, output_15_588;
mixer gate_output_15_588(.a(output_16_588), .b(output_16_13), .y(output_15_588));
wire output_1_589, output_1_14, output_0_589;
mixer gate_output_0_589(.a(output_1_589), .b(output_1_14), .y(output_0_589));
wire output_2_589, output_2_14, output_1_589;
mixer gate_output_1_589(.a(output_2_589), .b(output_2_14), .y(output_1_589));
wire output_3_589, output_3_14, output_2_589;
mixer gate_output_2_589(.a(output_3_589), .b(output_3_14), .y(output_2_589));
wire output_4_589, output_4_14, output_3_589;
mixer gate_output_3_589(.a(output_4_589), .b(output_4_14), .y(output_3_589));
wire output_5_589, output_5_14, output_4_589;
mixer gate_output_4_589(.a(output_5_589), .b(output_5_14), .y(output_4_589));
wire output_6_589, output_6_14, output_5_589;
mixer gate_output_5_589(.a(output_6_589), .b(output_6_14), .y(output_5_589));
wire output_7_589, output_7_14, output_6_589;
mixer gate_output_6_589(.a(output_7_589), .b(output_7_14), .y(output_6_589));
wire output_8_589, output_8_14, output_7_589;
mixer gate_output_7_589(.a(output_8_589), .b(output_8_14), .y(output_7_589));
wire output_9_589, output_9_14, output_8_589;
mixer gate_output_8_589(.a(output_9_589), .b(output_9_14), .y(output_8_589));
wire output_10_589, output_10_14, output_9_589;
mixer gate_output_9_589(.a(output_10_589), .b(output_10_14), .y(output_9_589));
wire output_11_589, output_11_14, output_10_589;
mixer gate_output_10_589(.a(output_11_589), .b(output_11_14), .y(output_10_589));
wire output_12_589, output_12_14, output_11_589;
mixer gate_output_11_589(.a(output_12_589), .b(output_12_14), .y(output_11_589));
wire output_13_589, output_13_14, output_12_589;
mixer gate_output_12_589(.a(output_13_589), .b(output_13_14), .y(output_12_589));
wire output_14_589, output_14_14, output_13_589;
mixer gate_output_13_589(.a(output_14_589), .b(output_14_14), .y(output_13_589));
wire output_15_589, output_15_14, output_14_589;
mixer gate_output_14_589(.a(output_15_589), .b(output_15_14), .y(output_14_589));
wire output_16_589, output_16_14, output_15_589;
mixer gate_output_15_589(.a(output_16_589), .b(output_16_14), .y(output_15_589));
wire output_1_590, output_1_15, output_0_590;
mixer gate_output_0_590(.a(output_1_590), .b(output_1_15), .y(output_0_590));
wire output_2_590, output_2_15, output_1_590;
mixer gate_output_1_590(.a(output_2_590), .b(output_2_15), .y(output_1_590));
wire output_3_590, output_3_15, output_2_590;
mixer gate_output_2_590(.a(output_3_590), .b(output_3_15), .y(output_2_590));
wire output_4_590, output_4_15, output_3_590;
mixer gate_output_3_590(.a(output_4_590), .b(output_4_15), .y(output_3_590));
wire output_5_590, output_5_15, output_4_590;
mixer gate_output_4_590(.a(output_5_590), .b(output_5_15), .y(output_4_590));
wire output_6_590, output_6_15, output_5_590;
mixer gate_output_5_590(.a(output_6_590), .b(output_6_15), .y(output_5_590));
wire output_7_590, output_7_15, output_6_590;
mixer gate_output_6_590(.a(output_7_590), .b(output_7_15), .y(output_6_590));
wire output_8_590, output_8_15, output_7_590;
mixer gate_output_7_590(.a(output_8_590), .b(output_8_15), .y(output_7_590));
wire output_9_590, output_9_15, output_8_590;
mixer gate_output_8_590(.a(output_9_590), .b(output_9_15), .y(output_8_590));
wire output_10_590, output_10_15, output_9_590;
mixer gate_output_9_590(.a(output_10_590), .b(output_10_15), .y(output_9_590));
wire output_11_590, output_11_15, output_10_590;
mixer gate_output_10_590(.a(output_11_590), .b(output_11_15), .y(output_10_590));
wire output_12_590, output_12_15, output_11_590;
mixer gate_output_11_590(.a(output_12_590), .b(output_12_15), .y(output_11_590));
wire output_13_590, output_13_15, output_12_590;
mixer gate_output_12_590(.a(output_13_590), .b(output_13_15), .y(output_12_590));
wire output_14_590, output_14_15, output_13_590;
mixer gate_output_13_590(.a(output_14_590), .b(output_14_15), .y(output_13_590));
wire output_15_590, output_15_15, output_14_590;
mixer gate_output_14_590(.a(output_15_590), .b(output_15_15), .y(output_14_590));
wire output_16_590, output_16_15, output_15_590;
mixer gate_output_15_590(.a(output_16_590), .b(output_16_15), .y(output_15_590));
wire output_1_591, output_1_0, output_0_591;
mixer gate_output_0_591(.a(output_1_591), .b(output_1_0), .y(output_0_591));
wire output_2_591, output_2_0, output_1_591;
mixer gate_output_1_591(.a(output_2_591), .b(output_2_0), .y(output_1_591));
wire output_3_591, output_3_0, output_2_591;
mixer gate_output_2_591(.a(output_3_591), .b(output_3_0), .y(output_2_591));
wire output_4_591, output_4_0, output_3_591;
mixer gate_output_3_591(.a(output_4_591), .b(output_4_0), .y(output_3_591));
wire output_5_591, output_5_0, output_4_591;
mixer gate_output_4_591(.a(output_5_591), .b(output_5_0), .y(output_4_591));
wire output_6_591, output_6_0, output_5_591;
mixer gate_output_5_591(.a(output_6_591), .b(output_6_0), .y(output_5_591));
wire output_7_591, output_7_0, output_6_591;
mixer gate_output_6_591(.a(output_7_591), .b(output_7_0), .y(output_6_591));
wire output_8_591, output_8_0, output_7_591;
mixer gate_output_7_591(.a(output_8_591), .b(output_8_0), .y(output_7_591));
wire output_9_591, output_9_0, output_8_591;
mixer gate_output_8_591(.a(output_9_591), .b(output_9_0), .y(output_8_591));
wire output_10_591, output_10_0, output_9_591;
mixer gate_output_9_591(.a(output_10_591), .b(output_10_0), .y(output_9_591));
wire output_11_591, output_11_0, output_10_591;
mixer gate_output_10_591(.a(output_11_591), .b(output_11_0), .y(output_10_591));
wire output_12_591, output_12_0, output_11_591;
mixer gate_output_11_591(.a(output_12_591), .b(output_12_0), .y(output_11_591));
wire output_13_591, output_13_0, output_12_591;
mixer gate_output_12_591(.a(output_13_591), .b(output_13_0), .y(output_12_591));
wire output_14_591, output_14_0, output_13_591;
mixer gate_output_13_591(.a(output_14_591), .b(output_14_0), .y(output_13_591));
wire output_15_591, output_15_0, output_14_591;
mixer gate_output_14_591(.a(output_15_591), .b(output_15_0), .y(output_14_591));
wire output_16_591, output_16_0, output_15_591;
mixer gate_output_15_591(.a(output_16_591), .b(output_16_0), .y(output_15_591));
wire output_1_592, output_1_1, output_0_592;
mixer gate_output_0_592(.a(output_1_592), .b(output_1_1), .y(output_0_592));
wire output_2_592, output_2_1, output_1_592;
mixer gate_output_1_592(.a(output_2_592), .b(output_2_1), .y(output_1_592));
wire output_3_592, output_3_1, output_2_592;
mixer gate_output_2_592(.a(output_3_592), .b(output_3_1), .y(output_2_592));
wire output_4_592, output_4_1, output_3_592;
mixer gate_output_3_592(.a(output_4_592), .b(output_4_1), .y(output_3_592));
wire output_5_592, output_5_1, output_4_592;
mixer gate_output_4_592(.a(output_5_592), .b(output_5_1), .y(output_4_592));
wire output_6_592, output_6_1, output_5_592;
mixer gate_output_5_592(.a(output_6_592), .b(output_6_1), .y(output_5_592));
wire output_7_592, output_7_1, output_6_592;
mixer gate_output_6_592(.a(output_7_592), .b(output_7_1), .y(output_6_592));
wire output_8_592, output_8_1, output_7_592;
mixer gate_output_7_592(.a(output_8_592), .b(output_8_1), .y(output_7_592));
wire output_9_592, output_9_1, output_8_592;
mixer gate_output_8_592(.a(output_9_592), .b(output_9_1), .y(output_8_592));
wire output_10_592, output_10_1, output_9_592;
mixer gate_output_9_592(.a(output_10_592), .b(output_10_1), .y(output_9_592));
wire output_11_592, output_11_1, output_10_592;
mixer gate_output_10_592(.a(output_11_592), .b(output_11_1), .y(output_10_592));
wire output_12_592, output_12_1, output_11_592;
mixer gate_output_11_592(.a(output_12_592), .b(output_12_1), .y(output_11_592));
wire output_13_592, output_13_1, output_12_592;
mixer gate_output_12_592(.a(output_13_592), .b(output_13_1), .y(output_12_592));
wire output_14_592, output_14_1, output_13_592;
mixer gate_output_13_592(.a(output_14_592), .b(output_14_1), .y(output_13_592));
wire output_15_592, output_15_1, output_14_592;
mixer gate_output_14_592(.a(output_15_592), .b(output_15_1), .y(output_14_592));
wire output_16_592, output_16_1, output_15_592;
mixer gate_output_15_592(.a(output_16_592), .b(output_16_1), .y(output_15_592));
wire output_1_593, output_1_2, output_0_593;
mixer gate_output_0_593(.a(output_1_593), .b(output_1_2), .y(output_0_593));
wire output_2_593, output_2_2, output_1_593;
mixer gate_output_1_593(.a(output_2_593), .b(output_2_2), .y(output_1_593));
wire output_3_593, output_3_2, output_2_593;
mixer gate_output_2_593(.a(output_3_593), .b(output_3_2), .y(output_2_593));
wire output_4_593, output_4_2, output_3_593;
mixer gate_output_3_593(.a(output_4_593), .b(output_4_2), .y(output_3_593));
wire output_5_593, output_5_2, output_4_593;
mixer gate_output_4_593(.a(output_5_593), .b(output_5_2), .y(output_4_593));
wire output_6_593, output_6_2, output_5_593;
mixer gate_output_5_593(.a(output_6_593), .b(output_6_2), .y(output_5_593));
wire output_7_593, output_7_2, output_6_593;
mixer gate_output_6_593(.a(output_7_593), .b(output_7_2), .y(output_6_593));
wire output_8_593, output_8_2, output_7_593;
mixer gate_output_7_593(.a(output_8_593), .b(output_8_2), .y(output_7_593));
wire output_9_593, output_9_2, output_8_593;
mixer gate_output_8_593(.a(output_9_593), .b(output_9_2), .y(output_8_593));
wire output_10_593, output_10_2, output_9_593;
mixer gate_output_9_593(.a(output_10_593), .b(output_10_2), .y(output_9_593));
wire output_11_593, output_11_2, output_10_593;
mixer gate_output_10_593(.a(output_11_593), .b(output_11_2), .y(output_10_593));
wire output_12_593, output_12_2, output_11_593;
mixer gate_output_11_593(.a(output_12_593), .b(output_12_2), .y(output_11_593));
wire output_13_593, output_13_2, output_12_593;
mixer gate_output_12_593(.a(output_13_593), .b(output_13_2), .y(output_12_593));
wire output_14_593, output_14_2, output_13_593;
mixer gate_output_13_593(.a(output_14_593), .b(output_14_2), .y(output_13_593));
wire output_15_593, output_15_2, output_14_593;
mixer gate_output_14_593(.a(output_15_593), .b(output_15_2), .y(output_14_593));
wire output_16_593, output_16_2, output_15_593;
mixer gate_output_15_593(.a(output_16_593), .b(output_16_2), .y(output_15_593));
wire output_1_594, output_1_3, output_0_594;
mixer gate_output_0_594(.a(output_1_594), .b(output_1_3), .y(output_0_594));
wire output_2_594, output_2_3, output_1_594;
mixer gate_output_1_594(.a(output_2_594), .b(output_2_3), .y(output_1_594));
wire output_3_594, output_3_3, output_2_594;
mixer gate_output_2_594(.a(output_3_594), .b(output_3_3), .y(output_2_594));
wire output_4_594, output_4_3, output_3_594;
mixer gate_output_3_594(.a(output_4_594), .b(output_4_3), .y(output_3_594));
wire output_5_594, output_5_3, output_4_594;
mixer gate_output_4_594(.a(output_5_594), .b(output_5_3), .y(output_4_594));
wire output_6_594, output_6_3, output_5_594;
mixer gate_output_5_594(.a(output_6_594), .b(output_6_3), .y(output_5_594));
wire output_7_594, output_7_3, output_6_594;
mixer gate_output_6_594(.a(output_7_594), .b(output_7_3), .y(output_6_594));
wire output_8_594, output_8_3, output_7_594;
mixer gate_output_7_594(.a(output_8_594), .b(output_8_3), .y(output_7_594));
wire output_9_594, output_9_3, output_8_594;
mixer gate_output_8_594(.a(output_9_594), .b(output_9_3), .y(output_8_594));
wire output_10_594, output_10_3, output_9_594;
mixer gate_output_9_594(.a(output_10_594), .b(output_10_3), .y(output_9_594));
wire output_11_594, output_11_3, output_10_594;
mixer gate_output_10_594(.a(output_11_594), .b(output_11_3), .y(output_10_594));
wire output_12_594, output_12_3, output_11_594;
mixer gate_output_11_594(.a(output_12_594), .b(output_12_3), .y(output_11_594));
wire output_13_594, output_13_3, output_12_594;
mixer gate_output_12_594(.a(output_13_594), .b(output_13_3), .y(output_12_594));
wire output_14_594, output_14_3, output_13_594;
mixer gate_output_13_594(.a(output_14_594), .b(output_14_3), .y(output_13_594));
wire output_15_594, output_15_3, output_14_594;
mixer gate_output_14_594(.a(output_15_594), .b(output_15_3), .y(output_14_594));
wire output_16_594, output_16_3, output_15_594;
mixer gate_output_15_594(.a(output_16_594), .b(output_16_3), .y(output_15_594));
wire output_1_595, output_1_4, output_0_595;
mixer gate_output_0_595(.a(output_1_595), .b(output_1_4), .y(output_0_595));
wire output_2_595, output_2_4, output_1_595;
mixer gate_output_1_595(.a(output_2_595), .b(output_2_4), .y(output_1_595));
wire output_3_595, output_3_4, output_2_595;
mixer gate_output_2_595(.a(output_3_595), .b(output_3_4), .y(output_2_595));
wire output_4_595, output_4_4, output_3_595;
mixer gate_output_3_595(.a(output_4_595), .b(output_4_4), .y(output_3_595));
wire output_5_595, output_5_4, output_4_595;
mixer gate_output_4_595(.a(output_5_595), .b(output_5_4), .y(output_4_595));
wire output_6_595, output_6_4, output_5_595;
mixer gate_output_5_595(.a(output_6_595), .b(output_6_4), .y(output_5_595));
wire output_7_595, output_7_4, output_6_595;
mixer gate_output_6_595(.a(output_7_595), .b(output_7_4), .y(output_6_595));
wire output_8_595, output_8_4, output_7_595;
mixer gate_output_7_595(.a(output_8_595), .b(output_8_4), .y(output_7_595));
wire output_9_595, output_9_4, output_8_595;
mixer gate_output_8_595(.a(output_9_595), .b(output_9_4), .y(output_8_595));
wire output_10_595, output_10_4, output_9_595;
mixer gate_output_9_595(.a(output_10_595), .b(output_10_4), .y(output_9_595));
wire output_11_595, output_11_4, output_10_595;
mixer gate_output_10_595(.a(output_11_595), .b(output_11_4), .y(output_10_595));
wire output_12_595, output_12_4, output_11_595;
mixer gate_output_11_595(.a(output_12_595), .b(output_12_4), .y(output_11_595));
wire output_13_595, output_13_4, output_12_595;
mixer gate_output_12_595(.a(output_13_595), .b(output_13_4), .y(output_12_595));
wire output_14_595, output_14_4, output_13_595;
mixer gate_output_13_595(.a(output_14_595), .b(output_14_4), .y(output_13_595));
wire output_15_595, output_15_4, output_14_595;
mixer gate_output_14_595(.a(output_15_595), .b(output_15_4), .y(output_14_595));
wire output_16_595, output_16_4, output_15_595;
mixer gate_output_15_595(.a(output_16_595), .b(output_16_4), .y(output_15_595));
wire output_1_596, output_1_5, output_0_596;
mixer gate_output_0_596(.a(output_1_596), .b(output_1_5), .y(output_0_596));
wire output_2_596, output_2_5, output_1_596;
mixer gate_output_1_596(.a(output_2_596), .b(output_2_5), .y(output_1_596));
wire output_3_596, output_3_5, output_2_596;
mixer gate_output_2_596(.a(output_3_596), .b(output_3_5), .y(output_2_596));
wire output_4_596, output_4_5, output_3_596;
mixer gate_output_3_596(.a(output_4_596), .b(output_4_5), .y(output_3_596));
wire output_5_596, output_5_5, output_4_596;
mixer gate_output_4_596(.a(output_5_596), .b(output_5_5), .y(output_4_596));
wire output_6_596, output_6_5, output_5_596;
mixer gate_output_5_596(.a(output_6_596), .b(output_6_5), .y(output_5_596));
wire output_7_596, output_7_5, output_6_596;
mixer gate_output_6_596(.a(output_7_596), .b(output_7_5), .y(output_6_596));
wire output_8_596, output_8_5, output_7_596;
mixer gate_output_7_596(.a(output_8_596), .b(output_8_5), .y(output_7_596));
wire output_9_596, output_9_5, output_8_596;
mixer gate_output_8_596(.a(output_9_596), .b(output_9_5), .y(output_8_596));
wire output_10_596, output_10_5, output_9_596;
mixer gate_output_9_596(.a(output_10_596), .b(output_10_5), .y(output_9_596));
wire output_11_596, output_11_5, output_10_596;
mixer gate_output_10_596(.a(output_11_596), .b(output_11_5), .y(output_10_596));
wire output_12_596, output_12_5, output_11_596;
mixer gate_output_11_596(.a(output_12_596), .b(output_12_5), .y(output_11_596));
wire output_13_596, output_13_5, output_12_596;
mixer gate_output_12_596(.a(output_13_596), .b(output_13_5), .y(output_12_596));
wire output_14_596, output_14_5, output_13_596;
mixer gate_output_13_596(.a(output_14_596), .b(output_14_5), .y(output_13_596));
wire output_15_596, output_15_5, output_14_596;
mixer gate_output_14_596(.a(output_15_596), .b(output_15_5), .y(output_14_596));
wire output_16_596, output_16_5, output_15_596;
mixer gate_output_15_596(.a(output_16_596), .b(output_16_5), .y(output_15_596));
wire output_1_597, output_1_6, output_0_597;
mixer gate_output_0_597(.a(output_1_597), .b(output_1_6), .y(output_0_597));
wire output_2_597, output_2_6, output_1_597;
mixer gate_output_1_597(.a(output_2_597), .b(output_2_6), .y(output_1_597));
wire output_3_597, output_3_6, output_2_597;
mixer gate_output_2_597(.a(output_3_597), .b(output_3_6), .y(output_2_597));
wire output_4_597, output_4_6, output_3_597;
mixer gate_output_3_597(.a(output_4_597), .b(output_4_6), .y(output_3_597));
wire output_5_597, output_5_6, output_4_597;
mixer gate_output_4_597(.a(output_5_597), .b(output_5_6), .y(output_4_597));
wire output_6_597, output_6_6, output_5_597;
mixer gate_output_5_597(.a(output_6_597), .b(output_6_6), .y(output_5_597));
wire output_7_597, output_7_6, output_6_597;
mixer gate_output_6_597(.a(output_7_597), .b(output_7_6), .y(output_6_597));
wire output_8_597, output_8_6, output_7_597;
mixer gate_output_7_597(.a(output_8_597), .b(output_8_6), .y(output_7_597));
wire output_9_597, output_9_6, output_8_597;
mixer gate_output_8_597(.a(output_9_597), .b(output_9_6), .y(output_8_597));
wire output_10_597, output_10_6, output_9_597;
mixer gate_output_9_597(.a(output_10_597), .b(output_10_6), .y(output_9_597));
wire output_11_597, output_11_6, output_10_597;
mixer gate_output_10_597(.a(output_11_597), .b(output_11_6), .y(output_10_597));
wire output_12_597, output_12_6, output_11_597;
mixer gate_output_11_597(.a(output_12_597), .b(output_12_6), .y(output_11_597));
wire output_13_597, output_13_6, output_12_597;
mixer gate_output_12_597(.a(output_13_597), .b(output_13_6), .y(output_12_597));
wire output_14_597, output_14_6, output_13_597;
mixer gate_output_13_597(.a(output_14_597), .b(output_14_6), .y(output_13_597));
wire output_15_597, output_15_6, output_14_597;
mixer gate_output_14_597(.a(output_15_597), .b(output_15_6), .y(output_14_597));
wire output_16_597, output_16_6, output_15_597;
mixer gate_output_15_597(.a(output_16_597), .b(output_16_6), .y(output_15_597));
wire output_1_598, output_1_7, output_0_598;
mixer gate_output_0_598(.a(output_1_598), .b(output_1_7), .y(output_0_598));
wire output_2_598, output_2_7, output_1_598;
mixer gate_output_1_598(.a(output_2_598), .b(output_2_7), .y(output_1_598));
wire output_3_598, output_3_7, output_2_598;
mixer gate_output_2_598(.a(output_3_598), .b(output_3_7), .y(output_2_598));
wire output_4_598, output_4_7, output_3_598;
mixer gate_output_3_598(.a(output_4_598), .b(output_4_7), .y(output_3_598));
wire output_5_598, output_5_7, output_4_598;
mixer gate_output_4_598(.a(output_5_598), .b(output_5_7), .y(output_4_598));
wire output_6_598, output_6_7, output_5_598;
mixer gate_output_5_598(.a(output_6_598), .b(output_6_7), .y(output_5_598));
wire output_7_598, output_7_7, output_6_598;
mixer gate_output_6_598(.a(output_7_598), .b(output_7_7), .y(output_6_598));
wire output_8_598, output_8_7, output_7_598;
mixer gate_output_7_598(.a(output_8_598), .b(output_8_7), .y(output_7_598));
wire output_9_598, output_9_7, output_8_598;
mixer gate_output_8_598(.a(output_9_598), .b(output_9_7), .y(output_8_598));
wire output_10_598, output_10_7, output_9_598;
mixer gate_output_9_598(.a(output_10_598), .b(output_10_7), .y(output_9_598));
wire output_11_598, output_11_7, output_10_598;
mixer gate_output_10_598(.a(output_11_598), .b(output_11_7), .y(output_10_598));
wire output_12_598, output_12_7, output_11_598;
mixer gate_output_11_598(.a(output_12_598), .b(output_12_7), .y(output_11_598));
wire output_13_598, output_13_7, output_12_598;
mixer gate_output_12_598(.a(output_13_598), .b(output_13_7), .y(output_12_598));
wire output_14_598, output_14_7, output_13_598;
mixer gate_output_13_598(.a(output_14_598), .b(output_14_7), .y(output_13_598));
wire output_15_598, output_15_7, output_14_598;
mixer gate_output_14_598(.a(output_15_598), .b(output_15_7), .y(output_14_598));
wire output_16_598, output_16_7, output_15_598;
mixer gate_output_15_598(.a(output_16_598), .b(output_16_7), .y(output_15_598));
wire output_1_599, output_1_8, output_0_599;
mixer gate_output_0_599(.a(output_1_599), .b(output_1_8), .y(output_0_599));
wire output_2_599, output_2_8, output_1_599;
mixer gate_output_1_599(.a(output_2_599), .b(output_2_8), .y(output_1_599));
wire output_3_599, output_3_8, output_2_599;
mixer gate_output_2_599(.a(output_3_599), .b(output_3_8), .y(output_2_599));
wire output_4_599, output_4_8, output_3_599;
mixer gate_output_3_599(.a(output_4_599), .b(output_4_8), .y(output_3_599));
wire output_5_599, output_5_8, output_4_599;
mixer gate_output_4_599(.a(output_5_599), .b(output_5_8), .y(output_4_599));
wire output_6_599, output_6_8, output_5_599;
mixer gate_output_5_599(.a(output_6_599), .b(output_6_8), .y(output_5_599));
wire output_7_599, output_7_8, output_6_599;
mixer gate_output_6_599(.a(output_7_599), .b(output_7_8), .y(output_6_599));
wire output_8_599, output_8_8, output_7_599;
mixer gate_output_7_599(.a(output_8_599), .b(output_8_8), .y(output_7_599));
wire output_9_599, output_9_8, output_8_599;
mixer gate_output_8_599(.a(output_9_599), .b(output_9_8), .y(output_8_599));
wire output_10_599, output_10_8, output_9_599;
mixer gate_output_9_599(.a(output_10_599), .b(output_10_8), .y(output_9_599));
wire output_11_599, output_11_8, output_10_599;
mixer gate_output_10_599(.a(output_11_599), .b(output_11_8), .y(output_10_599));
wire output_12_599, output_12_8, output_11_599;
mixer gate_output_11_599(.a(output_12_599), .b(output_12_8), .y(output_11_599));
wire output_13_599, output_13_8, output_12_599;
mixer gate_output_12_599(.a(output_13_599), .b(output_13_8), .y(output_12_599));
wire output_14_599, output_14_8, output_13_599;
mixer gate_output_13_599(.a(output_14_599), .b(output_14_8), .y(output_13_599));
wire output_15_599, output_15_8, output_14_599;
mixer gate_output_14_599(.a(output_15_599), .b(output_15_8), .y(output_14_599));
wire output_16_599, output_16_8, output_15_599;
mixer gate_output_15_599(.a(output_16_599), .b(output_16_8), .y(output_15_599));
wire output_1_600, output_1_9, output_0_600;
mixer gate_output_0_600(.a(output_1_600), .b(output_1_9), .y(output_0_600));
wire output_2_600, output_2_9, output_1_600;
mixer gate_output_1_600(.a(output_2_600), .b(output_2_9), .y(output_1_600));
wire output_3_600, output_3_9, output_2_600;
mixer gate_output_2_600(.a(output_3_600), .b(output_3_9), .y(output_2_600));
wire output_4_600, output_4_9, output_3_600;
mixer gate_output_3_600(.a(output_4_600), .b(output_4_9), .y(output_3_600));
wire output_5_600, output_5_9, output_4_600;
mixer gate_output_4_600(.a(output_5_600), .b(output_5_9), .y(output_4_600));
wire output_6_600, output_6_9, output_5_600;
mixer gate_output_5_600(.a(output_6_600), .b(output_6_9), .y(output_5_600));
wire output_7_600, output_7_9, output_6_600;
mixer gate_output_6_600(.a(output_7_600), .b(output_7_9), .y(output_6_600));
wire output_8_600, output_8_9, output_7_600;
mixer gate_output_7_600(.a(output_8_600), .b(output_8_9), .y(output_7_600));
wire output_9_600, output_9_9, output_8_600;
mixer gate_output_8_600(.a(output_9_600), .b(output_9_9), .y(output_8_600));
wire output_10_600, output_10_9, output_9_600;
mixer gate_output_9_600(.a(output_10_600), .b(output_10_9), .y(output_9_600));
wire output_11_600, output_11_9, output_10_600;
mixer gate_output_10_600(.a(output_11_600), .b(output_11_9), .y(output_10_600));
wire output_12_600, output_12_9, output_11_600;
mixer gate_output_11_600(.a(output_12_600), .b(output_12_9), .y(output_11_600));
wire output_13_600, output_13_9, output_12_600;
mixer gate_output_12_600(.a(output_13_600), .b(output_13_9), .y(output_12_600));
wire output_14_600, output_14_9, output_13_600;
mixer gate_output_13_600(.a(output_14_600), .b(output_14_9), .y(output_13_600));
wire output_15_600, output_15_9, output_14_600;
mixer gate_output_14_600(.a(output_15_600), .b(output_15_9), .y(output_14_600));
wire output_16_600, output_16_9, output_15_600;
mixer gate_output_15_600(.a(output_16_600), .b(output_16_9), .y(output_15_600));
wire output_1_601, output_1_10, output_0_601;
mixer gate_output_0_601(.a(output_1_601), .b(output_1_10), .y(output_0_601));
wire output_2_601, output_2_10, output_1_601;
mixer gate_output_1_601(.a(output_2_601), .b(output_2_10), .y(output_1_601));
wire output_3_601, output_3_10, output_2_601;
mixer gate_output_2_601(.a(output_3_601), .b(output_3_10), .y(output_2_601));
wire output_4_601, output_4_10, output_3_601;
mixer gate_output_3_601(.a(output_4_601), .b(output_4_10), .y(output_3_601));
wire output_5_601, output_5_10, output_4_601;
mixer gate_output_4_601(.a(output_5_601), .b(output_5_10), .y(output_4_601));
wire output_6_601, output_6_10, output_5_601;
mixer gate_output_5_601(.a(output_6_601), .b(output_6_10), .y(output_5_601));
wire output_7_601, output_7_10, output_6_601;
mixer gate_output_6_601(.a(output_7_601), .b(output_7_10), .y(output_6_601));
wire output_8_601, output_8_10, output_7_601;
mixer gate_output_7_601(.a(output_8_601), .b(output_8_10), .y(output_7_601));
wire output_9_601, output_9_10, output_8_601;
mixer gate_output_8_601(.a(output_9_601), .b(output_9_10), .y(output_8_601));
wire output_10_601, output_10_10, output_9_601;
mixer gate_output_9_601(.a(output_10_601), .b(output_10_10), .y(output_9_601));
wire output_11_601, output_11_10, output_10_601;
mixer gate_output_10_601(.a(output_11_601), .b(output_11_10), .y(output_10_601));
wire output_12_601, output_12_10, output_11_601;
mixer gate_output_11_601(.a(output_12_601), .b(output_12_10), .y(output_11_601));
wire output_13_601, output_13_10, output_12_601;
mixer gate_output_12_601(.a(output_13_601), .b(output_13_10), .y(output_12_601));
wire output_14_601, output_14_10, output_13_601;
mixer gate_output_13_601(.a(output_14_601), .b(output_14_10), .y(output_13_601));
wire output_15_601, output_15_10, output_14_601;
mixer gate_output_14_601(.a(output_15_601), .b(output_15_10), .y(output_14_601));
wire output_16_601, output_16_10, output_15_601;
mixer gate_output_15_601(.a(output_16_601), .b(output_16_10), .y(output_15_601));
wire output_1_602, output_1_11, output_0_602;
mixer gate_output_0_602(.a(output_1_602), .b(output_1_11), .y(output_0_602));
wire output_2_602, output_2_11, output_1_602;
mixer gate_output_1_602(.a(output_2_602), .b(output_2_11), .y(output_1_602));
wire output_3_602, output_3_11, output_2_602;
mixer gate_output_2_602(.a(output_3_602), .b(output_3_11), .y(output_2_602));
wire output_4_602, output_4_11, output_3_602;
mixer gate_output_3_602(.a(output_4_602), .b(output_4_11), .y(output_3_602));
wire output_5_602, output_5_11, output_4_602;
mixer gate_output_4_602(.a(output_5_602), .b(output_5_11), .y(output_4_602));
wire output_6_602, output_6_11, output_5_602;
mixer gate_output_5_602(.a(output_6_602), .b(output_6_11), .y(output_5_602));
wire output_7_602, output_7_11, output_6_602;
mixer gate_output_6_602(.a(output_7_602), .b(output_7_11), .y(output_6_602));
wire output_8_602, output_8_11, output_7_602;
mixer gate_output_7_602(.a(output_8_602), .b(output_8_11), .y(output_7_602));
wire output_9_602, output_9_11, output_8_602;
mixer gate_output_8_602(.a(output_9_602), .b(output_9_11), .y(output_8_602));
wire output_10_602, output_10_11, output_9_602;
mixer gate_output_9_602(.a(output_10_602), .b(output_10_11), .y(output_9_602));
wire output_11_602, output_11_11, output_10_602;
mixer gate_output_10_602(.a(output_11_602), .b(output_11_11), .y(output_10_602));
wire output_12_602, output_12_11, output_11_602;
mixer gate_output_11_602(.a(output_12_602), .b(output_12_11), .y(output_11_602));
wire output_13_602, output_13_11, output_12_602;
mixer gate_output_12_602(.a(output_13_602), .b(output_13_11), .y(output_12_602));
wire output_14_602, output_14_11, output_13_602;
mixer gate_output_13_602(.a(output_14_602), .b(output_14_11), .y(output_13_602));
wire output_15_602, output_15_11, output_14_602;
mixer gate_output_14_602(.a(output_15_602), .b(output_15_11), .y(output_14_602));
wire output_16_602, output_16_11, output_15_602;
mixer gate_output_15_602(.a(output_16_602), .b(output_16_11), .y(output_15_602));
wire output_1_603, output_1_12, output_0_603;
mixer gate_output_0_603(.a(output_1_603), .b(output_1_12), .y(output_0_603));
wire output_2_603, output_2_12, output_1_603;
mixer gate_output_1_603(.a(output_2_603), .b(output_2_12), .y(output_1_603));
wire output_3_603, output_3_12, output_2_603;
mixer gate_output_2_603(.a(output_3_603), .b(output_3_12), .y(output_2_603));
wire output_4_603, output_4_12, output_3_603;
mixer gate_output_3_603(.a(output_4_603), .b(output_4_12), .y(output_3_603));
wire output_5_603, output_5_12, output_4_603;
mixer gate_output_4_603(.a(output_5_603), .b(output_5_12), .y(output_4_603));
wire output_6_603, output_6_12, output_5_603;
mixer gate_output_5_603(.a(output_6_603), .b(output_6_12), .y(output_5_603));
wire output_7_603, output_7_12, output_6_603;
mixer gate_output_6_603(.a(output_7_603), .b(output_7_12), .y(output_6_603));
wire output_8_603, output_8_12, output_7_603;
mixer gate_output_7_603(.a(output_8_603), .b(output_8_12), .y(output_7_603));
wire output_9_603, output_9_12, output_8_603;
mixer gate_output_8_603(.a(output_9_603), .b(output_9_12), .y(output_8_603));
wire output_10_603, output_10_12, output_9_603;
mixer gate_output_9_603(.a(output_10_603), .b(output_10_12), .y(output_9_603));
wire output_11_603, output_11_12, output_10_603;
mixer gate_output_10_603(.a(output_11_603), .b(output_11_12), .y(output_10_603));
wire output_12_603, output_12_12, output_11_603;
mixer gate_output_11_603(.a(output_12_603), .b(output_12_12), .y(output_11_603));
wire output_13_603, output_13_12, output_12_603;
mixer gate_output_12_603(.a(output_13_603), .b(output_13_12), .y(output_12_603));
wire output_14_603, output_14_12, output_13_603;
mixer gate_output_13_603(.a(output_14_603), .b(output_14_12), .y(output_13_603));
wire output_15_603, output_15_12, output_14_603;
mixer gate_output_14_603(.a(output_15_603), .b(output_15_12), .y(output_14_603));
wire output_16_603, output_16_12, output_15_603;
mixer gate_output_15_603(.a(output_16_603), .b(output_16_12), .y(output_15_603));
wire output_1_604, output_1_13, output_0_604;
mixer gate_output_0_604(.a(output_1_604), .b(output_1_13), .y(output_0_604));
wire output_2_604, output_2_13, output_1_604;
mixer gate_output_1_604(.a(output_2_604), .b(output_2_13), .y(output_1_604));
wire output_3_604, output_3_13, output_2_604;
mixer gate_output_2_604(.a(output_3_604), .b(output_3_13), .y(output_2_604));
wire output_4_604, output_4_13, output_3_604;
mixer gate_output_3_604(.a(output_4_604), .b(output_4_13), .y(output_3_604));
wire output_5_604, output_5_13, output_4_604;
mixer gate_output_4_604(.a(output_5_604), .b(output_5_13), .y(output_4_604));
wire output_6_604, output_6_13, output_5_604;
mixer gate_output_5_604(.a(output_6_604), .b(output_6_13), .y(output_5_604));
wire output_7_604, output_7_13, output_6_604;
mixer gate_output_6_604(.a(output_7_604), .b(output_7_13), .y(output_6_604));
wire output_8_604, output_8_13, output_7_604;
mixer gate_output_7_604(.a(output_8_604), .b(output_8_13), .y(output_7_604));
wire output_9_604, output_9_13, output_8_604;
mixer gate_output_8_604(.a(output_9_604), .b(output_9_13), .y(output_8_604));
wire output_10_604, output_10_13, output_9_604;
mixer gate_output_9_604(.a(output_10_604), .b(output_10_13), .y(output_9_604));
wire output_11_604, output_11_13, output_10_604;
mixer gate_output_10_604(.a(output_11_604), .b(output_11_13), .y(output_10_604));
wire output_12_604, output_12_13, output_11_604;
mixer gate_output_11_604(.a(output_12_604), .b(output_12_13), .y(output_11_604));
wire output_13_604, output_13_13, output_12_604;
mixer gate_output_12_604(.a(output_13_604), .b(output_13_13), .y(output_12_604));
wire output_14_604, output_14_13, output_13_604;
mixer gate_output_13_604(.a(output_14_604), .b(output_14_13), .y(output_13_604));
wire output_15_604, output_15_13, output_14_604;
mixer gate_output_14_604(.a(output_15_604), .b(output_15_13), .y(output_14_604));
wire output_16_604, output_16_13, output_15_604;
mixer gate_output_15_604(.a(output_16_604), .b(output_16_13), .y(output_15_604));
wire output_1_605, output_1_14, output_0_605;
mixer gate_output_0_605(.a(output_1_605), .b(output_1_14), .y(output_0_605));
wire output_2_605, output_2_14, output_1_605;
mixer gate_output_1_605(.a(output_2_605), .b(output_2_14), .y(output_1_605));
wire output_3_605, output_3_14, output_2_605;
mixer gate_output_2_605(.a(output_3_605), .b(output_3_14), .y(output_2_605));
wire output_4_605, output_4_14, output_3_605;
mixer gate_output_3_605(.a(output_4_605), .b(output_4_14), .y(output_3_605));
wire output_5_605, output_5_14, output_4_605;
mixer gate_output_4_605(.a(output_5_605), .b(output_5_14), .y(output_4_605));
wire output_6_605, output_6_14, output_5_605;
mixer gate_output_5_605(.a(output_6_605), .b(output_6_14), .y(output_5_605));
wire output_7_605, output_7_14, output_6_605;
mixer gate_output_6_605(.a(output_7_605), .b(output_7_14), .y(output_6_605));
wire output_8_605, output_8_14, output_7_605;
mixer gate_output_7_605(.a(output_8_605), .b(output_8_14), .y(output_7_605));
wire output_9_605, output_9_14, output_8_605;
mixer gate_output_8_605(.a(output_9_605), .b(output_9_14), .y(output_8_605));
wire output_10_605, output_10_14, output_9_605;
mixer gate_output_9_605(.a(output_10_605), .b(output_10_14), .y(output_9_605));
wire output_11_605, output_11_14, output_10_605;
mixer gate_output_10_605(.a(output_11_605), .b(output_11_14), .y(output_10_605));
wire output_12_605, output_12_14, output_11_605;
mixer gate_output_11_605(.a(output_12_605), .b(output_12_14), .y(output_11_605));
wire output_13_605, output_13_14, output_12_605;
mixer gate_output_12_605(.a(output_13_605), .b(output_13_14), .y(output_12_605));
wire output_14_605, output_14_14, output_13_605;
mixer gate_output_13_605(.a(output_14_605), .b(output_14_14), .y(output_13_605));
wire output_15_605, output_15_14, output_14_605;
mixer gate_output_14_605(.a(output_15_605), .b(output_15_14), .y(output_14_605));
wire output_16_605, output_16_14, output_15_605;
mixer gate_output_15_605(.a(output_16_605), .b(output_16_14), .y(output_15_605));
wire output_1_606, output_1_15, output_0_606;
mixer gate_output_0_606(.a(output_1_606), .b(output_1_15), .y(output_0_606));
wire output_2_606, output_2_15, output_1_606;
mixer gate_output_1_606(.a(output_2_606), .b(output_2_15), .y(output_1_606));
wire output_3_606, output_3_15, output_2_606;
mixer gate_output_2_606(.a(output_3_606), .b(output_3_15), .y(output_2_606));
wire output_4_606, output_4_15, output_3_606;
mixer gate_output_3_606(.a(output_4_606), .b(output_4_15), .y(output_3_606));
wire output_5_606, output_5_15, output_4_606;
mixer gate_output_4_606(.a(output_5_606), .b(output_5_15), .y(output_4_606));
wire output_6_606, output_6_15, output_5_606;
mixer gate_output_5_606(.a(output_6_606), .b(output_6_15), .y(output_5_606));
wire output_7_606, output_7_15, output_6_606;
mixer gate_output_6_606(.a(output_7_606), .b(output_7_15), .y(output_6_606));
wire output_8_606, output_8_15, output_7_606;
mixer gate_output_7_606(.a(output_8_606), .b(output_8_15), .y(output_7_606));
wire output_9_606, output_9_15, output_8_606;
mixer gate_output_8_606(.a(output_9_606), .b(output_9_15), .y(output_8_606));
wire output_10_606, output_10_15, output_9_606;
mixer gate_output_9_606(.a(output_10_606), .b(output_10_15), .y(output_9_606));
wire output_11_606, output_11_15, output_10_606;
mixer gate_output_10_606(.a(output_11_606), .b(output_11_15), .y(output_10_606));
wire output_12_606, output_12_15, output_11_606;
mixer gate_output_11_606(.a(output_12_606), .b(output_12_15), .y(output_11_606));
wire output_13_606, output_13_15, output_12_606;
mixer gate_output_12_606(.a(output_13_606), .b(output_13_15), .y(output_12_606));
wire output_14_606, output_14_15, output_13_606;
mixer gate_output_13_606(.a(output_14_606), .b(output_14_15), .y(output_13_606));
wire output_15_606, output_15_15, output_14_606;
mixer gate_output_14_606(.a(output_15_606), .b(output_15_15), .y(output_14_606));
wire output_16_606, output_16_15, output_15_606;
mixer gate_output_15_606(.a(output_16_606), .b(output_16_15), .y(output_15_606));
wire output_1_607, output_1_0, output_0_607;
mixer gate_output_0_607(.a(output_1_607), .b(output_1_0), .y(output_0_607));
wire output_2_607, output_2_0, output_1_607;
mixer gate_output_1_607(.a(output_2_607), .b(output_2_0), .y(output_1_607));
wire output_3_607, output_3_0, output_2_607;
mixer gate_output_2_607(.a(output_3_607), .b(output_3_0), .y(output_2_607));
wire output_4_607, output_4_0, output_3_607;
mixer gate_output_3_607(.a(output_4_607), .b(output_4_0), .y(output_3_607));
wire output_5_607, output_5_0, output_4_607;
mixer gate_output_4_607(.a(output_5_607), .b(output_5_0), .y(output_4_607));
wire output_6_607, output_6_0, output_5_607;
mixer gate_output_5_607(.a(output_6_607), .b(output_6_0), .y(output_5_607));
wire output_7_607, output_7_0, output_6_607;
mixer gate_output_6_607(.a(output_7_607), .b(output_7_0), .y(output_6_607));
wire output_8_607, output_8_0, output_7_607;
mixer gate_output_7_607(.a(output_8_607), .b(output_8_0), .y(output_7_607));
wire output_9_607, output_9_0, output_8_607;
mixer gate_output_8_607(.a(output_9_607), .b(output_9_0), .y(output_8_607));
wire output_10_607, output_10_0, output_9_607;
mixer gate_output_9_607(.a(output_10_607), .b(output_10_0), .y(output_9_607));
wire output_11_607, output_11_0, output_10_607;
mixer gate_output_10_607(.a(output_11_607), .b(output_11_0), .y(output_10_607));
wire output_12_607, output_12_0, output_11_607;
mixer gate_output_11_607(.a(output_12_607), .b(output_12_0), .y(output_11_607));
wire output_13_607, output_13_0, output_12_607;
mixer gate_output_12_607(.a(output_13_607), .b(output_13_0), .y(output_12_607));
wire output_14_607, output_14_0, output_13_607;
mixer gate_output_13_607(.a(output_14_607), .b(output_14_0), .y(output_13_607));
wire output_15_607, output_15_0, output_14_607;
mixer gate_output_14_607(.a(output_15_607), .b(output_15_0), .y(output_14_607));
wire output_16_607, output_16_0, output_15_607;
mixer gate_output_15_607(.a(output_16_607), .b(output_16_0), .y(output_15_607));
wire output_1_608, output_1_1, output_0_608;
mixer gate_output_0_608(.a(output_1_608), .b(output_1_1), .y(output_0_608));
wire output_2_608, output_2_1, output_1_608;
mixer gate_output_1_608(.a(output_2_608), .b(output_2_1), .y(output_1_608));
wire output_3_608, output_3_1, output_2_608;
mixer gate_output_2_608(.a(output_3_608), .b(output_3_1), .y(output_2_608));
wire output_4_608, output_4_1, output_3_608;
mixer gate_output_3_608(.a(output_4_608), .b(output_4_1), .y(output_3_608));
wire output_5_608, output_5_1, output_4_608;
mixer gate_output_4_608(.a(output_5_608), .b(output_5_1), .y(output_4_608));
wire output_6_608, output_6_1, output_5_608;
mixer gate_output_5_608(.a(output_6_608), .b(output_6_1), .y(output_5_608));
wire output_7_608, output_7_1, output_6_608;
mixer gate_output_6_608(.a(output_7_608), .b(output_7_1), .y(output_6_608));
wire output_8_608, output_8_1, output_7_608;
mixer gate_output_7_608(.a(output_8_608), .b(output_8_1), .y(output_7_608));
wire output_9_608, output_9_1, output_8_608;
mixer gate_output_8_608(.a(output_9_608), .b(output_9_1), .y(output_8_608));
wire output_10_608, output_10_1, output_9_608;
mixer gate_output_9_608(.a(output_10_608), .b(output_10_1), .y(output_9_608));
wire output_11_608, output_11_1, output_10_608;
mixer gate_output_10_608(.a(output_11_608), .b(output_11_1), .y(output_10_608));
wire output_12_608, output_12_1, output_11_608;
mixer gate_output_11_608(.a(output_12_608), .b(output_12_1), .y(output_11_608));
wire output_13_608, output_13_1, output_12_608;
mixer gate_output_12_608(.a(output_13_608), .b(output_13_1), .y(output_12_608));
wire output_14_608, output_14_1, output_13_608;
mixer gate_output_13_608(.a(output_14_608), .b(output_14_1), .y(output_13_608));
wire output_15_608, output_15_1, output_14_608;
mixer gate_output_14_608(.a(output_15_608), .b(output_15_1), .y(output_14_608));
wire output_16_608, output_16_1, output_15_608;
mixer gate_output_15_608(.a(output_16_608), .b(output_16_1), .y(output_15_608));
wire output_1_609, output_1_2, output_0_609;
mixer gate_output_0_609(.a(output_1_609), .b(output_1_2), .y(output_0_609));
wire output_2_609, output_2_2, output_1_609;
mixer gate_output_1_609(.a(output_2_609), .b(output_2_2), .y(output_1_609));
wire output_3_609, output_3_2, output_2_609;
mixer gate_output_2_609(.a(output_3_609), .b(output_3_2), .y(output_2_609));
wire output_4_609, output_4_2, output_3_609;
mixer gate_output_3_609(.a(output_4_609), .b(output_4_2), .y(output_3_609));
wire output_5_609, output_5_2, output_4_609;
mixer gate_output_4_609(.a(output_5_609), .b(output_5_2), .y(output_4_609));
wire output_6_609, output_6_2, output_5_609;
mixer gate_output_5_609(.a(output_6_609), .b(output_6_2), .y(output_5_609));
wire output_7_609, output_7_2, output_6_609;
mixer gate_output_6_609(.a(output_7_609), .b(output_7_2), .y(output_6_609));
wire output_8_609, output_8_2, output_7_609;
mixer gate_output_7_609(.a(output_8_609), .b(output_8_2), .y(output_7_609));
wire output_9_609, output_9_2, output_8_609;
mixer gate_output_8_609(.a(output_9_609), .b(output_9_2), .y(output_8_609));
wire output_10_609, output_10_2, output_9_609;
mixer gate_output_9_609(.a(output_10_609), .b(output_10_2), .y(output_9_609));
wire output_11_609, output_11_2, output_10_609;
mixer gate_output_10_609(.a(output_11_609), .b(output_11_2), .y(output_10_609));
wire output_12_609, output_12_2, output_11_609;
mixer gate_output_11_609(.a(output_12_609), .b(output_12_2), .y(output_11_609));
wire output_13_609, output_13_2, output_12_609;
mixer gate_output_12_609(.a(output_13_609), .b(output_13_2), .y(output_12_609));
wire output_14_609, output_14_2, output_13_609;
mixer gate_output_13_609(.a(output_14_609), .b(output_14_2), .y(output_13_609));
wire output_15_609, output_15_2, output_14_609;
mixer gate_output_14_609(.a(output_15_609), .b(output_15_2), .y(output_14_609));
wire output_16_609, output_16_2, output_15_609;
mixer gate_output_15_609(.a(output_16_609), .b(output_16_2), .y(output_15_609));
wire output_1_610, output_1_3, output_0_610;
mixer gate_output_0_610(.a(output_1_610), .b(output_1_3), .y(output_0_610));
wire output_2_610, output_2_3, output_1_610;
mixer gate_output_1_610(.a(output_2_610), .b(output_2_3), .y(output_1_610));
wire output_3_610, output_3_3, output_2_610;
mixer gate_output_2_610(.a(output_3_610), .b(output_3_3), .y(output_2_610));
wire output_4_610, output_4_3, output_3_610;
mixer gate_output_3_610(.a(output_4_610), .b(output_4_3), .y(output_3_610));
wire output_5_610, output_5_3, output_4_610;
mixer gate_output_4_610(.a(output_5_610), .b(output_5_3), .y(output_4_610));
wire output_6_610, output_6_3, output_5_610;
mixer gate_output_5_610(.a(output_6_610), .b(output_6_3), .y(output_5_610));
wire output_7_610, output_7_3, output_6_610;
mixer gate_output_6_610(.a(output_7_610), .b(output_7_3), .y(output_6_610));
wire output_8_610, output_8_3, output_7_610;
mixer gate_output_7_610(.a(output_8_610), .b(output_8_3), .y(output_7_610));
wire output_9_610, output_9_3, output_8_610;
mixer gate_output_8_610(.a(output_9_610), .b(output_9_3), .y(output_8_610));
wire output_10_610, output_10_3, output_9_610;
mixer gate_output_9_610(.a(output_10_610), .b(output_10_3), .y(output_9_610));
wire output_11_610, output_11_3, output_10_610;
mixer gate_output_10_610(.a(output_11_610), .b(output_11_3), .y(output_10_610));
wire output_12_610, output_12_3, output_11_610;
mixer gate_output_11_610(.a(output_12_610), .b(output_12_3), .y(output_11_610));
wire output_13_610, output_13_3, output_12_610;
mixer gate_output_12_610(.a(output_13_610), .b(output_13_3), .y(output_12_610));
wire output_14_610, output_14_3, output_13_610;
mixer gate_output_13_610(.a(output_14_610), .b(output_14_3), .y(output_13_610));
wire output_15_610, output_15_3, output_14_610;
mixer gate_output_14_610(.a(output_15_610), .b(output_15_3), .y(output_14_610));
wire output_16_610, output_16_3, output_15_610;
mixer gate_output_15_610(.a(output_16_610), .b(output_16_3), .y(output_15_610));
wire output_1_611, output_1_4, output_0_611;
mixer gate_output_0_611(.a(output_1_611), .b(output_1_4), .y(output_0_611));
wire output_2_611, output_2_4, output_1_611;
mixer gate_output_1_611(.a(output_2_611), .b(output_2_4), .y(output_1_611));
wire output_3_611, output_3_4, output_2_611;
mixer gate_output_2_611(.a(output_3_611), .b(output_3_4), .y(output_2_611));
wire output_4_611, output_4_4, output_3_611;
mixer gate_output_3_611(.a(output_4_611), .b(output_4_4), .y(output_3_611));
wire output_5_611, output_5_4, output_4_611;
mixer gate_output_4_611(.a(output_5_611), .b(output_5_4), .y(output_4_611));
wire output_6_611, output_6_4, output_5_611;
mixer gate_output_5_611(.a(output_6_611), .b(output_6_4), .y(output_5_611));
wire output_7_611, output_7_4, output_6_611;
mixer gate_output_6_611(.a(output_7_611), .b(output_7_4), .y(output_6_611));
wire output_8_611, output_8_4, output_7_611;
mixer gate_output_7_611(.a(output_8_611), .b(output_8_4), .y(output_7_611));
wire output_9_611, output_9_4, output_8_611;
mixer gate_output_8_611(.a(output_9_611), .b(output_9_4), .y(output_8_611));
wire output_10_611, output_10_4, output_9_611;
mixer gate_output_9_611(.a(output_10_611), .b(output_10_4), .y(output_9_611));
wire output_11_611, output_11_4, output_10_611;
mixer gate_output_10_611(.a(output_11_611), .b(output_11_4), .y(output_10_611));
wire output_12_611, output_12_4, output_11_611;
mixer gate_output_11_611(.a(output_12_611), .b(output_12_4), .y(output_11_611));
wire output_13_611, output_13_4, output_12_611;
mixer gate_output_12_611(.a(output_13_611), .b(output_13_4), .y(output_12_611));
wire output_14_611, output_14_4, output_13_611;
mixer gate_output_13_611(.a(output_14_611), .b(output_14_4), .y(output_13_611));
wire output_15_611, output_15_4, output_14_611;
mixer gate_output_14_611(.a(output_15_611), .b(output_15_4), .y(output_14_611));
wire output_16_611, output_16_4, output_15_611;
mixer gate_output_15_611(.a(output_16_611), .b(output_16_4), .y(output_15_611));
wire output_1_612, output_1_5, output_0_612;
mixer gate_output_0_612(.a(output_1_612), .b(output_1_5), .y(output_0_612));
wire output_2_612, output_2_5, output_1_612;
mixer gate_output_1_612(.a(output_2_612), .b(output_2_5), .y(output_1_612));
wire output_3_612, output_3_5, output_2_612;
mixer gate_output_2_612(.a(output_3_612), .b(output_3_5), .y(output_2_612));
wire output_4_612, output_4_5, output_3_612;
mixer gate_output_3_612(.a(output_4_612), .b(output_4_5), .y(output_3_612));
wire output_5_612, output_5_5, output_4_612;
mixer gate_output_4_612(.a(output_5_612), .b(output_5_5), .y(output_4_612));
wire output_6_612, output_6_5, output_5_612;
mixer gate_output_5_612(.a(output_6_612), .b(output_6_5), .y(output_5_612));
wire output_7_612, output_7_5, output_6_612;
mixer gate_output_6_612(.a(output_7_612), .b(output_7_5), .y(output_6_612));
wire output_8_612, output_8_5, output_7_612;
mixer gate_output_7_612(.a(output_8_612), .b(output_8_5), .y(output_7_612));
wire output_9_612, output_9_5, output_8_612;
mixer gate_output_8_612(.a(output_9_612), .b(output_9_5), .y(output_8_612));
wire output_10_612, output_10_5, output_9_612;
mixer gate_output_9_612(.a(output_10_612), .b(output_10_5), .y(output_9_612));
wire output_11_612, output_11_5, output_10_612;
mixer gate_output_10_612(.a(output_11_612), .b(output_11_5), .y(output_10_612));
wire output_12_612, output_12_5, output_11_612;
mixer gate_output_11_612(.a(output_12_612), .b(output_12_5), .y(output_11_612));
wire output_13_612, output_13_5, output_12_612;
mixer gate_output_12_612(.a(output_13_612), .b(output_13_5), .y(output_12_612));
wire output_14_612, output_14_5, output_13_612;
mixer gate_output_13_612(.a(output_14_612), .b(output_14_5), .y(output_13_612));
wire output_15_612, output_15_5, output_14_612;
mixer gate_output_14_612(.a(output_15_612), .b(output_15_5), .y(output_14_612));
wire output_16_612, output_16_5, output_15_612;
mixer gate_output_15_612(.a(output_16_612), .b(output_16_5), .y(output_15_612));
wire output_1_613, output_1_6, output_0_613;
mixer gate_output_0_613(.a(output_1_613), .b(output_1_6), .y(output_0_613));
wire output_2_613, output_2_6, output_1_613;
mixer gate_output_1_613(.a(output_2_613), .b(output_2_6), .y(output_1_613));
wire output_3_613, output_3_6, output_2_613;
mixer gate_output_2_613(.a(output_3_613), .b(output_3_6), .y(output_2_613));
wire output_4_613, output_4_6, output_3_613;
mixer gate_output_3_613(.a(output_4_613), .b(output_4_6), .y(output_3_613));
wire output_5_613, output_5_6, output_4_613;
mixer gate_output_4_613(.a(output_5_613), .b(output_5_6), .y(output_4_613));
wire output_6_613, output_6_6, output_5_613;
mixer gate_output_5_613(.a(output_6_613), .b(output_6_6), .y(output_5_613));
wire output_7_613, output_7_6, output_6_613;
mixer gate_output_6_613(.a(output_7_613), .b(output_7_6), .y(output_6_613));
wire output_8_613, output_8_6, output_7_613;
mixer gate_output_7_613(.a(output_8_613), .b(output_8_6), .y(output_7_613));
wire output_9_613, output_9_6, output_8_613;
mixer gate_output_8_613(.a(output_9_613), .b(output_9_6), .y(output_8_613));
wire output_10_613, output_10_6, output_9_613;
mixer gate_output_9_613(.a(output_10_613), .b(output_10_6), .y(output_9_613));
wire output_11_613, output_11_6, output_10_613;
mixer gate_output_10_613(.a(output_11_613), .b(output_11_6), .y(output_10_613));
wire output_12_613, output_12_6, output_11_613;
mixer gate_output_11_613(.a(output_12_613), .b(output_12_6), .y(output_11_613));
wire output_13_613, output_13_6, output_12_613;
mixer gate_output_12_613(.a(output_13_613), .b(output_13_6), .y(output_12_613));
wire output_14_613, output_14_6, output_13_613;
mixer gate_output_13_613(.a(output_14_613), .b(output_14_6), .y(output_13_613));
wire output_15_613, output_15_6, output_14_613;
mixer gate_output_14_613(.a(output_15_613), .b(output_15_6), .y(output_14_613));
wire output_16_613, output_16_6, output_15_613;
mixer gate_output_15_613(.a(output_16_613), .b(output_16_6), .y(output_15_613));
wire output_1_614, output_1_7, output_0_614;
mixer gate_output_0_614(.a(output_1_614), .b(output_1_7), .y(output_0_614));
wire output_2_614, output_2_7, output_1_614;
mixer gate_output_1_614(.a(output_2_614), .b(output_2_7), .y(output_1_614));
wire output_3_614, output_3_7, output_2_614;
mixer gate_output_2_614(.a(output_3_614), .b(output_3_7), .y(output_2_614));
wire output_4_614, output_4_7, output_3_614;
mixer gate_output_3_614(.a(output_4_614), .b(output_4_7), .y(output_3_614));
wire output_5_614, output_5_7, output_4_614;
mixer gate_output_4_614(.a(output_5_614), .b(output_5_7), .y(output_4_614));
wire output_6_614, output_6_7, output_5_614;
mixer gate_output_5_614(.a(output_6_614), .b(output_6_7), .y(output_5_614));
wire output_7_614, output_7_7, output_6_614;
mixer gate_output_6_614(.a(output_7_614), .b(output_7_7), .y(output_6_614));
wire output_8_614, output_8_7, output_7_614;
mixer gate_output_7_614(.a(output_8_614), .b(output_8_7), .y(output_7_614));
wire output_9_614, output_9_7, output_8_614;
mixer gate_output_8_614(.a(output_9_614), .b(output_9_7), .y(output_8_614));
wire output_10_614, output_10_7, output_9_614;
mixer gate_output_9_614(.a(output_10_614), .b(output_10_7), .y(output_9_614));
wire output_11_614, output_11_7, output_10_614;
mixer gate_output_10_614(.a(output_11_614), .b(output_11_7), .y(output_10_614));
wire output_12_614, output_12_7, output_11_614;
mixer gate_output_11_614(.a(output_12_614), .b(output_12_7), .y(output_11_614));
wire output_13_614, output_13_7, output_12_614;
mixer gate_output_12_614(.a(output_13_614), .b(output_13_7), .y(output_12_614));
wire output_14_614, output_14_7, output_13_614;
mixer gate_output_13_614(.a(output_14_614), .b(output_14_7), .y(output_13_614));
wire output_15_614, output_15_7, output_14_614;
mixer gate_output_14_614(.a(output_15_614), .b(output_15_7), .y(output_14_614));
wire output_16_614, output_16_7, output_15_614;
mixer gate_output_15_614(.a(output_16_614), .b(output_16_7), .y(output_15_614));
wire output_1_615, output_1_8, output_0_615;
mixer gate_output_0_615(.a(output_1_615), .b(output_1_8), .y(output_0_615));
wire output_2_615, output_2_8, output_1_615;
mixer gate_output_1_615(.a(output_2_615), .b(output_2_8), .y(output_1_615));
wire output_3_615, output_3_8, output_2_615;
mixer gate_output_2_615(.a(output_3_615), .b(output_3_8), .y(output_2_615));
wire output_4_615, output_4_8, output_3_615;
mixer gate_output_3_615(.a(output_4_615), .b(output_4_8), .y(output_3_615));
wire output_5_615, output_5_8, output_4_615;
mixer gate_output_4_615(.a(output_5_615), .b(output_5_8), .y(output_4_615));
wire output_6_615, output_6_8, output_5_615;
mixer gate_output_5_615(.a(output_6_615), .b(output_6_8), .y(output_5_615));
wire output_7_615, output_7_8, output_6_615;
mixer gate_output_6_615(.a(output_7_615), .b(output_7_8), .y(output_6_615));
wire output_8_615, output_8_8, output_7_615;
mixer gate_output_7_615(.a(output_8_615), .b(output_8_8), .y(output_7_615));
wire output_9_615, output_9_8, output_8_615;
mixer gate_output_8_615(.a(output_9_615), .b(output_9_8), .y(output_8_615));
wire output_10_615, output_10_8, output_9_615;
mixer gate_output_9_615(.a(output_10_615), .b(output_10_8), .y(output_9_615));
wire output_11_615, output_11_8, output_10_615;
mixer gate_output_10_615(.a(output_11_615), .b(output_11_8), .y(output_10_615));
wire output_12_615, output_12_8, output_11_615;
mixer gate_output_11_615(.a(output_12_615), .b(output_12_8), .y(output_11_615));
wire output_13_615, output_13_8, output_12_615;
mixer gate_output_12_615(.a(output_13_615), .b(output_13_8), .y(output_12_615));
wire output_14_615, output_14_8, output_13_615;
mixer gate_output_13_615(.a(output_14_615), .b(output_14_8), .y(output_13_615));
wire output_15_615, output_15_8, output_14_615;
mixer gate_output_14_615(.a(output_15_615), .b(output_15_8), .y(output_14_615));
wire output_16_615, output_16_8, output_15_615;
mixer gate_output_15_615(.a(output_16_615), .b(output_16_8), .y(output_15_615));
wire output_1_616, output_1_9, output_0_616;
mixer gate_output_0_616(.a(output_1_616), .b(output_1_9), .y(output_0_616));
wire output_2_616, output_2_9, output_1_616;
mixer gate_output_1_616(.a(output_2_616), .b(output_2_9), .y(output_1_616));
wire output_3_616, output_3_9, output_2_616;
mixer gate_output_2_616(.a(output_3_616), .b(output_3_9), .y(output_2_616));
wire output_4_616, output_4_9, output_3_616;
mixer gate_output_3_616(.a(output_4_616), .b(output_4_9), .y(output_3_616));
wire output_5_616, output_5_9, output_4_616;
mixer gate_output_4_616(.a(output_5_616), .b(output_5_9), .y(output_4_616));
wire output_6_616, output_6_9, output_5_616;
mixer gate_output_5_616(.a(output_6_616), .b(output_6_9), .y(output_5_616));
wire output_7_616, output_7_9, output_6_616;
mixer gate_output_6_616(.a(output_7_616), .b(output_7_9), .y(output_6_616));
wire output_8_616, output_8_9, output_7_616;
mixer gate_output_7_616(.a(output_8_616), .b(output_8_9), .y(output_7_616));
wire output_9_616, output_9_9, output_8_616;
mixer gate_output_8_616(.a(output_9_616), .b(output_9_9), .y(output_8_616));
wire output_10_616, output_10_9, output_9_616;
mixer gate_output_9_616(.a(output_10_616), .b(output_10_9), .y(output_9_616));
wire output_11_616, output_11_9, output_10_616;
mixer gate_output_10_616(.a(output_11_616), .b(output_11_9), .y(output_10_616));
wire output_12_616, output_12_9, output_11_616;
mixer gate_output_11_616(.a(output_12_616), .b(output_12_9), .y(output_11_616));
wire output_13_616, output_13_9, output_12_616;
mixer gate_output_12_616(.a(output_13_616), .b(output_13_9), .y(output_12_616));
wire output_14_616, output_14_9, output_13_616;
mixer gate_output_13_616(.a(output_14_616), .b(output_14_9), .y(output_13_616));
wire output_15_616, output_15_9, output_14_616;
mixer gate_output_14_616(.a(output_15_616), .b(output_15_9), .y(output_14_616));
wire output_16_616, output_16_9, output_15_616;
mixer gate_output_15_616(.a(output_16_616), .b(output_16_9), .y(output_15_616));
wire output_1_617, output_1_10, output_0_617;
mixer gate_output_0_617(.a(output_1_617), .b(output_1_10), .y(output_0_617));
wire output_2_617, output_2_10, output_1_617;
mixer gate_output_1_617(.a(output_2_617), .b(output_2_10), .y(output_1_617));
wire output_3_617, output_3_10, output_2_617;
mixer gate_output_2_617(.a(output_3_617), .b(output_3_10), .y(output_2_617));
wire output_4_617, output_4_10, output_3_617;
mixer gate_output_3_617(.a(output_4_617), .b(output_4_10), .y(output_3_617));
wire output_5_617, output_5_10, output_4_617;
mixer gate_output_4_617(.a(output_5_617), .b(output_5_10), .y(output_4_617));
wire output_6_617, output_6_10, output_5_617;
mixer gate_output_5_617(.a(output_6_617), .b(output_6_10), .y(output_5_617));
wire output_7_617, output_7_10, output_6_617;
mixer gate_output_6_617(.a(output_7_617), .b(output_7_10), .y(output_6_617));
wire output_8_617, output_8_10, output_7_617;
mixer gate_output_7_617(.a(output_8_617), .b(output_8_10), .y(output_7_617));
wire output_9_617, output_9_10, output_8_617;
mixer gate_output_8_617(.a(output_9_617), .b(output_9_10), .y(output_8_617));
wire output_10_617, output_10_10, output_9_617;
mixer gate_output_9_617(.a(output_10_617), .b(output_10_10), .y(output_9_617));
wire output_11_617, output_11_10, output_10_617;
mixer gate_output_10_617(.a(output_11_617), .b(output_11_10), .y(output_10_617));
wire output_12_617, output_12_10, output_11_617;
mixer gate_output_11_617(.a(output_12_617), .b(output_12_10), .y(output_11_617));
wire output_13_617, output_13_10, output_12_617;
mixer gate_output_12_617(.a(output_13_617), .b(output_13_10), .y(output_12_617));
wire output_14_617, output_14_10, output_13_617;
mixer gate_output_13_617(.a(output_14_617), .b(output_14_10), .y(output_13_617));
wire output_15_617, output_15_10, output_14_617;
mixer gate_output_14_617(.a(output_15_617), .b(output_15_10), .y(output_14_617));
wire output_16_617, output_16_10, output_15_617;
mixer gate_output_15_617(.a(output_16_617), .b(output_16_10), .y(output_15_617));
wire output_1_618, output_1_11, output_0_618;
mixer gate_output_0_618(.a(output_1_618), .b(output_1_11), .y(output_0_618));
wire output_2_618, output_2_11, output_1_618;
mixer gate_output_1_618(.a(output_2_618), .b(output_2_11), .y(output_1_618));
wire output_3_618, output_3_11, output_2_618;
mixer gate_output_2_618(.a(output_3_618), .b(output_3_11), .y(output_2_618));
wire output_4_618, output_4_11, output_3_618;
mixer gate_output_3_618(.a(output_4_618), .b(output_4_11), .y(output_3_618));
wire output_5_618, output_5_11, output_4_618;
mixer gate_output_4_618(.a(output_5_618), .b(output_5_11), .y(output_4_618));
wire output_6_618, output_6_11, output_5_618;
mixer gate_output_5_618(.a(output_6_618), .b(output_6_11), .y(output_5_618));
wire output_7_618, output_7_11, output_6_618;
mixer gate_output_6_618(.a(output_7_618), .b(output_7_11), .y(output_6_618));
wire output_8_618, output_8_11, output_7_618;
mixer gate_output_7_618(.a(output_8_618), .b(output_8_11), .y(output_7_618));
wire output_9_618, output_9_11, output_8_618;
mixer gate_output_8_618(.a(output_9_618), .b(output_9_11), .y(output_8_618));
wire output_10_618, output_10_11, output_9_618;
mixer gate_output_9_618(.a(output_10_618), .b(output_10_11), .y(output_9_618));
wire output_11_618, output_11_11, output_10_618;
mixer gate_output_10_618(.a(output_11_618), .b(output_11_11), .y(output_10_618));
wire output_12_618, output_12_11, output_11_618;
mixer gate_output_11_618(.a(output_12_618), .b(output_12_11), .y(output_11_618));
wire output_13_618, output_13_11, output_12_618;
mixer gate_output_12_618(.a(output_13_618), .b(output_13_11), .y(output_12_618));
wire output_14_618, output_14_11, output_13_618;
mixer gate_output_13_618(.a(output_14_618), .b(output_14_11), .y(output_13_618));
wire output_15_618, output_15_11, output_14_618;
mixer gate_output_14_618(.a(output_15_618), .b(output_15_11), .y(output_14_618));
wire output_16_618, output_16_11, output_15_618;
mixer gate_output_15_618(.a(output_16_618), .b(output_16_11), .y(output_15_618));
wire output_1_619, output_1_12, output_0_619;
mixer gate_output_0_619(.a(output_1_619), .b(output_1_12), .y(output_0_619));
wire output_2_619, output_2_12, output_1_619;
mixer gate_output_1_619(.a(output_2_619), .b(output_2_12), .y(output_1_619));
wire output_3_619, output_3_12, output_2_619;
mixer gate_output_2_619(.a(output_3_619), .b(output_3_12), .y(output_2_619));
wire output_4_619, output_4_12, output_3_619;
mixer gate_output_3_619(.a(output_4_619), .b(output_4_12), .y(output_3_619));
wire output_5_619, output_5_12, output_4_619;
mixer gate_output_4_619(.a(output_5_619), .b(output_5_12), .y(output_4_619));
wire output_6_619, output_6_12, output_5_619;
mixer gate_output_5_619(.a(output_6_619), .b(output_6_12), .y(output_5_619));
wire output_7_619, output_7_12, output_6_619;
mixer gate_output_6_619(.a(output_7_619), .b(output_7_12), .y(output_6_619));
wire output_8_619, output_8_12, output_7_619;
mixer gate_output_7_619(.a(output_8_619), .b(output_8_12), .y(output_7_619));
wire output_9_619, output_9_12, output_8_619;
mixer gate_output_8_619(.a(output_9_619), .b(output_9_12), .y(output_8_619));
wire output_10_619, output_10_12, output_9_619;
mixer gate_output_9_619(.a(output_10_619), .b(output_10_12), .y(output_9_619));
wire output_11_619, output_11_12, output_10_619;
mixer gate_output_10_619(.a(output_11_619), .b(output_11_12), .y(output_10_619));
wire output_12_619, output_12_12, output_11_619;
mixer gate_output_11_619(.a(output_12_619), .b(output_12_12), .y(output_11_619));
wire output_13_619, output_13_12, output_12_619;
mixer gate_output_12_619(.a(output_13_619), .b(output_13_12), .y(output_12_619));
wire output_14_619, output_14_12, output_13_619;
mixer gate_output_13_619(.a(output_14_619), .b(output_14_12), .y(output_13_619));
wire output_15_619, output_15_12, output_14_619;
mixer gate_output_14_619(.a(output_15_619), .b(output_15_12), .y(output_14_619));
wire output_16_619, output_16_12, output_15_619;
mixer gate_output_15_619(.a(output_16_619), .b(output_16_12), .y(output_15_619));
wire output_1_620, output_1_13, output_0_620;
mixer gate_output_0_620(.a(output_1_620), .b(output_1_13), .y(output_0_620));
wire output_2_620, output_2_13, output_1_620;
mixer gate_output_1_620(.a(output_2_620), .b(output_2_13), .y(output_1_620));
wire output_3_620, output_3_13, output_2_620;
mixer gate_output_2_620(.a(output_3_620), .b(output_3_13), .y(output_2_620));
wire output_4_620, output_4_13, output_3_620;
mixer gate_output_3_620(.a(output_4_620), .b(output_4_13), .y(output_3_620));
wire output_5_620, output_5_13, output_4_620;
mixer gate_output_4_620(.a(output_5_620), .b(output_5_13), .y(output_4_620));
wire output_6_620, output_6_13, output_5_620;
mixer gate_output_5_620(.a(output_6_620), .b(output_6_13), .y(output_5_620));
wire output_7_620, output_7_13, output_6_620;
mixer gate_output_6_620(.a(output_7_620), .b(output_7_13), .y(output_6_620));
wire output_8_620, output_8_13, output_7_620;
mixer gate_output_7_620(.a(output_8_620), .b(output_8_13), .y(output_7_620));
wire output_9_620, output_9_13, output_8_620;
mixer gate_output_8_620(.a(output_9_620), .b(output_9_13), .y(output_8_620));
wire output_10_620, output_10_13, output_9_620;
mixer gate_output_9_620(.a(output_10_620), .b(output_10_13), .y(output_9_620));
wire output_11_620, output_11_13, output_10_620;
mixer gate_output_10_620(.a(output_11_620), .b(output_11_13), .y(output_10_620));
wire output_12_620, output_12_13, output_11_620;
mixer gate_output_11_620(.a(output_12_620), .b(output_12_13), .y(output_11_620));
wire output_13_620, output_13_13, output_12_620;
mixer gate_output_12_620(.a(output_13_620), .b(output_13_13), .y(output_12_620));
wire output_14_620, output_14_13, output_13_620;
mixer gate_output_13_620(.a(output_14_620), .b(output_14_13), .y(output_13_620));
wire output_15_620, output_15_13, output_14_620;
mixer gate_output_14_620(.a(output_15_620), .b(output_15_13), .y(output_14_620));
wire output_16_620, output_16_13, output_15_620;
mixer gate_output_15_620(.a(output_16_620), .b(output_16_13), .y(output_15_620));
wire output_1_621, output_1_14, output_0_621;
mixer gate_output_0_621(.a(output_1_621), .b(output_1_14), .y(output_0_621));
wire output_2_621, output_2_14, output_1_621;
mixer gate_output_1_621(.a(output_2_621), .b(output_2_14), .y(output_1_621));
wire output_3_621, output_3_14, output_2_621;
mixer gate_output_2_621(.a(output_3_621), .b(output_3_14), .y(output_2_621));
wire output_4_621, output_4_14, output_3_621;
mixer gate_output_3_621(.a(output_4_621), .b(output_4_14), .y(output_3_621));
wire output_5_621, output_5_14, output_4_621;
mixer gate_output_4_621(.a(output_5_621), .b(output_5_14), .y(output_4_621));
wire output_6_621, output_6_14, output_5_621;
mixer gate_output_5_621(.a(output_6_621), .b(output_6_14), .y(output_5_621));
wire output_7_621, output_7_14, output_6_621;
mixer gate_output_6_621(.a(output_7_621), .b(output_7_14), .y(output_6_621));
wire output_8_621, output_8_14, output_7_621;
mixer gate_output_7_621(.a(output_8_621), .b(output_8_14), .y(output_7_621));
wire output_9_621, output_9_14, output_8_621;
mixer gate_output_8_621(.a(output_9_621), .b(output_9_14), .y(output_8_621));
wire output_10_621, output_10_14, output_9_621;
mixer gate_output_9_621(.a(output_10_621), .b(output_10_14), .y(output_9_621));
wire output_11_621, output_11_14, output_10_621;
mixer gate_output_10_621(.a(output_11_621), .b(output_11_14), .y(output_10_621));
wire output_12_621, output_12_14, output_11_621;
mixer gate_output_11_621(.a(output_12_621), .b(output_12_14), .y(output_11_621));
wire output_13_621, output_13_14, output_12_621;
mixer gate_output_12_621(.a(output_13_621), .b(output_13_14), .y(output_12_621));
wire output_14_621, output_14_14, output_13_621;
mixer gate_output_13_621(.a(output_14_621), .b(output_14_14), .y(output_13_621));
wire output_15_621, output_15_14, output_14_621;
mixer gate_output_14_621(.a(output_15_621), .b(output_15_14), .y(output_14_621));
wire output_16_621, output_16_14, output_15_621;
mixer gate_output_15_621(.a(output_16_621), .b(output_16_14), .y(output_15_621));
wire output_1_622, output_1_15, output_0_622;
mixer gate_output_0_622(.a(output_1_622), .b(output_1_15), .y(output_0_622));
wire output_2_622, output_2_15, output_1_622;
mixer gate_output_1_622(.a(output_2_622), .b(output_2_15), .y(output_1_622));
wire output_3_622, output_3_15, output_2_622;
mixer gate_output_2_622(.a(output_3_622), .b(output_3_15), .y(output_2_622));
wire output_4_622, output_4_15, output_3_622;
mixer gate_output_3_622(.a(output_4_622), .b(output_4_15), .y(output_3_622));
wire output_5_622, output_5_15, output_4_622;
mixer gate_output_4_622(.a(output_5_622), .b(output_5_15), .y(output_4_622));
wire output_6_622, output_6_15, output_5_622;
mixer gate_output_5_622(.a(output_6_622), .b(output_6_15), .y(output_5_622));
wire output_7_622, output_7_15, output_6_622;
mixer gate_output_6_622(.a(output_7_622), .b(output_7_15), .y(output_6_622));
wire output_8_622, output_8_15, output_7_622;
mixer gate_output_7_622(.a(output_8_622), .b(output_8_15), .y(output_7_622));
wire output_9_622, output_9_15, output_8_622;
mixer gate_output_8_622(.a(output_9_622), .b(output_9_15), .y(output_8_622));
wire output_10_622, output_10_15, output_9_622;
mixer gate_output_9_622(.a(output_10_622), .b(output_10_15), .y(output_9_622));
wire output_11_622, output_11_15, output_10_622;
mixer gate_output_10_622(.a(output_11_622), .b(output_11_15), .y(output_10_622));
wire output_12_622, output_12_15, output_11_622;
mixer gate_output_11_622(.a(output_12_622), .b(output_12_15), .y(output_11_622));
wire output_13_622, output_13_15, output_12_622;
mixer gate_output_12_622(.a(output_13_622), .b(output_13_15), .y(output_12_622));
wire output_14_622, output_14_15, output_13_622;
mixer gate_output_13_622(.a(output_14_622), .b(output_14_15), .y(output_13_622));
wire output_15_622, output_15_15, output_14_622;
mixer gate_output_14_622(.a(output_15_622), .b(output_15_15), .y(output_14_622));
wire output_16_622, output_16_15, output_15_622;
mixer gate_output_15_622(.a(output_16_622), .b(output_16_15), .y(output_15_622));
wire output_1_623, output_1_0, output_0_623;
mixer gate_output_0_623(.a(output_1_623), .b(output_1_0), .y(output_0_623));
wire output_2_623, output_2_0, output_1_623;
mixer gate_output_1_623(.a(output_2_623), .b(output_2_0), .y(output_1_623));
wire output_3_623, output_3_0, output_2_623;
mixer gate_output_2_623(.a(output_3_623), .b(output_3_0), .y(output_2_623));
wire output_4_623, output_4_0, output_3_623;
mixer gate_output_3_623(.a(output_4_623), .b(output_4_0), .y(output_3_623));
wire output_5_623, output_5_0, output_4_623;
mixer gate_output_4_623(.a(output_5_623), .b(output_5_0), .y(output_4_623));
wire output_6_623, output_6_0, output_5_623;
mixer gate_output_5_623(.a(output_6_623), .b(output_6_0), .y(output_5_623));
wire output_7_623, output_7_0, output_6_623;
mixer gate_output_6_623(.a(output_7_623), .b(output_7_0), .y(output_6_623));
wire output_8_623, output_8_0, output_7_623;
mixer gate_output_7_623(.a(output_8_623), .b(output_8_0), .y(output_7_623));
wire output_9_623, output_9_0, output_8_623;
mixer gate_output_8_623(.a(output_9_623), .b(output_9_0), .y(output_8_623));
wire output_10_623, output_10_0, output_9_623;
mixer gate_output_9_623(.a(output_10_623), .b(output_10_0), .y(output_9_623));
wire output_11_623, output_11_0, output_10_623;
mixer gate_output_10_623(.a(output_11_623), .b(output_11_0), .y(output_10_623));
wire output_12_623, output_12_0, output_11_623;
mixer gate_output_11_623(.a(output_12_623), .b(output_12_0), .y(output_11_623));
wire output_13_623, output_13_0, output_12_623;
mixer gate_output_12_623(.a(output_13_623), .b(output_13_0), .y(output_12_623));
wire output_14_623, output_14_0, output_13_623;
mixer gate_output_13_623(.a(output_14_623), .b(output_14_0), .y(output_13_623));
wire output_15_623, output_15_0, output_14_623;
mixer gate_output_14_623(.a(output_15_623), .b(output_15_0), .y(output_14_623));
wire output_16_623, output_16_0, output_15_623;
mixer gate_output_15_623(.a(output_16_623), .b(output_16_0), .y(output_15_623));
wire output_1_624, output_1_1, output_0_624;
mixer gate_output_0_624(.a(output_1_624), .b(output_1_1), .y(output_0_624));
wire output_2_624, output_2_1, output_1_624;
mixer gate_output_1_624(.a(output_2_624), .b(output_2_1), .y(output_1_624));
wire output_3_624, output_3_1, output_2_624;
mixer gate_output_2_624(.a(output_3_624), .b(output_3_1), .y(output_2_624));
wire output_4_624, output_4_1, output_3_624;
mixer gate_output_3_624(.a(output_4_624), .b(output_4_1), .y(output_3_624));
wire output_5_624, output_5_1, output_4_624;
mixer gate_output_4_624(.a(output_5_624), .b(output_5_1), .y(output_4_624));
wire output_6_624, output_6_1, output_5_624;
mixer gate_output_5_624(.a(output_6_624), .b(output_6_1), .y(output_5_624));
wire output_7_624, output_7_1, output_6_624;
mixer gate_output_6_624(.a(output_7_624), .b(output_7_1), .y(output_6_624));
wire output_8_624, output_8_1, output_7_624;
mixer gate_output_7_624(.a(output_8_624), .b(output_8_1), .y(output_7_624));
wire output_9_624, output_9_1, output_8_624;
mixer gate_output_8_624(.a(output_9_624), .b(output_9_1), .y(output_8_624));
wire output_10_624, output_10_1, output_9_624;
mixer gate_output_9_624(.a(output_10_624), .b(output_10_1), .y(output_9_624));
wire output_11_624, output_11_1, output_10_624;
mixer gate_output_10_624(.a(output_11_624), .b(output_11_1), .y(output_10_624));
wire output_12_624, output_12_1, output_11_624;
mixer gate_output_11_624(.a(output_12_624), .b(output_12_1), .y(output_11_624));
wire output_13_624, output_13_1, output_12_624;
mixer gate_output_12_624(.a(output_13_624), .b(output_13_1), .y(output_12_624));
wire output_14_624, output_14_1, output_13_624;
mixer gate_output_13_624(.a(output_14_624), .b(output_14_1), .y(output_13_624));
wire output_15_624, output_15_1, output_14_624;
mixer gate_output_14_624(.a(output_15_624), .b(output_15_1), .y(output_14_624));
wire output_16_624, output_16_1, output_15_624;
mixer gate_output_15_624(.a(output_16_624), .b(output_16_1), .y(output_15_624));
wire output_1_625, output_1_2, output_0_625;
mixer gate_output_0_625(.a(output_1_625), .b(output_1_2), .y(output_0_625));
wire output_2_625, output_2_2, output_1_625;
mixer gate_output_1_625(.a(output_2_625), .b(output_2_2), .y(output_1_625));
wire output_3_625, output_3_2, output_2_625;
mixer gate_output_2_625(.a(output_3_625), .b(output_3_2), .y(output_2_625));
wire output_4_625, output_4_2, output_3_625;
mixer gate_output_3_625(.a(output_4_625), .b(output_4_2), .y(output_3_625));
wire output_5_625, output_5_2, output_4_625;
mixer gate_output_4_625(.a(output_5_625), .b(output_5_2), .y(output_4_625));
wire output_6_625, output_6_2, output_5_625;
mixer gate_output_5_625(.a(output_6_625), .b(output_6_2), .y(output_5_625));
wire output_7_625, output_7_2, output_6_625;
mixer gate_output_6_625(.a(output_7_625), .b(output_7_2), .y(output_6_625));
wire output_8_625, output_8_2, output_7_625;
mixer gate_output_7_625(.a(output_8_625), .b(output_8_2), .y(output_7_625));
wire output_9_625, output_9_2, output_8_625;
mixer gate_output_8_625(.a(output_9_625), .b(output_9_2), .y(output_8_625));
wire output_10_625, output_10_2, output_9_625;
mixer gate_output_9_625(.a(output_10_625), .b(output_10_2), .y(output_9_625));
wire output_11_625, output_11_2, output_10_625;
mixer gate_output_10_625(.a(output_11_625), .b(output_11_2), .y(output_10_625));
wire output_12_625, output_12_2, output_11_625;
mixer gate_output_11_625(.a(output_12_625), .b(output_12_2), .y(output_11_625));
wire output_13_625, output_13_2, output_12_625;
mixer gate_output_12_625(.a(output_13_625), .b(output_13_2), .y(output_12_625));
wire output_14_625, output_14_2, output_13_625;
mixer gate_output_13_625(.a(output_14_625), .b(output_14_2), .y(output_13_625));
wire output_15_625, output_15_2, output_14_625;
mixer gate_output_14_625(.a(output_15_625), .b(output_15_2), .y(output_14_625));
wire output_16_625, output_16_2, output_15_625;
mixer gate_output_15_625(.a(output_16_625), .b(output_16_2), .y(output_15_625));
wire output_1_626, output_1_3, output_0_626;
mixer gate_output_0_626(.a(output_1_626), .b(output_1_3), .y(output_0_626));
wire output_2_626, output_2_3, output_1_626;
mixer gate_output_1_626(.a(output_2_626), .b(output_2_3), .y(output_1_626));
wire output_3_626, output_3_3, output_2_626;
mixer gate_output_2_626(.a(output_3_626), .b(output_3_3), .y(output_2_626));
wire output_4_626, output_4_3, output_3_626;
mixer gate_output_3_626(.a(output_4_626), .b(output_4_3), .y(output_3_626));
wire output_5_626, output_5_3, output_4_626;
mixer gate_output_4_626(.a(output_5_626), .b(output_5_3), .y(output_4_626));
wire output_6_626, output_6_3, output_5_626;
mixer gate_output_5_626(.a(output_6_626), .b(output_6_3), .y(output_5_626));
wire output_7_626, output_7_3, output_6_626;
mixer gate_output_6_626(.a(output_7_626), .b(output_7_3), .y(output_6_626));
wire output_8_626, output_8_3, output_7_626;
mixer gate_output_7_626(.a(output_8_626), .b(output_8_3), .y(output_7_626));
wire output_9_626, output_9_3, output_8_626;
mixer gate_output_8_626(.a(output_9_626), .b(output_9_3), .y(output_8_626));
wire output_10_626, output_10_3, output_9_626;
mixer gate_output_9_626(.a(output_10_626), .b(output_10_3), .y(output_9_626));
wire output_11_626, output_11_3, output_10_626;
mixer gate_output_10_626(.a(output_11_626), .b(output_11_3), .y(output_10_626));
wire output_12_626, output_12_3, output_11_626;
mixer gate_output_11_626(.a(output_12_626), .b(output_12_3), .y(output_11_626));
wire output_13_626, output_13_3, output_12_626;
mixer gate_output_12_626(.a(output_13_626), .b(output_13_3), .y(output_12_626));
wire output_14_626, output_14_3, output_13_626;
mixer gate_output_13_626(.a(output_14_626), .b(output_14_3), .y(output_13_626));
wire output_15_626, output_15_3, output_14_626;
mixer gate_output_14_626(.a(output_15_626), .b(output_15_3), .y(output_14_626));
wire output_16_626, output_16_3, output_15_626;
mixer gate_output_15_626(.a(output_16_626), .b(output_16_3), .y(output_15_626));
wire output_1_627, output_1_4, output_0_627;
mixer gate_output_0_627(.a(output_1_627), .b(output_1_4), .y(output_0_627));
wire output_2_627, output_2_4, output_1_627;
mixer gate_output_1_627(.a(output_2_627), .b(output_2_4), .y(output_1_627));
wire output_3_627, output_3_4, output_2_627;
mixer gate_output_2_627(.a(output_3_627), .b(output_3_4), .y(output_2_627));
wire output_4_627, output_4_4, output_3_627;
mixer gate_output_3_627(.a(output_4_627), .b(output_4_4), .y(output_3_627));
wire output_5_627, output_5_4, output_4_627;
mixer gate_output_4_627(.a(output_5_627), .b(output_5_4), .y(output_4_627));
wire output_6_627, output_6_4, output_5_627;
mixer gate_output_5_627(.a(output_6_627), .b(output_6_4), .y(output_5_627));
wire output_7_627, output_7_4, output_6_627;
mixer gate_output_6_627(.a(output_7_627), .b(output_7_4), .y(output_6_627));
wire output_8_627, output_8_4, output_7_627;
mixer gate_output_7_627(.a(output_8_627), .b(output_8_4), .y(output_7_627));
wire output_9_627, output_9_4, output_8_627;
mixer gate_output_8_627(.a(output_9_627), .b(output_9_4), .y(output_8_627));
wire output_10_627, output_10_4, output_9_627;
mixer gate_output_9_627(.a(output_10_627), .b(output_10_4), .y(output_9_627));
wire output_11_627, output_11_4, output_10_627;
mixer gate_output_10_627(.a(output_11_627), .b(output_11_4), .y(output_10_627));
wire output_12_627, output_12_4, output_11_627;
mixer gate_output_11_627(.a(output_12_627), .b(output_12_4), .y(output_11_627));
wire output_13_627, output_13_4, output_12_627;
mixer gate_output_12_627(.a(output_13_627), .b(output_13_4), .y(output_12_627));
wire output_14_627, output_14_4, output_13_627;
mixer gate_output_13_627(.a(output_14_627), .b(output_14_4), .y(output_13_627));
wire output_15_627, output_15_4, output_14_627;
mixer gate_output_14_627(.a(output_15_627), .b(output_15_4), .y(output_14_627));
wire output_16_627, output_16_4, output_15_627;
mixer gate_output_15_627(.a(output_16_627), .b(output_16_4), .y(output_15_627));
wire output_1_628, output_1_5, output_0_628;
mixer gate_output_0_628(.a(output_1_628), .b(output_1_5), .y(output_0_628));
wire output_2_628, output_2_5, output_1_628;
mixer gate_output_1_628(.a(output_2_628), .b(output_2_5), .y(output_1_628));
wire output_3_628, output_3_5, output_2_628;
mixer gate_output_2_628(.a(output_3_628), .b(output_3_5), .y(output_2_628));
wire output_4_628, output_4_5, output_3_628;
mixer gate_output_3_628(.a(output_4_628), .b(output_4_5), .y(output_3_628));
wire output_5_628, output_5_5, output_4_628;
mixer gate_output_4_628(.a(output_5_628), .b(output_5_5), .y(output_4_628));
wire output_6_628, output_6_5, output_5_628;
mixer gate_output_5_628(.a(output_6_628), .b(output_6_5), .y(output_5_628));
wire output_7_628, output_7_5, output_6_628;
mixer gate_output_6_628(.a(output_7_628), .b(output_7_5), .y(output_6_628));
wire output_8_628, output_8_5, output_7_628;
mixer gate_output_7_628(.a(output_8_628), .b(output_8_5), .y(output_7_628));
wire output_9_628, output_9_5, output_8_628;
mixer gate_output_8_628(.a(output_9_628), .b(output_9_5), .y(output_8_628));
wire output_10_628, output_10_5, output_9_628;
mixer gate_output_9_628(.a(output_10_628), .b(output_10_5), .y(output_9_628));
wire output_11_628, output_11_5, output_10_628;
mixer gate_output_10_628(.a(output_11_628), .b(output_11_5), .y(output_10_628));
wire output_12_628, output_12_5, output_11_628;
mixer gate_output_11_628(.a(output_12_628), .b(output_12_5), .y(output_11_628));
wire output_13_628, output_13_5, output_12_628;
mixer gate_output_12_628(.a(output_13_628), .b(output_13_5), .y(output_12_628));
wire output_14_628, output_14_5, output_13_628;
mixer gate_output_13_628(.a(output_14_628), .b(output_14_5), .y(output_13_628));
wire output_15_628, output_15_5, output_14_628;
mixer gate_output_14_628(.a(output_15_628), .b(output_15_5), .y(output_14_628));
wire output_16_628, output_16_5, output_15_628;
mixer gate_output_15_628(.a(output_16_628), .b(output_16_5), .y(output_15_628));
wire output_1_629, output_1_6, output_0_629;
mixer gate_output_0_629(.a(output_1_629), .b(output_1_6), .y(output_0_629));
wire output_2_629, output_2_6, output_1_629;
mixer gate_output_1_629(.a(output_2_629), .b(output_2_6), .y(output_1_629));
wire output_3_629, output_3_6, output_2_629;
mixer gate_output_2_629(.a(output_3_629), .b(output_3_6), .y(output_2_629));
wire output_4_629, output_4_6, output_3_629;
mixer gate_output_3_629(.a(output_4_629), .b(output_4_6), .y(output_3_629));
wire output_5_629, output_5_6, output_4_629;
mixer gate_output_4_629(.a(output_5_629), .b(output_5_6), .y(output_4_629));
wire output_6_629, output_6_6, output_5_629;
mixer gate_output_5_629(.a(output_6_629), .b(output_6_6), .y(output_5_629));
wire output_7_629, output_7_6, output_6_629;
mixer gate_output_6_629(.a(output_7_629), .b(output_7_6), .y(output_6_629));
wire output_8_629, output_8_6, output_7_629;
mixer gate_output_7_629(.a(output_8_629), .b(output_8_6), .y(output_7_629));
wire output_9_629, output_9_6, output_8_629;
mixer gate_output_8_629(.a(output_9_629), .b(output_9_6), .y(output_8_629));
wire output_10_629, output_10_6, output_9_629;
mixer gate_output_9_629(.a(output_10_629), .b(output_10_6), .y(output_9_629));
wire output_11_629, output_11_6, output_10_629;
mixer gate_output_10_629(.a(output_11_629), .b(output_11_6), .y(output_10_629));
wire output_12_629, output_12_6, output_11_629;
mixer gate_output_11_629(.a(output_12_629), .b(output_12_6), .y(output_11_629));
wire output_13_629, output_13_6, output_12_629;
mixer gate_output_12_629(.a(output_13_629), .b(output_13_6), .y(output_12_629));
wire output_14_629, output_14_6, output_13_629;
mixer gate_output_13_629(.a(output_14_629), .b(output_14_6), .y(output_13_629));
wire output_15_629, output_15_6, output_14_629;
mixer gate_output_14_629(.a(output_15_629), .b(output_15_6), .y(output_14_629));
wire output_16_629, output_16_6, output_15_629;
mixer gate_output_15_629(.a(output_16_629), .b(output_16_6), .y(output_15_629));
wire output_1_630, output_1_7, output_0_630;
mixer gate_output_0_630(.a(output_1_630), .b(output_1_7), .y(output_0_630));
wire output_2_630, output_2_7, output_1_630;
mixer gate_output_1_630(.a(output_2_630), .b(output_2_7), .y(output_1_630));
wire output_3_630, output_3_7, output_2_630;
mixer gate_output_2_630(.a(output_3_630), .b(output_3_7), .y(output_2_630));
wire output_4_630, output_4_7, output_3_630;
mixer gate_output_3_630(.a(output_4_630), .b(output_4_7), .y(output_3_630));
wire output_5_630, output_5_7, output_4_630;
mixer gate_output_4_630(.a(output_5_630), .b(output_5_7), .y(output_4_630));
wire output_6_630, output_6_7, output_5_630;
mixer gate_output_5_630(.a(output_6_630), .b(output_6_7), .y(output_5_630));
wire output_7_630, output_7_7, output_6_630;
mixer gate_output_6_630(.a(output_7_630), .b(output_7_7), .y(output_6_630));
wire output_8_630, output_8_7, output_7_630;
mixer gate_output_7_630(.a(output_8_630), .b(output_8_7), .y(output_7_630));
wire output_9_630, output_9_7, output_8_630;
mixer gate_output_8_630(.a(output_9_630), .b(output_9_7), .y(output_8_630));
wire output_10_630, output_10_7, output_9_630;
mixer gate_output_9_630(.a(output_10_630), .b(output_10_7), .y(output_9_630));
wire output_11_630, output_11_7, output_10_630;
mixer gate_output_10_630(.a(output_11_630), .b(output_11_7), .y(output_10_630));
wire output_12_630, output_12_7, output_11_630;
mixer gate_output_11_630(.a(output_12_630), .b(output_12_7), .y(output_11_630));
wire output_13_630, output_13_7, output_12_630;
mixer gate_output_12_630(.a(output_13_630), .b(output_13_7), .y(output_12_630));
wire output_14_630, output_14_7, output_13_630;
mixer gate_output_13_630(.a(output_14_630), .b(output_14_7), .y(output_13_630));
wire output_15_630, output_15_7, output_14_630;
mixer gate_output_14_630(.a(output_15_630), .b(output_15_7), .y(output_14_630));
wire output_16_630, output_16_7, output_15_630;
mixer gate_output_15_630(.a(output_16_630), .b(output_16_7), .y(output_15_630));
wire output_1_631, output_1_8, output_0_631;
mixer gate_output_0_631(.a(output_1_631), .b(output_1_8), .y(output_0_631));
wire output_2_631, output_2_8, output_1_631;
mixer gate_output_1_631(.a(output_2_631), .b(output_2_8), .y(output_1_631));
wire output_3_631, output_3_8, output_2_631;
mixer gate_output_2_631(.a(output_3_631), .b(output_3_8), .y(output_2_631));
wire output_4_631, output_4_8, output_3_631;
mixer gate_output_3_631(.a(output_4_631), .b(output_4_8), .y(output_3_631));
wire output_5_631, output_5_8, output_4_631;
mixer gate_output_4_631(.a(output_5_631), .b(output_5_8), .y(output_4_631));
wire output_6_631, output_6_8, output_5_631;
mixer gate_output_5_631(.a(output_6_631), .b(output_6_8), .y(output_5_631));
wire output_7_631, output_7_8, output_6_631;
mixer gate_output_6_631(.a(output_7_631), .b(output_7_8), .y(output_6_631));
wire output_8_631, output_8_8, output_7_631;
mixer gate_output_7_631(.a(output_8_631), .b(output_8_8), .y(output_7_631));
wire output_9_631, output_9_8, output_8_631;
mixer gate_output_8_631(.a(output_9_631), .b(output_9_8), .y(output_8_631));
wire output_10_631, output_10_8, output_9_631;
mixer gate_output_9_631(.a(output_10_631), .b(output_10_8), .y(output_9_631));
wire output_11_631, output_11_8, output_10_631;
mixer gate_output_10_631(.a(output_11_631), .b(output_11_8), .y(output_10_631));
wire output_12_631, output_12_8, output_11_631;
mixer gate_output_11_631(.a(output_12_631), .b(output_12_8), .y(output_11_631));
wire output_13_631, output_13_8, output_12_631;
mixer gate_output_12_631(.a(output_13_631), .b(output_13_8), .y(output_12_631));
wire output_14_631, output_14_8, output_13_631;
mixer gate_output_13_631(.a(output_14_631), .b(output_14_8), .y(output_13_631));
wire output_15_631, output_15_8, output_14_631;
mixer gate_output_14_631(.a(output_15_631), .b(output_15_8), .y(output_14_631));
wire output_16_631, output_16_8, output_15_631;
mixer gate_output_15_631(.a(output_16_631), .b(output_16_8), .y(output_15_631));
wire output_1_632, output_1_9, output_0_632;
mixer gate_output_0_632(.a(output_1_632), .b(output_1_9), .y(output_0_632));
wire output_2_632, output_2_9, output_1_632;
mixer gate_output_1_632(.a(output_2_632), .b(output_2_9), .y(output_1_632));
wire output_3_632, output_3_9, output_2_632;
mixer gate_output_2_632(.a(output_3_632), .b(output_3_9), .y(output_2_632));
wire output_4_632, output_4_9, output_3_632;
mixer gate_output_3_632(.a(output_4_632), .b(output_4_9), .y(output_3_632));
wire output_5_632, output_5_9, output_4_632;
mixer gate_output_4_632(.a(output_5_632), .b(output_5_9), .y(output_4_632));
wire output_6_632, output_6_9, output_5_632;
mixer gate_output_5_632(.a(output_6_632), .b(output_6_9), .y(output_5_632));
wire output_7_632, output_7_9, output_6_632;
mixer gate_output_6_632(.a(output_7_632), .b(output_7_9), .y(output_6_632));
wire output_8_632, output_8_9, output_7_632;
mixer gate_output_7_632(.a(output_8_632), .b(output_8_9), .y(output_7_632));
wire output_9_632, output_9_9, output_8_632;
mixer gate_output_8_632(.a(output_9_632), .b(output_9_9), .y(output_8_632));
wire output_10_632, output_10_9, output_9_632;
mixer gate_output_9_632(.a(output_10_632), .b(output_10_9), .y(output_9_632));
wire output_11_632, output_11_9, output_10_632;
mixer gate_output_10_632(.a(output_11_632), .b(output_11_9), .y(output_10_632));
wire output_12_632, output_12_9, output_11_632;
mixer gate_output_11_632(.a(output_12_632), .b(output_12_9), .y(output_11_632));
wire output_13_632, output_13_9, output_12_632;
mixer gate_output_12_632(.a(output_13_632), .b(output_13_9), .y(output_12_632));
wire output_14_632, output_14_9, output_13_632;
mixer gate_output_13_632(.a(output_14_632), .b(output_14_9), .y(output_13_632));
wire output_15_632, output_15_9, output_14_632;
mixer gate_output_14_632(.a(output_15_632), .b(output_15_9), .y(output_14_632));
wire output_16_632, output_16_9, output_15_632;
mixer gate_output_15_632(.a(output_16_632), .b(output_16_9), .y(output_15_632));
wire output_1_633, output_1_10, output_0_633;
mixer gate_output_0_633(.a(output_1_633), .b(output_1_10), .y(output_0_633));
wire output_2_633, output_2_10, output_1_633;
mixer gate_output_1_633(.a(output_2_633), .b(output_2_10), .y(output_1_633));
wire output_3_633, output_3_10, output_2_633;
mixer gate_output_2_633(.a(output_3_633), .b(output_3_10), .y(output_2_633));
wire output_4_633, output_4_10, output_3_633;
mixer gate_output_3_633(.a(output_4_633), .b(output_4_10), .y(output_3_633));
wire output_5_633, output_5_10, output_4_633;
mixer gate_output_4_633(.a(output_5_633), .b(output_5_10), .y(output_4_633));
wire output_6_633, output_6_10, output_5_633;
mixer gate_output_5_633(.a(output_6_633), .b(output_6_10), .y(output_5_633));
wire output_7_633, output_7_10, output_6_633;
mixer gate_output_6_633(.a(output_7_633), .b(output_7_10), .y(output_6_633));
wire output_8_633, output_8_10, output_7_633;
mixer gate_output_7_633(.a(output_8_633), .b(output_8_10), .y(output_7_633));
wire output_9_633, output_9_10, output_8_633;
mixer gate_output_8_633(.a(output_9_633), .b(output_9_10), .y(output_8_633));
wire output_10_633, output_10_10, output_9_633;
mixer gate_output_9_633(.a(output_10_633), .b(output_10_10), .y(output_9_633));
wire output_11_633, output_11_10, output_10_633;
mixer gate_output_10_633(.a(output_11_633), .b(output_11_10), .y(output_10_633));
wire output_12_633, output_12_10, output_11_633;
mixer gate_output_11_633(.a(output_12_633), .b(output_12_10), .y(output_11_633));
wire output_13_633, output_13_10, output_12_633;
mixer gate_output_12_633(.a(output_13_633), .b(output_13_10), .y(output_12_633));
wire output_14_633, output_14_10, output_13_633;
mixer gate_output_13_633(.a(output_14_633), .b(output_14_10), .y(output_13_633));
wire output_15_633, output_15_10, output_14_633;
mixer gate_output_14_633(.a(output_15_633), .b(output_15_10), .y(output_14_633));
wire output_16_633, output_16_10, output_15_633;
mixer gate_output_15_633(.a(output_16_633), .b(output_16_10), .y(output_15_633));
wire output_1_634, output_1_11, output_0_634;
mixer gate_output_0_634(.a(output_1_634), .b(output_1_11), .y(output_0_634));
wire output_2_634, output_2_11, output_1_634;
mixer gate_output_1_634(.a(output_2_634), .b(output_2_11), .y(output_1_634));
wire output_3_634, output_3_11, output_2_634;
mixer gate_output_2_634(.a(output_3_634), .b(output_3_11), .y(output_2_634));
wire output_4_634, output_4_11, output_3_634;
mixer gate_output_3_634(.a(output_4_634), .b(output_4_11), .y(output_3_634));
wire output_5_634, output_5_11, output_4_634;
mixer gate_output_4_634(.a(output_5_634), .b(output_5_11), .y(output_4_634));
wire output_6_634, output_6_11, output_5_634;
mixer gate_output_5_634(.a(output_6_634), .b(output_6_11), .y(output_5_634));
wire output_7_634, output_7_11, output_6_634;
mixer gate_output_6_634(.a(output_7_634), .b(output_7_11), .y(output_6_634));
wire output_8_634, output_8_11, output_7_634;
mixer gate_output_7_634(.a(output_8_634), .b(output_8_11), .y(output_7_634));
wire output_9_634, output_9_11, output_8_634;
mixer gate_output_8_634(.a(output_9_634), .b(output_9_11), .y(output_8_634));
wire output_10_634, output_10_11, output_9_634;
mixer gate_output_9_634(.a(output_10_634), .b(output_10_11), .y(output_9_634));
wire output_11_634, output_11_11, output_10_634;
mixer gate_output_10_634(.a(output_11_634), .b(output_11_11), .y(output_10_634));
wire output_12_634, output_12_11, output_11_634;
mixer gate_output_11_634(.a(output_12_634), .b(output_12_11), .y(output_11_634));
wire output_13_634, output_13_11, output_12_634;
mixer gate_output_12_634(.a(output_13_634), .b(output_13_11), .y(output_12_634));
wire output_14_634, output_14_11, output_13_634;
mixer gate_output_13_634(.a(output_14_634), .b(output_14_11), .y(output_13_634));
wire output_15_634, output_15_11, output_14_634;
mixer gate_output_14_634(.a(output_15_634), .b(output_15_11), .y(output_14_634));
wire output_16_634, output_16_11, output_15_634;
mixer gate_output_15_634(.a(output_16_634), .b(output_16_11), .y(output_15_634));
wire output_1_635, output_1_12, output_0_635;
mixer gate_output_0_635(.a(output_1_635), .b(output_1_12), .y(output_0_635));
wire output_2_635, output_2_12, output_1_635;
mixer gate_output_1_635(.a(output_2_635), .b(output_2_12), .y(output_1_635));
wire output_3_635, output_3_12, output_2_635;
mixer gate_output_2_635(.a(output_3_635), .b(output_3_12), .y(output_2_635));
wire output_4_635, output_4_12, output_3_635;
mixer gate_output_3_635(.a(output_4_635), .b(output_4_12), .y(output_3_635));
wire output_5_635, output_5_12, output_4_635;
mixer gate_output_4_635(.a(output_5_635), .b(output_5_12), .y(output_4_635));
wire output_6_635, output_6_12, output_5_635;
mixer gate_output_5_635(.a(output_6_635), .b(output_6_12), .y(output_5_635));
wire output_7_635, output_7_12, output_6_635;
mixer gate_output_6_635(.a(output_7_635), .b(output_7_12), .y(output_6_635));
wire output_8_635, output_8_12, output_7_635;
mixer gate_output_7_635(.a(output_8_635), .b(output_8_12), .y(output_7_635));
wire output_9_635, output_9_12, output_8_635;
mixer gate_output_8_635(.a(output_9_635), .b(output_9_12), .y(output_8_635));
wire output_10_635, output_10_12, output_9_635;
mixer gate_output_9_635(.a(output_10_635), .b(output_10_12), .y(output_9_635));
wire output_11_635, output_11_12, output_10_635;
mixer gate_output_10_635(.a(output_11_635), .b(output_11_12), .y(output_10_635));
wire output_12_635, output_12_12, output_11_635;
mixer gate_output_11_635(.a(output_12_635), .b(output_12_12), .y(output_11_635));
wire output_13_635, output_13_12, output_12_635;
mixer gate_output_12_635(.a(output_13_635), .b(output_13_12), .y(output_12_635));
wire output_14_635, output_14_12, output_13_635;
mixer gate_output_13_635(.a(output_14_635), .b(output_14_12), .y(output_13_635));
wire output_15_635, output_15_12, output_14_635;
mixer gate_output_14_635(.a(output_15_635), .b(output_15_12), .y(output_14_635));
wire output_16_635, output_16_12, output_15_635;
mixer gate_output_15_635(.a(output_16_635), .b(output_16_12), .y(output_15_635));
wire output_1_636, output_1_13, output_0_636;
mixer gate_output_0_636(.a(output_1_636), .b(output_1_13), .y(output_0_636));
wire output_2_636, output_2_13, output_1_636;
mixer gate_output_1_636(.a(output_2_636), .b(output_2_13), .y(output_1_636));
wire output_3_636, output_3_13, output_2_636;
mixer gate_output_2_636(.a(output_3_636), .b(output_3_13), .y(output_2_636));
wire output_4_636, output_4_13, output_3_636;
mixer gate_output_3_636(.a(output_4_636), .b(output_4_13), .y(output_3_636));
wire output_5_636, output_5_13, output_4_636;
mixer gate_output_4_636(.a(output_5_636), .b(output_5_13), .y(output_4_636));
wire output_6_636, output_6_13, output_5_636;
mixer gate_output_5_636(.a(output_6_636), .b(output_6_13), .y(output_5_636));
wire output_7_636, output_7_13, output_6_636;
mixer gate_output_6_636(.a(output_7_636), .b(output_7_13), .y(output_6_636));
wire output_8_636, output_8_13, output_7_636;
mixer gate_output_7_636(.a(output_8_636), .b(output_8_13), .y(output_7_636));
wire output_9_636, output_9_13, output_8_636;
mixer gate_output_8_636(.a(output_9_636), .b(output_9_13), .y(output_8_636));
wire output_10_636, output_10_13, output_9_636;
mixer gate_output_9_636(.a(output_10_636), .b(output_10_13), .y(output_9_636));
wire output_11_636, output_11_13, output_10_636;
mixer gate_output_10_636(.a(output_11_636), .b(output_11_13), .y(output_10_636));
wire output_12_636, output_12_13, output_11_636;
mixer gate_output_11_636(.a(output_12_636), .b(output_12_13), .y(output_11_636));
wire output_13_636, output_13_13, output_12_636;
mixer gate_output_12_636(.a(output_13_636), .b(output_13_13), .y(output_12_636));
wire output_14_636, output_14_13, output_13_636;
mixer gate_output_13_636(.a(output_14_636), .b(output_14_13), .y(output_13_636));
wire output_15_636, output_15_13, output_14_636;
mixer gate_output_14_636(.a(output_15_636), .b(output_15_13), .y(output_14_636));
wire output_16_636, output_16_13, output_15_636;
mixer gate_output_15_636(.a(output_16_636), .b(output_16_13), .y(output_15_636));
wire output_1_637, output_1_14, output_0_637;
mixer gate_output_0_637(.a(output_1_637), .b(output_1_14), .y(output_0_637));
wire output_2_637, output_2_14, output_1_637;
mixer gate_output_1_637(.a(output_2_637), .b(output_2_14), .y(output_1_637));
wire output_3_637, output_3_14, output_2_637;
mixer gate_output_2_637(.a(output_3_637), .b(output_3_14), .y(output_2_637));
wire output_4_637, output_4_14, output_3_637;
mixer gate_output_3_637(.a(output_4_637), .b(output_4_14), .y(output_3_637));
wire output_5_637, output_5_14, output_4_637;
mixer gate_output_4_637(.a(output_5_637), .b(output_5_14), .y(output_4_637));
wire output_6_637, output_6_14, output_5_637;
mixer gate_output_5_637(.a(output_6_637), .b(output_6_14), .y(output_5_637));
wire output_7_637, output_7_14, output_6_637;
mixer gate_output_6_637(.a(output_7_637), .b(output_7_14), .y(output_6_637));
wire output_8_637, output_8_14, output_7_637;
mixer gate_output_7_637(.a(output_8_637), .b(output_8_14), .y(output_7_637));
wire output_9_637, output_9_14, output_8_637;
mixer gate_output_8_637(.a(output_9_637), .b(output_9_14), .y(output_8_637));
wire output_10_637, output_10_14, output_9_637;
mixer gate_output_9_637(.a(output_10_637), .b(output_10_14), .y(output_9_637));
wire output_11_637, output_11_14, output_10_637;
mixer gate_output_10_637(.a(output_11_637), .b(output_11_14), .y(output_10_637));
wire output_12_637, output_12_14, output_11_637;
mixer gate_output_11_637(.a(output_12_637), .b(output_12_14), .y(output_11_637));
wire output_13_637, output_13_14, output_12_637;
mixer gate_output_12_637(.a(output_13_637), .b(output_13_14), .y(output_12_637));
wire output_14_637, output_14_14, output_13_637;
mixer gate_output_13_637(.a(output_14_637), .b(output_14_14), .y(output_13_637));
wire output_15_637, output_15_14, output_14_637;
mixer gate_output_14_637(.a(output_15_637), .b(output_15_14), .y(output_14_637));
wire output_16_637, output_16_14, output_15_637;
mixer gate_output_15_637(.a(output_16_637), .b(output_16_14), .y(output_15_637));
wire output_1_638, output_1_15, output_0_638;
mixer gate_output_0_638(.a(output_1_638), .b(output_1_15), .y(output_0_638));
wire output_2_638, output_2_15, output_1_638;
mixer gate_output_1_638(.a(output_2_638), .b(output_2_15), .y(output_1_638));
wire output_3_638, output_3_15, output_2_638;
mixer gate_output_2_638(.a(output_3_638), .b(output_3_15), .y(output_2_638));
wire output_4_638, output_4_15, output_3_638;
mixer gate_output_3_638(.a(output_4_638), .b(output_4_15), .y(output_3_638));
wire output_5_638, output_5_15, output_4_638;
mixer gate_output_4_638(.a(output_5_638), .b(output_5_15), .y(output_4_638));
wire output_6_638, output_6_15, output_5_638;
mixer gate_output_5_638(.a(output_6_638), .b(output_6_15), .y(output_5_638));
wire output_7_638, output_7_15, output_6_638;
mixer gate_output_6_638(.a(output_7_638), .b(output_7_15), .y(output_6_638));
wire output_8_638, output_8_15, output_7_638;
mixer gate_output_7_638(.a(output_8_638), .b(output_8_15), .y(output_7_638));
wire output_9_638, output_9_15, output_8_638;
mixer gate_output_8_638(.a(output_9_638), .b(output_9_15), .y(output_8_638));
wire output_10_638, output_10_15, output_9_638;
mixer gate_output_9_638(.a(output_10_638), .b(output_10_15), .y(output_9_638));
wire output_11_638, output_11_15, output_10_638;
mixer gate_output_10_638(.a(output_11_638), .b(output_11_15), .y(output_10_638));
wire output_12_638, output_12_15, output_11_638;
mixer gate_output_11_638(.a(output_12_638), .b(output_12_15), .y(output_11_638));
wire output_13_638, output_13_15, output_12_638;
mixer gate_output_12_638(.a(output_13_638), .b(output_13_15), .y(output_12_638));
wire output_14_638, output_14_15, output_13_638;
mixer gate_output_13_638(.a(output_14_638), .b(output_14_15), .y(output_13_638));
wire output_15_638, output_15_15, output_14_638;
mixer gate_output_14_638(.a(output_15_638), .b(output_15_15), .y(output_14_638));
wire output_16_638, output_16_15, output_15_638;
mixer gate_output_15_638(.a(output_16_638), .b(output_16_15), .y(output_15_638));
wire output_1_639, output_1_0, output_0_639;
mixer gate_output_0_639(.a(output_1_639), .b(output_1_0), .y(output_0_639));
wire output_2_639, output_2_0, output_1_639;
mixer gate_output_1_639(.a(output_2_639), .b(output_2_0), .y(output_1_639));
wire output_3_639, output_3_0, output_2_639;
mixer gate_output_2_639(.a(output_3_639), .b(output_3_0), .y(output_2_639));
wire output_4_639, output_4_0, output_3_639;
mixer gate_output_3_639(.a(output_4_639), .b(output_4_0), .y(output_3_639));
wire output_5_639, output_5_0, output_4_639;
mixer gate_output_4_639(.a(output_5_639), .b(output_5_0), .y(output_4_639));
wire output_6_639, output_6_0, output_5_639;
mixer gate_output_5_639(.a(output_6_639), .b(output_6_0), .y(output_5_639));
wire output_7_639, output_7_0, output_6_639;
mixer gate_output_6_639(.a(output_7_639), .b(output_7_0), .y(output_6_639));
wire output_8_639, output_8_0, output_7_639;
mixer gate_output_7_639(.a(output_8_639), .b(output_8_0), .y(output_7_639));
wire output_9_639, output_9_0, output_8_639;
mixer gate_output_8_639(.a(output_9_639), .b(output_9_0), .y(output_8_639));
wire output_10_639, output_10_0, output_9_639;
mixer gate_output_9_639(.a(output_10_639), .b(output_10_0), .y(output_9_639));
wire output_11_639, output_11_0, output_10_639;
mixer gate_output_10_639(.a(output_11_639), .b(output_11_0), .y(output_10_639));
wire output_12_639, output_12_0, output_11_639;
mixer gate_output_11_639(.a(output_12_639), .b(output_12_0), .y(output_11_639));
wire output_13_639, output_13_0, output_12_639;
mixer gate_output_12_639(.a(output_13_639), .b(output_13_0), .y(output_12_639));
wire output_14_639, output_14_0, output_13_639;
mixer gate_output_13_639(.a(output_14_639), .b(output_14_0), .y(output_13_639));
wire output_15_639, output_15_0, output_14_639;
mixer gate_output_14_639(.a(output_15_639), .b(output_15_0), .y(output_14_639));
wire output_16_639, output_16_0, output_15_639;
mixer gate_output_15_639(.a(output_16_639), .b(output_16_0), .y(output_15_639));
wire output_1_640, output_1_1, output_0_640;
mixer gate_output_0_640(.a(output_1_640), .b(output_1_1), .y(output_0_640));
wire output_2_640, output_2_1, output_1_640;
mixer gate_output_1_640(.a(output_2_640), .b(output_2_1), .y(output_1_640));
wire output_3_640, output_3_1, output_2_640;
mixer gate_output_2_640(.a(output_3_640), .b(output_3_1), .y(output_2_640));
wire output_4_640, output_4_1, output_3_640;
mixer gate_output_3_640(.a(output_4_640), .b(output_4_1), .y(output_3_640));
wire output_5_640, output_5_1, output_4_640;
mixer gate_output_4_640(.a(output_5_640), .b(output_5_1), .y(output_4_640));
wire output_6_640, output_6_1, output_5_640;
mixer gate_output_5_640(.a(output_6_640), .b(output_6_1), .y(output_5_640));
wire output_7_640, output_7_1, output_6_640;
mixer gate_output_6_640(.a(output_7_640), .b(output_7_1), .y(output_6_640));
wire output_8_640, output_8_1, output_7_640;
mixer gate_output_7_640(.a(output_8_640), .b(output_8_1), .y(output_7_640));
wire output_9_640, output_9_1, output_8_640;
mixer gate_output_8_640(.a(output_9_640), .b(output_9_1), .y(output_8_640));
wire output_10_640, output_10_1, output_9_640;
mixer gate_output_9_640(.a(output_10_640), .b(output_10_1), .y(output_9_640));
wire output_11_640, output_11_1, output_10_640;
mixer gate_output_10_640(.a(output_11_640), .b(output_11_1), .y(output_10_640));
wire output_12_640, output_12_1, output_11_640;
mixer gate_output_11_640(.a(output_12_640), .b(output_12_1), .y(output_11_640));
wire output_13_640, output_13_1, output_12_640;
mixer gate_output_12_640(.a(output_13_640), .b(output_13_1), .y(output_12_640));
wire output_14_640, output_14_1, output_13_640;
mixer gate_output_13_640(.a(output_14_640), .b(output_14_1), .y(output_13_640));
wire output_15_640, output_15_1, output_14_640;
mixer gate_output_14_640(.a(output_15_640), .b(output_15_1), .y(output_14_640));
wire output_16_640, output_16_1, output_15_640;
mixer gate_output_15_640(.a(output_16_640), .b(output_16_1), .y(output_15_640));
wire output_1_641, output_1_2, output_0_641;
mixer gate_output_0_641(.a(output_1_641), .b(output_1_2), .y(output_0_641));
wire output_2_641, output_2_2, output_1_641;
mixer gate_output_1_641(.a(output_2_641), .b(output_2_2), .y(output_1_641));
wire output_3_641, output_3_2, output_2_641;
mixer gate_output_2_641(.a(output_3_641), .b(output_3_2), .y(output_2_641));
wire output_4_641, output_4_2, output_3_641;
mixer gate_output_3_641(.a(output_4_641), .b(output_4_2), .y(output_3_641));
wire output_5_641, output_5_2, output_4_641;
mixer gate_output_4_641(.a(output_5_641), .b(output_5_2), .y(output_4_641));
wire output_6_641, output_6_2, output_5_641;
mixer gate_output_5_641(.a(output_6_641), .b(output_6_2), .y(output_5_641));
wire output_7_641, output_7_2, output_6_641;
mixer gate_output_6_641(.a(output_7_641), .b(output_7_2), .y(output_6_641));
wire output_8_641, output_8_2, output_7_641;
mixer gate_output_7_641(.a(output_8_641), .b(output_8_2), .y(output_7_641));
wire output_9_641, output_9_2, output_8_641;
mixer gate_output_8_641(.a(output_9_641), .b(output_9_2), .y(output_8_641));
wire output_10_641, output_10_2, output_9_641;
mixer gate_output_9_641(.a(output_10_641), .b(output_10_2), .y(output_9_641));
wire output_11_641, output_11_2, output_10_641;
mixer gate_output_10_641(.a(output_11_641), .b(output_11_2), .y(output_10_641));
wire output_12_641, output_12_2, output_11_641;
mixer gate_output_11_641(.a(output_12_641), .b(output_12_2), .y(output_11_641));
wire output_13_641, output_13_2, output_12_641;
mixer gate_output_12_641(.a(output_13_641), .b(output_13_2), .y(output_12_641));
wire output_14_641, output_14_2, output_13_641;
mixer gate_output_13_641(.a(output_14_641), .b(output_14_2), .y(output_13_641));
wire output_15_641, output_15_2, output_14_641;
mixer gate_output_14_641(.a(output_15_641), .b(output_15_2), .y(output_14_641));
wire output_16_641, output_16_2, output_15_641;
mixer gate_output_15_641(.a(output_16_641), .b(output_16_2), .y(output_15_641));
wire output_1_642, output_1_3, output_0_642;
mixer gate_output_0_642(.a(output_1_642), .b(output_1_3), .y(output_0_642));
wire output_2_642, output_2_3, output_1_642;
mixer gate_output_1_642(.a(output_2_642), .b(output_2_3), .y(output_1_642));
wire output_3_642, output_3_3, output_2_642;
mixer gate_output_2_642(.a(output_3_642), .b(output_3_3), .y(output_2_642));
wire output_4_642, output_4_3, output_3_642;
mixer gate_output_3_642(.a(output_4_642), .b(output_4_3), .y(output_3_642));
wire output_5_642, output_5_3, output_4_642;
mixer gate_output_4_642(.a(output_5_642), .b(output_5_3), .y(output_4_642));
wire output_6_642, output_6_3, output_5_642;
mixer gate_output_5_642(.a(output_6_642), .b(output_6_3), .y(output_5_642));
wire output_7_642, output_7_3, output_6_642;
mixer gate_output_6_642(.a(output_7_642), .b(output_7_3), .y(output_6_642));
wire output_8_642, output_8_3, output_7_642;
mixer gate_output_7_642(.a(output_8_642), .b(output_8_3), .y(output_7_642));
wire output_9_642, output_9_3, output_8_642;
mixer gate_output_8_642(.a(output_9_642), .b(output_9_3), .y(output_8_642));
wire output_10_642, output_10_3, output_9_642;
mixer gate_output_9_642(.a(output_10_642), .b(output_10_3), .y(output_9_642));
wire output_11_642, output_11_3, output_10_642;
mixer gate_output_10_642(.a(output_11_642), .b(output_11_3), .y(output_10_642));
wire output_12_642, output_12_3, output_11_642;
mixer gate_output_11_642(.a(output_12_642), .b(output_12_3), .y(output_11_642));
wire output_13_642, output_13_3, output_12_642;
mixer gate_output_12_642(.a(output_13_642), .b(output_13_3), .y(output_12_642));
wire output_14_642, output_14_3, output_13_642;
mixer gate_output_13_642(.a(output_14_642), .b(output_14_3), .y(output_13_642));
wire output_15_642, output_15_3, output_14_642;
mixer gate_output_14_642(.a(output_15_642), .b(output_15_3), .y(output_14_642));
wire output_16_642, output_16_3, output_15_642;
mixer gate_output_15_642(.a(output_16_642), .b(output_16_3), .y(output_15_642));
wire output_1_643, output_1_4, output_0_643;
mixer gate_output_0_643(.a(output_1_643), .b(output_1_4), .y(output_0_643));
wire output_2_643, output_2_4, output_1_643;
mixer gate_output_1_643(.a(output_2_643), .b(output_2_4), .y(output_1_643));
wire output_3_643, output_3_4, output_2_643;
mixer gate_output_2_643(.a(output_3_643), .b(output_3_4), .y(output_2_643));
wire output_4_643, output_4_4, output_3_643;
mixer gate_output_3_643(.a(output_4_643), .b(output_4_4), .y(output_3_643));
wire output_5_643, output_5_4, output_4_643;
mixer gate_output_4_643(.a(output_5_643), .b(output_5_4), .y(output_4_643));
wire output_6_643, output_6_4, output_5_643;
mixer gate_output_5_643(.a(output_6_643), .b(output_6_4), .y(output_5_643));
wire output_7_643, output_7_4, output_6_643;
mixer gate_output_6_643(.a(output_7_643), .b(output_7_4), .y(output_6_643));
wire output_8_643, output_8_4, output_7_643;
mixer gate_output_7_643(.a(output_8_643), .b(output_8_4), .y(output_7_643));
wire output_9_643, output_9_4, output_8_643;
mixer gate_output_8_643(.a(output_9_643), .b(output_9_4), .y(output_8_643));
wire output_10_643, output_10_4, output_9_643;
mixer gate_output_9_643(.a(output_10_643), .b(output_10_4), .y(output_9_643));
wire output_11_643, output_11_4, output_10_643;
mixer gate_output_10_643(.a(output_11_643), .b(output_11_4), .y(output_10_643));
wire output_12_643, output_12_4, output_11_643;
mixer gate_output_11_643(.a(output_12_643), .b(output_12_4), .y(output_11_643));
wire output_13_643, output_13_4, output_12_643;
mixer gate_output_12_643(.a(output_13_643), .b(output_13_4), .y(output_12_643));
wire output_14_643, output_14_4, output_13_643;
mixer gate_output_13_643(.a(output_14_643), .b(output_14_4), .y(output_13_643));
wire output_15_643, output_15_4, output_14_643;
mixer gate_output_14_643(.a(output_15_643), .b(output_15_4), .y(output_14_643));
wire output_16_643, output_16_4, output_15_643;
mixer gate_output_15_643(.a(output_16_643), .b(output_16_4), .y(output_15_643));
wire output_1_644, output_1_5, output_0_644;
mixer gate_output_0_644(.a(output_1_644), .b(output_1_5), .y(output_0_644));
wire output_2_644, output_2_5, output_1_644;
mixer gate_output_1_644(.a(output_2_644), .b(output_2_5), .y(output_1_644));
wire output_3_644, output_3_5, output_2_644;
mixer gate_output_2_644(.a(output_3_644), .b(output_3_5), .y(output_2_644));
wire output_4_644, output_4_5, output_3_644;
mixer gate_output_3_644(.a(output_4_644), .b(output_4_5), .y(output_3_644));
wire output_5_644, output_5_5, output_4_644;
mixer gate_output_4_644(.a(output_5_644), .b(output_5_5), .y(output_4_644));
wire output_6_644, output_6_5, output_5_644;
mixer gate_output_5_644(.a(output_6_644), .b(output_6_5), .y(output_5_644));
wire output_7_644, output_7_5, output_6_644;
mixer gate_output_6_644(.a(output_7_644), .b(output_7_5), .y(output_6_644));
wire output_8_644, output_8_5, output_7_644;
mixer gate_output_7_644(.a(output_8_644), .b(output_8_5), .y(output_7_644));
wire output_9_644, output_9_5, output_8_644;
mixer gate_output_8_644(.a(output_9_644), .b(output_9_5), .y(output_8_644));
wire output_10_644, output_10_5, output_9_644;
mixer gate_output_9_644(.a(output_10_644), .b(output_10_5), .y(output_9_644));
wire output_11_644, output_11_5, output_10_644;
mixer gate_output_10_644(.a(output_11_644), .b(output_11_5), .y(output_10_644));
wire output_12_644, output_12_5, output_11_644;
mixer gate_output_11_644(.a(output_12_644), .b(output_12_5), .y(output_11_644));
wire output_13_644, output_13_5, output_12_644;
mixer gate_output_12_644(.a(output_13_644), .b(output_13_5), .y(output_12_644));
wire output_14_644, output_14_5, output_13_644;
mixer gate_output_13_644(.a(output_14_644), .b(output_14_5), .y(output_13_644));
wire output_15_644, output_15_5, output_14_644;
mixer gate_output_14_644(.a(output_15_644), .b(output_15_5), .y(output_14_644));
wire output_16_644, output_16_5, output_15_644;
mixer gate_output_15_644(.a(output_16_644), .b(output_16_5), .y(output_15_644));
wire output_1_645, output_1_6, output_0_645;
mixer gate_output_0_645(.a(output_1_645), .b(output_1_6), .y(output_0_645));
wire output_2_645, output_2_6, output_1_645;
mixer gate_output_1_645(.a(output_2_645), .b(output_2_6), .y(output_1_645));
wire output_3_645, output_3_6, output_2_645;
mixer gate_output_2_645(.a(output_3_645), .b(output_3_6), .y(output_2_645));
wire output_4_645, output_4_6, output_3_645;
mixer gate_output_3_645(.a(output_4_645), .b(output_4_6), .y(output_3_645));
wire output_5_645, output_5_6, output_4_645;
mixer gate_output_4_645(.a(output_5_645), .b(output_5_6), .y(output_4_645));
wire output_6_645, output_6_6, output_5_645;
mixer gate_output_5_645(.a(output_6_645), .b(output_6_6), .y(output_5_645));
wire output_7_645, output_7_6, output_6_645;
mixer gate_output_6_645(.a(output_7_645), .b(output_7_6), .y(output_6_645));
wire output_8_645, output_8_6, output_7_645;
mixer gate_output_7_645(.a(output_8_645), .b(output_8_6), .y(output_7_645));
wire output_9_645, output_9_6, output_8_645;
mixer gate_output_8_645(.a(output_9_645), .b(output_9_6), .y(output_8_645));
wire output_10_645, output_10_6, output_9_645;
mixer gate_output_9_645(.a(output_10_645), .b(output_10_6), .y(output_9_645));
wire output_11_645, output_11_6, output_10_645;
mixer gate_output_10_645(.a(output_11_645), .b(output_11_6), .y(output_10_645));
wire output_12_645, output_12_6, output_11_645;
mixer gate_output_11_645(.a(output_12_645), .b(output_12_6), .y(output_11_645));
wire output_13_645, output_13_6, output_12_645;
mixer gate_output_12_645(.a(output_13_645), .b(output_13_6), .y(output_12_645));
wire output_14_645, output_14_6, output_13_645;
mixer gate_output_13_645(.a(output_14_645), .b(output_14_6), .y(output_13_645));
wire output_15_645, output_15_6, output_14_645;
mixer gate_output_14_645(.a(output_15_645), .b(output_15_6), .y(output_14_645));
wire output_16_645, output_16_6, output_15_645;
mixer gate_output_15_645(.a(output_16_645), .b(output_16_6), .y(output_15_645));
wire output_1_646, output_1_7, output_0_646;
mixer gate_output_0_646(.a(output_1_646), .b(output_1_7), .y(output_0_646));
wire output_2_646, output_2_7, output_1_646;
mixer gate_output_1_646(.a(output_2_646), .b(output_2_7), .y(output_1_646));
wire output_3_646, output_3_7, output_2_646;
mixer gate_output_2_646(.a(output_3_646), .b(output_3_7), .y(output_2_646));
wire output_4_646, output_4_7, output_3_646;
mixer gate_output_3_646(.a(output_4_646), .b(output_4_7), .y(output_3_646));
wire output_5_646, output_5_7, output_4_646;
mixer gate_output_4_646(.a(output_5_646), .b(output_5_7), .y(output_4_646));
wire output_6_646, output_6_7, output_5_646;
mixer gate_output_5_646(.a(output_6_646), .b(output_6_7), .y(output_5_646));
wire output_7_646, output_7_7, output_6_646;
mixer gate_output_6_646(.a(output_7_646), .b(output_7_7), .y(output_6_646));
wire output_8_646, output_8_7, output_7_646;
mixer gate_output_7_646(.a(output_8_646), .b(output_8_7), .y(output_7_646));
wire output_9_646, output_9_7, output_8_646;
mixer gate_output_8_646(.a(output_9_646), .b(output_9_7), .y(output_8_646));
wire output_10_646, output_10_7, output_9_646;
mixer gate_output_9_646(.a(output_10_646), .b(output_10_7), .y(output_9_646));
wire output_11_646, output_11_7, output_10_646;
mixer gate_output_10_646(.a(output_11_646), .b(output_11_7), .y(output_10_646));
wire output_12_646, output_12_7, output_11_646;
mixer gate_output_11_646(.a(output_12_646), .b(output_12_7), .y(output_11_646));
wire output_13_646, output_13_7, output_12_646;
mixer gate_output_12_646(.a(output_13_646), .b(output_13_7), .y(output_12_646));
wire output_14_646, output_14_7, output_13_646;
mixer gate_output_13_646(.a(output_14_646), .b(output_14_7), .y(output_13_646));
wire output_15_646, output_15_7, output_14_646;
mixer gate_output_14_646(.a(output_15_646), .b(output_15_7), .y(output_14_646));
wire output_16_646, output_16_7, output_15_646;
mixer gate_output_15_646(.a(output_16_646), .b(output_16_7), .y(output_15_646));
wire output_1_647, output_1_8, output_0_647;
mixer gate_output_0_647(.a(output_1_647), .b(output_1_8), .y(output_0_647));
wire output_2_647, output_2_8, output_1_647;
mixer gate_output_1_647(.a(output_2_647), .b(output_2_8), .y(output_1_647));
wire output_3_647, output_3_8, output_2_647;
mixer gate_output_2_647(.a(output_3_647), .b(output_3_8), .y(output_2_647));
wire output_4_647, output_4_8, output_3_647;
mixer gate_output_3_647(.a(output_4_647), .b(output_4_8), .y(output_3_647));
wire output_5_647, output_5_8, output_4_647;
mixer gate_output_4_647(.a(output_5_647), .b(output_5_8), .y(output_4_647));
wire output_6_647, output_6_8, output_5_647;
mixer gate_output_5_647(.a(output_6_647), .b(output_6_8), .y(output_5_647));
wire output_7_647, output_7_8, output_6_647;
mixer gate_output_6_647(.a(output_7_647), .b(output_7_8), .y(output_6_647));
wire output_8_647, output_8_8, output_7_647;
mixer gate_output_7_647(.a(output_8_647), .b(output_8_8), .y(output_7_647));
wire output_9_647, output_9_8, output_8_647;
mixer gate_output_8_647(.a(output_9_647), .b(output_9_8), .y(output_8_647));
wire output_10_647, output_10_8, output_9_647;
mixer gate_output_9_647(.a(output_10_647), .b(output_10_8), .y(output_9_647));
wire output_11_647, output_11_8, output_10_647;
mixer gate_output_10_647(.a(output_11_647), .b(output_11_8), .y(output_10_647));
wire output_12_647, output_12_8, output_11_647;
mixer gate_output_11_647(.a(output_12_647), .b(output_12_8), .y(output_11_647));
wire output_13_647, output_13_8, output_12_647;
mixer gate_output_12_647(.a(output_13_647), .b(output_13_8), .y(output_12_647));
wire output_14_647, output_14_8, output_13_647;
mixer gate_output_13_647(.a(output_14_647), .b(output_14_8), .y(output_13_647));
wire output_15_647, output_15_8, output_14_647;
mixer gate_output_14_647(.a(output_15_647), .b(output_15_8), .y(output_14_647));
wire output_16_647, output_16_8, output_15_647;
mixer gate_output_15_647(.a(output_16_647), .b(output_16_8), .y(output_15_647));
wire output_1_648, output_1_9, output_0_648;
mixer gate_output_0_648(.a(output_1_648), .b(output_1_9), .y(output_0_648));
wire output_2_648, output_2_9, output_1_648;
mixer gate_output_1_648(.a(output_2_648), .b(output_2_9), .y(output_1_648));
wire output_3_648, output_3_9, output_2_648;
mixer gate_output_2_648(.a(output_3_648), .b(output_3_9), .y(output_2_648));
wire output_4_648, output_4_9, output_3_648;
mixer gate_output_3_648(.a(output_4_648), .b(output_4_9), .y(output_3_648));
wire output_5_648, output_5_9, output_4_648;
mixer gate_output_4_648(.a(output_5_648), .b(output_5_9), .y(output_4_648));
wire output_6_648, output_6_9, output_5_648;
mixer gate_output_5_648(.a(output_6_648), .b(output_6_9), .y(output_5_648));
wire output_7_648, output_7_9, output_6_648;
mixer gate_output_6_648(.a(output_7_648), .b(output_7_9), .y(output_6_648));
wire output_8_648, output_8_9, output_7_648;
mixer gate_output_7_648(.a(output_8_648), .b(output_8_9), .y(output_7_648));
wire output_9_648, output_9_9, output_8_648;
mixer gate_output_8_648(.a(output_9_648), .b(output_9_9), .y(output_8_648));
wire output_10_648, output_10_9, output_9_648;
mixer gate_output_9_648(.a(output_10_648), .b(output_10_9), .y(output_9_648));
wire output_11_648, output_11_9, output_10_648;
mixer gate_output_10_648(.a(output_11_648), .b(output_11_9), .y(output_10_648));
wire output_12_648, output_12_9, output_11_648;
mixer gate_output_11_648(.a(output_12_648), .b(output_12_9), .y(output_11_648));
wire output_13_648, output_13_9, output_12_648;
mixer gate_output_12_648(.a(output_13_648), .b(output_13_9), .y(output_12_648));
wire output_14_648, output_14_9, output_13_648;
mixer gate_output_13_648(.a(output_14_648), .b(output_14_9), .y(output_13_648));
wire output_15_648, output_15_9, output_14_648;
mixer gate_output_14_648(.a(output_15_648), .b(output_15_9), .y(output_14_648));
wire output_16_648, output_16_9, output_15_648;
mixer gate_output_15_648(.a(output_16_648), .b(output_16_9), .y(output_15_648));
wire output_1_649, output_1_10, output_0_649;
mixer gate_output_0_649(.a(output_1_649), .b(output_1_10), .y(output_0_649));
wire output_2_649, output_2_10, output_1_649;
mixer gate_output_1_649(.a(output_2_649), .b(output_2_10), .y(output_1_649));
wire output_3_649, output_3_10, output_2_649;
mixer gate_output_2_649(.a(output_3_649), .b(output_3_10), .y(output_2_649));
wire output_4_649, output_4_10, output_3_649;
mixer gate_output_3_649(.a(output_4_649), .b(output_4_10), .y(output_3_649));
wire output_5_649, output_5_10, output_4_649;
mixer gate_output_4_649(.a(output_5_649), .b(output_5_10), .y(output_4_649));
wire output_6_649, output_6_10, output_5_649;
mixer gate_output_5_649(.a(output_6_649), .b(output_6_10), .y(output_5_649));
wire output_7_649, output_7_10, output_6_649;
mixer gate_output_6_649(.a(output_7_649), .b(output_7_10), .y(output_6_649));
wire output_8_649, output_8_10, output_7_649;
mixer gate_output_7_649(.a(output_8_649), .b(output_8_10), .y(output_7_649));
wire output_9_649, output_9_10, output_8_649;
mixer gate_output_8_649(.a(output_9_649), .b(output_9_10), .y(output_8_649));
wire output_10_649, output_10_10, output_9_649;
mixer gate_output_9_649(.a(output_10_649), .b(output_10_10), .y(output_9_649));
wire output_11_649, output_11_10, output_10_649;
mixer gate_output_10_649(.a(output_11_649), .b(output_11_10), .y(output_10_649));
wire output_12_649, output_12_10, output_11_649;
mixer gate_output_11_649(.a(output_12_649), .b(output_12_10), .y(output_11_649));
wire output_13_649, output_13_10, output_12_649;
mixer gate_output_12_649(.a(output_13_649), .b(output_13_10), .y(output_12_649));
wire output_14_649, output_14_10, output_13_649;
mixer gate_output_13_649(.a(output_14_649), .b(output_14_10), .y(output_13_649));
wire output_15_649, output_15_10, output_14_649;
mixer gate_output_14_649(.a(output_15_649), .b(output_15_10), .y(output_14_649));
wire output_16_649, output_16_10, output_15_649;
mixer gate_output_15_649(.a(output_16_649), .b(output_16_10), .y(output_15_649));
wire output_1_650, output_1_11, output_0_650;
mixer gate_output_0_650(.a(output_1_650), .b(output_1_11), .y(output_0_650));
wire output_2_650, output_2_11, output_1_650;
mixer gate_output_1_650(.a(output_2_650), .b(output_2_11), .y(output_1_650));
wire output_3_650, output_3_11, output_2_650;
mixer gate_output_2_650(.a(output_3_650), .b(output_3_11), .y(output_2_650));
wire output_4_650, output_4_11, output_3_650;
mixer gate_output_3_650(.a(output_4_650), .b(output_4_11), .y(output_3_650));
wire output_5_650, output_5_11, output_4_650;
mixer gate_output_4_650(.a(output_5_650), .b(output_5_11), .y(output_4_650));
wire output_6_650, output_6_11, output_5_650;
mixer gate_output_5_650(.a(output_6_650), .b(output_6_11), .y(output_5_650));
wire output_7_650, output_7_11, output_6_650;
mixer gate_output_6_650(.a(output_7_650), .b(output_7_11), .y(output_6_650));
wire output_8_650, output_8_11, output_7_650;
mixer gate_output_7_650(.a(output_8_650), .b(output_8_11), .y(output_7_650));
wire output_9_650, output_9_11, output_8_650;
mixer gate_output_8_650(.a(output_9_650), .b(output_9_11), .y(output_8_650));
wire output_10_650, output_10_11, output_9_650;
mixer gate_output_9_650(.a(output_10_650), .b(output_10_11), .y(output_9_650));
wire output_11_650, output_11_11, output_10_650;
mixer gate_output_10_650(.a(output_11_650), .b(output_11_11), .y(output_10_650));
wire output_12_650, output_12_11, output_11_650;
mixer gate_output_11_650(.a(output_12_650), .b(output_12_11), .y(output_11_650));
wire output_13_650, output_13_11, output_12_650;
mixer gate_output_12_650(.a(output_13_650), .b(output_13_11), .y(output_12_650));
wire output_14_650, output_14_11, output_13_650;
mixer gate_output_13_650(.a(output_14_650), .b(output_14_11), .y(output_13_650));
wire output_15_650, output_15_11, output_14_650;
mixer gate_output_14_650(.a(output_15_650), .b(output_15_11), .y(output_14_650));
wire output_16_650, output_16_11, output_15_650;
mixer gate_output_15_650(.a(output_16_650), .b(output_16_11), .y(output_15_650));
wire output_1_651, output_1_12, output_0_651;
mixer gate_output_0_651(.a(output_1_651), .b(output_1_12), .y(output_0_651));
wire output_2_651, output_2_12, output_1_651;
mixer gate_output_1_651(.a(output_2_651), .b(output_2_12), .y(output_1_651));
wire output_3_651, output_3_12, output_2_651;
mixer gate_output_2_651(.a(output_3_651), .b(output_3_12), .y(output_2_651));
wire output_4_651, output_4_12, output_3_651;
mixer gate_output_3_651(.a(output_4_651), .b(output_4_12), .y(output_3_651));
wire output_5_651, output_5_12, output_4_651;
mixer gate_output_4_651(.a(output_5_651), .b(output_5_12), .y(output_4_651));
wire output_6_651, output_6_12, output_5_651;
mixer gate_output_5_651(.a(output_6_651), .b(output_6_12), .y(output_5_651));
wire output_7_651, output_7_12, output_6_651;
mixer gate_output_6_651(.a(output_7_651), .b(output_7_12), .y(output_6_651));
wire output_8_651, output_8_12, output_7_651;
mixer gate_output_7_651(.a(output_8_651), .b(output_8_12), .y(output_7_651));
wire output_9_651, output_9_12, output_8_651;
mixer gate_output_8_651(.a(output_9_651), .b(output_9_12), .y(output_8_651));
wire output_10_651, output_10_12, output_9_651;
mixer gate_output_9_651(.a(output_10_651), .b(output_10_12), .y(output_9_651));
wire output_11_651, output_11_12, output_10_651;
mixer gate_output_10_651(.a(output_11_651), .b(output_11_12), .y(output_10_651));
wire output_12_651, output_12_12, output_11_651;
mixer gate_output_11_651(.a(output_12_651), .b(output_12_12), .y(output_11_651));
wire output_13_651, output_13_12, output_12_651;
mixer gate_output_12_651(.a(output_13_651), .b(output_13_12), .y(output_12_651));
wire output_14_651, output_14_12, output_13_651;
mixer gate_output_13_651(.a(output_14_651), .b(output_14_12), .y(output_13_651));
wire output_15_651, output_15_12, output_14_651;
mixer gate_output_14_651(.a(output_15_651), .b(output_15_12), .y(output_14_651));
wire output_16_651, output_16_12, output_15_651;
mixer gate_output_15_651(.a(output_16_651), .b(output_16_12), .y(output_15_651));
wire output_1_652, output_1_13, output_0_652;
mixer gate_output_0_652(.a(output_1_652), .b(output_1_13), .y(output_0_652));
wire output_2_652, output_2_13, output_1_652;
mixer gate_output_1_652(.a(output_2_652), .b(output_2_13), .y(output_1_652));
wire output_3_652, output_3_13, output_2_652;
mixer gate_output_2_652(.a(output_3_652), .b(output_3_13), .y(output_2_652));
wire output_4_652, output_4_13, output_3_652;
mixer gate_output_3_652(.a(output_4_652), .b(output_4_13), .y(output_3_652));
wire output_5_652, output_5_13, output_4_652;
mixer gate_output_4_652(.a(output_5_652), .b(output_5_13), .y(output_4_652));
wire output_6_652, output_6_13, output_5_652;
mixer gate_output_5_652(.a(output_6_652), .b(output_6_13), .y(output_5_652));
wire output_7_652, output_7_13, output_6_652;
mixer gate_output_6_652(.a(output_7_652), .b(output_7_13), .y(output_6_652));
wire output_8_652, output_8_13, output_7_652;
mixer gate_output_7_652(.a(output_8_652), .b(output_8_13), .y(output_7_652));
wire output_9_652, output_9_13, output_8_652;
mixer gate_output_8_652(.a(output_9_652), .b(output_9_13), .y(output_8_652));
wire output_10_652, output_10_13, output_9_652;
mixer gate_output_9_652(.a(output_10_652), .b(output_10_13), .y(output_9_652));
wire output_11_652, output_11_13, output_10_652;
mixer gate_output_10_652(.a(output_11_652), .b(output_11_13), .y(output_10_652));
wire output_12_652, output_12_13, output_11_652;
mixer gate_output_11_652(.a(output_12_652), .b(output_12_13), .y(output_11_652));
wire output_13_652, output_13_13, output_12_652;
mixer gate_output_12_652(.a(output_13_652), .b(output_13_13), .y(output_12_652));
wire output_14_652, output_14_13, output_13_652;
mixer gate_output_13_652(.a(output_14_652), .b(output_14_13), .y(output_13_652));
wire output_15_652, output_15_13, output_14_652;
mixer gate_output_14_652(.a(output_15_652), .b(output_15_13), .y(output_14_652));
wire output_16_652, output_16_13, output_15_652;
mixer gate_output_15_652(.a(output_16_652), .b(output_16_13), .y(output_15_652));
wire output_1_653, output_1_14, output_0_653;
mixer gate_output_0_653(.a(output_1_653), .b(output_1_14), .y(output_0_653));
wire output_2_653, output_2_14, output_1_653;
mixer gate_output_1_653(.a(output_2_653), .b(output_2_14), .y(output_1_653));
wire output_3_653, output_3_14, output_2_653;
mixer gate_output_2_653(.a(output_3_653), .b(output_3_14), .y(output_2_653));
wire output_4_653, output_4_14, output_3_653;
mixer gate_output_3_653(.a(output_4_653), .b(output_4_14), .y(output_3_653));
wire output_5_653, output_5_14, output_4_653;
mixer gate_output_4_653(.a(output_5_653), .b(output_5_14), .y(output_4_653));
wire output_6_653, output_6_14, output_5_653;
mixer gate_output_5_653(.a(output_6_653), .b(output_6_14), .y(output_5_653));
wire output_7_653, output_7_14, output_6_653;
mixer gate_output_6_653(.a(output_7_653), .b(output_7_14), .y(output_6_653));
wire output_8_653, output_8_14, output_7_653;
mixer gate_output_7_653(.a(output_8_653), .b(output_8_14), .y(output_7_653));
wire output_9_653, output_9_14, output_8_653;
mixer gate_output_8_653(.a(output_9_653), .b(output_9_14), .y(output_8_653));
wire output_10_653, output_10_14, output_9_653;
mixer gate_output_9_653(.a(output_10_653), .b(output_10_14), .y(output_9_653));
wire output_11_653, output_11_14, output_10_653;
mixer gate_output_10_653(.a(output_11_653), .b(output_11_14), .y(output_10_653));
wire output_12_653, output_12_14, output_11_653;
mixer gate_output_11_653(.a(output_12_653), .b(output_12_14), .y(output_11_653));
wire output_13_653, output_13_14, output_12_653;
mixer gate_output_12_653(.a(output_13_653), .b(output_13_14), .y(output_12_653));
wire output_14_653, output_14_14, output_13_653;
mixer gate_output_13_653(.a(output_14_653), .b(output_14_14), .y(output_13_653));
wire output_15_653, output_15_14, output_14_653;
mixer gate_output_14_653(.a(output_15_653), .b(output_15_14), .y(output_14_653));
wire output_16_653, output_16_14, output_15_653;
mixer gate_output_15_653(.a(output_16_653), .b(output_16_14), .y(output_15_653));
wire output_1_654, output_1_15, output_0_654;
mixer gate_output_0_654(.a(output_1_654), .b(output_1_15), .y(output_0_654));
wire output_2_654, output_2_15, output_1_654;
mixer gate_output_1_654(.a(output_2_654), .b(output_2_15), .y(output_1_654));
wire output_3_654, output_3_15, output_2_654;
mixer gate_output_2_654(.a(output_3_654), .b(output_3_15), .y(output_2_654));
wire output_4_654, output_4_15, output_3_654;
mixer gate_output_3_654(.a(output_4_654), .b(output_4_15), .y(output_3_654));
wire output_5_654, output_5_15, output_4_654;
mixer gate_output_4_654(.a(output_5_654), .b(output_5_15), .y(output_4_654));
wire output_6_654, output_6_15, output_5_654;
mixer gate_output_5_654(.a(output_6_654), .b(output_6_15), .y(output_5_654));
wire output_7_654, output_7_15, output_6_654;
mixer gate_output_6_654(.a(output_7_654), .b(output_7_15), .y(output_6_654));
wire output_8_654, output_8_15, output_7_654;
mixer gate_output_7_654(.a(output_8_654), .b(output_8_15), .y(output_7_654));
wire output_9_654, output_9_15, output_8_654;
mixer gate_output_8_654(.a(output_9_654), .b(output_9_15), .y(output_8_654));
wire output_10_654, output_10_15, output_9_654;
mixer gate_output_9_654(.a(output_10_654), .b(output_10_15), .y(output_9_654));
wire output_11_654, output_11_15, output_10_654;
mixer gate_output_10_654(.a(output_11_654), .b(output_11_15), .y(output_10_654));
wire output_12_654, output_12_15, output_11_654;
mixer gate_output_11_654(.a(output_12_654), .b(output_12_15), .y(output_11_654));
wire output_13_654, output_13_15, output_12_654;
mixer gate_output_12_654(.a(output_13_654), .b(output_13_15), .y(output_12_654));
wire output_14_654, output_14_15, output_13_654;
mixer gate_output_13_654(.a(output_14_654), .b(output_14_15), .y(output_13_654));
wire output_15_654, output_15_15, output_14_654;
mixer gate_output_14_654(.a(output_15_654), .b(output_15_15), .y(output_14_654));
wire output_16_654, output_16_15, output_15_654;
mixer gate_output_15_654(.a(output_16_654), .b(output_16_15), .y(output_15_654));
wire output_1_655, output_1_0, output_0_655;
mixer gate_output_0_655(.a(output_1_655), .b(output_1_0), .y(output_0_655));
wire output_2_655, output_2_0, output_1_655;
mixer gate_output_1_655(.a(output_2_655), .b(output_2_0), .y(output_1_655));
wire output_3_655, output_3_0, output_2_655;
mixer gate_output_2_655(.a(output_3_655), .b(output_3_0), .y(output_2_655));
wire output_4_655, output_4_0, output_3_655;
mixer gate_output_3_655(.a(output_4_655), .b(output_4_0), .y(output_3_655));
wire output_5_655, output_5_0, output_4_655;
mixer gate_output_4_655(.a(output_5_655), .b(output_5_0), .y(output_4_655));
wire output_6_655, output_6_0, output_5_655;
mixer gate_output_5_655(.a(output_6_655), .b(output_6_0), .y(output_5_655));
wire output_7_655, output_7_0, output_6_655;
mixer gate_output_6_655(.a(output_7_655), .b(output_7_0), .y(output_6_655));
wire output_8_655, output_8_0, output_7_655;
mixer gate_output_7_655(.a(output_8_655), .b(output_8_0), .y(output_7_655));
wire output_9_655, output_9_0, output_8_655;
mixer gate_output_8_655(.a(output_9_655), .b(output_9_0), .y(output_8_655));
wire output_10_655, output_10_0, output_9_655;
mixer gate_output_9_655(.a(output_10_655), .b(output_10_0), .y(output_9_655));
wire output_11_655, output_11_0, output_10_655;
mixer gate_output_10_655(.a(output_11_655), .b(output_11_0), .y(output_10_655));
wire output_12_655, output_12_0, output_11_655;
mixer gate_output_11_655(.a(output_12_655), .b(output_12_0), .y(output_11_655));
wire output_13_655, output_13_0, output_12_655;
mixer gate_output_12_655(.a(output_13_655), .b(output_13_0), .y(output_12_655));
wire output_14_655, output_14_0, output_13_655;
mixer gate_output_13_655(.a(output_14_655), .b(output_14_0), .y(output_13_655));
wire output_15_655, output_15_0, output_14_655;
mixer gate_output_14_655(.a(output_15_655), .b(output_15_0), .y(output_14_655));
wire output_16_655, output_16_0, output_15_655;
mixer gate_output_15_655(.a(output_16_655), .b(output_16_0), .y(output_15_655));
wire output_1_656, output_1_1, output_0_656;
mixer gate_output_0_656(.a(output_1_656), .b(output_1_1), .y(output_0_656));
wire output_2_656, output_2_1, output_1_656;
mixer gate_output_1_656(.a(output_2_656), .b(output_2_1), .y(output_1_656));
wire output_3_656, output_3_1, output_2_656;
mixer gate_output_2_656(.a(output_3_656), .b(output_3_1), .y(output_2_656));
wire output_4_656, output_4_1, output_3_656;
mixer gate_output_3_656(.a(output_4_656), .b(output_4_1), .y(output_3_656));
wire output_5_656, output_5_1, output_4_656;
mixer gate_output_4_656(.a(output_5_656), .b(output_5_1), .y(output_4_656));
wire output_6_656, output_6_1, output_5_656;
mixer gate_output_5_656(.a(output_6_656), .b(output_6_1), .y(output_5_656));
wire output_7_656, output_7_1, output_6_656;
mixer gate_output_6_656(.a(output_7_656), .b(output_7_1), .y(output_6_656));
wire output_8_656, output_8_1, output_7_656;
mixer gate_output_7_656(.a(output_8_656), .b(output_8_1), .y(output_7_656));
wire output_9_656, output_9_1, output_8_656;
mixer gate_output_8_656(.a(output_9_656), .b(output_9_1), .y(output_8_656));
wire output_10_656, output_10_1, output_9_656;
mixer gate_output_9_656(.a(output_10_656), .b(output_10_1), .y(output_9_656));
wire output_11_656, output_11_1, output_10_656;
mixer gate_output_10_656(.a(output_11_656), .b(output_11_1), .y(output_10_656));
wire output_12_656, output_12_1, output_11_656;
mixer gate_output_11_656(.a(output_12_656), .b(output_12_1), .y(output_11_656));
wire output_13_656, output_13_1, output_12_656;
mixer gate_output_12_656(.a(output_13_656), .b(output_13_1), .y(output_12_656));
wire output_14_656, output_14_1, output_13_656;
mixer gate_output_13_656(.a(output_14_656), .b(output_14_1), .y(output_13_656));
wire output_15_656, output_15_1, output_14_656;
mixer gate_output_14_656(.a(output_15_656), .b(output_15_1), .y(output_14_656));
wire output_16_656, output_16_1, output_15_656;
mixer gate_output_15_656(.a(output_16_656), .b(output_16_1), .y(output_15_656));
wire output_1_657, output_1_2, output_0_657;
mixer gate_output_0_657(.a(output_1_657), .b(output_1_2), .y(output_0_657));
wire output_2_657, output_2_2, output_1_657;
mixer gate_output_1_657(.a(output_2_657), .b(output_2_2), .y(output_1_657));
wire output_3_657, output_3_2, output_2_657;
mixer gate_output_2_657(.a(output_3_657), .b(output_3_2), .y(output_2_657));
wire output_4_657, output_4_2, output_3_657;
mixer gate_output_3_657(.a(output_4_657), .b(output_4_2), .y(output_3_657));
wire output_5_657, output_5_2, output_4_657;
mixer gate_output_4_657(.a(output_5_657), .b(output_5_2), .y(output_4_657));
wire output_6_657, output_6_2, output_5_657;
mixer gate_output_5_657(.a(output_6_657), .b(output_6_2), .y(output_5_657));
wire output_7_657, output_7_2, output_6_657;
mixer gate_output_6_657(.a(output_7_657), .b(output_7_2), .y(output_6_657));
wire output_8_657, output_8_2, output_7_657;
mixer gate_output_7_657(.a(output_8_657), .b(output_8_2), .y(output_7_657));
wire output_9_657, output_9_2, output_8_657;
mixer gate_output_8_657(.a(output_9_657), .b(output_9_2), .y(output_8_657));
wire output_10_657, output_10_2, output_9_657;
mixer gate_output_9_657(.a(output_10_657), .b(output_10_2), .y(output_9_657));
wire output_11_657, output_11_2, output_10_657;
mixer gate_output_10_657(.a(output_11_657), .b(output_11_2), .y(output_10_657));
wire output_12_657, output_12_2, output_11_657;
mixer gate_output_11_657(.a(output_12_657), .b(output_12_2), .y(output_11_657));
wire output_13_657, output_13_2, output_12_657;
mixer gate_output_12_657(.a(output_13_657), .b(output_13_2), .y(output_12_657));
wire output_14_657, output_14_2, output_13_657;
mixer gate_output_13_657(.a(output_14_657), .b(output_14_2), .y(output_13_657));
wire output_15_657, output_15_2, output_14_657;
mixer gate_output_14_657(.a(output_15_657), .b(output_15_2), .y(output_14_657));
wire output_16_657, output_16_2, output_15_657;
mixer gate_output_15_657(.a(output_16_657), .b(output_16_2), .y(output_15_657));
wire output_1_658, output_1_3, output_0_658;
mixer gate_output_0_658(.a(output_1_658), .b(output_1_3), .y(output_0_658));
wire output_2_658, output_2_3, output_1_658;
mixer gate_output_1_658(.a(output_2_658), .b(output_2_3), .y(output_1_658));
wire output_3_658, output_3_3, output_2_658;
mixer gate_output_2_658(.a(output_3_658), .b(output_3_3), .y(output_2_658));
wire output_4_658, output_4_3, output_3_658;
mixer gate_output_3_658(.a(output_4_658), .b(output_4_3), .y(output_3_658));
wire output_5_658, output_5_3, output_4_658;
mixer gate_output_4_658(.a(output_5_658), .b(output_5_3), .y(output_4_658));
wire output_6_658, output_6_3, output_5_658;
mixer gate_output_5_658(.a(output_6_658), .b(output_6_3), .y(output_5_658));
wire output_7_658, output_7_3, output_6_658;
mixer gate_output_6_658(.a(output_7_658), .b(output_7_3), .y(output_6_658));
wire output_8_658, output_8_3, output_7_658;
mixer gate_output_7_658(.a(output_8_658), .b(output_8_3), .y(output_7_658));
wire output_9_658, output_9_3, output_8_658;
mixer gate_output_8_658(.a(output_9_658), .b(output_9_3), .y(output_8_658));
wire output_10_658, output_10_3, output_9_658;
mixer gate_output_9_658(.a(output_10_658), .b(output_10_3), .y(output_9_658));
wire output_11_658, output_11_3, output_10_658;
mixer gate_output_10_658(.a(output_11_658), .b(output_11_3), .y(output_10_658));
wire output_12_658, output_12_3, output_11_658;
mixer gate_output_11_658(.a(output_12_658), .b(output_12_3), .y(output_11_658));
wire output_13_658, output_13_3, output_12_658;
mixer gate_output_12_658(.a(output_13_658), .b(output_13_3), .y(output_12_658));
wire output_14_658, output_14_3, output_13_658;
mixer gate_output_13_658(.a(output_14_658), .b(output_14_3), .y(output_13_658));
wire output_15_658, output_15_3, output_14_658;
mixer gate_output_14_658(.a(output_15_658), .b(output_15_3), .y(output_14_658));
wire output_16_658, output_16_3, output_15_658;
mixer gate_output_15_658(.a(output_16_658), .b(output_16_3), .y(output_15_658));
wire output_1_659, output_1_4, output_0_659;
mixer gate_output_0_659(.a(output_1_659), .b(output_1_4), .y(output_0_659));
wire output_2_659, output_2_4, output_1_659;
mixer gate_output_1_659(.a(output_2_659), .b(output_2_4), .y(output_1_659));
wire output_3_659, output_3_4, output_2_659;
mixer gate_output_2_659(.a(output_3_659), .b(output_3_4), .y(output_2_659));
wire output_4_659, output_4_4, output_3_659;
mixer gate_output_3_659(.a(output_4_659), .b(output_4_4), .y(output_3_659));
wire output_5_659, output_5_4, output_4_659;
mixer gate_output_4_659(.a(output_5_659), .b(output_5_4), .y(output_4_659));
wire output_6_659, output_6_4, output_5_659;
mixer gate_output_5_659(.a(output_6_659), .b(output_6_4), .y(output_5_659));
wire output_7_659, output_7_4, output_6_659;
mixer gate_output_6_659(.a(output_7_659), .b(output_7_4), .y(output_6_659));
wire output_8_659, output_8_4, output_7_659;
mixer gate_output_7_659(.a(output_8_659), .b(output_8_4), .y(output_7_659));
wire output_9_659, output_9_4, output_8_659;
mixer gate_output_8_659(.a(output_9_659), .b(output_9_4), .y(output_8_659));
wire output_10_659, output_10_4, output_9_659;
mixer gate_output_9_659(.a(output_10_659), .b(output_10_4), .y(output_9_659));
wire output_11_659, output_11_4, output_10_659;
mixer gate_output_10_659(.a(output_11_659), .b(output_11_4), .y(output_10_659));
wire output_12_659, output_12_4, output_11_659;
mixer gate_output_11_659(.a(output_12_659), .b(output_12_4), .y(output_11_659));
wire output_13_659, output_13_4, output_12_659;
mixer gate_output_12_659(.a(output_13_659), .b(output_13_4), .y(output_12_659));
wire output_14_659, output_14_4, output_13_659;
mixer gate_output_13_659(.a(output_14_659), .b(output_14_4), .y(output_13_659));
wire output_15_659, output_15_4, output_14_659;
mixer gate_output_14_659(.a(output_15_659), .b(output_15_4), .y(output_14_659));
wire output_16_659, output_16_4, output_15_659;
mixer gate_output_15_659(.a(output_16_659), .b(output_16_4), .y(output_15_659));
wire output_1_660, output_1_5, output_0_660;
mixer gate_output_0_660(.a(output_1_660), .b(output_1_5), .y(output_0_660));
wire output_2_660, output_2_5, output_1_660;
mixer gate_output_1_660(.a(output_2_660), .b(output_2_5), .y(output_1_660));
wire output_3_660, output_3_5, output_2_660;
mixer gate_output_2_660(.a(output_3_660), .b(output_3_5), .y(output_2_660));
wire output_4_660, output_4_5, output_3_660;
mixer gate_output_3_660(.a(output_4_660), .b(output_4_5), .y(output_3_660));
wire output_5_660, output_5_5, output_4_660;
mixer gate_output_4_660(.a(output_5_660), .b(output_5_5), .y(output_4_660));
wire output_6_660, output_6_5, output_5_660;
mixer gate_output_5_660(.a(output_6_660), .b(output_6_5), .y(output_5_660));
wire output_7_660, output_7_5, output_6_660;
mixer gate_output_6_660(.a(output_7_660), .b(output_7_5), .y(output_6_660));
wire output_8_660, output_8_5, output_7_660;
mixer gate_output_7_660(.a(output_8_660), .b(output_8_5), .y(output_7_660));
wire output_9_660, output_9_5, output_8_660;
mixer gate_output_8_660(.a(output_9_660), .b(output_9_5), .y(output_8_660));
wire output_10_660, output_10_5, output_9_660;
mixer gate_output_9_660(.a(output_10_660), .b(output_10_5), .y(output_9_660));
wire output_11_660, output_11_5, output_10_660;
mixer gate_output_10_660(.a(output_11_660), .b(output_11_5), .y(output_10_660));
wire output_12_660, output_12_5, output_11_660;
mixer gate_output_11_660(.a(output_12_660), .b(output_12_5), .y(output_11_660));
wire output_13_660, output_13_5, output_12_660;
mixer gate_output_12_660(.a(output_13_660), .b(output_13_5), .y(output_12_660));
wire output_14_660, output_14_5, output_13_660;
mixer gate_output_13_660(.a(output_14_660), .b(output_14_5), .y(output_13_660));
wire output_15_660, output_15_5, output_14_660;
mixer gate_output_14_660(.a(output_15_660), .b(output_15_5), .y(output_14_660));
wire output_16_660, output_16_5, output_15_660;
mixer gate_output_15_660(.a(output_16_660), .b(output_16_5), .y(output_15_660));
wire output_1_661, output_1_6, output_0_661;
mixer gate_output_0_661(.a(output_1_661), .b(output_1_6), .y(output_0_661));
wire output_2_661, output_2_6, output_1_661;
mixer gate_output_1_661(.a(output_2_661), .b(output_2_6), .y(output_1_661));
wire output_3_661, output_3_6, output_2_661;
mixer gate_output_2_661(.a(output_3_661), .b(output_3_6), .y(output_2_661));
wire output_4_661, output_4_6, output_3_661;
mixer gate_output_3_661(.a(output_4_661), .b(output_4_6), .y(output_3_661));
wire output_5_661, output_5_6, output_4_661;
mixer gate_output_4_661(.a(output_5_661), .b(output_5_6), .y(output_4_661));
wire output_6_661, output_6_6, output_5_661;
mixer gate_output_5_661(.a(output_6_661), .b(output_6_6), .y(output_5_661));
wire output_7_661, output_7_6, output_6_661;
mixer gate_output_6_661(.a(output_7_661), .b(output_7_6), .y(output_6_661));
wire output_8_661, output_8_6, output_7_661;
mixer gate_output_7_661(.a(output_8_661), .b(output_8_6), .y(output_7_661));
wire output_9_661, output_9_6, output_8_661;
mixer gate_output_8_661(.a(output_9_661), .b(output_9_6), .y(output_8_661));
wire output_10_661, output_10_6, output_9_661;
mixer gate_output_9_661(.a(output_10_661), .b(output_10_6), .y(output_9_661));
wire output_11_661, output_11_6, output_10_661;
mixer gate_output_10_661(.a(output_11_661), .b(output_11_6), .y(output_10_661));
wire output_12_661, output_12_6, output_11_661;
mixer gate_output_11_661(.a(output_12_661), .b(output_12_6), .y(output_11_661));
wire output_13_661, output_13_6, output_12_661;
mixer gate_output_12_661(.a(output_13_661), .b(output_13_6), .y(output_12_661));
wire output_14_661, output_14_6, output_13_661;
mixer gate_output_13_661(.a(output_14_661), .b(output_14_6), .y(output_13_661));
wire output_15_661, output_15_6, output_14_661;
mixer gate_output_14_661(.a(output_15_661), .b(output_15_6), .y(output_14_661));
wire output_16_661, output_16_6, output_15_661;
mixer gate_output_15_661(.a(output_16_661), .b(output_16_6), .y(output_15_661));
wire output_1_662, output_1_7, output_0_662;
mixer gate_output_0_662(.a(output_1_662), .b(output_1_7), .y(output_0_662));
wire output_2_662, output_2_7, output_1_662;
mixer gate_output_1_662(.a(output_2_662), .b(output_2_7), .y(output_1_662));
wire output_3_662, output_3_7, output_2_662;
mixer gate_output_2_662(.a(output_3_662), .b(output_3_7), .y(output_2_662));
wire output_4_662, output_4_7, output_3_662;
mixer gate_output_3_662(.a(output_4_662), .b(output_4_7), .y(output_3_662));
wire output_5_662, output_5_7, output_4_662;
mixer gate_output_4_662(.a(output_5_662), .b(output_5_7), .y(output_4_662));
wire output_6_662, output_6_7, output_5_662;
mixer gate_output_5_662(.a(output_6_662), .b(output_6_7), .y(output_5_662));
wire output_7_662, output_7_7, output_6_662;
mixer gate_output_6_662(.a(output_7_662), .b(output_7_7), .y(output_6_662));
wire output_8_662, output_8_7, output_7_662;
mixer gate_output_7_662(.a(output_8_662), .b(output_8_7), .y(output_7_662));
wire output_9_662, output_9_7, output_8_662;
mixer gate_output_8_662(.a(output_9_662), .b(output_9_7), .y(output_8_662));
wire output_10_662, output_10_7, output_9_662;
mixer gate_output_9_662(.a(output_10_662), .b(output_10_7), .y(output_9_662));
wire output_11_662, output_11_7, output_10_662;
mixer gate_output_10_662(.a(output_11_662), .b(output_11_7), .y(output_10_662));
wire output_12_662, output_12_7, output_11_662;
mixer gate_output_11_662(.a(output_12_662), .b(output_12_7), .y(output_11_662));
wire output_13_662, output_13_7, output_12_662;
mixer gate_output_12_662(.a(output_13_662), .b(output_13_7), .y(output_12_662));
wire output_14_662, output_14_7, output_13_662;
mixer gate_output_13_662(.a(output_14_662), .b(output_14_7), .y(output_13_662));
wire output_15_662, output_15_7, output_14_662;
mixer gate_output_14_662(.a(output_15_662), .b(output_15_7), .y(output_14_662));
wire output_16_662, output_16_7, output_15_662;
mixer gate_output_15_662(.a(output_16_662), .b(output_16_7), .y(output_15_662));
wire output_1_663, output_1_8, output_0_663;
mixer gate_output_0_663(.a(output_1_663), .b(output_1_8), .y(output_0_663));
wire output_2_663, output_2_8, output_1_663;
mixer gate_output_1_663(.a(output_2_663), .b(output_2_8), .y(output_1_663));
wire output_3_663, output_3_8, output_2_663;
mixer gate_output_2_663(.a(output_3_663), .b(output_3_8), .y(output_2_663));
wire output_4_663, output_4_8, output_3_663;
mixer gate_output_3_663(.a(output_4_663), .b(output_4_8), .y(output_3_663));
wire output_5_663, output_5_8, output_4_663;
mixer gate_output_4_663(.a(output_5_663), .b(output_5_8), .y(output_4_663));
wire output_6_663, output_6_8, output_5_663;
mixer gate_output_5_663(.a(output_6_663), .b(output_6_8), .y(output_5_663));
wire output_7_663, output_7_8, output_6_663;
mixer gate_output_6_663(.a(output_7_663), .b(output_7_8), .y(output_6_663));
wire output_8_663, output_8_8, output_7_663;
mixer gate_output_7_663(.a(output_8_663), .b(output_8_8), .y(output_7_663));
wire output_9_663, output_9_8, output_8_663;
mixer gate_output_8_663(.a(output_9_663), .b(output_9_8), .y(output_8_663));
wire output_10_663, output_10_8, output_9_663;
mixer gate_output_9_663(.a(output_10_663), .b(output_10_8), .y(output_9_663));
wire output_11_663, output_11_8, output_10_663;
mixer gate_output_10_663(.a(output_11_663), .b(output_11_8), .y(output_10_663));
wire output_12_663, output_12_8, output_11_663;
mixer gate_output_11_663(.a(output_12_663), .b(output_12_8), .y(output_11_663));
wire output_13_663, output_13_8, output_12_663;
mixer gate_output_12_663(.a(output_13_663), .b(output_13_8), .y(output_12_663));
wire output_14_663, output_14_8, output_13_663;
mixer gate_output_13_663(.a(output_14_663), .b(output_14_8), .y(output_13_663));
wire output_15_663, output_15_8, output_14_663;
mixer gate_output_14_663(.a(output_15_663), .b(output_15_8), .y(output_14_663));
wire output_16_663, output_16_8, output_15_663;
mixer gate_output_15_663(.a(output_16_663), .b(output_16_8), .y(output_15_663));
wire output_1_664, output_1_9, output_0_664;
mixer gate_output_0_664(.a(output_1_664), .b(output_1_9), .y(output_0_664));
wire output_2_664, output_2_9, output_1_664;
mixer gate_output_1_664(.a(output_2_664), .b(output_2_9), .y(output_1_664));
wire output_3_664, output_3_9, output_2_664;
mixer gate_output_2_664(.a(output_3_664), .b(output_3_9), .y(output_2_664));
wire output_4_664, output_4_9, output_3_664;
mixer gate_output_3_664(.a(output_4_664), .b(output_4_9), .y(output_3_664));
wire output_5_664, output_5_9, output_4_664;
mixer gate_output_4_664(.a(output_5_664), .b(output_5_9), .y(output_4_664));
wire output_6_664, output_6_9, output_5_664;
mixer gate_output_5_664(.a(output_6_664), .b(output_6_9), .y(output_5_664));
wire output_7_664, output_7_9, output_6_664;
mixer gate_output_6_664(.a(output_7_664), .b(output_7_9), .y(output_6_664));
wire output_8_664, output_8_9, output_7_664;
mixer gate_output_7_664(.a(output_8_664), .b(output_8_9), .y(output_7_664));
wire output_9_664, output_9_9, output_8_664;
mixer gate_output_8_664(.a(output_9_664), .b(output_9_9), .y(output_8_664));
wire output_10_664, output_10_9, output_9_664;
mixer gate_output_9_664(.a(output_10_664), .b(output_10_9), .y(output_9_664));
wire output_11_664, output_11_9, output_10_664;
mixer gate_output_10_664(.a(output_11_664), .b(output_11_9), .y(output_10_664));
wire output_12_664, output_12_9, output_11_664;
mixer gate_output_11_664(.a(output_12_664), .b(output_12_9), .y(output_11_664));
wire output_13_664, output_13_9, output_12_664;
mixer gate_output_12_664(.a(output_13_664), .b(output_13_9), .y(output_12_664));
wire output_14_664, output_14_9, output_13_664;
mixer gate_output_13_664(.a(output_14_664), .b(output_14_9), .y(output_13_664));
wire output_15_664, output_15_9, output_14_664;
mixer gate_output_14_664(.a(output_15_664), .b(output_15_9), .y(output_14_664));
wire output_16_664, output_16_9, output_15_664;
mixer gate_output_15_664(.a(output_16_664), .b(output_16_9), .y(output_15_664));
wire output_1_665, output_1_10, output_0_665;
mixer gate_output_0_665(.a(output_1_665), .b(output_1_10), .y(output_0_665));
wire output_2_665, output_2_10, output_1_665;
mixer gate_output_1_665(.a(output_2_665), .b(output_2_10), .y(output_1_665));
wire output_3_665, output_3_10, output_2_665;
mixer gate_output_2_665(.a(output_3_665), .b(output_3_10), .y(output_2_665));
wire output_4_665, output_4_10, output_3_665;
mixer gate_output_3_665(.a(output_4_665), .b(output_4_10), .y(output_3_665));
wire output_5_665, output_5_10, output_4_665;
mixer gate_output_4_665(.a(output_5_665), .b(output_5_10), .y(output_4_665));
wire output_6_665, output_6_10, output_5_665;
mixer gate_output_5_665(.a(output_6_665), .b(output_6_10), .y(output_5_665));
wire output_7_665, output_7_10, output_6_665;
mixer gate_output_6_665(.a(output_7_665), .b(output_7_10), .y(output_6_665));
wire output_8_665, output_8_10, output_7_665;
mixer gate_output_7_665(.a(output_8_665), .b(output_8_10), .y(output_7_665));
wire output_9_665, output_9_10, output_8_665;
mixer gate_output_8_665(.a(output_9_665), .b(output_9_10), .y(output_8_665));
wire output_10_665, output_10_10, output_9_665;
mixer gate_output_9_665(.a(output_10_665), .b(output_10_10), .y(output_9_665));
wire output_11_665, output_11_10, output_10_665;
mixer gate_output_10_665(.a(output_11_665), .b(output_11_10), .y(output_10_665));
wire output_12_665, output_12_10, output_11_665;
mixer gate_output_11_665(.a(output_12_665), .b(output_12_10), .y(output_11_665));
wire output_13_665, output_13_10, output_12_665;
mixer gate_output_12_665(.a(output_13_665), .b(output_13_10), .y(output_12_665));
wire output_14_665, output_14_10, output_13_665;
mixer gate_output_13_665(.a(output_14_665), .b(output_14_10), .y(output_13_665));
wire output_15_665, output_15_10, output_14_665;
mixer gate_output_14_665(.a(output_15_665), .b(output_15_10), .y(output_14_665));
wire output_16_665, output_16_10, output_15_665;
mixer gate_output_15_665(.a(output_16_665), .b(output_16_10), .y(output_15_665));
wire output_1_666, output_1_11, output_0_666;
mixer gate_output_0_666(.a(output_1_666), .b(output_1_11), .y(output_0_666));
wire output_2_666, output_2_11, output_1_666;
mixer gate_output_1_666(.a(output_2_666), .b(output_2_11), .y(output_1_666));
wire output_3_666, output_3_11, output_2_666;
mixer gate_output_2_666(.a(output_3_666), .b(output_3_11), .y(output_2_666));
wire output_4_666, output_4_11, output_3_666;
mixer gate_output_3_666(.a(output_4_666), .b(output_4_11), .y(output_3_666));
wire output_5_666, output_5_11, output_4_666;
mixer gate_output_4_666(.a(output_5_666), .b(output_5_11), .y(output_4_666));
wire output_6_666, output_6_11, output_5_666;
mixer gate_output_5_666(.a(output_6_666), .b(output_6_11), .y(output_5_666));
wire output_7_666, output_7_11, output_6_666;
mixer gate_output_6_666(.a(output_7_666), .b(output_7_11), .y(output_6_666));
wire output_8_666, output_8_11, output_7_666;
mixer gate_output_7_666(.a(output_8_666), .b(output_8_11), .y(output_7_666));
wire output_9_666, output_9_11, output_8_666;
mixer gate_output_8_666(.a(output_9_666), .b(output_9_11), .y(output_8_666));
wire output_10_666, output_10_11, output_9_666;
mixer gate_output_9_666(.a(output_10_666), .b(output_10_11), .y(output_9_666));
wire output_11_666, output_11_11, output_10_666;
mixer gate_output_10_666(.a(output_11_666), .b(output_11_11), .y(output_10_666));
wire output_12_666, output_12_11, output_11_666;
mixer gate_output_11_666(.a(output_12_666), .b(output_12_11), .y(output_11_666));
wire output_13_666, output_13_11, output_12_666;
mixer gate_output_12_666(.a(output_13_666), .b(output_13_11), .y(output_12_666));
wire output_14_666, output_14_11, output_13_666;
mixer gate_output_13_666(.a(output_14_666), .b(output_14_11), .y(output_13_666));
wire output_15_666, output_15_11, output_14_666;
mixer gate_output_14_666(.a(output_15_666), .b(output_15_11), .y(output_14_666));
wire output_16_666, output_16_11, output_15_666;
mixer gate_output_15_666(.a(output_16_666), .b(output_16_11), .y(output_15_666));
wire output_1_667, output_1_12, output_0_667;
mixer gate_output_0_667(.a(output_1_667), .b(output_1_12), .y(output_0_667));
wire output_2_667, output_2_12, output_1_667;
mixer gate_output_1_667(.a(output_2_667), .b(output_2_12), .y(output_1_667));
wire output_3_667, output_3_12, output_2_667;
mixer gate_output_2_667(.a(output_3_667), .b(output_3_12), .y(output_2_667));
wire output_4_667, output_4_12, output_3_667;
mixer gate_output_3_667(.a(output_4_667), .b(output_4_12), .y(output_3_667));
wire output_5_667, output_5_12, output_4_667;
mixer gate_output_4_667(.a(output_5_667), .b(output_5_12), .y(output_4_667));
wire output_6_667, output_6_12, output_5_667;
mixer gate_output_5_667(.a(output_6_667), .b(output_6_12), .y(output_5_667));
wire output_7_667, output_7_12, output_6_667;
mixer gate_output_6_667(.a(output_7_667), .b(output_7_12), .y(output_6_667));
wire output_8_667, output_8_12, output_7_667;
mixer gate_output_7_667(.a(output_8_667), .b(output_8_12), .y(output_7_667));
wire output_9_667, output_9_12, output_8_667;
mixer gate_output_8_667(.a(output_9_667), .b(output_9_12), .y(output_8_667));
wire output_10_667, output_10_12, output_9_667;
mixer gate_output_9_667(.a(output_10_667), .b(output_10_12), .y(output_9_667));
wire output_11_667, output_11_12, output_10_667;
mixer gate_output_10_667(.a(output_11_667), .b(output_11_12), .y(output_10_667));
wire output_12_667, output_12_12, output_11_667;
mixer gate_output_11_667(.a(output_12_667), .b(output_12_12), .y(output_11_667));
wire output_13_667, output_13_12, output_12_667;
mixer gate_output_12_667(.a(output_13_667), .b(output_13_12), .y(output_12_667));
wire output_14_667, output_14_12, output_13_667;
mixer gate_output_13_667(.a(output_14_667), .b(output_14_12), .y(output_13_667));
wire output_15_667, output_15_12, output_14_667;
mixer gate_output_14_667(.a(output_15_667), .b(output_15_12), .y(output_14_667));
wire output_16_667, output_16_12, output_15_667;
mixer gate_output_15_667(.a(output_16_667), .b(output_16_12), .y(output_15_667));
wire output_1_668, output_1_13, output_0_668;
mixer gate_output_0_668(.a(output_1_668), .b(output_1_13), .y(output_0_668));
wire output_2_668, output_2_13, output_1_668;
mixer gate_output_1_668(.a(output_2_668), .b(output_2_13), .y(output_1_668));
wire output_3_668, output_3_13, output_2_668;
mixer gate_output_2_668(.a(output_3_668), .b(output_3_13), .y(output_2_668));
wire output_4_668, output_4_13, output_3_668;
mixer gate_output_3_668(.a(output_4_668), .b(output_4_13), .y(output_3_668));
wire output_5_668, output_5_13, output_4_668;
mixer gate_output_4_668(.a(output_5_668), .b(output_5_13), .y(output_4_668));
wire output_6_668, output_6_13, output_5_668;
mixer gate_output_5_668(.a(output_6_668), .b(output_6_13), .y(output_5_668));
wire output_7_668, output_7_13, output_6_668;
mixer gate_output_6_668(.a(output_7_668), .b(output_7_13), .y(output_6_668));
wire output_8_668, output_8_13, output_7_668;
mixer gate_output_7_668(.a(output_8_668), .b(output_8_13), .y(output_7_668));
wire output_9_668, output_9_13, output_8_668;
mixer gate_output_8_668(.a(output_9_668), .b(output_9_13), .y(output_8_668));
wire output_10_668, output_10_13, output_9_668;
mixer gate_output_9_668(.a(output_10_668), .b(output_10_13), .y(output_9_668));
wire output_11_668, output_11_13, output_10_668;
mixer gate_output_10_668(.a(output_11_668), .b(output_11_13), .y(output_10_668));
wire output_12_668, output_12_13, output_11_668;
mixer gate_output_11_668(.a(output_12_668), .b(output_12_13), .y(output_11_668));
wire output_13_668, output_13_13, output_12_668;
mixer gate_output_12_668(.a(output_13_668), .b(output_13_13), .y(output_12_668));
wire output_14_668, output_14_13, output_13_668;
mixer gate_output_13_668(.a(output_14_668), .b(output_14_13), .y(output_13_668));
wire output_15_668, output_15_13, output_14_668;
mixer gate_output_14_668(.a(output_15_668), .b(output_15_13), .y(output_14_668));
wire output_16_668, output_16_13, output_15_668;
mixer gate_output_15_668(.a(output_16_668), .b(output_16_13), .y(output_15_668));
wire output_1_669, output_1_14, output_0_669;
mixer gate_output_0_669(.a(output_1_669), .b(output_1_14), .y(output_0_669));
wire output_2_669, output_2_14, output_1_669;
mixer gate_output_1_669(.a(output_2_669), .b(output_2_14), .y(output_1_669));
wire output_3_669, output_3_14, output_2_669;
mixer gate_output_2_669(.a(output_3_669), .b(output_3_14), .y(output_2_669));
wire output_4_669, output_4_14, output_3_669;
mixer gate_output_3_669(.a(output_4_669), .b(output_4_14), .y(output_3_669));
wire output_5_669, output_5_14, output_4_669;
mixer gate_output_4_669(.a(output_5_669), .b(output_5_14), .y(output_4_669));
wire output_6_669, output_6_14, output_5_669;
mixer gate_output_5_669(.a(output_6_669), .b(output_6_14), .y(output_5_669));
wire output_7_669, output_7_14, output_6_669;
mixer gate_output_6_669(.a(output_7_669), .b(output_7_14), .y(output_6_669));
wire output_8_669, output_8_14, output_7_669;
mixer gate_output_7_669(.a(output_8_669), .b(output_8_14), .y(output_7_669));
wire output_9_669, output_9_14, output_8_669;
mixer gate_output_8_669(.a(output_9_669), .b(output_9_14), .y(output_8_669));
wire output_10_669, output_10_14, output_9_669;
mixer gate_output_9_669(.a(output_10_669), .b(output_10_14), .y(output_9_669));
wire output_11_669, output_11_14, output_10_669;
mixer gate_output_10_669(.a(output_11_669), .b(output_11_14), .y(output_10_669));
wire output_12_669, output_12_14, output_11_669;
mixer gate_output_11_669(.a(output_12_669), .b(output_12_14), .y(output_11_669));
wire output_13_669, output_13_14, output_12_669;
mixer gate_output_12_669(.a(output_13_669), .b(output_13_14), .y(output_12_669));
wire output_14_669, output_14_14, output_13_669;
mixer gate_output_13_669(.a(output_14_669), .b(output_14_14), .y(output_13_669));
wire output_15_669, output_15_14, output_14_669;
mixer gate_output_14_669(.a(output_15_669), .b(output_15_14), .y(output_14_669));
wire output_16_669, output_16_14, output_15_669;
mixer gate_output_15_669(.a(output_16_669), .b(output_16_14), .y(output_15_669));
wire output_1_670, output_1_15, output_0_670;
mixer gate_output_0_670(.a(output_1_670), .b(output_1_15), .y(output_0_670));
wire output_2_670, output_2_15, output_1_670;
mixer gate_output_1_670(.a(output_2_670), .b(output_2_15), .y(output_1_670));
wire output_3_670, output_3_15, output_2_670;
mixer gate_output_2_670(.a(output_3_670), .b(output_3_15), .y(output_2_670));
wire output_4_670, output_4_15, output_3_670;
mixer gate_output_3_670(.a(output_4_670), .b(output_4_15), .y(output_3_670));
wire output_5_670, output_5_15, output_4_670;
mixer gate_output_4_670(.a(output_5_670), .b(output_5_15), .y(output_4_670));
wire output_6_670, output_6_15, output_5_670;
mixer gate_output_5_670(.a(output_6_670), .b(output_6_15), .y(output_5_670));
wire output_7_670, output_7_15, output_6_670;
mixer gate_output_6_670(.a(output_7_670), .b(output_7_15), .y(output_6_670));
wire output_8_670, output_8_15, output_7_670;
mixer gate_output_7_670(.a(output_8_670), .b(output_8_15), .y(output_7_670));
wire output_9_670, output_9_15, output_8_670;
mixer gate_output_8_670(.a(output_9_670), .b(output_9_15), .y(output_8_670));
wire output_10_670, output_10_15, output_9_670;
mixer gate_output_9_670(.a(output_10_670), .b(output_10_15), .y(output_9_670));
wire output_11_670, output_11_15, output_10_670;
mixer gate_output_10_670(.a(output_11_670), .b(output_11_15), .y(output_10_670));
wire output_12_670, output_12_15, output_11_670;
mixer gate_output_11_670(.a(output_12_670), .b(output_12_15), .y(output_11_670));
wire output_13_670, output_13_15, output_12_670;
mixer gate_output_12_670(.a(output_13_670), .b(output_13_15), .y(output_12_670));
wire output_14_670, output_14_15, output_13_670;
mixer gate_output_13_670(.a(output_14_670), .b(output_14_15), .y(output_13_670));
wire output_15_670, output_15_15, output_14_670;
mixer gate_output_14_670(.a(output_15_670), .b(output_15_15), .y(output_14_670));
wire output_16_670, output_16_15, output_15_670;
mixer gate_output_15_670(.a(output_16_670), .b(output_16_15), .y(output_15_670));
wire output_1_671, output_1_0, output_0_671;
mixer gate_output_0_671(.a(output_1_671), .b(output_1_0), .y(output_0_671));
wire output_2_671, output_2_0, output_1_671;
mixer gate_output_1_671(.a(output_2_671), .b(output_2_0), .y(output_1_671));
wire output_3_671, output_3_0, output_2_671;
mixer gate_output_2_671(.a(output_3_671), .b(output_3_0), .y(output_2_671));
wire output_4_671, output_4_0, output_3_671;
mixer gate_output_3_671(.a(output_4_671), .b(output_4_0), .y(output_3_671));
wire output_5_671, output_5_0, output_4_671;
mixer gate_output_4_671(.a(output_5_671), .b(output_5_0), .y(output_4_671));
wire output_6_671, output_6_0, output_5_671;
mixer gate_output_5_671(.a(output_6_671), .b(output_6_0), .y(output_5_671));
wire output_7_671, output_7_0, output_6_671;
mixer gate_output_6_671(.a(output_7_671), .b(output_7_0), .y(output_6_671));
wire output_8_671, output_8_0, output_7_671;
mixer gate_output_7_671(.a(output_8_671), .b(output_8_0), .y(output_7_671));
wire output_9_671, output_9_0, output_8_671;
mixer gate_output_8_671(.a(output_9_671), .b(output_9_0), .y(output_8_671));
wire output_10_671, output_10_0, output_9_671;
mixer gate_output_9_671(.a(output_10_671), .b(output_10_0), .y(output_9_671));
wire output_11_671, output_11_0, output_10_671;
mixer gate_output_10_671(.a(output_11_671), .b(output_11_0), .y(output_10_671));
wire output_12_671, output_12_0, output_11_671;
mixer gate_output_11_671(.a(output_12_671), .b(output_12_0), .y(output_11_671));
wire output_13_671, output_13_0, output_12_671;
mixer gate_output_12_671(.a(output_13_671), .b(output_13_0), .y(output_12_671));
wire output_14_671, output_14_0, output_13_671;
mixer gate_output_13_671(.a(output_14_671), .b(output_14_0), .y(output_13_671));
wire output_15_671, output_15_0, output_14_671;
mixer gate_output_14_671(.a(output_15_671), .b(output_15_0), .y(output_14_671));
wire output_16_671, output_16_0, output_15_671;
mixer gate_output_15_671(.a(output_16_671), .b(output_16_0), .y(output_15_671));
wire output_1_672, output_1_1, output_0_672;
mixer gate_output_0_672(.a(output_1_672), .b(output_1_1), .y(output_0_672));
wire output_2_672, output_2_1, output_1_672;
mixer gate_output_1_672(.a(output_2_672), .b(output_2_1), .y(output_1_672));
wire output_3_672, output_3_1, output_2_672;
mixer gate_output_2_672(.a(output_3_672), .b(output_3_1), .y(output_2_672));
wire output_4_672, output_4_1, output_3_672;
mixer gate_output_3_672(.a(output_4_672), .b(output_4_1), .y(output_3_672));
wire output_5_672, output_5_1, output_4_672;
mixer gate_output_4_672(.a(output_5_672), .b(output_5_1), .y(output_4_672));
wire output_6_672, output_6_1, output_5_672;
mixer gate_output_5_672(.a(output_6_672), .b(output_6_1), .y(output_5_672));
wire output_7_672, output_7_1, output_6_672;
mixer gate_output_6_672(.a(output_7_672), .b(output_7_1), .y(output_6_672));
wire output_8_672, output_8_1, output_7_672;
mixer gate_output_7_672(.a(output_8_672), .b(output_8_1), .y(output_7_672));
wire output_9_672, output_9_1, output_8_672;
mixer gate_output_8_672(.a(output_9_672), .b(output_9_1), .y(output_8_672));
wire output_10_672, output_10_1, output_9_672;
mixer gate_output_9_672(.a(output_10_672), .b(output_10_1), .y(output_9_672));
wire output_11_672, output_11_1, output_10_672;
mixer gate_output_10_672(.a(output_11_672), .b(output_11_1), .y(output_10_672));
wire output_12_672, output_12_1, output_11_672;
mixer gate_output_11_672(.a(output_12_672), .b(output_12_1), .y(output_11_672));
wire output_13_672, output_13_1, output_12_672;
mixer gate_output_12_672(.a(output_13_672), .b(output_13_1), .y(output_12_672));
wire output_14_672, output_14_1, output_13_672;
mixer gate_output_13_672(.a(output_14_672), .b(output_14_1), .y(output_13_672));
wire output_15_672, output_15_1, output_14_672;
mixer gate_output_14_672(.a(output_15_672), .b(output_15_1), .y(output_14_672));
wire output_16_672, output_16_1, output_15_672;
mixer gate_output_15_672(.a(output_16_672), .b(output_16_1), .y(output_15_672));
wire output_1_673, output_1_2, output_0_673;
mixer gate_output_0_673(.a(output_1_673), .b(output_1_2), .y(output_0_673));
wire output_2_673, output_2_2, output_1_673;
mixer gate_output_1_673(.a(output_2_673), .b(output_2_2), .y(output_1_673));
wire output_3_673, output_3_2, output_2_673;
mixer gate_output_2_673(.a(output_3_673), .b(output_3_2), .y(output_2_673));
wire output_4_673, output_4_2, output_3_673;
mixer gate_output_3_673(.a(output_4_673), .b(output_4_2), .y(output_3_673));
wire output_5_673, output_5_2, output_4_673;
mixer gate_output_4_673(.a(output_5_673), .b(output_5_2), .y(output_4_673));
wire output_6_673, output_6_2, output_5_673;
mixer gate_output_5_673(.a(output_6_673), .b(output_6_2), .y(output_5_673));
wire output_7_673, output_7_2, output_6_673;
mixer gate_output_6_673(.a(output_7_673), .b(output_7_2), .y(output_6_673));
wire output_8_673, output_8_2, output_7_673;
mixer gate_output_7_673(.a(output_8_673), .b(output_8_2), .y(output_7_673));
wire output_9_673, output_9_2, output_8_673;
mixer gate_output_8_673(.a(output_9_673), .b(output_9_2), .y(output_8_673));
wire output_10_673, output_10_2, output_9_673;
mixer gate_output_9_673(.a(output_10_673), .b(output_10_2), .y(output_9_673));
wire output_11_673, output_11_2, output_10_673;
mixer gate_output_10_673(.a(output_11_673), .b(output_11_2), .y(output_10_673));
wire output_12_673, output_12_2, output_11_673;
mixer gate_output_11_673(.a(output_12_673), .b(output_12_2), .y(output_11_673));
wire output_13_673, output_13_2, output_12_673;
mixer gate_output_12_673(.a(output_13_673), .b(output_13_2), .y(output_12_673));
wire output_14_673, output_14_2, output_13_673;
mixer gate_output_13_673(.a(output_14_673), .b(output_14_2), .y(output_13_673));
wire output_15_673, output_15_2, output_14_673;
mixer gate_output_14_673(.a(output_15_673), .b(output_15_2), .y(output_14_673));
wire output_16_673, output_16_2, output_15_673;
mixer gate_output_15_673(.a(output_16_673), .b(output_16_2), .y(output_15_673));
wire output_1_674, output_1_3, output_0_674;
mixer gate_output_0_674(.a(output_1_674), .b(output_1_3), .y(output_0_674));
wire output_2_674, output_2_3, output_1_674;
mixer gate_output_1_674(.a(output_2_674), .b(output_2_3), .y(output_1_674));
wire output_3_674, output_3_3, output_2_674;
mixer gate_output_2_674(.a(output_3_674), .b(output_3_3), .y(output_2_674));
wire output_4_674, output_4_3, output_3_674;
mixer gate_output_3_674(.a(output_4_674), .b(output_4_3), .y(output_3_674));
wire output_5_674, output_5_3, output_4_674;
mixer gate_output_4_674(.a(output_5_674), .b(output_5_3), .y(output_4_674));
wire output_6_674, output_6_3, output_5_674;
mixer gate_output_5_674(.a(output_6_674), .b(output_6_3), .y(output_5_674));
wire output_7_674, output_7_3, output_6_674;
mixer gate_output_6_674(.a(output_7_674), .b(output_7_3), .y(output_6_674));
wire output_8_674, output_8_3, output_7_674;
mixer gate_output_7_674(.a(output_8_674), .b(output_8_3), .y(output_7_674));
wire output_9_674, output_9_3, output_8_674;
mixer gate_output_8_674(.a(output_9_674), .b(output_9_3), .y(output_8_674));
wire output_10_674, output_10_3, output_9_674;
mixer gate_output_9_674(.a(output_10_674), .b(output_10_3), .y(output_9_674));
wire output_11_674, output_11_3, output_10_674;
mixer gate_output_10_674(.a(output_11_674), .b(output_11_3), .y(output_10_674));
wire output_12_674, output_12_3, output_11_674;
mixer gate_output_11_674(.a(output_12_674), .b(output_12_3), .y(output_11_674));
wire output_13_674, output_13_3, output_12_674;
mixer gate_output_12_674(.a(output_13_674), .b(output_13_3), .y(output_12_674));
wire output_14_674, output_14_3, output_13_674;
mixer gate_output_13_674(.a(output_14_674), .b(output_14_3), .y(output_13_674));
wire output_15_674, output_15_3, output_14_674;
mixer gate_output_14_674(.a(output_15_674), .b(output_15_3), .y(output_14_674));
wire output_16_674, output_16_3, output_15_674;
mixer gate_output_15_674(.a(output_16_674), .b(output_16_3), .y(output_15_674));
wire output_1_675, output_1_4, output_0_675;
mixer gate_output_0_675(.a(output_1_675), .b(output_1_4), .y(output_0_675));
wire output_2_675, output_2_4, output_1_675;
mixer gate_output_1_675(.a(output_2_675), .b(output_2_4), .y(output_1_675));
wire output_3_675, output_3_4, output_2_675;
mixer gate_output_2_675(.a(output_3_675), .b(output_3_4), .y(output_2_675));
wire output_4_675, output_4_4, output_3_675;
mixer gate_output_3_675(.a(output_4_675), .b(output_4_4), .y(output_3_675));
wire output_5_675, output_5_4, output_4_675;
mixer gate_output_4_675(.a(output_5_675), .b(output_5_4), .y(output_4_675));
wire output_6_675, output_6_4, output_5_675;
mixer gate_output_5_675(.a(output_6_675), .b(output_6_4), .y(output_5_675));
wire output_7_675, output_7_4, output_6_675;
mixer gate_output_6_675(.a(output_7_675), .b(output_7_4), .y(output_6_675));
wire output_8_675, output_8_4, output_7_675;
mixer gate_output_7_675(.a(output_8_675), .b(output_8_4), .y(output_7_675));
wire output_9_675, output_9_4, output_8_675;
mixer gate_output_8_675(.a(output_9_675), .b(output_9_4), .y(output_8_675));
wire output_10_675, output_10_4, output_9_675;
mixer gate_output_9_675(.a(output_10_675), .b(output_10_4), .y(output_9_675));
wire output_11_675, output_11_4, output_10_675;
mixer gate_output_10_675(.a(output_11_675), .b(output_11_4), .y(output_10_675));
wire output_12_675, output_12_4, output_11_675;
mixer gate_output_11_675(.a(output_12_675), .b(output_12_4), .y(output_11_675));
wire output_13_675, output_13_4, output_12_675;
mixer gate_output_12_675(.a(output_13_675), .b(output_13_4), .y(output_12_675));
wire output_14_675, output_14_4, output_13_675;
mixer gate_output_13_675(.a(output_14_675), .b(output_14_4), .y(output_13_675));
wire output_15_675, output_15_4, output_14_675;
mixer gate_output_14_675(.a(output_15_675), .b(output_15_4), .y(output_14_675));
wire output_16_675, output_16_4, output_15_675;
mixer gate_output_15_675(.a(output_16_675), .b(output_16_4), .y(output_15_675));
wire output_1_676, output_1_5, output_0_676;
mixer gate_output_0_676(.a(output_1_676), .b(output_1_5), .y(output_0_676));
wire output_2_676, output_2_5, output_1_676;
mixer gate_output_1_676(.a(output_2_676), .b(output_2_5), .y(output_1_676));
wire output_3_676, output_3_5, output_2_676;
mixer gate_output_2_676(.a(output_3_676), .b(output_3_5), .y(output_2_676));
wire output_4_676, output_4_5, output_3_676;
mixer gate_output_3_676(.a(output_4_676), .b(output_4_5), .y(output_3_676));
wire output_5_676, output_5_5, output_4_676;
mixer gate_output_4_676(.a(output_5_676), .b(output_5_5), .y(output_4_676));
wire output_6_676, output_6_5, output_5_676;
mixer gate_output_5_676(.a(output_6_676), .b(output_6_5), .y(output_5_676));
wire output_7_676, output_7_5, output_6_676;
mixer gate_output_6_676(.a(output_7_676), .b(output_7_5), .y(output_6_676));
wire output_8_676, output_8_5, output_7_676;
mixer gate_output_7_676(.a(output_8_676), .b(output_8_5), .y(output_7_676));
wire output_9_676, output_9_5, output_8_676;
mixer gate_output_8_676(.a(output_9_676), .b(output_9_5), .y(output_8_676));
wire output_10_676, output_10_5, output_9_676;
mixer gate_output_9_676(.a(output_10_676), .b(output_10_5), .y(output_9_676));
wire output_11_676, output_11_5, output_10_676;
mixer gate_output_10_676(.a(output_11_676), .b(output_11_5), .y(output_10_676));
wire output_12_676, output_12_5, output_11_676;
mixer gate_output_11_676(.a(output_12_676), .b(output_12_5), .y(output_11_676));
wire output_13_676, output_13_5, output_12_676;
mixer gate_output_12_676(.a(output_13_676), .b(output_13_5), .y(output_12_676));
wire output_14_676, output_14_5, output_13_676;
mixer gate_output_13_676(.a(output_14_676), .b(output_14_5), .y(output_13_676));
wire output_15_676, output_15_5, output_14_676;
mixer gate_output_14_676(.a(output_15_676), .b(output_15_5), .y(output_14_676));
wire output_16_676, output_16_5, output_15_676;
mixer gate_output_15_676(.a(output_16_676), .b(output_16_5), .y(output_15_676));
wire output_1_677, output_1_6, output_0_677;
mixer gate_output_0_677(.a(output_1_677), .b(output_1_6), .y(output_0_677));
wire output_2_677, output_2_6, output_1_677;
mixer gate_output_1_677(.a(output_2_677), .b(output_2_6), .y(output_1_677));
wire output_3_677, output_3_6, output_2_677;
mixer gate_output_2_677(.a(output_3_677), .b(output_3_6), .y(output_2_677));
wire output_4_677, output_4_6, output_3_677;
mixer gate_output_3_677(.a(output_4_677), .b(output_4_6), .y(output_3_677));
wire output_5_677, output_5_6, output_4_677;
mixer gate_output_4_677(.a(output_5_677), .b(output_5_6), .y(output_4_677));
wire output_6_677, output_6_6, output_5_677;
mixer gate_output_5_677(.a(output_6_677), .b(output_6_6), .y(output_5_677));
wire output_7_677, output_7_6, output_6_677;
mixer gate_output_6_677(.a(output_7_677), .b(output_7_6), .y(output_6_677));
wire output_8_677, output_8_6, output_7_677;
mixer gate_output_7_677(.a(output_8_677), .b(output_8_6), .y(output_7_677));
wire output_9_677, output_9_6, output_8_677;
mixer gate_output_8_677(.a(output_9_677), .b(output_9_6), .y(output_8_677));
wire output_10_677, output_10_6, output_9_677;
mixer gate_output_9_677(.a(output_10_677), .b(output_10_6), .y(output_9_677));
wire output_11_677, output_11_6, output_10_677;
mixer gate_output_10_677(.a(output_11_677), .b(output_11_6), .y(output_10_677));
wire output_12_677, output_12_6, output_11_677;
mixer gate_output_11_677(.a(output_12_677), .b(output_12_6), .y(output_11_677));
wire output_13_677, output_13_6, output_12_677;
mixer gate_output_12_677(.a(output_13_677), .b(output_13_6), .y(output_12_677));
wire output_14_677, output_14_6, output_13_677;
mixer gate_output_13_677(.a(output_14_677), .b(output_14_6), .y(output_13_677));
wire output_15_677, output_15_6, output_14_677;
mixer gate_output_14_677(.a(output_15_677), .b(output_15_6), .y(output_14_677));
wire output_16_677, output_16_6, output_15_677;
mixer gate_output_15_677(.a(output_16_677), .b(output_16_6), .y(output_15_677));
wire output_1_678, output_1_7, output_0_678;
mixer gate_output_0_678(.a(output_1_678), .b(output_1_7), .y(output_0_678));
wire output_2_678, output_2_7, output_1_678;
mixer gate_output_1_678(.a(output_2_678), .b(output_2_7), .y(output_1_678));
wire output_3_678, output_3_7, output_2_678;
mixer gate_output_2_678(.a(output_3_678), .b(output_3_7), .y(output_2_678));
wire output_4_678, output_4_7, output_3_678;
mixer gate_output_3_678(.a(output_4_678), .b(output_4_7), .y(output_3_678));
wire output_5_678, output_5_7, output_4_678;
mixer gate_output_4_678(.a(output_5_678), .b(output_5_7), .y(output_4_678));
wire output_6_678, output_6_7, output_5_678;
mixer gate_output_5_678(.a(output_6_678), .b(output_6_7), .y(output_5_678));
wire output_7_678, output_7_7, output_6_678;
mixer gate_output_6_678(.a(output_7_678), .b(output_7_7), .y(output_6_678));
wire output_8_678, output_8_7, output_7_678;
mixer gate_output_7_678(.a(output_8_678), .b(output_8_7), .y(output_7_678));
wire output_9_678, output_9_7, output_8_678;
mixer gate_output_8_678(.a(output_9_678), .b(output_9_7), .y(output_8_678));
wire output_10_678, output_10_7, output_9_678;
mixer gate_output_9_678(.a(output_10_678), .b(output_10_7), .y(output_9_678));
wire output_11_678, output_11_7, output_10_678;
mixer gate_output_10_678(.a(output_11_678), .b(output_11_7), .y(output_10_678));
wire output_12_678, output_12_7, output_11_678;
mixer gate_output_11_678(.a(output_12_678), .b(output_12_7), .y(output_11_678));
wire output_13_678, output_13_7, output_12_678;
mixer gate_output_12_678(.a(output_13_678), .b(output_13_7), .y(output_12_678));
wire output_14_678, output_14_7, output_13_678;
mixer gate_output_13_678(.a(output_14_678), .b(output_14_7), .y(output_13_678));
wire output_15_678, output_15_7, output_14_678;
mixer gate_output_14_678(.a(output_15_678), .b(output_15_7), .y(output_14_678));
wire output_16_678, output_16_7, output_15_678;
mixer gate_output_15_678(.a(output_16_678), .b(output_16_7), .y(output_15_678));
wire output_1_679, output_1_8, output_0_679;
mixer gate_output_0_679(.a(output_1_679), .b(output_1_8), .y(output_0_679));
wire output_2_679, output_2_8, output_1_679;
mixer gate_output_1_679(.a(output_2_679), .b(output_2_8), .y(output_1_679));
wire output_3_679, output_3_8, output_2_679;
mixer gate_output_2_679(.a(output_3_679), .b(output_3_8), .y(output_2_679));
wire output_4_679, output_4_8, output_3_679;
mixer gate_output_3_679(.a(output_4_679), .b(output_4_8), .y(output_3_679));
wire output_5_679, output_5_8, output_4_679;
mixer gate_output_4_679(.a(output_5_679), .b(output_5_8), .y(output_4_679));
wire output_6_679, output_6_8, output_5_679;
mixer gate_output_5_679(.a(output_6_679), .b(output_6_8), .y(output_5_679));
wire output_7_679, output_7_8, output_6_679;
mixer gate_output_6_679(.a(output_7_679), .b(output_7_8), .y(output_6_679));
wire output_8_679, output_8_8, output_7_679;
mixer gate_output_7_679(.a(output_8_679), .b(output_8_8), .y(output_7_679));
wire output_9_679, output_9_8, output_8_679;
mixer gate_output_8_679(.a(output_9_679), .b(output_9_8), .y(output_8_679));
wire output_10_679, output_10_8, output_9_679;
mixer gate_output_9_679(.a(output_10_679), .b(output_10_8), .y(output_9_679));
wire output_11_679, output_11_8, output_10_679;
mixer gate_output_10_679(.a(output_11_679), .b(output_11_8), .y(output_10_679));
wire output_12_679, output_12_8, output_11_679;
mixer gate_output_11_679(.a(output_12_679), .b(output_12_8), .y(output_11_679));
wire output_13_679, output_13_8, output_12_679;
mixer gate_output_12_679(.a(output_13_679), .b(output_13_8), .y(output_12_679));
wire output_14_679, output_14_8, output_13_679;
mixer gate_output_13_679(.a(output_14_679), .b(output_14_8), .y(output_13_679));
wire output_15_679, output_15_8, output_14_679;
mixer gate_output_14_679(.a(output_15_679), .b(output_15_8), .y(output_14_679));
wire output_16_679, output_16_8, output_15_679;
mixer gate_output_15_679(.a(output_16_679), .b(output_16_8), .y(output_15_679));
wire output_1_680, output_1_9, output_0_680;
mixer gate_output_0_680(.a(output_1_680), .b(output_1_9), .y(output_0_680));
wire output_2_680, output_2_9, output_1_680;
mixer gate_output_1_680(.a(output_2_680), .b(output_2_9), .y(output_1_680));
wire output_3_680, output_3_9, output_2_680;
mixer gate_output_2_680(.a(output_3_680), .b(output_3_9), .y(output_2_680));
wire output_4_680, output_4_9, output_3_680;
mixer gate_output_3_680(.a(output_4_680), .b(output_4_9), .y(output_3_680));
wire output_5_680, output_5_9, output_4_680;
mixer gate_output_4_680(.a(output_5_680), .b(output_5_9), .y(output_4_680));
wire output_6_680, output_6_9, output_5_680;
mixer gate_output_5_680(.a(output_6_680), .b(output_6_9), .y(output_5_680));
wire output_7_680, output_7_9, output_6_680;
mixer gate_output_6_680(.a(output_7_680), .b(output_7_9), .y(output_6_680));
wire output_8_680, output_8_9, output_7_680;
mixer gate_output_7_680(.a(output_8_680), .b(output_8_9), .y(output_7_680));
wire output_9_680, output_9_9, output_8_680;
mixer gate_output_8_680(.a(output_9_680), .b(output_9_9), .y(output_8_680));
wire output_10_680, output_10_9, output_9_680;
mixer gate_output_9_680(.a(output_10_680), .b(output_10_9), .y(output_9_680));
wire output_11_680, output_11_9, output_10_680;
mixer gate_output_10_680(.a(output_11_680), .b(output_11_9), .y(output_10_680));
wire output_12_680, output_12_9, output_11_680;
mixer gate_output_11_680(.a(output_12_680), .b(output_12_9), .y(output_11_680));
wire output_13_680, output_13_9, output_12_680;
mixer gate_output_12_680(.a(output_13_680), .b(output_13_9), .y(output_12_680));
wire output_14_680, output_14_9, output_13_680;
mixer gate_output_13_680(.a(output_14_680), .b(output_14_9), .y(output_13_680));
wire output_15_680, output_15_9, output_14_680;
mixer gate_output_14_680(.a(output_15_680), .b(output_15_9), .y(output_14_680));
wire output_16_680, output_16_9, output_15_680;
mixer gate_output_15_680(.a(output_16_680), .b(output_16_9), .y(output_15_680));
wire output_1_681, output_1_10, output_0_681;
mixer gate_output_0_681(.a(output_1_681), .b(output_1_10), .y(output_0_681));
wire output_2_681, output_2_10, output_1_681;
mixer gate_output_1_681(.a(output_2_681), .b(output_2_10), .y(output_1_681));
wire output_3_681, output_3_10, output_2_681;
mixer gate_output_2_681(.a(output_3_681), .b(output_3_10), .y(output_2_681));
wire output_4_681, output_4_10, output_3_681;
mixer gate_output_3_681(.a(output_4_681), .b(output_4_10), .y(output_3_681));
wire output_5_681, output_5_10, output_4_681;
mixer gate_output_4_681(.a(output_5_681), .b(output_5_10), .y(output_4_681));
wire output_6_681, output_6_10, output_5_681;
mixer gate_output_5_681(.a(output_6_681), .b(output_6_10), .y(output_5_681));
wire output_7_681, output_7_10, output_6_681;
mixer gate_output_6_681(.a(output_7_681), .b(output_7_10), .y(output_6_681));
wire output_8_681, output_8_10, output_7_681;
mixer gate_output_7_681(.a(output_8_681), .b(output_8_10), .y(output_7_681));
wire output_9_681, output_9_10, output_8_681;
mixer gate_output_8_681(.a(output_9_681), .b(output_9_10), .y(output_8_681));
wire output_10_681, output_10_10, output_9_681;
mixer gate_output_9_681(.a(output_10_681), .b(output_10_10), .y(output_9_681));
wire output_11_681, output_11_10, output_10_681;
mixer gate_output_10_681(.a(output_11_681), .b(output_11_10), .y(output_10_681));
wire output_12_681, output_12_10, output_11_681;
mixer gate_output_11_681(.a(output_12_681), .b(output_12_10), .y(output_11_681));
wire output_13_681, output_13_10, output_12_681;
mixer gate_output_12_681(.a(output_13_681), .b(output_13_10), .y(output_12_681));
wire output_14_681, output_14_10, output_13_681;
mixer gate_output_13_681(.a(output_14_681), .b(output_14_10), .y(output_13_681));
wire output_15_681, output_15_10, output_14_681;
mixer gate_output_14_681(.a(output_15_681), .b(output_15_10), .y(output_14_681));
wire output_16_681, output_16_10, output_15_681;
mixer gate_output_15_681(.a(output_16_681), .b(output_16_10), .y(output_15_681));
wire output_1_682, output_1_11, output_0_682;
mixer gate_output_0_682(.a(output_1_682), .b(output_1_11), .y(output_0_682));
wire output_2_682, output_2_11, output_1_682;
mixer gate_output_1_682(.a(output_2_682), .b(output_2_11), .y(output_1_682));
wire output_3_682, output_3_11, output_2_682;
mixer gate_output_2_682(.a(output_3_682), .b(output_3_11), .y(output_2_682));
wire output_4_682, output_4_11, output_3_682;
mixer gate_output_3_682(.a(output_4_682), .b(output_4_11), .y(output_3_682));
wire output_5_682, output_5_11, output_4_682;
mixer gate_output_4_682(.a(output_5_682), .b(output_5_11), .y(output_4_682));
wire output_6_682, output_6_11, output_5_682;
mixer gate_output_5_682(.a(output_6_682), .b(output_6_11), .y(output_5_682));
wire output_7_682, output_7_11, output_6_682;
mixer gate_output_6_682(.a(output_7_682), .b(output_7_11), .y(output_6_682));
wire output_8_682, output_8_11, output_7_682;
mixer gate_output_7_682(.a(output_8_682), .b(output_8_11), .y(output_7_682));
wire output_9_682, output_9_11, output_8_682;
mixer gate_output_8_682(.a(output_9_682), .b(output_9_11), .y(output_8_682));
wire output_10_682, output_10_11, output_9_682;
mixer gate_output_9_682(.a(output_10_682), .b(output_10_11), .y(output_9_682));
wire output_11_682, output_11_11, output_10_682;
mixer gate_output_10_682(.a(output_11_682), .b(output_11_11), .y(output_10_682));
wire output_12_682, output_12_11, output_11_682;
mixer gate_output_11_682(.a(output_12_682), .b(output_12_11), .y(output_11_682));
wire output_13_682, output_13_11, output_12_682;
mixer gate_output_12_682(.a(output_13_682), .b(output_13_11), .y(output_12_682));
wire output_14_682, output_14_11, output_13_682;
mixer gate_output_13_682(.a(output_14_682), .b(output_14_11), .y(output_13_682));
wire output_15_682, output_15_11, output_14_682;
mixer gate_output_14_682(.a(output_15_682), .b(output_15_11), .y(output_14_682));
wire output_16_682, output_16_11, output_15_682;
mixer gate_output_15_682(.a(output_16_682), .b(output_16_11), .y(output_15_682));
wire output_1_683, output_1_12, output_0_683;
mixer gate_output_0_683(.a(output_1_683), .b(output_1_12), .y(output_0_683));
wire output_2_683, output_2_12, output_1_683;
mixer gate_output_1_683(.a(output_2_683), .b(output_2_12), .y(output_1_683));
wire output_3_683, output_3_12, output_2_683;
mixer gate_output_2_683(.a(output_3_683), .b(output_3_12), .y(output_2_683));
wire output_4_683, output_4_12, output_3_683;
mixer gate_output_3_683(.a(output_4_683), .b(output_4_12), .y(output_3_683));
wire output_5_683, output_5_12, output_4_683;
mixer gate_output_4_683(.a(output_5_683), .b(output_5_12), .y(output_4_683));
wire output_6_683, output_6_12, output_5_683;
mixer gate_output_5_683(.a(output_6_683), .b(output_6_12), .y(output_5_683));
wire output_7_683, output_7_12, output_6_683;
mixer gate_output_6_683(.a(output_7_683), .b(output_7_12), .y(output_6_683));
wire output_8_683, output_8_12, output_7_683;
mixer gate_output_7_683(.a(output_8_683), .b(output_8_12), .y(output_7_683));
wire output_9_683, output_9_12, output_8_683;
mixer gate_output_8_683(.a(output_9_683), .b(output_9_12), .y(output_8_683));
wire output_10_683, output_10_12, output_9_683;
mixer gate_output_9_683(.a(output_10_683), .b(output_10_12), .y(output_9_683));
wire output_11_683, output_11_12, output_10_683;
mixer gate_output_10_683(.a(output_11_683), .b(output_11_12), .y(output_10_683));
wire output_12_683, output_12_12, output_11_683;
mixer gate_output_11_683(.a(output_12_683), .b(output_12_12), .y(output_11_683));
wire output_13_683, output_13_12, output_12_683;
mixer gate_output_12_683(.a(output_13_683), .b(output_13_12), .y(output_12_683));
wire output_14_683, output_14_12, output_13_683;
mixer gate_output_13_683(.a(output_14_683), .b(output_14_12), .y(output_13_683));
wire output_15_683, output_15_12, output_14_683;
mixer gate_output_14_683(.a(output_15_683), .b(output_15_12), .y(output_14_683));
wire output_16_683, output_16_12, output_15_683;
mixer gate_output_15_683(.a(output_16_683), .b(output_16_12), .y(output_15_683));
wire output_1_684, output_1_13, output_0_684;
mixer gate_output_0_684(.a(output_1_684), .b(output_1_13), .y(output_0_684));
wire output_2_684, output_2_13, output_1_684;
mixer gate_output_1_684(.a(output_2_684), .b(output_2_13), .y(output_1_684));
wire output_3_684, output_3_13, output_2_684;
mixer gate_output_2_684(.a(output_3_684), .b(output_3_13), .y(output_2_684));
wire output_4_684, output_4_13, output_3_684;
mixer gate_output_3_684(.a(output_4_684), .b(output_4_13), .y(output_3_684));
wire output_5_684, output_5_13, output_4_684;
mixer gate_output_4_684(.a(output_5_684), .b(output_5_13), .y(output_4_684));
wire output_6_684, output_6_13, output_5_684;
mixer gate_output_5_684(.a(output_6_684), .b(output_6_13), .y(output_5_684));
wire output_7_684, output_7_13, output_6_684;
mixer gate_output_6_684(.a(output_7_684), .b(output_7_13), .y(output_6_684));
wire output_8_684, output_8_13, output_7_684;
mixer gate_output_7_684(.a(output_8_684), .b(output_8_13), .y(output_7_684));
wire output_9_684, output_9_13, output_8_684;
mixer gate_output_8_684(.a(output_9_684), .b(output_9_13), .y(output_8_684));
wire output_10_684, output_10_13, output_9_684;
mixer gate_output_9_684(.a(output_10_684), .b(output_10_13), .y(output_9_684));
wire output_11_684, output_11_13, output_10_684;
mixer gate_output_10_684(.a(output_11_684), .b(output_11_13), .y(output_10_684));
wire output_12_684, output_12_13, output_11_684;
mixer gate_output_11_684(.a(output_12_684), .b(output_12_13), .y(output_11_684));
wire output_13_684, output_13_13, output_12_684;
mixer gate_output_12_684(.a(output_13_684), .b(output_13_13), .y(output_12_684));
wire output_14_684, output_14_13, output_13_684;
mixer gate_output_13_684(.a(output_14_684), .b(output_14_13), .y(output_13_684));
wire output_15_684, output_15_13, output_14_684;
mixer gate_output_14_684(.a(output_15_684), .b(output_15_13), .y(output_14_684));
wire output_16_684, output_16_13, output_15_684;
mixer gate_output_15_684(.a(output_16_684), .b(output_16_13), .y(output_15_684));
wire output_1_685, output_1_14, output_0_685;
mixer gate_output_0_685(.a(output_1_685), .b(output_1_14), .y(output_0_685));
wire output_2_685, output_2_14, output_1_685;
mixer gate_output_1_685(.a(output_2_685), .b(output_2_14), .y(output_1_685));
wire output_3_685, output_3_14, output_2_685;
mixer gate_output_2_685(.a(output_3_685), .b(output_3_14), .y(output_2_685));
wire output_4_685, output_4_14, output_3_685;
mixer gate_output_3_685(.a(output_4_685), .b(output_4_14), .y(output_3_685));
wire output_5_685, output_5_14, output_4_685;
mixer gate_output_4_685(.a(output_5_685), .b(output_5_14), .y(output_4_685));
wire output_6_685, output_6_14, output_5_685;
mixer gate_output_5_685(.a(output_6_685), .b(output_6_14), .y(output_5_685));
wire output_7_685, output_7_14, output_6_685;
mixer gate_output_6_685(.a(output_7_685), .b(output_7_14), .y(output_6_685));
wire output_8_685, output_8_14, output_7_685;
mixer gate_output_7_685(.a(output_8_685), .b(output_8_14), .y(output_7_685));
wire output_9_685, output_9_14, output_8_685;
mixer gate_output_8_685(.a(output_9_685), .b(output_9_14), .y(output_8_685));
wire output_10_685, output_10_14, output_9_685;
mixer gate_output_9_685(.a(output_10_685), .b(output_10_14), .y(output_9_685));
wire output_11_685, output_11_14, output_10_685;
mixer gate_output_10_685(.a(output_11_685), .b(output_11_14), .y(output_10_685));
wire output_12_685, output_12_14, output_11_685;
mixer gate_output_11_685(.a(output_12_685), .b(output_12_14), .y(output_11_685));
wire output_13_685, output_13_14, output_12_685;
mixer gate_output_12_685(.a(output_13_685), .b(output_13_14), .y(output_12_685));
wire output_14_685, output_14_14, output_13_685;
mixer gate_output_13_685(.a(output_14_685), .b(output_14_14), .y(output_13_685));
wire output_15_685, output_15_14, output_14_685;
mixer gate_output_14_685(.a(output_15_685), .b(output_15_14), .y(output_14_685));
wire output_16_685, output_16_14, output_15_685;
mixer gate_output_15_685(.a(output_16_685), .b(output_16_14), .y(output_15_685));
wire output_1_686, output_1_15, output_0_686;
mixer gate_output_0_686(.a(output_1_686), .b(output_1_15), .y(output_0_686));
wire output_2_686, output_2_15, output_1_686;
mixer gate_output_1_686(.a(output_2_686), .b(output_2_15), .y(output_1_686));
wire output_3_686, output_3_15, output_2_686;
mixer gate_output_2_686(.a(output_3_686), .b(output_3_15), .y(output_2_686));
wire output_4_686, output_4_15, output_3_686;
mixer gate_output_3_686(.a(output_4_686), .b(output_4_15), .y(output_3_686));
wire output_5_686, output_5_15, output_4_686;
mixer gate_output_4_686(.a(output_5_686), .b(output_5_15), .y(output_4_686));
wire output_6_686, output_6_15, output_5_686;
mixer gate_output_5_686(.a(output_6_686), .b(output_6_15), .y(output_5_686));
wire output_7_686, output_7_15, output_6_686;
mixer gate_output_6_686(.a(output_7_686), .b(output_7_15), .y(output_6_686));
wire output_8_686, output_8_15, output_7_686;
mixer gate_output_7_686(.a(output_8_686), .b(output_8_15), .y(output_7_686));
wire output_9_686, output_9_15, output_8_686;
mixer gate_output_8_686(.a(output_9_686), .b(output_9_15), .y(output_8_686));
wire output_10_686, output_10_15, output_9_686;
mixer gate_output_9_686(.a(output_10_686), .b(output_10_15), .y(output_9_686));
wire output_11_686, output_11_15, output_10_686;
mixer gate_output_10_686(.a(output_11_686), .b(output_11_15), .y(output_10_686));
wire output_12_686, output_12_15, output_11_686;
mixer gate_output_11_686(.a(output_12_686), .b(output_12_15), .y(output_11_686));
wire output_13_686, output_13_15, output_12_686;
mixer gate_output_12_686(.a(output_13_686), .b(output_13_15), .y(output_12_686));
wire output_14_686, output_14_15, output_13_686;
mixer gate_output_13_686(.a(output_14_686), .b(output_14_15), .y(output_13_686));
wire output_15_686, output_15_15, output_14_686;
mixer gate_output_14_686(.a(output_15_686), .b(output_15_15), .y(output_14_686));
wire output_16_686, output_16_15, output_15_686;
mixer gate_output_15_686(.a(output_16_686), .b(output_16_15), .y(output_15_686));
wire output_1_687, output_1_0, output_0_687;
mixer gate_output_0_687(.a(output_1_687), .b(output_1_0), .y(output_0_687));
wire output_2_687, output_2_0, output_1_687;
mixer gate_output_1_687(.a(output_2_687), .b(output_2_0), .y(output_1_687));
wire output_3_687, output_3_0, output_2_687;
mixer gate_output_2_687(.a(output_3_687), .b(output_3_0), .y(output_2_687));
wire output_4_687, output_4_0, output_3_687;
mixer gate_output_3_687(.a(output_4_687), .b(output_4_0), .y(output_3_687));
wire output_5_687, output_5_0, output_4_687;
mixer gate_output_4_687(.a(output_5_687), .b(output_5_0), .y(output_4_687));
wire output_6_687, output_6_0, output_5_687;
mixer gate_output_5_687(.a(output_6_687), .b(output_6_0), .y(output_5_687));
wire output_7_687, output_7_0, output_6_687;
mixer gate_output_6_687(.a(output_7_687), .b(output_7_0), .y(output_6_687));
wire output_8_687, output_8_0, output_7_687;
mixer gate_output_7_687(.a(output_8_687), .b(output_8_0), .y(output_7_687));
wire output_9_687, output_9_0, output_8_687;
mixer gate_output_8_687(.a(output_9_687), .b(output_9_0), .y(output_8_687));
wire output_10_687, output_10_0, output_9_687;
mixer gate_output_9_687(.a(output_10_687), .b(output_10_0), .y(output_9_687));
wire output_11_687, output_11_0, output_10_687;
mixer gate_output_10_687(.a(output_11_687), .b(output_11_0), .y(output_10_687));
wire output_12_687, output_12_0, output_11_687;
mixer gate_output_11_687(.a(output_12_687), .b(output_12_0), .y(output_11_687));
wire output_13_687, output_13_0, output_12_687;
mixer gate_output_12_687(.a(output_13_687), .b(output_13_0), .y(output_12_687));
wire output_14_687, output_14_0, output_13_687;
mixer gate_output_13_687(.a(output_14_687), .b(output_14_0), .y(output_13_687));
wire output_15_687, output_15_0, output_14_687;
mixer gate_output_14_687(.a(output_15_687), .b(output_15_0), .y(output_14_687));
wire output_16_687, output_16_0, output_15_687;
mixer gate_output_15_687(.a(output_16_687), .b(output_16_0), .y(output_15_687));
wire output_1_688, output_1_1, output_0_688;
mixer gate_output_0_688(.a(output_1_688), .b(output_1_1), .y(output_0_688));
wire output_2_688, output_2_1, output_1_688;
mixer gate_output_1_688(.a(output_2_688), .b(output_2_1), .y(output_1_688));
wire output_3_688, output_3_1, output_2_688;
mixer gate_output_2_688(.a(output_3_688), .b(output_3_1), .y(output_2_688));
wire output_4_688, output_4_1, output_3_688;
mixer gate_output_3_688(.a(output_4_688), .b(output_4_1), .y(output_3_688));
wire output_5_688, output_5_1, output_4_688;
mixer gate_output_4_688(.a(output_5_688), .b(output_5_1), .y(output_4_688));
wire output_6_688, output_6_1, output_5_688;
mixer gate_output_5_688(.a(output_6_688), .b(output_6_1), .y(output_5_688));
wire output_7_688, output_7_1, output_6_688;
mixer gate_output_6_688(.a(output_7_688), .b(output_7_1), .y(output_6_688));
wire output_8_688, output_8_1, output_7_688;
mixer gate_output_7_688(.a(output_8_688), .b(output_8_1), .y(output_7_688));
wire output_9_688, output_9_1, output_8_688;
mixer gate_output_8_688(.a(output_9_688), .b(output_9_1), .y(output_8_688));
wire output_10_688, output_10_1, output_9_688;
mixer gate_output_9_688(.a(output_10_688), .b(output_10_1), .y(output_9_688));
wire output_11_688, output_11_1, output_10_688;
mixer gate_output_10_688(.a(output_11_688), .b(output_11_1), .y(output_10_688));
wire output_12_688, output_12_1, output_11_688;
mixer gate_output_11_688(.a(output_12_688), .b(output_12_1), .y(output_11_688));
wire output_13_688, output_13_1, output_12_688;
mixer gate_output_12_688(.a(output_13_688), .b(output_13_1), .y(output_12_688));
wire output_14_688, output_14_1, output_13_688;
mixer gate_output_13_688(.a(output_14_688), .b(output_14_1), .y(output_13_688));
wire output_15_688, output_15_1, output_14_688;
mixer gate_output_14_688(.a(output_15_688), .b(output_15_1), .y(output_14_688));
wire output_16_688, output_16_1, output_15_688;
mixer gate_output_15_688(.a(output_16_688), .b(output_16_1), .y(output_15_688));
wire output_1_689, output_1_2, output_0_689;
mixer gate_output_0_689(.a(output_1_689), .b(output_1_2), .y(output_0_689));
wire output_2_689, output_2_2, output_1_689;
mixer gate_output_1_689(.a(output_2_689), .b(output_2_2), .y(output_1_689));
wire output_3_689, output_3_2, output_2_689;
mixer gate_output_2_689(.a(output_3_689), .b(output_3_2), .y(output_2_689));
wire output_4_689, output_4_2, output_3_689;
mixer gate_output_3_689(.a(output_4_689), .b(output_4_2), .y(output_3_689));
wire output_5_689, output_5_2, output_4_689;
mixer gate_output_4_689(.a(output_5_689), .b(output_5_2), .y(output_4_689));
wire output_6_689, output_6_2, output_5_689;
mixer gate_output_5_689(.a(output_6_689), .b(output_6_2), .y(output_5_689));
wire output_7_689, output_7_2, output_6_689;
mixer gate_output_6_689(.a(output_7_689), .b(output_7_2), .y(output_6_689));
wire output_8_689, output_8_2, output_7_689;
mixer gate_output_7_689(.a(output_8_689), .b(output_8_2), .y(output_7_689));
wire output_9_689, output_9_2, output_8_689;
mixer gate_output_8_689(.a(output_9_689), .b(output_9_2), .y(output_8_689));
wire output_10_689, output_10_2, output_9_689;
mixer gate_output_9_689(.a(output_10_689), .b(output_10_2), .y(output_9_689));
wire output_11_689, output_11_2, output_10_689;
mixer gate_output_10_689(.a(output_11_689), .b(output_11_2), .y(output_10_689));
wire output_12_689, output_12_2, output_11_689;
mixer gate_output_11_689(.a(output_12_689), .b(output_12_2), .y(output_11_689));
wire output_13_689, output_13_2, output_12_689;
mixer gate_output_12_689(.a(output_13_689), .b(output_13_2), .y(output_12_689));
wire output_14_689, output_14_2, output_13_689;
mixer gate_output_13_689(.a(output_14_689), .b(output_14_2), .y(output_13_689));
wire output_15_689, output_15_2, output_14_689;
mixer gate_output_14_689(.a(output_15_689), .b(output_15_2), .y(output_14_689));
wire output_16_689, output_16_2, output_15_689;
mixer gate_output_15_689(.a(output_16_689), .b(output_16_2), .y(output_15_689));
wire output_1_690, output_1_3, output_0_690;
mixer gate_output_0_690(.a(output_1_690), .b(output_1_3), .y(output_0_690));
wire output_2_690, output_2_3, output_1_690;
mixer gate_output_1_690(.a(output_2_690), .b(output_2_3), .y(output_1_690));
wire output_3_690, output_3_3, output_2_690;
mixer gate_output_2_690(.a(output_3_690), .b(output_3_3), .y(output_2_690));
wire output_4_690, output_4_3, output_3_690;
mixer gate_output_3_690(.a(output_4_690), .b(output_4_3), .y(output_3_690));
wire output_5_690, output_5_3, output_4_690;
mixer gate_output_4_690(.a(output_5_690), .b(output_5_3), .y(output_4_690));
wire output_6_690, output_6_3, output_5_690;
mixer gate_output_5_690(.a(output_6_690), .b(output_6_3), .y(output_5_690));
wire output_7_690, output_7_3, output_6_690;
mixer gate_output_6_690(.a(output_7_690), .b(output_7_3), .y(output_6_690));
wire output_8_690, output_8_3, output_7_690;
mixer gate_output_7_690(.a(output_8_690), .b(output_8_3), .y(output_7_690));
wire output_9_690, output_9_3, output_8_690;
mixer gate_output_8_690(.a(output_9_690), .b(output_9_3), .y(output_8_690));
wire output_10_690, output_10_3, output_9_690;
mixer gate_output_9_690(.a(output_10_690), .b(output_10_3), .y(output_9_690));
wire output_11_690, output_11_3, output_10_690;
mixer gate_output_10_690(.a(output_11_690), .b(output_11_3), .y(output_10_690));
wire output_12_690, output_12_3, output_11_690;
mixer gate_output_11_690(.a(output_12_690), .b(output_12_3), .y(output_11_690));
wire output_13_690, output_13_3, output_12_690;
mixer gate_output_12_690(.a(output_13_690), .b(output_13_3), .y(output_12_690));
wire output_14_690, output_14_3, output_13_690;
mixer gate_output_13_690(.a(output_14_690), .b(output_14_3), .y(output_13_690));
wire output_15_690, output_15_3, output_14_690;
mixer gate_output_14_690(.a(output_15_690), .b(output_15_3), .y(output_14_690));
wire output_16_690, output_16_3, output_15_690;
mixer gate_output_15_690(.a(output_16_690), .b(output_16_3), .y(output_15_690));
wire output_1_691, output_1_4, output_0_691;
mixer gate_output_0_691(.a(output_1_691), .b(output_1_4), .y(output_0_691));
wire output_2_691, output_2_4, output_1_691;
mixer gate_output_1_691(.a(output_2_691), .b(output_2_4), .y(output_1_691));
wire output_3_691, output_3_4, output_2_691;
mixer gate_output_2_691(.a(output_3_691), .b(output_3_4), .y(output_2_691));
wire output_4_691, output_4_4, output_3_691;
mixer gate_output_3_691(.a(output_4_691), .b(output_4_4), .y(output_3_691));
wire output_5_691, output_5_4, output_4_691;
mixer gate_output_4_691(.a(output_5_691), .b(output_5_4), .y(output_4_691));
wire output_6_691, output_6_4, output_5_691;
mixer gate_output_5_691(.a(output_6_691), .b(output_6_4), .y(output_5_691));
wire output_7_691, output_7_4, output_6_691;
mixer gate_output_6_691(.a(output_7_691), .b(output_7_4), .y(output_6_691));
wire output_8_691, output_8_4, output_7_691;
mixer gate_output_7_691(.a(output_8_691), .b(output_8_4), .y(output_7_691));
wire output_9_691, output_9_4, output_8_691;
mixer gate_output_8_691(.a(output_9_691), .b(output_9_4), .y(output_8_691));
wire output_10_691, output_10_4, output_9_691;
mixer gate_output_9_691(.a(output_10_691), .b(output_10_4), .y(output_9_691));
wire output_11_691, output_11_4, output_10_691;
mixer gate_output_10_691(.a(output_11_691), .b(output_11_4), .y(output_10_691));
wire output_12_691, output_12_4, output_11_691;
mixer gate_output_11_691(.a(output_12_691), .b(output_12_4), .y(output_11_691));
wire output_13_691, output_13_4, output_12_691;
mixer gate_output_12_691(.a(output_13_691), .b(output_13_4), .y(output_12_691));
wire output_14_691, output_14_4, output_13_691;
mixer gate_output_13_691(.a(output_14_691), .b(output_14_4), .y(output_13_691));
wire output_15_691, output_15_4, output_14_691;
mixer gate_output_14_691(.a(output_15_691), .b(output_15_4), .y(output_14_691));
wire output_16_691, output_16_4, output_15_691;
mixer gate_output_15_691(.a(output_16_691), .b(output_16_4), .y(output_15_691));
wire output_1_692, output_1_5, output_0_692;
mixer gate_output_0_692(.a(output_1_692), .b(output_1_5), .y(output_0_692));
wire output_2_692, output_2_5, output_1_692;
mixer gate_output_1_692(.a(output_2_692), .b(output_2_5), .y(output_1_692));
wire output_3_692, output_3_5, output_2_692;
mixer gate_output_2_692(.a(output_3_692), .b(output_3_5), .y(output_2_692));
wire output_4_692, output_4_5, output_3_692;
mixer gate_output_3_692(.a(output_4_692), .b(output_4_5), .y(output_3_692));
wire output_5_692, output_5_5, output_4_692;
mixer gate_output_4_692(.a(output_5_692), .b(output_5_5), .y(output_4_692));
wire output_6_692, output_6_5, output_5_692;
mixer gate_output_5_692(.a(output_6_692), .b(output_6_5), .y(output_5_692));
wire output_7_692, output_7_5, output_6_692;
mixer gate_output_6_692(.a(output_7_692), .b(output_7_5), .y(output_6_692));
wire output_8_692, output_8_5, output_7_692;
mixer gate_output_7_692(.a(output_8_692), .b(output_8_5), .y(output_7_692));
wire output_9_692, output_9_5, output_8_692;
mixer gate_output_8_692(.a(output_9_692), .b(output_9_5), .y(output_8_692));
wire output_10_692, output_10_5, output_9_692;
mixer gate_output_9_692(.a(output_10_692), .b(output_10_5), .y(output_9_692));
wire output_11_692, output_11_5, output_10_692;
mixer gate_output_10_692(.a(output_11_692), .b(output_11_5), .y(output_10_692));
wire output_12_692, output_12_5, output_11_692;
mixer gate_output_11_692(.a(output_12_692), .b(output_12_5), .y(output_11_692));
wire output_13_692, output_13_5, output_12_692;
mixer gate_output_12_692(.a(output_13_692), .b(output_13_5), .y(output_12_692));
wire output_14_692, output_14_5, output_13_692;
mixer gate_output_13_692(.a(output_14_692), .b(output_14_5), .y(output_13_692));
wire output_15_692, output_15_5, output_14_692;
mixer gate_output_14_692(.a(output_15_692), .b(output_15_5), .y(output_14_692));
wire output_16_692, output_16_5, output_15_692;
mixer gate_output_15_692(.a(output_16_692), .b(output_16_5), .y(output_15_692));
wire output_1_693, output_1_6, output_0_693;
mixer gate_output_0_693(.a(output_1_693), .b(output_1_6), .y(output_0_693));
wire output_2_693, output_2_6, output_1_693;
mixer gate_output_1_693(.a(output_2_693), .b(output_2_6), .y(output_1_693));
wire output_3_693, output_3_6, output_2_693;
mixer gate_output_2_693(.a(output_3_693), .b(output_3_6), .y(output_2_693));
wire output_4_693, output_4_6, output_3_693;
mixer gate_output_3_693(.a(output_4_693), .b(output_4_6), .y(output_3_693));
wire output_5_693, output_5_6, output_4_693;
mixer gate_output_4_693(.a(output_5_693), .b(output_5_6), .y(output_4_693));
wire output_6_693, output_6_6, output_5_693;
mixer gate_output_5_693(.a(output_6_693), .b(output_6_6), .y(output_5_693));
wire output_7_693, output_7_6, output_6_693;
mixer gate_output_6_693(.a(output_7_693), .b(output_7_6), .y(output_6_693));
wire output_8_693, output_8_6, output_7_693;
mixer gate_output_7_693(.a(output_8_693), .b(output_8_6), .y(output_7_693));
wire output_9_693, output_9_6, output_8_693;
mixer gate_output_8_693(.a(output_9_693), .b(output_9_6), .y(output_8_693));
wire output_10_693, output_10_6, output_9_693;
mixer gate_output_9_693(.a(output_10_693), .b(output_10_6), .y(output_9_693));
wire output_11_693, output_11_6, output_10_693;
mixer gate_output_10_693(.a(output_11_693), .b(output_11_6), .y(output_10_693));
wire output_12_693, output_12_6, output_11_693;
mixer gate_output_11_693(.a(output_12_693), .b(output_12_6), .y(output_11_693));
wire output_13_693, output_13_6, output_12_693;
mixer gate_output_12_693(.a(output_13_693), .b(output_13_6), .y(output_12_693));
wire output_14_693, output_14_6, output_13_693;
mixer gate_output_13_693(.a(output_14_693), .b(output_14_6), .y(output_13_693));
wire output_15_693, output_15_6, output_14_693;
mixer gate_output_14_693(.a(output_15_693), .b(output_15_6), .y(output_14_693));
wire output_16_693, output_16_6, output_15_693;
mixer gate_output_15_693(.a(output_16_693), .b(output_16_6), .y(output_15_693));
wire output_1_694, output_1_7, output_0_694;
mixer gate_output_0_694(.a(output_1_694), .b(output_1_7), .y(output_0_694));
wire output_2_694, output_2_7, output_1_694;
mixer gate_output_1_694(.a(output_2_694), .b(output_2_7), .y(output_1_694));
wire output_3_694, output_3_7, output_2_694;
mixer gate_output_2_694(.a(output_3_694), .b(output_3_7), .y(output_2_694));
wire output_4_694, output_4_7, output_3_694;
mixer gate_output_3_694(.a(output_4_694), .b(output_4_7), .y(output_3_694));
wire output_5_694, output_5_7, output_4_694;
mixer gate_output_4_694(.a(output_5_694), .b(output_5_7), .y(output_4_694));
wire output_6_694, output_6_7, output_5_694;
mixer gate_output_5_694(.a(output_6_694), .b(output_6_7), .y(output_5_694));
wire output_7_694, output_7_7, output_6_694;
mixer gate_output_6_694(.a(output_7_694), .b(output_7_7), .y(output_6_694));
wire output_8_694, output_8_7, output_7_694;
mixer gate_output_7_694(.a(output_8_694), .b(output_8_7), .y(output_7_694));
wire output_9_694, output_9_7, output_8_694;
mixer gate_output_8_694(.a(output_9_694), .b(output_9_7), .y(output_8_694));
wire output_10_694, output_10_7, output_9_694;
mixer gate_output_9_694(.a(output_10_694), .b(output_10_7), .y(output_9_694));
wire output_11_694, output_11_7, output_10_694;
mixer gate_output_10_694(.a(output_11_694), .b(output_11_7), .y(output_10_694));
wire output_12_694, output_12_7, output_11_694;
mixer gate_output_11_694(.a(output_12_694), .b(output_12_7), .y(output_11_694));
wire output_13_694, output_13_7, output_12_694;
mixer gate_output_12_694(.a(output_13_694), .b(output_13_7), .y(output_12_694));
wire output_14_694, output_14_7, output_13_694;
mixer gate_output_13_694(.a(output_14_694), .b(output_14_7), .y(output_13_694));
wire output_15_694, output_15_7, output_14_694;
mixer gate_output_14_694(.a(output_15_694), .b(output_15_7), .y(output_14_694));
wire output_16_694, output_16_7, output_15_694;
mixer gate_output_15_694(.a(output_16_694), .b(output_16_7), .y(output_15_694));
wire output_1_695, output_1_8, output_0_695;
mixer gate_output_0_695(.a(output_1_695), .b(output_1_8), .y(output_0_695));
wire output_2_695, output_2_8, output_1_695;
mixer gate_output_1_695(.a(output_2_695), .b(output_2_8), .y(output_1_695));
wire output_3_695, output_3_8, output_2_695;
mixer gate_output_2_695(.a(output_3_695), .b(output_3_8), .y(output_2_695));
wire output_4_695, output_4_8, output_3_695;
mixer gate_output_3_695(.a(output_4_695), .b(output_4_8), .y(output_3_695));
wire output_5_695, output_5_8, output_4_695;
mixer gate_output_4_695(.a(output_5_695), .b(output_5_8), .y(output_4_695));
wire output_6_695, output_6_8, output_5_695;
mixer gate_output_5_695(.a(output_6_695), .b(output_6_8), .y(output_5_695));
wire output_7_695, output_7_8, output_6_695;
mixer gate_output_6_695(.a(output_7_695), .b(output_7_8), .y(output_6_695));
wire output_8_695, output_8_8, output_7_695;
mixer gate_output_7_695(.a(output_8_695), .b(output_8_8), .y(output_7_695));
wire output_9_695, output_9_8, output_8_695;
mixer gate_output_8_695(.a(output_9_695), .b(output_9_8), .y(output_8_695));
wire output_10_695, output_10_8, output_9_695;
mixer gate_output_9_695(.a(output_10_695), .b(output_10_8), .y(output_9_695));
wire output_11_695, output_11_8, output_10_695;
mixer gate_output_10_695(.a(output_11_695), .b(output_11_8), .y(output_10_695));
wire output_12_695, output_12_8, output_11_695;
mixer gate_output_11_695(.a(output_12_695), .b(output_12_8), .y(output_11_695));
wire output_13_695, output_13_8, output_12_695;
mixer gate_output_12_695(.a(output_13_695), .b(output_13_8), .y(output_12_695));
wire output_14_695, output_14_8, output_13_695;
mixer gate_output_13_695(.a(output_14_695), .b(output_14_8), .y(output_13_695));
wire output_15_695, output_15_8, output_14_695;
mixer gate_output_14_695(.a(output_15_695), .b(output_15_8), .y(output_14_695));
wire output_16_695, output_16_8, output_15_695;
mixer gate_output_15_695(.a(output_16_695), .b(output_16_8), .y(output_15_695));
wire output_1_696, output_1_9, output_0_696;
mixer gate_output_0_696(.a(output_1_696), .b(output_1_9), .y(output_0_696));
wire output_2_696, output_2_9, output_1_696;
mixer gate_output_1_696(.a(output_2_696), .b(output_2_9), .y(output_1_696));
wire output_3_696, output_3_9, output_2_696;
mixer gate_output_2_696(.a(output_3_696), .b(output_3_9), .y(output_2_696));
wire output_4_696, output_4_9, output_3_696;
mixer gate_output_3_696(.a(output_4_696), .b(output_4_9), .y(output_3_696));
wire output_5_696, output_5_9, output_4_696;
mixer gate_output_4_696(.a(output_5_696), .b(output_5_9), .y(output_4_696));
wire output_6_696, output_6_9, output_5_696;
mixer gate_output_5_696(.a(output_6_696), .b(output_6_9), .y(output_5_696));
wire output_7_696, output_7_9, output_6_696;
mixer gate_output_6_696(.a(output_7_696), .b(output_7_9), .y(output_6_696));
wire output_8_696, output_8_9, output_7_696;
mixer gate_output_7_696(.a(output_8_696), .b(output_8_9), .y(output_7_696));
wire output_9_696, output_9_9, output_8_696;
mixer gate_output_8_696(.a(output_9_696), .b(output_9_9), .y(output_8_696));
wire output_10_696, output_10_9, output_9_696;
mixer gate_output_9_696(.a(output_10_696), .b(output_10_9), .y(output_9_696));
wire output_11_696, output_11_9, output_10_696;
mixer gate_output_10_696(.a(output_11_696), .b(output_11_9), .y(output_10_696));
wire output_12_696, output_12_9, output_11_696;
mixer gate_output_11_696(.a(output_12_696), .b(output_12_9), .y(output_11_696));
wire output_13_696, output_13_9, output_12_696;
mixer gate_output_12_696(.a(output_13_696), .b(output_13_9), .y(output_12_696));
wire output_14_696, output_14_9, output_13_696;
mixer gate_output_13_696(.a(output_14_696), .b(output_14_9), .y(output_13_696));
wire output_15_696, output_15_9, output_14_696;
mixer gate_output_14_696(.a(output_15_696), .b(output_15_9), .y(output_14_696));
wire output_16_696, output_16_9, output_15_696;
mixer gate_output_15_696(.a(output_16_696), .b(output_16_9), .y(output_15_696));
wire output_1_697, output_1_10, output_0_697;
mixer gate_output_0_697(.a(output_1_697), .b(output_1_10), .y(output_0_697));
wire output_2_697, output_2_10, output_1_697;
mixer gate_output_1_697(.a(output_2_697), .b(output_2_10), .y(output_1_697));
wire output_3_697, output_3_10, output_2_697;
mixer gate_output_2_697(.a(output_3_697), .b(output_3_10), .y(output_2_697));
wire output_4_697, output_4_10, output_3_697;
mixer gate_output_3_697(.a(output_4_697), .b(output_4_10), .y(output_3_697));
wire output_5_697, output_5_10, output_4_697;
mixer gate_output_4_697(.a(output_5_697), .b(output_5_10), .y(output_4_697));
wire output_6_697, output_6_10, output_5_697;
mixer gate_output_5_697(.a(output_6_697), .b(output_6_10), .y(output_5_697));
wire output_7_697, output_7_10, output_6_697;
mixer gate_output_6_697(.a(output_7_697), .b(output_7_10), .y(output_6_697));
wire output_8_697, output_8_10, output_7_697;
mixer gate_output_7_697(.a(output_8_697), .b(output_8_10), .y(output_7_697));
wire output_9_697, output_9_10, output_8_697;
mixer gate_output_8_697(.a(output_9_697), .b(output_9_10), .y(output_8_697));
wire output_10_697, output_10_10, output_9_697;
mixer gate_output_9_697(.a(output_10_697), .b(output_10_10), .y(output_9_697));
wire output_11_697, output_11_10, output_10_697;
mixer gate_output_10_697(.a(output_11_697), .b(output_11_10), .y(output_10_697));
wire output_12_697, output_12_10, output_11_697;
mixer gate_output_11_697(.a(output_12_697), .b(output_12_10), .y(output_11_697));
wire output_13_697, output_13_10, output_12_697;
mixer gate_output_12_697(.a(output_13_697), .b(output_13_10), .y(output_12_697));
wire output_14_697, output_14_10, output_13_697;
mixer gate_output_13_697(.a(output_14_697), .b(output_14_10), .y(output_13_697));
wire output_15_697, output_15_10, output_14_697;
mixer gate_output_14_697(.a(output_15_697), .b(output_15_10), .y(output_14_697));
wire output_16_697, output_16_10, output_15_697;
mixer gate_output_15_697(.a(output_16_697), .b(output_16_10), .y(output_15_697));
wire output_1_698, output_1_11, output_0_698;
mixer gate_output_0_698(.a(output_1_698), .b(output_1_11), .y(output_0_698));
wire output_2_698, output_2_11, output_1_698;
mixer gate_output_1_698(.a(output_2_698), .b(output_2_11), .y(output_1_698));
wire output_3_698, output_3_11, output_2_698;
mixer gate_output_2_698(.a(output_3_698), .b(output_3_11), .y(output_2_698));
wire output_4_698, output_4_11, output_3_698;
mixer gate_output_3_698(.a(output_4_698), .b(output_4_11), .y(output_3_698));
wire output_5_698, output_5_11, output_4_698;
mixer gate_output_4_698(.a(output_5_698), .b(output_5_11), .y(output_4_698));
wire output_6_698, output_6_11, output_5_698;
mixer gate_output_5_698(.a(output_6_698), .b(output_6_11), .y(output_5_698));
wire output_7_698, output_7_11, output_6_698;
mixer gate_output_6_698(.a(output_7_698), .b(output_7_11), .y(output_6_698));
wire output_8_698, output_8_11, output_7_698;
mixer gate_output_7_698(.a(output_8_698), .b(output_8_11), .y(output_7_698));
wire output_9_698, output_9_11, output_8_698;
mixer gate_output_8_698(.a(output_9_698), .b(output_9_11), .y(output_8_698));
wire output_10_698, output_10_11, output_9_698;
mixer gate_output_9_698(.a(output_10_698), .b(output_10_11), .y(output_9_698));
wire output_11_698, output_11_11, output_10_698;
mixer gate_output_10_698(.a(output_11_698), .b(output_11_11), .y(output_10_698));
wire output_12_698, output_12_11, output_11_698;
mixer gate_output_11_698(.a(output_12_698), .b(output_12_11), .y(output_11_698));
wire output_13_698, output_13_11, output_12_698;
mixer gate_output_12_698(.a(output_13_698), .b(output_13_11), .y(output_12_698));
wire output_14_698, output_14_11, output_13_698;
mixer gate_output_13_698(.a(output_14_698), .b(output_14_11), .y(output_13_698));
wire output_15_698, output_15_11, output_14_698;
mixer gate_output_14_698(.a(output_15_698), .b(output_15_11), .y(output_14_698));
wire output_16_698, output_16_11, output_15_698;
mixer gate_output_15_698(.a(output_16_698), .b(output_16_11), .y(output_15_698));
wire output_1_699, output_1_12, output_0_699;
mixer gate_output_0_699(.a(output_1_699), .b(output_1_12), .y(output_0_699));
wire output_2_699, output_2_12, output_1_699;
mixer gate_output_1_699(.a(output_2_699), .b(output_2_12), .y(output_1_699));
wire output_3_699, output_3_12, output_2_699;
mixer gate_output_2_699(.a(output_3_699), .b(output_3_12), .y(output_2_699));
wire output_4_699, output_4_12, output_3_699;
mixer gate_output_3_699(.a(output_4_699), .b(output_4_12), .y(output_3_699));
wire output_5_699, output_5_12, output_4_699;
mixer gate_output_4_699(.a(output_5_699), .b(output_5_12), .y(output_4_699));
wire output_6_699, output_6_12, output_5_699;
mixer gate_output_5_699(.a(output_6_699), .b(output_6_12), .y(output_5_699));
wire output_7_699, output_7_12, output_6_699;
mixer gate_output_6_699(.a(output_7_699), .b(output_7_12), .y(output_6_699));
wire output_8_699, output_8_12, output_7_699;
mixer gate_output_7_699(.a(output_8_699), .b(output_8_12), .y(output_7_699));
wire output_9_699, output_9_12, output_8_699;
mixer gate_output_8_699(.a(output_9_699), .b(output_9_12), .y(output_8_699));
wire output_10_699, output_10_12, output_9_699;
mixer gate_output_9_699(.a(output_10_699), .b(output_10_12), .y(output_9_699));
wire output_11_699, output_11_12, output_10_699;
mixer gate_output_10_699(.a(output_11_699), .b(output_11_12), .y(output_10_699));
wire output_12_699, output_12_12, output_11_699;
mixer gate_output_11_699(.a(output_12_699), .b(output_12_12), .y(output_11_699));
wire output_13_699, output_13_12, output_12_699;
mixer gate_output_12_699(.a(output_13_699), .b(output_13_12), .y(output_12_699));
wire output_14_699, output_14_12, output_13_699;
mixer gate_output_13_699(.a(output_14_699), .b(output_14_12), .y(output_13_699));
wire output_15_699, output_15_12, output_14_699;
mixer gate_output_14_699(.a(output_15_699), .b(output_15_12), .y(output_14_699));
wire output_16_699, output_16_12, output_15_699;
mixer gate_output_15_699(.a(output_16_699), .b(output_16_12), .y(output_15_699));
wire output_1_700, output_1_13, output_0_700;
mixer gate_output_0_700(.a(output_1_700), .b(output_1_13), .y(output_0_700));
wire output_2_700, output_2_13, output_1_700;
mixer gate_output_1_700(.a(output_2_700), .b(output_2_13), .y(output_1_700));
wire output_3_700, output_3_13, output_2_700;
mixer gate_output_2_700(.a(output_3_700), .b(output_3_13), .y(output_2_700));
wire output_4_700, output_4_13, output_3_700;
mixer gate_output_3_700(.a(output_4_700), .b(output_4_13), .y(output_3_700));
wire output_5_700, output_5_13, output_4_700;
mixer gate_output_4_700(.a(output_5_700), .b(output_5_13), .y(output_4_700));
wire output_6_700, output_6_13, output_5_700;
mixer gate_output_5_700(.a(output_6_700), .b(output_6_13), .y(output_5_700));
wire output_7_700, output_7_13, output_6_700;
mixer gate_output_6_700(.a(output_7_700), .b(output_7_13), .y(output_6_700));
wire output_8_700, output_8_13, output_7_700;
mixer gate_output_7_700(.a(output_8_700), .b(output_8_13), .y(output_7_700));
wire output_9_700, output_9_13, output_8_700;
mixer gate_output_8_700(.a(output_9_700), .b(output_9_13), .y(output_8_700));
wire output_10_700, output_10_13, output_9_700;
mixer gate_output_9_700(.a(output_10_700), .b(output_10_13), .y(output_9_700));
wire output_11_700, output_11_13, output_10_700;
mixer gate_output_10_700(.a(output_11_700), .b(output_11_13), .y(output_10_700));
wire output_12_700, output_12_13, output_11_700;
mixer gate_output_11_700(.a(output_12_700), .b(output_12_13), .y(output_11_700));
wire output_13_700, output_13_13, output_12_700;
mixer gate_output_12_700(.a(output_13_700), .b(output_13_13), .y(output_12_700));
wire output_14_700, output_14_13, output_13_700;
mixer gate_output_13_700(.a(output_14_700), .b(output_14_13), .y(output_13_700));
wire output_15_700, output_15_13, output_14_700;
mixer gate_output_14_700(.a(output_15_700), .b(output_15_13), .y(output_14_700));
wire output_16_700, output_16_13, output_15_700;
mixer gate_output_15_700(.a(output_16_700), .b(output_16_13), .y(output_15_700));
wire output_1_701, output_1_14, output_0_701;
mixer gate_output_0_701(.a(output_1_701), .b(output_1_14), .y(output_0_701));
wire output_2_701, output_2_14, output_1_701;
mixer gate_output_1_701(.a(output_2_701), .b(output_2_14), .y(output_1_701));
wire output_3_701, output_3_14, output_2_701;
mixer gate_output_2_701(.a(output_3_701), .b(output_3_14), .y(output_2_701));
wire output_4_701, output_4_14, output_3_701;
mixer gate_output_3_701(.a(output_4_701), .b(output_4_14), .y(output_3_701));
wire output_5_701, output_5_14, output_4_701;
mixer gate_output_4_701(.a(output_5_701), .b(output_5_14), .y(output_4_701));
wire output_6_701, output_6_14, output_5_701;
mixer gate_output_5_701(.a(output_6_701), .b(output_6_14), .y(output_5_701));
wire output_7_701, output_7_14, output_6_701;
mixer gate_output_6_701(.a(output_7_701), .b(output_7_14), .y(output_6_701));
wire output_8_701, output_8_14, output_7_701;
mixer gate_output_7_701(.a(output_8_701), .b(output_8_14), .y(output_7_701));
wire output_9_701, output_9_14, output_8_701;
mixer gate_output_8_701(.a(output_9_701), .b(output_9_14), .y(output_8_701));
wire output_10_701, output_10_14, output_9_701;
mixer gate_output_9_701(.a(output_10_701), .b(output_10_14), .y(output_9_701));
wire output_11_701, output_11_14, output_10_701;
mixer gate_output_10_701(.a(output_11_701), .b(output_11_14), .y(output_10_701));
wire output_12_701, output_12_14, output_11_701;
mixer gate_output_11_701(.a(output_12_701), .b(output_12_14), .y(output_11_701));
wire output_13_701, output_13_14, output_12_701;
mixer gate_output_12_701(.a(output_13_701), .b(output_13_14), .y(output_12_701));
wire output_14_701, output_14_14, output_13_701;
mixer gate_output_13_701(.a(output_14_701), .b(output_14_14), .y(output_13_701));
wire output_15_701, output_15_14, output_14_701;
mixer gate_output_14_701(.a(output_15_701), .b(output_15_14), .y(output_14_701));
wire output_16_701, output_16_14, output_15_701;
mixer gate_output_15_701(.a(output_16_701), .b(output_16_14), .y(output_15_701));
wire output_1_702, output_1_15, output_0_702;
mixer gate_output_0_702(.a(output_1_702), .b(output_1_15), .y(output_0_702));
wire output_2_702, output_2_15, output_1_702;
mixer gate_output_1_702(.a(output_2_702), .b(output_2_15), .y(output_1_702));
wire output_3_702, output_3_15, output_2_702;
mixer gate_output_2_702(.a(output_3_702), .b(output_3_15), .y(output_2_702));
wire output_4_702, output_4_15, output_3_702;
mixer gate_output_3_702(.a(output_4_702), .b(output_4_15), .y(output_3_702));
wire output_5_702, output_5_15, output_4_702;
mixer gate_output_4_702(.a(output_5_702), .b(output_5_15), .y(output_4_702));
wire output_6_702, output_6_15, output_5_702;
mixer gate_output_5_702(.a(output_6_702), .b(output_6_15), .y(output_5_702));
wire output_7_702, output_7_15, output_6_702;
mixer gate_output_6_702(.a(output_7_702), .b(output_7_15), .y(output_6_702));
wire output_8_702, output_8_15, output_7_702;
mixer gate_output_7_702(.a(output_8_702), .b(output_8_15), .y(output_7_702));
wire output_9_702, output_9_15, output_8_702;
mixer gate_output_8_702(.a(output_9_702), .b(output_9_15), .y(output_8_702));
wire output_10_702, output_10_15, output_9_702;
mixer gate_output_9_702(.a(output_10_702), .b(output_10_15), .y(output_9_702));
wire output_11_702, output_11_15, output_10_702;
mixer gate_output_10_702(.a(output_11_702), .b(output_11_15), .y(output_10_702));
wire output_12_702, output_12_15, output_11_702;
mixer gate_output_11_702(.a(output_12_702), .b(output_12_15), .y(output_11_702));
wire output_13_702, output_13_15, output_12_702;
mixer gate_output_12_702(.a(output_13_702), .b(output_13_15), .y(output_12_702));
wire output_14_702, output_14_15, output_13_702;
mixer gate_output_13_702(.a(output_14_702), .b(output_14_15), .y(output_13_702));
wire output_15_702, output_15_15, output_14_702;
mixer gate_output_14_702(.a(output_15_702), .b(output_15_15), .y(output_14_702));
wire output_16_702, output_16_15, output_15_702;
mixer gate_output_15_702(.a(output_16_702), .b(output_16_15), .y(output_15_702));
wire output_1_703, output_1_0, output_0_703;
mixer gate_output_0_703(.a(output_1_703), .b(output_1_0), .y(output_0_703));
wire output_2_703, output_2_0, output_1_703;
mixer gate_output_1_703(.a(output_2_703), .b(output_2_0), .y(output_1_703));
wire output_3_703, output_3_0, output_2_703;
mixer gate_output_2_703(.a(output_3_703), .b(output_3_0), .y(output_2_703));
wire output_4_703, output_4_0, output_3_703;
mixer gate_output_3_703(.a(output_4_703), .b(output_4_0), .y(output_3_703));
wire output_5_703, output_5_0, output_4_703;
mixer gate_output_4_703(.a(output_5_703), .b(output_5_0), .y(output_4_703));
wire output_6_703, output_6_0, output_5_703;
mixer gate_output_5_703(.a(output_6_703), .b(output_6_0), .y(output_5_703));
wire output_7_703, output_7_0, output_6_703;
mixer gate_output_6_703(.a(output_7_703), .b(output_7_0), .y(output_6_703));
wire output_8_703, output_8_0, output_7_703;
mixer gate_output_7_703(.a(output_8_703), .b(output_8_0), .y(output_7_703));
wire output_9_703, output_9_0, output_8_703;
mixer gate_output_8_703(.a(output_9_703), .b(output_9_0), .y(output_8_703));
wire output_10_703, output_10_0, output_9_703;
mixer gate_output_9_703(.a(output_10_703), .b(output_10_0), .y(output_9_703));
wire output_11_703, output_11_0, output_10_703;
mixer gate_output_10_703(.a(output_11_703), .b(output_11_0), .y(output_10_703));
wire output_12_703, output_12_0, output_11_703;
mixer gate_output_11_703(.a(output_12_703), .b(output_12_0), .y(output_11_703));
wire output_13_703, output_13_0, output_12_703;
mixer gate_output_12_703(.a(output_13_703), .b(output_13_0), .y(output_12_703));
wire output_14_703, output_14_0, output_13_703;
mixer gate_output_13_703(.a(output_14_703), .b(output_14_0), .y(output_13_703));
wire output_15_703, output_15_0, output_14_703;
mixer gate_output_14_703(.a(output_15_703), .b(output_15_0), .y(output_14_703));
wire output_16_703, output_16_0, output_15_703;
mixer gate_output_15_703(.a(output_16_703), .b(output_16_0), .y(output_15_703));
wire output_1_704, output_1_1, output_0_704;
mixer gate_output_0_704(.a(output_1_704), .b(output_1_1), .y(output_0_704));
wire output_2_704, output_2_1, output_1_704;
mixer gate_output_1_704(.a(output_2_704), .b(output_2_1), .y(output_1_704));
wire output_3_704, output_3_1, output_2_704;
mixer gate_output_2_704(.a(output_3_704), .b(output_3_1), .y(output_2_704));
wire output_4_704, output_4_1, output_3_704;
mixer gate_output_3_704(.a(output_4_704), .b(output_4_1), .y(output_3_704));
wire output_5_704, output_5_1, output_4_704;
mixer gate_output_4_704(.a(output_5_704), .b(output_5_1), .y(output_4_704));
wire output_6_704, output_6_1, output_5_704;
mixer gate_output_5_704(.a(output_6_704), .b(output_6_1), .y(output_5_704));
wire output_7_704, output_7_1, output_6_704;
mixer gate_output_6_704(.a(output_7_704), .b(output_7_1), .y(output_6_704));
wire output_8_704, output_8_1, output_7_704;
mixer gate_output_7_704(.a(output_8_704), .b(output_8_1), .y(output_7_704));
wire output_9_704, output_9_1, output_8_704;
mixer gate_output_8_704(.a(output_9_704), .b(output_9_1), .y(output_8_704));
wire output_10_704, output_10_1, output_9_704;
mixer gate_output_9_704(.a(output_10_704), .b(output_10_1), .y(output_9_704));
wire output_11_704, output_11_1, output_10_704;
mixer gate_output_10_704(.a(output_11_704), .b(output_11_1), .y(output_10_704));
wire output_12_704, output_12_1, output_11_704;
mixer gate_output_11_704(.a(output_12_704), .b(output_12_1), .y(output_11_704));
wire output_13_704, output_13_1, output_12_704;
mixer gate_output_12_704(.a(output_13_704), .b(output_13_1), .y(output_12_704));
wire output_14_704, output_14_1, output_13_704;
mixer gate_output_13_704(.a(output_14_704), .b(output_14_1), .y(output_13_704));
wire output_15_704, output_15_1, output_14_704;
mixer gate_output_14_704(.a(output_15_704), .b(output_15_1), .y(output_14_704));
wire output_16_704, output_16_1, output_15_704;
mixer gate_output_15_704(.a(output_16_704), .b(output_16_1), .y(output_15_704));
wire output_1_705, output_1_2, output_0_705;
mixer gate_output_0_705(.a(output_1_705), .b(output_1_2), .y(output_0_705));
wire output_2_705, output_2_2, output_1_705;
mixer gate_output_1_705(.a(output_2_705), .b(output_2_2), .y(output_1_705));
wire output_3_705, output_3_2, output_2_705;
mixer gate_output_2_705(.a(output_3_705), .b(output_3_2), .y(output_2_705));
wire output_4_705, output_4_2, output_3_705;
mixer gate_output_3_705(.a(output_4_705), .b(output_4_2), .y(output_3_705));
wire output_5_705, output_5_2, output_4_705;
mixer gate_output_4_705(.a(output_5_705), .b(output_5_2), .y(output_4_705));
wire output_6_705, output_6_2, output_5_705;
mixer gate_output_5_705(.a(output_6_705), .b(output_6_2), .y(output_5_705));
wire output_7_705, output_7_2, output_6_705;
mixer gate_output_6_705(.a(output_7_705), .b(output_7_2), .y(output_6_705));
wire output_8_705, output_8_2, output_7_705;
mixer gate_output_7_705(.a(output_8_705), .b(output_8_2), .y(output_7_705));
wire output_9_705, output_9_2, output_8_705;
mixer gate_output_8_705(.a(output_9_705), .b(output_9_2), .y(output_8_705));
wire output_10_705, output_10_2, output_9_705;
mixer gate_output_9_705(.a(output_10_705), .b(output_10_2), .y(output_9_705));
wire output_11_705, output_11_2, output_10_705;
mixer gate_output_10_705(.a(output_11_705), .b(output_11_2), .y(output_10_705));
wire output_12_705, output_12_2, output_11_705;
mixer gate_output_11_705(.a(output_12_705), .b(output_12_2), .y(output_11_705));
wire output_13_705, output_13_2, output_12_705;
mixer gate_output_12_705(.a(output_13_705), .b(output_13_2), .y(output_12_705));
wire output_14_705, output_14_2, output_13_705;
mixer gate_output_13_705(.a(output_14_705), .b(output_14_2), .y(output_13_705));
wire output_15_705, output_15_2, output_14_705;
mixer gate_output_14_705(.a(output_15_705), .b(output_15_2), .y(output_14_705));
wire output_16_705, output_16_2, output_15_705;
mixer gate_output_15_705(.a(output_16_705), .b(output_16_2), .y(output_15_705));
wire output_1_706, output_1_3, output_0_706;
mixer gate_output_0_706(.a(output_1_706), .b(output_1_3), .y(output_0_706));
wire output_2_706, output_2_3, output_1_706;
mixer gate_output_1_706(.a(output_2_706), .b(output_2_3), .y(output_1_706));
wire output_3_706, output_3_3, output_2_706;
mixer gate_output_2_706(.a(output_3_706), .b(output_3_3), .y(output_2_706));
wire output_4_706, output_4_3, output_3_706;
mixer gate_output_3_706(.a(output_4_706), .b(output_4_3), .y(output_3_706));
wire output_5_706, output_5_3, output_4_706;
mixer gate_output_4_706(.a(output_5_706), .b(output_5_3), .y(output_4_706));
wire output_6_706, output_6_3, output_5_706;
mixer gate_output_5_706(.a(output_6_706), .b(output_6_3), .y(output_5_706));
wire output_7_706, output_7_3, output_6_706;
mixer gate_output_6_706(.a(output_7_706), .b(output_7_3), .y(output_6_706));
wire output_8_706, output_8_3, output_7_706;
mixer gate_output_7_706(.a(output_8_706), .b(output_8_3), .y(output_7_706));
wire output_9_706, output_9_3, output_8_706;
mixer gate_output_8_706(.a(output_9_706), .b(output_9_3), .y(output_8_706));
wire output_10_706, output_10_3, output_9_706;
mixer gate_output_9_706(.a(output_10_706), .b(output_10_3), .y(output_9_706));
wire output_11_706, output_11_3, output_10_706;
mixer gate_output_10_706(.a(output_11_706), .b(output_11_3), .y(output_10_706));
wire output_12_706, output_12_3, output_11_706;
mixer gate_output_11_706(.a(output_12_706), .b(output_12_3), .y(output_11_706));
wire output_13_706, output_13_3, output_12_706;
mixer gate_output_12_706(.a(output_13_706), .b(output_13_3), .y(output_12_706));
wire output_14_706, output_14_3, output_13_706;
mixer gate_output_13_706(.a(output_14_706), .b(output_14_3), .y(output_13_706));
wire output_15_706, output_15_3, output_14_706;
mixer gate_output_14_706(.a(output_15_706), .b(output_15_3), .y(output_14_706));
wire output_16_706, output_16_3, output_15_706;
mixer gate_output_15_706(.a(output_16_706), .b(output_16_3), .y(output_15_706));
wire output_1_707, output_1_4, output_0_707;
mixer gate_output_0_707(.a(output_1_707), .b(output_1_4), .y(output_0_707));
wire output_2_707, output_2_4, output_1_707;
mixer gate_output_1_707(.a(output_2_707), .b(output_2_4), .y(output_1_707));
wire output_3_707, output_3_4, output_2_707;
mixer gate_output_2_707(.a(output_3_707), .b(output_3_4), .y(output_2_707));
wire output_4_707, output_4_4, output_3_707;
mixer gate_output_3_707(.a(output_4_707), .b(output_4_4), .y(output_3_707));
wire output_5_707, output_5_4, output_4_707;
mixer gate_output_4_707(.a(output_5_707), .b(output_5_4), .y(output_4_707));
wire output_6_707, output_6_4, output_5_707;
mixer gate_output_5_707(.a(output_6_707), .b(output_6_4), .y(output_5_707));
wire output_7_707, output_7_4, output_6_707;
mixer gate_output_6_707(.a(output_7_707), .b(output_7_4), .y(output_6_707));
wire output_8_707, output_8_4, output_7_707;
mixer gate_output_7_707(.a(output_8_707), .b(output_8_4), .y(output_7_707));
wire output_9_707, output_9_4, output_8_707;
mixer gate_output_8_707(.a(output_9_707), .b(output_9_4), .y(output_8_707));
wire output_10_707, output_10_4, output_9_707;
mixer gate_output_9_707(.a(output_10_707), .b(output_10_4), .y(output_9_707));
wire output_11_707, output_11_4, output_10_707;
mixer gate_output_10_707(.a(output_11_707), .b(output_11_4), .y(output_10_707));
wire output_12_707, output_12_4, output_11_707;
mixer gate_output_11_707(.a(output_12_707), .b(output_12_4), .y(output_11_707));
wire output_13_707, output_13_4, output_12_707;
mixer gate_output_12_707(.a(output_13_707), .b(output_13_4), .y(output_12_707));
wire output_14_707, output_14_4, output_13_707;
mixer gate_output_13_707(.a(output_14_707), .b(output_14_4), .y(output_13_707));
wire output_15_707, output_15_4, output_14_707;
mixer gate_output_14_707(.a(output_15_707), .b(output_15_4), .y(output_14_707));
wire output_16_707, output_16_4, output_15_707;
mixer gate_output_15_707(.a(output_16_707), .b(output_16_4), .y(output_15_707));
wire output_1_708, output_1_5, output_0_708;
mixer gate_output_0_708(.a(output_1_708), .b(output_1_5), .y(output_0_708));
wire output_2_708, output_2_5, output_1_708;
mixer gate_output_1_708(.a(output_2_708), .b(output_2_5), .y(output_1_708));
wire output_3_708, output_3_5, output_2_708;
mixer gate_output_2_708(.a(output_3_708), .b(output_3_5), .y(output_2_708));
wire output_4_708, output_4_5, output_3_708;
mixer gate_output_3_708(.a(output_4_708), .b(output_4_5), .y(output_3_708));
wire output_5_708, output_5_5, output_4_708;
mixer gate_output_4_708(.a(output_5_708), .b(output_5_5), .y(output_4_708));
wire output_6_708, output_6_5, output_5_708;
mixer gate_output_5_708(.a(output_6_708), .b(output_6_5), .y(output_5_708));
wire output_7_708, output_7_5, output_6_708;
mixer gate_output_6_708(.a(output_7_708), .b(output_7_5), .y(output_6_708));
wire output_8_708, output_8_5, output_7_708;
mixer gate_output_7_708(.a(output_8_708), .b(output_8_5), .y(output_7_708));
wire output_9_708, output_9_5, output_8_708;
mixer gate_output_8_708(.a(output_9_708), .b(output_9_5), .y(output_8_708));
wire output_10_708, output_10_5, output_9_708;
mixer gate_output_9_708(.a(output_10_708), .b(output_10_5), .y(output_9_708));
wire output_11_708, output_11_5, output_10_708;
mixer gate_output_10_708(.a(output_11_708), .b(output_11_5), .y(output_10_708));
wire output_12_708, output_12_5, output_11_708;
mixer gate_output_11_708(.a(output_12_708), .b(output_12_5), .y(output_11_708));
wire output_13_708, output_13_5, output_12_708;
mixer gate_output_12_708(.a(output_13_708), .b(output_13_5), .y(output_12_708));
wire output_14_708, output_14_5, output_13_708;
mixer gate_output_13_708(.a(output_14_708), .b(output_14_5), .y(output_13_708));
wire output_15_708, output_15_5, output_14_708;
mixer gate_output_14_708(.a(output_15_708), .b(output_15_5), .y(output_14_708));
wire output_16_708, output_16_5, output_15_708;
mixer gate_output_15_708(.a(output_16_708), .b(output_16_5), .y(output_15_708));
wire output_1_709, output_1_6, output_0_709;
mixer gate_output_0_709(.a(output_1_709), .b(output_1_6), .y(output_0_709));
wire output_2_709, output_2_6, output_1_709;
mixer gate_output_1_709(.a(output_2_709), .b(output_2_6), .y(output_1_709));
wire output_3_709, output_3_6, output_2_709;
mixer gate_output_2_709(.a(output_3_709), .b(output_3_6), .y(output_2_709));
wire output_4_709, output_4_6, output_3_709;
mixer gate_output_3_709(.a(output_4_709), .b(output_4_6), .y(output_3_709));
wire output_5_709, output_5_6, output_4_709;
mixer gate_output_4_709(.a(output_5_709), .b(output_5_6), .y(output_4_709));
wire output_6_709, output_6_6, output_5_709;
mixer gate_output_5_709(.a(output_6_709), .b(output_6_6), .y(output_5_709));
wire output_7_709, output_7_6, output_6_709;
mixer gate_output_6_709(.a(output_7_709), .b(output_7_6), .y(output_6_709));
wire output_8_709, output_8_6, output_7_709;
mixer gate_output_7_709(.a(output_8_709), .b(output_8_6), .y(output_7_709));
wire output_9_709, output_9_6, output_8_709;
mixer gate_output_8_709(.a(output_9_709), .b(output_9_6), .y(output_8_709));
wire output_10_709, output_10_6, output_9_709;
mixer gate_output_9_709(.a(output_10_709), .b(output_10_6), .y(output_9_709));
wire output_11_709, output_11_6, output_10_709;
mixer gate_output_10_709(.a(output_11_709), .b(output_11_6), .y(output_10_709));
wire output_12_709, output_12_6, output_11_709;
mixer gate_output_11_709(.a(output_12_709), .b(output_12_6), .y(output_11_709));
wire output_13_709, output_13_6, output_12_709;
mixer gate_output_12_709(.a(output_13_709), .b(output_13_6), .y(output_12_709));
wire output_14_709, output_14_6, output_13_709;
mixer gate_output_13_709(.a(output_14_709), .b(output_14_6), .y(output_13_709));
wire output_15_709, output_15_6, output_14_709;
mixer gate_output_14_709(.a(output_15_709), .b(output_15_6), .y(output_14_709));
wire output_16_709, output_16_6, output_15_709;
mixer gate_output_15_709(.a(output_16_709), .b(output_16_6), .y(output_15_709));
wire output_1_710, output_1_7, output_0_710;
mixer gate_output_0_710(.a(output_1_710), .b(output_1_7), .y(output_0_710));
wire output_2_710, output_2_7, output_1_710;
mixer gate_output_1_710(.a(output_2_710), .b(output_2_7), .y(output_1_710));
wire output_3_710, output_3_7, output_2_710;
mixer gate_output_2_710(.a(output_3_710), .b(output_3_7), .y(output_2_710));
wire output_4_710, output_4_7, output_3_710;
mixer gate_output_3_710(.a(output_4_710), .b(output_4_7), .y(output_3_710));
wire output_5_710, output_5_7, output_4_710;
mixer gate_output_4_710(.a(output_5_710), .b(output_5_7), .y(output_4_710));
wire output_6_710, output_6_7, output_5_710;
mixer gate_output_5_710(.a(output_6_710), .b(output_6_7), .y(output_5_710));
wire output_7_710, output_7_7, output_6_710;
mixer gate_output_6_710(.a(output_7_710), .b(output_7_7), .y(output_6_710));
wire output_8_710, output_8_7, output_7_710;
mixer gate_output_7_710(.a(output_8_710), .b(output_8_7), .y(output_7_710));
wire output_9_710, output_9_7, output_8_710;
mixer gate_output_8_710(.a(output_9_710), .b(output_9_7), .y(output_8_710));
wire output_10_710, output_10_7, output_9_710;
mixer gate_output_9_710(.a(output_10_710), .b(output_10_7), .y(output_9_710));
wire output_11_710, output_11_7, output_10_710;
mixer gate_output_10_710(.a(output_11_710), .b(output_11_7), .y(output_10_710));
wire output_12_710, output_12_7, output_11_710;
mixer gate_output_11_710(.a(output_12_710), .b(output_12_7), .y(output_11_710));
wire output_13_710, output_13_7, output_12_710;
mixer gate_output_12_710(.a(output_13_710), .b(output_13_7), .y(output_12_710));
wire output_14_710, output_14_7, output_13_710;
mixer gate_output_13_710(.a(output_14_710), .b(output_14_7), .y(output_13_710));
wire output_15_710, output_15_7, output_14_710;
mixer gate_output_14_710(.a(output_15_710), .b(output_15_7), .y(output_14_710));
wire output_16_710, output_16_7, output_15_710;
mixer gate_output_15_710(.a(output_16_710), .b(output_16_7), .y(output_15_710));
wire output_1_711, output_1_8, output_0_711;
mixer gate_output_0_711(.a(output_1_711), .b(output_1_8), .y(output_0_711));
wire output_2_711, output_2_8, output_1_711;
mixer gate_output_1_711(.a(output_2_711), .b(output_2_8), .y(output_1_711));
wire output_3_711, output_3_8, output_2_711;
mixer gate_output_2_711(.a(output_3_711), .b(output_3_8), .y(output_2_711));
wire output_4_711, output_4_8, output_3_711;
mixer gate_output_3_711(.a(output_4_711), .b(output_4_8), .y(output_3_711));
wire output_5_711, output_5_8, output_4_711;
mixer gate_output_4_711(.a(output_5_711), .b(output_5_8), .y(output_4_711));
wire output_6_711, output_6_8, output_5_711;
mixer gate_output_5_711(.a(output_6_711), .b(output_6_8), .y(output_5_711));
wire output_7_711, output_7_8, output_6_711;
mixer gate_output_6_711(.a(output_7_711), .b(output_7_8), .y(output_6_711));
wire output_8_711, output_8_8, output_7_711;
mixer gate_output_7_711(.a(output_8_711), .b(output_8_8), .y(output_7_711));
wire output_9_711, output_9_8, output_8_711;
mixer gate_output_8_711(.a(output_9_711), .b(output_9_8), .y(output_8_711));
wire output_10_711, output_10_8, output_9_711;
mixer gate_output_9_711(.a(output_10_711), .b(output_10_8), .y(output_9_711));
wire output_11_711, output_11_8, output_10_711;
mixer gate_output_10_711(.a(output_11_711), .b(output_11_8), .y(output_10_711));
wire output_12_711, output_12_8, output_11_711;
mixer gate_output_11_711(.a(output_12_711), .b(output_12_8), .y(output_11_711));
wire output_13_711, output_13_8, output_12_711;
mixer gate_output_12_711(.a(output_13_711), .b(output_13_8), .y(output_12_711));
wire output_14_711, output_14_8, output_13_711;
mixer gate_output_13_711(.a(output_14_711), .b(output_14_8), .y(output_13_711));
wire output_15_711, output_15_8, output_14_711;
mixer gate_output_14_711(.a(output_15_711), .b(output_15_8), .y(output_14_711));
wire output_16_711, output_16_8, output_15_711;
mixer gate_output_15_711(.a(output_16_711), .b(output_16_8), .y(output_15_711));
wire output_1_712, output_1_9, output_0_712;
mixer gate_output_0_712(.a(output_1_712), .b(output_1_9), .y(output_0_712));
wire output_2_712, output_2_9, output_1_712;
mixer gate_output_1_712(.a(output_2_712), .b(output_2_9), .y(output_1_712));
wire output_3_712, output_3_9, output_2_712;
mixer gate_output_2_712(.a(output_3_712), .b(output_3_9), .y(output_2_712));
wire output_4_712, output_4_9, output_3_712;
mixer gate_output_3_712(.a(output_4_712), .b(output_4_9), .y(output_3_712));
wire output_5_712, output_5_9, output_4_712;
mixer gate_output_4_712(.a(output_5_712), .b(output_5_9), .y(output_4_712));
wire output_6_712, output_6_9, output_5_712;
mixer gate_output_5_712(.a(output_6_712), .b(output_6_9), .y(output_5_712));
wire output_7_712, output_7_9, output_6_712;
mixer gate_output_6_712(.a(output_7_712), .b(output_7_9), .y(output_6_712));
wire output_8_712, output_8_9, output_7_712;
mixer gate_output_7_712(.a(output_8_712), .b(output_8_9), .y(output_7_712));
wire output_9_712, output_9_9, output_8_712;
mixer gate_output_8_712(.a(output_9_712), .b(output_9_9), .y(output_8_712));
wire output_10_712, output_10_9, output_9_712;
mixer gate_output_9_712(.a(output_10_712), .b(output_10_9), .y(output_9_712));
wire output_11_712, output_11_9, output_10_712;
mixer gate_output_10_712(.a(output_11_712), .b(output_11_9), .y(output_10_712));
wire output_12_712, output_12_9, output_11_712;
mixer gate_output_11_712(.a(output_12_712), .b(output_12_9), .y(output_11_712));
wire output_13_712, output_13_9, output_12_712;
mixer gate_output_12_712(.a(output_13_712), .b(output_13_9), .y(output_12_712));
wire output_14_712, output_14_9, output_13_712;
mixer gate_output_13_712(.a(output_14_712), .b(output_14_9), .y(output_13_712));
wire output_15_712, output_15_9, output_14_712;
mixer gate_output_14_712(.a(output_15_712), .b(output_15_9), .y(output_14_712));
wire output_16_712, output_16_9, output_15_712;
mixer gate_output_15_712(.a(output_16_712), .b(output_16_9), .y(output_15_712));
wire output_1_713, output_1_10, output_0_713;
mixer gate_output_0_713(.a(output_1_713), .b(output_1_10), .y(output_0_713));
wire output_2_713, output_2_10, output_1_713;
mixer gate_output_1_713(.a(output_2_713), .b(output_2_10), .y(output_1_713));
wire output_3_713, output_3_10, output_2_713;
mixer gate_output_2_713(.a(output_3_713), .b(output_3_10), .y(output_2_713));
wire output_4_713, output_4_10, output_3_713;
mixer gate_output_3_713(.a(output_4_713), .b(output_4_10), .y(output_3_713));
wire output_5_713, output_5_10, output_4_713;
mixer gate_output_4_713(.a(output_5_713), .b(output_5_10), .y(output_4_713));
wire output_6_713, output_6_10, output_5_713;
mixer gate_output_5_713(.a(output_6_713), .b(output_6_10), .y(output_5_713));
wire output_7_713, output_7_10, output_6_713;
mixer gate_output_6_713(.a(output_7_713), .b(output_7_10), .y(output_6_713));
wire output_8_713, output_8_10, output_7_713;
mixer gate_output_7_713(.a(output_8_713), .b(output_8_10), .y(output_7_713));
wire output_9_713, output_9_10, output_8_713;
mixer gate_output_8_713(.a(output_9_713), .b(output_9_10), .y(output_8_713));
wire output_10_713, output_10_10, output_9_713;
mixer gate_output_9_713(.a(output_10_713), .b(output_10_10), .y(output_9_713));
wire output_11_713, output_11_10, output_10_713;
mixer gate_output_10_713(.a(output_11_713), .b(output_11_10), .y(output_10_713));
wire output_12_713, output_12_10, output_11_713;
mixer gate_output_11_713(.a(output_12_713), .b(output_12_10), .y(output_11_713));
wire output_13_713, output_13_10, output_12_713;
mixer gate_output_12_713(.a(output_13_713), .b(output_13_10), .y(output_12_713));
wire output_14_713, output_14_10, output_13_713;
mixer gate_output_13_713(.a(output_14_713), .b(output_14_10), .y(output_13_713));
wire output_15_713, output_15_10, output_14_713;
mixer gate_output_14_713(.a(output_15_713), .b(output_15_10), .y(output_14_713));
wire output_16_713, output_16_10, output_15_713;
mixer gate_output_15_713(.a(output_16_713), .b(output_16_10), .y(output_15_713));
wire output_1_714, output_1_11, output_0_714;
mixer gate_output_0_714(.a(output_1_714), .b(output_1_11), .y(output_0_714));
wire output_2_714, output_2_11, output_1_714;
mixer gate_output_1_714(.a(output_2_714), .b(output_2_11), .y(output_1_714));
wire output_3_714, output_3_11, output_2_714;
mixer gate_output_2_714(.a(output_3_714), .b(output_3_11), .y(output_2_714));
wire output_4_714, output_4_11, output_3_714;
mixer gate_output_3_714(.a(output_4_714), .b(output_4_11), .y(output_3_714));
wire output_5_714, output_5_11, output_4_714;
mixer gate_output_4_714(.a(output_5_714), .b(output_5_11), .y(output_4_714));
wire output_6_714, output_6_11, output_5_714;
mixer gate_output_5_714(.a(output_6_714), .b(output_6_11), .y(output_5_714));
wire output_7_714, output_7_11, output_6_714;
mixer gate_output_6_714(.a(output_7_714), .b(output_7_11), .y(output_6_714));
wire output_8_714, output_8_11, output_7_714;
mixer gate_output_7_714(.a(output_8_714), .b(output_8_11), .y(output_7_714));
wire output_9_714, output_9_11, output_8_714;
mixer gate_output_8_714(.a(output_9_714), .b(output_9_11), .y(output_8_714));
wire output_10_714, output_10_11, output_9_714;
mixer gate_output_9_714(.a(output_10_714), .b(output_10_11), .y(output_9_714));
wire output_11_714, output_11_11, output_10_714;
mixer gate_output_10_714(.a(output_11_714), .b(output_11_11), .y(output_10_714));
wire output_12_714, output_12_11, output_11_714;
mixer gate_output_11_714(.a(output_12_714), .b(output_12_11), .y(output_11_714));
wire output_13_714, output_13_11, output_12_714;
mixer gate_output_12_714(.a(output_13_714), .b(output_13_11), .y(output_12_714));
wire output_14_714, output_14_11, output_13_714;
mixer gate_output_13_714(.a(output_14_714), .b(output_14_11), .y(output_13_714));
wire output_15_714, output_15_11, output_14_714;
mixer gate_output_14_714(.a(output_15_714), .b(output_15_11), .y(output_14_714));
wire output_16_714, output_16_11, output_15_714;
mixer gate_output_15_714(.a(output_16_714), .b(output_16_11), .y(output_15_714));
wire output_1_715, output_1_12, output_0_715;
mixer gate_output_0_715(.a(output_1_715), .b(output_1_12), .y(output_0_715));
wire output_2_715, output_2_12, output_1_715;
mixer gate_output_1_715(.a(output_2_715), .b(output_2_12), .y(output_1_715));
wire output_3_715, output_3_12, output_2_715;
mixer gate_output_2_715(.a(output_3_715), .b(output_3_12), .y(output_2_715));
wire output_4_715, output_4_12, output_3_715;
mixer gate_output_3_715(.a(output_4_715), .b(output_4_12), .y(output_3_715));
wire output_5_715, output_5_12, output_4_715;
mixer gate_output_4_715(.a(output_5_715), .b(output_5_12), .y(output_4_715));
wire output_6_715, output_6_12, output_5_715;
mixer gate_output_5_715(.a(output_6_715), .b(output_6_12), .y(output_5_715));
wire output_7_715, output_7_12, output_6_715;
mixer gate_output_6_715(.a(output_7_715), .b(output_7_12), .y(output_6_715));
wire output_8_715, output_8_12, output_7_715;
mixer gate_output_7_715(.a(output_8_715), .b(output_8_12), .y(output_7_715));
wire output_9_715, output_9_12, output_8_715;
mixer gate_output_8_715(.a(output_9_715), .b(output_9_12), .y(output_8_715));
wire output_10_715, output_10_12, output_9_715;
mixer gate_output_9_715(.a(output_10_715), .b(output_10_12), .y(output_9_715));
wire output_11_715, output_11_12, output_10_715;
mixer gate_output_10_715(.a(output_11_715), .b(output_11_12), .y(output_10_715));
wire output_12_715, output_12_12, output_11_715;
mixer gate_output_11_715(.a(output_12_715), .b(output_12_12), .y(output_11_715));
wire output_13_715, output_13_12, output_12_715;
mixer gate_output_12_715(.a(output_13_715), .b(output_13_12), .y(output_12_715));
wire output_14_715, output_14_12, output_13_715;
mixer gate_output_13_715(.a(output_14_715), .b(output_14_12), .y(output_13_715));
wire output_15_715, output_15_12, output_14_715;
mixer gate_output_14_715(.a(output_15_715), .b(output_15_12), .y(output_14_715));
wire output_16_715, output_16_12, output_15_715;
mixer gate_output_15_715(.a(output_16_715), .b(output_16_12), .y(output_15_715));
wire output_1_716, output_1_13, output_0_716;
mixer gate_output_0_716(.a(output_1_716), .b(output_1_13), .y(output_0_716));
wire output_2_716, output_2_13, output_1_716;
mixer gate_output_1_716(.a(output_2_716), .b(output_2_13), .y(output_1_716));
wire output_3_716, output_3_13, output_2_716;
mixer gate_output_2_716(.a(output_3_716), .b(output_3_13), .y(output_2_716));
wire output_4_716, output_4_13, output_3_716;
mixer gate_output_3_716(.a(output_4_716), .b(output_4_13), .y(output_3_716));
wire output_5_716, output_5_13, output_4_716;
mixer gate_output_4_716(.a(output_5_716), .b(output_5_13), .y(output_4_716));
wire output_6_716, output_6_13, output_5_716;
mixer gate_output_5_716(.a(output_6_716), .b(output_6_13), .y(output_5_716));
wire output_7_716, output_7_13, output_6_716;
mixer gate_output_6_716(.a(output_7_716), .b(output_7_13), .y(output_6_716));
wire output_8_716, output_8_13, output_7_716;
mixer gate_output_7_716(.a(output_8_716), .b(output_8_13), .y(output_7_716));
wire output_9_716, output_9_13, output_8_716;
mixer gate_output_8_716(.a(output_9_716), .b(output_9_13), .y(output_8_716));
wire output_10_716, output_10_13, output_9_716;
mixer gate_output_9_716(.a(output_10_716), .b(output_10_13), .y(output_9_716));
wire output_11_716, output_11_13, output_10_716;
mixer gate_output_10_716(.a(output_11_716), .b(output_11_13), .y(output_10_716));
wire output_12_716, output_12_13, output_11_716;
mixer gate_output_11_716(.a(output_12_716), .b(output_12_13), .y(output_11_716));
wire output_13_716, output_13_13, output_12_716;
mixer gate_output_12_716(.a(output_13_716), .b(output_13_13), .y(output_12_716));
wire output_14_716, output_14_13, output_13_716;
mixer gate_output_13_716(.a(output_14_716), .b(output_14_13), .y(output_13_716));
wire output_15_716, output_15_13, output_14_716;
mixer gate_output_14_716(.a(output_15_716), .b(output_15_13), .y(output_14_716));
wire output_16_716, output_16_13, output_15_716;
mixer gate_output_15_716(.a(output_16_716), .b(output_16_13), .y(output_15_716));
wire output_1_717, output_1_14, output_0_717;
mixer gate_output_0_717(.a(output_1_717), .b(output_1_14), .y(output_0_717));
wire output_2_717, output_2_14, output_1_717;
mixer gate_output_1_717(.a(output_2_717), .b(output_2_14), .y(output_1_717));
wire output_3_717, output_3_14, output_2_717;
mixer gate_output_2_717(.a(output_3_717), .b(output_3_14), .y(output_2_717));
wire output_4_717, output_4_14, output_3_717;
mixer gate_output_3_717(.a(output_4_717), .b(output_4_14), .y(output_3_717));
wire output_5_717, output_5_14, output_4_717;
mixer gate_output_4_717(.a(output_5_717), .b(output_5_14), .y(output_4_717));
wire output_6_717, output_6_14, output_5_717;
mixer gate_output_5_717(.a(output_6_717), .b(output_6_14), .y(output_5_717));
wire output_7_717, output_7_14, output_6_717;
mixer gate_output_6_717(.a(output_7_717), .b(output_7_14), .y(output_6_717));
wire output_8_717, output_8_14, output_7_717;
mixer gate_output_7_717(.a(output_8_717), .b(output_8_14), .y(output_7_717));
wire output_9_717, output_9_14, output_8_717;
mixer gate_output_8_717(.a(output_9_717), .b(output_9_14), .y(output_8_717));
wire output_10_717, output_10_14, output_9_717;
mixer gate_output_9_717(.a(output_10_717), .b(output_10_14), .y(output_9_717));
wire output_11_717, output_11_14, output_10_717;
mixer gate_output_10_717(.a(output_11_717), .b(output_11_14), .y(output_10_717));
wire output_12_717, output_12_14, output_11_717;
mixer gate_output_11_717(.a(output_12_717), .b(output_12_14), .y(output_11_717));
wire output_13_717, output_13_14, output_12_717;
mixer gate_output_12_717(.a(output_13_717), .b(output_13_14), .y(output_12_717));
wire output_14_717, output_14_14, output_13_717;
mixer gate_output_13_717(.a(output_14_717), .b(output_14_14), .y(output_13_717));
wire output_15_717, output_15_14, output_14_717;
mixer gate_output_14_717(.a(output_15_717), .b(output_15_14), .y(output_14_717));
wire output_16_717, output_16_14, output_15_717;
mixer gate_output_15_717(.a(output_16_717), .b(output_16_14), .y(output_15_717));
wire output_1_718, output_1_15, output_0_718;
mixer gate_output_0_718(.a(output_1_718), .b(output_1_15), .y(output_0_718));
wire output_2_718, output_2_15, output_1_718;
mixer gate_output_1_718(.a(output_2_718), .b(output_2_15), .y(output_1_718));
wire output_3_718, output_3_15, output_2_718;
mixer gate_output_2_718(.a(output_3_718), .b(output_3_15), .y(output_2_718));
wire output_4_718, output_4_15, output_3_718;
mixer gate_output_3_718(.a(output_4_718), .b(output_4_15), .y(output_3_718));
wire output_5_718, output_5_15, output_4_718;
mixer gate_output_4_718(.a(output_5_718), .b(output_5_15), .y(output_4_718));
wire output_6_718, output_6_15, output_5_718;
mixer gate_output_5_718(.a(output_6_718), .b(output_6_15), .y(output_5_718));
wire output_7_718, output_7_15, output_6_718;
mixer gate_output_6_718(.a(output_7_718), .b(output_7_15), .y(output_6_718));
wire output_8_718, output_8_15, output_7_718;
mixer gate_output_7_718(.a(output_8_718), .b(output_8_15), .y(output_7_718));
wire output_9_718, output_9_15, output_8_718;
mixer gate_output_8_718(.a(output_9_718), .b(output_9_15), .y(output_8_718));
wire output_10_718, output_10_15, output_9_718;
mixer gate_output_9_718(.a(output_10_718), .b(output_10_15), .y(output_9_718));
wire output_11_718, output_11_15, output_10_718;
mixer gate_output_10_718(.a(output_11_718), .b(output_11_15), .y(output_10_718));
wire output_12_718, output_12_15, output_11_718;
mixer gate_output_11_718(.a(output_12_718), .b(output_12_15), .y(output_11_718));
wire output_13_718, output_13_15, output_12_718;
mixer gate_output_12_718(.a(output_13_718), .b(output_13_15), .y(output_12_718));
wire output_14_718, output_14_15, output_13_718;
mixer gate_output_13_718(.a(output_14_718), .b(output_14_15), .y(output_13_718));
wire output_15_718, output_15_15, output_14_718;
mixer gate_output_14_718(.a(output_15_718), .b(output_15_15), .y(output_14_718));
wire output_16_718, output_16_15, output_15_718;
mixer gate_output_15_718(.a(output_16_718), .b(output_16_15), .y(output_15_718));
wire output_1_719, output_1_0, output_0_719;
mixer gate_output_0_719(.a(output_1_719), .b(output_1_0), .y(output_0_719));
wire output_2_719, output_2_0, output_1_719;
mixer gate_output_1_719(.a(output_2_719), .b(output_2_0), .y(output_1_719));
wire output_3_719, output_3_0, output_2_719;
mixer gate_output_2_719(.a(output_3_719), .b(output_3_0), .y(output_2_719));
wire output_4_719, output_4_0, output_3_719;
mixer gate_output_3_719(.a(output_4_719), .b(output_4_0), .y(output_3_719));
wire output_5_719, output_5_0, output_4_719;
mixer gate_output_4_719(.a(output_5_719), .b(output_5_0), .y(output_4_719));
wire output_6_719, output_6_0, output_5_719;
mixer gate_output_5_719(.a(output_6_719), .b(output_6_0), .y(output_5_719));
wire output_7_719, output_7_0, output_6_719;
mixer gate_output_6_719(.a(output_7_719), .b(output_7_0), .y(output_6_719));
wire output_8_719, output_8_0, output_7_719;
mixer gate_output_7_719(.a(output_8_719), .b(output_8_0), .y(output_7_719));
wire output_9_719, output_9_0, output_8_719;
mixer gate_output_8_719(.a(output_9_719), .b(output_9_0), .y(output_8_719));
wire output_10_719, output_10_0, output_9_719;
mixer gate_output_9_719(.a(output_10_719), .b(output_10_0), .y(output_9_719));
wire output_11_719, output_11_0, output_10_719;
mixer gate_output_10_719(.a(output_11_719), .b(output_11_0), .y(output_10_719));
wire output_12_719, output_12_0, output_11_719;
mixer gate_output_11_719(.a(output_12_719), .b(output_12_0), .y(output_11_719));
wire output_13_719, output_13_0, output_12_719;
mixer gate_output_12_719(.a(output_13_719), .b(output_13_0), .y(output_12_719));
wire output_14_719, output_14_0, output_13_719;
mixer gate_output_13_719(.a(output_14_719), .b(output_14_0), .y(output_13_719));
wire output_15_719, output_15_0, output_14_719;
mixer gate_output_14_719(.a(output_15_719), .b(output_15_0), .y(output_14_719));
wire output_16_719, output_16_0, output_15_719;
mixer gate_output_15_719(.a(output_16_719), .b(output_16_0), .y(output_15_719));
wire output_1_720, output_1_1, output_0_720;
mixer gate_output_0_720(.a(output_1_720), .b(output_1_1), .y(output_0_720));
wire output_2_720, output_2_1, output_1_720;
mixer gate_output_1_720(.a(output_2_720), .b(output_2_1), .y(output_1_720));
wire output_3_720, output_3_1, output_2_720;
mixer gate_output_2_720(.a(output_3_720), .b(output_3_1), .y(output_2_720));
wire output_4_720, output_4_1, output_3_720;
mixer gate_output_3_720(.a(output_4_720), .b(output_4_1), .y(output_3_720));
wire output_5_720, output_5_1, output_4_720;
mixer gate_output_4_720(.a(output_5_720), .b(output_5_1), .y(output_4_720));
wire output_6_720, output_6_1, output_5_720;
mixer gate_output_5_720(.a(output_6_720), .b(output_6_1), .y(output_5_720));
wire output_7_720, output_7_1, output_6_720;
mixer gate_output_6_720(.a(output_7_720), .b(output_7_1), .y(output_6_720));
wire output_8_720, output_8_1, output_7_720;
mixer gate_output_7_720(.a(output_8_720), .b(output_8_1), .y(output_7_720));
wire output_9_720, output_9_1, output_8_720;
mixer gate_output_8_720(.a(output_9_720), .b(output_9_1), .y(output_8_720));
wire output_10_720, output_10_1, output_9_720;
mixer gate_output_9_720(.a(output_10_720), .b(output_10_1), .y(output_9_720));
wire output_11_720, output_11_1, output_10_720;
mixer gate_output_10_720(.a(output_11_720), .b(output_11_1), .y(output_10_720));
wire output_12_720, output_12_1, output_11_720;
mixer gate_output_11_720(.a(output_12_720), .b(output_12_1), .y(output_11_720));
wire output_13_720, output_13_1, output_12_720;
mixer gate_output_12_720(.a(output_13_720), .b(output_13_1), .y(output_12_720));
wire output_14_720, output_14_1, output_13_720;
mixer gate_output_13_720(.a(output_14_720), .b(output_14_1), .y(output_13_720));
wire output_15_720, output_15_1, output_14_720;
mixer gate_output_14_720(.a(output_15_720), .b(output_15_1), .y(output_14_720));
wire output_16_720, output_16_1, output_15_720;
mixer gate_output_15_720(.a(output_16_720), .b(output_16_1), .y(output_15_720));
wire output_1_721, output_1_2, output_0_721;
mixer gate_output_0_721(.a(output_1_721), .b(output_1_2), .y(output_0_721));
wire output_2_721, output_2_2, output_1_721;
mixer gate_output_1_721(.a(output_2_721), .b(output_2_2), .y(output_1_721));
wire output_3_721, output_3_2, output_2_721;
mixer gate_output_2_721(.a(output_3_721), .b(output_3_2), .y(output_2_721));
wire output_4_721, output_4_2, output_3_721;
mixer gate_output_3_721(.a(output_4_721), .b(output_4_2), .y(output_3_721));
wire output_5_721, output_5_2, output_4_721;
mixer gate_output_4_721(.a(output_5_721), .b(output_5_2), .y(output_4_721));
wire output_6_721, output_6_2, output_5_721;
mixer gate_output_5_721(.a(output_6_721), .b(output_6_2), .y(output_5_721));
wire output_7_721, output_7_2, output_6_721;
mixer gate_output_6_721(.a(output_7_721), .b(output_7_2), .y(output_6_721));
wire output_8_721, output_8_2, output_7_721;
mixer gate_output_7_721(.a(output_8_721), .b(output_8_2), .y(output_7_721));
wire output_9_721, output_9_2, output_8_721;
mixer gate_output_8_721(.a(output_9_721), .b(output_9_2), .y(output_8_721));
wire output_10_721, output_10_2, output_9_721;
mixer gate_output_9_721(.a(output_10_721), .b(output_10_2), .y(output_9_721));
wire output_11_721, output_11_2, output_10_721;
mixer gate_output_10_721(.a(output_11_721), .b(output_11_2), .y(output_10_721));
wire output_12_721, output_12_2, output_11_721;
mixer gate_output_11_721(.a(output_12_721), .b(output_12_2), .y(output_11_721));
wire output_13_721, output_13_2, output_12_721;
mixer gate_output_12_721(.a(output_13_721), .b(output_13_2), .y(output_12_721));
wire output_14_721, output_14_2, output_13_721;
mixer gate_output_13_721(.a(output_14_721), .b(output_14_2), .y(output_13_721));
wire output_15_721, output_15_2, output_14_721;
mixer gate_output_14_721(.a(output_15_721), .b(output_15_2), .y(output_14_721));
wire output_16_721, output_16_2, output_15_721;
mixer gate_output_15_721(.a(output_16_721), .b(output_16_2), .y(output_15_721));
wire output_1_722, output_1_3, output_0_722;
mixer gate_output_0_722(.a(output_1_722), .b(output_1_3), .y(output_0_722));
wire output_2_722, output_2_3, output_1_722;
mixer gate_output_1_722(.a(output_2_722), .b(output_2_3), .y(output_1_722));
wire output_3_722, output_3_3, output_2_722;
mixer gate_output_2_722(.a(output_3_722), .b(output_3_3), .y(output_2_722));
wire output_4_722, output_4_3, output_3_722;
mixer gate_output_3_722(.a(output_4_722), .b(output_4_3), .y(output_3_722));
wire output_5_722, output_5_3, output_4_722;
mixer gate_output_4_722(.a(output_5_722), .b(output_5_3), .y(output_4_722));
wire output_6_722, output_6_3, output_5_722;
mixer gate_output_5_722(.a(output_6_722), .b(output_6_3), .y(output_5_722));
wire output_7_722, output_7_3, output_6_722;
mixer gate_output_6_722(.a(output_7_722), .b(output_7_3), .y(output_6_722));
wire output_8_722, output_8_3, output_7_722;
mixer gate_output_7_722(.a(output_8_722), .b(output_8_3), .y(output_7_722));
wire output_9_722, output_9_3, output_8_722;
mixer gate_output_8_722(.a(output_9_722), .b(output_9_3), .y(output_8_722));
wire output_10_722, output_10_3, output_9_722;
mixer gate_output_9_722(.a(output_10_722), .b(output_10_3), .y(output_9_722));
wire output_11_722, output_11_3, output_10_722;
mixer gate_output_10_722(.a(output_11_722), .b(output_11_3), .y(output_10_722));
wire output_12_722, output_12_3, output_11_722;
mixer gate_output_11_722(.a(output_12_722), .b(output_12_3), .y(output_11_722));
wire output_13_722, output_13_3, output_12_722;
mixer gate_output_12_722(.a(output_13_722), .b(output_13_3), .y(output_12_722));
wire output_14_722, output_14_3, output_13_722;
mixer gate_output_13_722(.a(output_14_722), .b(output_14_3), .y(output_13_722));
wire output_15_722, output_15_3, output_14_722;
mixer gate_output_14_722(.a(output_15_722), .b(output_15_3), .y(output_14_722));
wire output_16_722, output_16_3, output_15_722;
mixer gate_output_15_722(.a(output_16_722), .b(output_16_3), .y(output_15_722));
wire output_1_723, output_1_4, output_0_723;
mixer gate_output_0_723(.a(output_1_723), .b(output_1_4), .y(output_0_723));
wire output_2_723, output_2_4, output_1_723;
mixer gate_output_1_723(.a(output_2_723), .b(output_2_4), .y(output_1_723));
wire output_3_723, output_3_4, output_2_723;
mixer gate_output_2_723(.a(output_3_723), .b(output_3_4), .y(output_2_723));
wire output_4_723, output_4_4, output_3_723;
mixer gate_output_3_723(.a(output_4_723), .b(output_4_4), .y(output_3_723));
wire output_5_723, output_5_4, output_4_723;
mixer gate_output_4_723(.a(output_5_723), .b(output_5_4), .y(output_4_723));
wire output_6_723, output_6_4, output_5_723;
mixer gate_output_5_723(.a(output_6_723), .b(output_6_4), .y(output_5_723));
wire output_7_723, output_7_4, output_6_723;
mixer gate_output_6_723(.a(output_7_723), .b(output_7_4), .y(output_6_723));
wire output_8_723, output_8_4, output_7_723;
mixer gate_output_7_723(.a(output_8_723), .b(output_8_4), .y(output_7_723));
wire output_9_723, output_9_4, output_8_723;
mixer gate_output_8_723(.a(output_9_723), .b(output_9_4), .y(output_8_723));
wire output_10_723, output_10_4, output_9_723;
mixer gate_output_9_723(.a(output_10_723), .b(output_10_4), .y(output_9_723));
wire output_11_723, output_11_4, output_10_723;
mixer gate_output_10_723(.a(output_11_723), .b(output_11_4), .y(output_10_723));
wire output_12_723, output_12_4, output_11_723;
mixer gate_output_11_723(.a(output_12_723), .b(output_12_4), .y(output_11_723));
wire output_13_723, output_13_4, output_12_723;
mixer gate_output_12_723(.a(output_13_723), .b(output_13_4), .y(output_12_723));
wire output_14_723, output_14_4, output_13_723;
mixer gate_output_13_723(.a(output_14_723), .b(output_14_4), .y(output_13_723));
wire output_15_723, output_15_4, output_14_723;
mixer gate_output_14_723(.a(output_15_723), .b(output_15_4), .y(output_14_723));
wire output_16_723, output_16_4, output_15_723;
mixer gate_output_15_723(.a(output_16_723), .b(output_16_4), .y(output_15_723));
wire output_1_724, output_1_5, output_0_724;
mixer gate_output_0_724(.a(output_1_724), .b(output_1_5), .y(output_0_724));
wire output_2_724, output_2_5, output_1_724;
mixer gate_output_1_724(.a(output_2_724), .b(output_2_5), .y(output_1_724));
wire output_3_724, output_3_5, output_2_724;
mixer gate_output_2_724(.a(output_3_724), .b(output_3_5), .y(output_2_724));
wire output_4_724, output_4_5, output_3_724;
mixer gate_output_3_724(.a(output_4_724), .b(output_4_5), .y(output_3_724));
wire output_5_724, output_5_5, output_4_724;
mixer gate_output_4_724(.a(output_5_724), .b(output_5_5), .y(output_4_724));
wire output_6_724, output_6_5, output_5_724;
mixer gate_output_5_724(.a(output_6_724), .b(output_6_5), .y(output_5_724));
wire output_7_724, output_7_5, output_6_724;
mixer gate_output_6_724(.a(output_7_724), .b(output_7_5), .y(output_6_724));
wire output_8_724, output_8_5, output_7_724;
mixer gate_output_7_724(.a(output_8_724), .b(output_8_5), .y(output_7_724));
wire output_9_724, output_9_5, output_8_724;
mixer gate_output_8_724(.a(output_9_724), .b(output_9_5), .y(output_8_724));
wire output_10_724, output_10_5, output_9_724;
mixer gate_output_9_724(.a(output_10_724), .b(output_10_5), .y(output_9_724));
wire output_11_724, output_11_5, output_10_724;
mixer gate_output_10_724(.a(output_11_724), .b(output_11_5), .y(output_10_724));
wire output_12_724, output_12_5, output_11_724;
mixer gate_output_11_724(.a(output_12_724), .b(output_12_5), .y(output_11_724));
wire output_13_724, output_13_5, output_12_724;
mixer gate_output_12_724(.a(output_13_724), .b(output_13_5), .y(output_12_724));
wire output_14_724, output_14_5, output_13_724;
mixer gate_output_13_724(.a(output_14_724), .b(output_14_5), .y(output_13_724));
wire output_15_724, output_15_5, output_14_724;
mixer gate_output_14_724(.a(output_15_724), .b(output_15_5), .y(output_14_724));
wire output_16_724, output_16_5, output_15_724;
mixer gate_output_15_724(.a(output_16_724), .b(output_16_5), .y(output_15_724));
wire output_1_725, output_1_6, output_0_725;
mixer gate_output_0_725(.a(output_1_725), .b(output_1_6), .y(output_0_725));
wire output_2_725, output_2_6, output_1_725;
mixer gate_output_1_725(.a(output_2_725), .b(output_2_6), .y(output_1_725));
wire output_3_725, output_3_6, output_2_725;
mixer gate_output_2_725(.a(output_3_725), .b(output_3_6), .y(output_2_725));
wire output_4_725, output_4_6, output_3_725;
mixer gate_output_3_725(.a(output_4_725), .b(output_4_6), .y(output_3_725));
wire output_5_725, output_5_6, output_4_725;
mixer gate_output_4_725(.a(output_5_725), .b(output_5_6), .y(output_4_725));
wire output_6_725, output_6_6, output_5_725;
mixer gate_output_5_725(.a(output_6_725), .b(output_6_6), .y(output_5_725));
wire output_7_725, output_7_6, output_6_725;
mixer gate_output_6_725(.a(output_7_725), .b(output_7_6), .y(output_6_725));
wire output_8_725, output_8_6, output_7_725;
mixer gate_output_7_725(.a(output_8_725), .b(output_8_6), .y(output_7_725));
wire output_9_725, output_9_6, output_8_725;
mixer gate_output_8_725(.a(output_9_725), .b(output_9_6), .y(output_8_725));
wire output_10_725, output_10_6, output_9_725;
mixer gate_output_9_725(.a(output_10_725), .b(output_10_6), .y(output_9_725));
wire output_11_725, output_11_6, output_10_725;
mixer gate_output_10_725(.a(output_11_725), .b(output_11_6), .y(output_10_725));
wire output_12_725, output_12_6, output_11_725;
mixer gate_output_11_725(.a(output_12_725), .b(output_12_6), .y(output_11_725));
wire output_13_725, output_13_6, output_12_725;
mixer gate_output_12_725(.a(output_13_725), .b(output_13_6), .y(output_12_725));
wire output_14_725, output_14_6, output_13_725;
mixer gate_output_13_725(.a(output_14_725), .b(output_14_6), .y(output_13_725));
wire output_15_725, output_15_6, output_14_725;
mixer gate_output_14_725(.a(output_15_725), .b(output_15_6), .y(output_14_725));
wire output_16_725, output_16_6, output_15_725;
mixer gate_output_15_725(.a(output_16_725), .b(output_16_6), .y(output_15_725));
wire output_1_726, output_1_7, output_0_726;
mixer gate_output_0_726(.a(output_1_726), .b(output_1_7), .y(output_0_726));
wire output_2_726, output_2_7, output_1_726;
mixer gate_output_1_726(.a(output_2_726), .b(output_2_7), .y(output_1_726));
wire output_3_726, output_3_7, output_2_726;
mixer gate_output_2_726(.a(output_3_726), .b(output_3_7), .y(output_2_726));
wire output_4_726, output_4_7, output_3_726;
mixer gate_output_3_726(.a(output_4_726), .b(output_4_7), .y(output_3_726));
wire output_5_726, output_5_7, output_4_726;
mixer gate_output_4_726(.a(output_5_726), .b(output_5_7), .y(output_4_726));
wire output_6_726, output_6_7, output_5_726;
mixer gate_output_5_726(.a(output_6_726), .b(output_6_7), .y(output_5_726));
wire output_7_726, output_7_7, output_6_726;
mixer gate_output_6_726(.a(output_7_726), .b(output_7_7), .y(output_6_726));
wire output_8_726, output_8_7, output_7_726;
mixer gate_output_7_726(.a(output_8_726), .b(output_8_7), .y(output_7_726));
wire output_9_726, output_9_7, output_8_726;
mixer gate_output_8_726(.a(output_9_726), .b(output_9_7), .y(output_8_726));
wire output_10_726, output_10_7, output_9_726;
mixer gate_output_9_726(.a(output_10_726), .b(output_10_7), .y(output_9_726));
wire output_11_726, output_11_7, output_10_726;
mixer gate_output_10_726(.a(output_11_726), .b(output_11_7), .y(output_10_726));
wire output_12_726, output_12_7, output_11_726;
mixer gate_output_11_726(.a(output_12_726), .b(output_12_7), .y(output_11_726));
wire output_13_726, output_13_7, output_12_726;
mixer gate_output_12_726(.a(output_13_726), .b(output_13_7), .y(output_12_726));
wire output_14_726, output_14_7, output_13_726;
mixer gate_output_13_726(.a(output_14_726), .b(output_14_7), .y(output_13_726));
wire output_15_726, output_15_7, output_14_726;
mixer gate_output_14_726(.a(output_15_726), .b(output_15_7), .y(output_14_726));
wire output_16_726, output_16_7, output_15_726;
mixer gate_output_15_726(.a(output_16_726), .b(output_16_7), .y(output_15_726));
wire output_1_727, output_1_8, output_0_727;
mixer gate_output_0_727(.a(output_1_727), .b(output_1_8), .y(output_0_727));
wire output_2_727, output_2_8, output_1_727;
mixer gate_output_1_727(.a(output_2_727), .b(output_2_8), .y(output_1_727));
wire output_3_727, output_3_8, output_2_727;
mixer gate_output_2_727(.a(output_3_727), .b(output_3_8), .y(output_2_727));
wire output_4_727, output_4_8, output_3_727;
mixer gate_output_3_727(.a(output_4_727), .b(output_4_8), .y(output_3_727));
wire output_5_727, output_5_8, output_4_727;
mixer gate_output_4_727(.a(output_5_727), .b(output_5_8), .y(output_4_727));
wire output_6_727, output_6_8, output_5_727;
mixer gate_output_5_727(.a(output_6_727), .b(output_6_8), .y(output_5_727));
wire output_7_727, output_7_8, output_6_727;
mixer gate_output_6_727(.a(output_7_727), .b(output_7_8), .y(output_6_727));
wire output_8_727, output_8_8, output_7_727;
mixer gate_output_7_727(.a(output_8_727), .b(output_8_8), .y(output_7_727));
wire output_9_727, output_9_8, output_8_727;
mixer gate_output_8_727(.a(output_9_727), .b(output_9_8), .y(output_8_727));
wire output_10_727, output_10_8, output_9_727;
mixer gate_output_9_727(.a(output_10_727), .b(output_10_8), .y(output_9_727));
wire output_11_727, output_11_8, output_10_727;
mixer gate_output_10_727(.a(output_11_727), .b(output_11_8), .y(output_10_727));
wire output_12_727, output_12_8, output_11_727;
mixer gate_output_11_727(.a(output_12_727), .b(output_12_8), .y(output_11_727));
wire output_13_727, output_13_8, output_12_727;
mixer gate_output_12_727(.a(output_13_727), .b(output_13_8), .y(output_12_727));
wire output_14_727, output_14_8, output_13_727;
mixer gate_output_13_727(.a(output_14_727), .b(output_14_8), .y(output_13_727));
wire output_15_727, output_15_8, output_14_727;
mixer gate_output_14_727(.a(output_15_727), .b(output_15_8), .y(output_14_727));
wire output_16_727, output_16_8, output_15_727;
mixer gate_output_15_727(.a(output_16_727), .b(output_16_8), .y(output_15_727));
wire output_1_728, output_1_9, output_0_728;
mixer gate_output_0_728(.a(output_1_728), .b(output_1_9), .y(output_0_728));
wire output_2_728, output_2_9, output_1_728;
mixer gate_output_1_728(.a(output_2_728), .b(output_2_9), .y(output_1_728));
wire output_3_728, output_3_9, output_2_728;
mixer gate_output_2_728(.a(output_3_728), .b(output_3_9), .y(output_2_728));
wire output_4_728, output_4_9, output_3_728;
mixer gate_output_3_728(.a(output_4_728), .b(output_4_9), .y(output_3_728));
wire output_5_728, output_5_9, output_4_728;
mixer gate_output_4_728(.a(output_5_728), .b(output_5_9), .y(output_4_728));
wire output_6_728, output_6_9, output_5_728;
mixer gate_output_5_728(.a(output_6_728), .b(output_6_9), .y(output_5_728));
wire output_7_728, output_7_9, output_6_728;
mixer gate_output_6_728(.a(output_7_728), .b(output_7_9), .y(output_6_728));
wire output_8_728, output_8_9, output_7_728;
mixer gate_output_7_728(.a(output_8_728), .b(output_8_9), .y(output_7_728));
wire output_9_728, output_9_9, output_8_728;
mixer gate_output_8_728(.a(output_9_728), .b(output_9_9), .y(output_8_728));
wire output_10_728, output_10_9, output_9_728;
mixer gate_output_9_728(.a(output_10_728), .b(output_10_9), .y(output_9_728));
wire output_11_728, output_11_9, output_10_728;
mixer gate_output_10_728(.a(output_11_728), .b(output_11_9), .y(output_10_728));
wire output_12_728, output_12_9, output_11_728;
mixer gate_output_11_728(.a(output_12_728), .b(output_12_9), .y(output_11_728));
wire output_13_728, output_13_9, output_12_728;
mixer gate_output_12_728(.a(output_13_728), .b(output_13_9), .y(output_12_728));
wire output_14_728, output_14_9, output_13_728;
mixer gate_output_13_728(.a(output_14_728), .b(output_14_9), .y(output_13_728));
wire output_15_728, output_15_9, output_14_728;
mixer gate_output_14_728(.a(output_15_728), .b(output_15_9), .y(output_14_728));
wire output_16_728, output_16_9, output_15_728;
mixer gate_output_15_728(.a(output_16_728), .b(output_16_9), .y(output_15_728));
wire output_1_729, output_1_10, output_0_729;
mixer gate_output_0_729(.a(output_1_729), .b(output_1_10), .y(output_0_729));
wire output_2_729, output_2_10, output_1_729;
mixer gate_output_1_729(.a(output_2_729), .b(output_2_10), .y(output_1_729));
wire output_3_729, output_3_10, output_2_729;
mixer gate_output_2_729(.a(output_3_729), .b(output_3_10), .y(output_2_729));
wire output_4_729, output_4_10, output_3_729;
mixer gate_output_3_729(.a(output_4_729), .b(output_4_10), .y(output_3_729));
wire output_5_729, output_5_10, output_4_729;
mixer gate_output_4_729(.a(output_5_729), .b(output_5_10), .y(output_4_729));
wire output_6_729, output_6_10, output_5_729;
mixer gate_output_5_729(.a(output_6_729), .b(output_6_10), .y(output_5_729));
wire output_7_729, output_7_10, output_6_729;
mixer gate_output_6_729(.a(output_7_729), .b(output_7_10), .y(output_6_729));
wire output_8_729, output_8_10, output_7_729;
mixer gate_output_7_729(.a(output_8_729), .b(output_8_10), .y(output_7_729));
wire output_9_729, output_9_10, output_8_729;
mixer gate_output_8_729(.a(output_9_729), .b(output_9_10), .y(output_8_729));
wire output_10_729, output_10_10, output_9_729;
mixer gate_output_9_729(.a(output_10_729), .b(output_10_10), .y(output_9_729));
wire output_11_729, output_11_10, output_10_729;
mixer gate_output_10_729(.a(output_11_729), .b(output_11_10), .y(output_10_729));
wire output_12_729, output_12_10, output_11_729;
mixer gate_output_11_729(.a(output_12_729), .b(output_12_10), .y(output_11_729));
wire output_13_729, output_13_10, output_12_729;
mixer gate_output_12_729(.a(output_13_729), .b(output_13_10), .y(output_12_729));
wire output_14_729, output_14_10, output_13_729;
mixer gate_output_13_729(.a(output_14_729), .b(output_14_10), .y(output_13_729));
wire output_15_729, output_15_10, output_14_729;
mixer gate_output_14_729(.a(output_15_729), .b(output_15_10), .y(output_14_729));
wire output_16_729, output_16_10, output_15_729;
mixer gate_output_15_729(.a(output_16_729), .b(output_16_10), .y(output_15_729));
wire output_1_730, output_1_11, output_0_730;
mixer gate_output_0_730(.a(output_1_730), .b(output_1_11), .y(output_0_730));
wire output_2_730, output_2_11, output_1_730;
mixer gate_output_1_730(.a(output_2_730), .b(output_2_11), .y(output_1_730));
wire output_3_730, output_3_11, output_2_730;
mixer gate_output_2_730(.a(output_3_730), .b(output_3_11), .y(output_2_730));
wire output_4_730, output_4_11, output_3_730;
mixer gate_output_3_730(.a(output_4_730), .b(output_4_11), .y(output_3_730));
wire output_5_730, output_5_11, output_4_730;
mixer gate_output_4_730(.a(output_5_730), .b(output_5_11), .y(output_4_730));
wire output_6_730, output_6_11, output_5_730;
mixer gate_output_5_730(.a(output_6_730), .b(output_6_11), .y(output_5_730));
wire output_7_730, output_7_11, output_6_730;
mixer gate_output_6_730(.a(output_7_730), .b(output_7_11), .y(output_6_730));
wire output_8_730, output_8_11, output_7_730;
mixer gate_output_7_730(.a(output_8_730), .b(output_8_11), .y(output_7_730));
wire output_9_730, output_9_11, output_8_730;
mixer gate_output_8_730(.a(output_9_730), .b(output_9_11), .y(output_8_730));
wire output_10_730, output_10_11, output_9_730;
mixer gate_output_9_730(.a(output_10_730), .b(output_10_11), .y(output_9_730));
wire output_11_730, output_11_11, output_10_730;
mixer gate_output_10_730(.a(output_11_730), .b(output_11_11), .y(output_10_730));
wire output_12_730, output_12_11, output_11_730;
mixer gate_output_11_730(.a(output_12_730), .b(output_12_11), .y(output_11_730));
wire output_13_730, output_13_11, output_12_730;
mixer gate_output_12_730(.a(output_13_730), .b(output_13_11), .y(output_12_730));
wire output_14_730, output_14_11, output_13_730;
mixer gate_output_13_730(.a(output_14_730), .b(output_14_11), .y(output_13_730));
wire output_15_730, output_15_11, output_14_730;
mixer gate_output_14_730(.a(output_15_730), .b(output_15_11), .y(output_14_730));
wire output_16_730, output_16_11, output_15_730;
mixer gate_output_15_730(.a(output_16_730), .b(output_16_11), .y(output_15_730));
wire output_1_731, output_1_12, output_0_731;
mixer gate_output_0_731(.a(output_1_731), .b(output_1_12), .y(output_0_731));
wire output_2_731, output_2_12, output_1_731;
mixer gate_output_1_731(.a(output_2_731), .b(output_2_12), .y(output_1_731));
wire output_3_731, output_3_12, output_2_731;
mixer gate_output_2_731(.a(output_3_731), .b(output_3_12), .y(output_2_731));
wire output_4_731, output_4_12, output_3_731;
mixer gate_output_3_731(.a(output_4_731), .b(output_4_12), .y(output_3_731));
wire output_5_731, output_5_12, output_4_731;
mixer gate_output_4_731(.a(output_5_731), .b(output_5_12), .y(output_4_731));
wire output_6_731, output_6_12, output_5_731;
mixer gate_output_5_731(.a(output_6_731), .b(output_6_12), .y(output_5_731));
wire output_7_731, output_7_12, output_6_731;
mixer gate_output_6_731(.a(output_7_731), .b(output_7_12), .y(output_6_731));
wire output_8_731, output_8_12, output_7_731;
mixer gate_output_7_731(.a(output_8_731), .b(output_8_12), .y(output_7_731));
wire output_9_731, output_9_12, output_8_731;
mixer gate_output_8_731(.a(output_9_731), .b(output_9_12), .y(output_8_731));
wire output_10_731, output_10_12, output_9_731;
mixer gate_output_9_731(.a(output_10_731), .b(output_10_12), .y(output_9_731));
wire output_11_731, output_11_12, output_10_731;
mixer gate_output_10_731(.a(output_11_731), .b(output_11_12), .y(output_10_731));
wire output_12_731, output_12_12, output_11_731;
mixer gate_output_11_731(.a(output_12_731), .b(output_12_12), .y(output_11_731));
wire output_13_731, output_13_12, output_12_731;
mixer gate_output_12_731(.a(output_13_731), .b(output_13_12), .y(output_12_731));
wire output_14_731, output_14_12, output_13_731;
mixer gate_output_13_731(.a(output_14_731), .b(output_14_12), .y(output_13_731));
wire output_15_731, output_15_12, output_14_731;
mixer gate_output_14_731(.a(output_15_731), .b(output_15_12), .y(output_14_731));
wire output_16_731, output_16_12, output_15_731;
mixer gate_output_15_731(.a(output_16_731), .b(output_16_12), .y(output_15_731));
wire output_1_732, output_1_13, output_0_732;
mixer gate_output_0_732(.a(output_1_732), .b(output_1_13), .y(output_0_732));
wire output_2_732, output_2_13, output_1_732;
mixer gate_output_1_732(.a(output_2_732), .b(output_2_13), .y(output_1_732));
wire output_3_732, output_3_13, output_2_732;
mixer gate_output_2_732(.a(output_3_732), .b(output_3_13), .y(output_2_732));
wire output_4_732, output_4_13, output_3_732;
mixer gate_output_3_732(.a(output_4_732), .b(output_4_13), .y(output_3_732));
wire output_5_732, output_5_13, output_4_732;
mixer gate_output_4_732(.a(output_5_732), .b(output_5_13), .y(output_4_732));
wire output_6_732, output_6_13, output_5_732;
mixer gate_output_5_732(.a(output_6_732), .b(output_6_13), .y(output_5_732));
wire output_7_732, output_7_13, output_6_732;
mixer gate_output_6_732(.a(output_7_732), .b(output_7_13), .y(output_6_732));
wire output_8_732, output_8_13, output_7_732;
mixer gate_output_7_732(.a(output_8_732), .b(output_8_13), .y(output_7_732));
wire output_9_732, output_9_13, output_8_732;
mixer gate_output_8_732(.a(output_9_732), .b(output_9_13), .y(output_8_732));
wire output_10_732, output_10_13, output_9_732;
mixer gate_output_9_732(.a(output_10_732), .b(output_10_13), .y(output_9_732));
wire output_11_732, output_11_13, output_10_732;
mixer gate_output_10_732(.a(output_11_732), .b(output_11_13), .y(output_10_732));
wire output_12_732, output_12_13, output_11_732;
mixer gate_output_11_732(.a(output_12_732), .b(output_12_13), .y(output_11_732));
wire output_13_732, output_13_13, output_12_732;
mixer gate_output_12_732(.a(output_13_732), .b(output_13_13), .y(output_12_732));
wire output_14_732, output_14_13, output_13_732;
mixer gate_output_13_732(.a(output_14_732), .b(output_14_13), .y(output_13_732));
wire output_15_732, output_15_13, output_14_732;
mixer gate_output_14_732(.a(output_15_732), .b(output_15_13), .y(output_14_732));
wire output_16_732, output_16_13, output_15_732;
mixer gate_output_15_732(.a(output_16_732), .b(output_16_13), .y(output_15_732));
wire output_1_733, output_1_14, output_0_733;
mixer gate_output_0_733(.a(output_1_733), .b(output_1_14), .y(output_0_733));
wire output_2_733, output_2_14, output_1_733;
mixer gate_output_1_733(.a(output_2_733), .b(output_2_14), .y(output_1_733));
wire output_3_733, output_3_14, output_2_733;
mixer gate_output_2_733(.a(output_3_733), .b(output_3_14), .y(output_2_733));
wire output_4_733, output_4_14, output_3_733;
mixer gate_output_3_733(.a(output_4_733), .b(output_4_14), .y(output_3_733));
wire output_5_733, output_5_14, output_4_733;
mixer gate_output_4_733(.a(output_5_733), .b(output_5_14), .y(output_4_733));
wire output_6_733, output_6_14, output_5_733;
mixer gate_output_5_733(.a(output_6_733), .b(output_6_14), .y(output_5_733));
wire output_7_733, output_7_14, output_6_733;
mixer gate_output_6_733(.a(output_7_733), .b(output_7_14), .y(output_6_733));
wire output_8_733, output_8_14, output_7_733;
mixer gate_output_7_733(.a(output_8_733), .b(output_8_14), .y(output_7_733));
wire output_9_733, output_9_14, output_8_733;
mixer gate_output_8_733(.a(output_9_733), .b(output_9_14), .y(output_8_733));
wire output_10_733, output_10_14, output_9_733;
mixer gate_output_9_733(.a(output_10_733), .b(output_10_14), .y(output_9_733));
wire output_11_733, output_11_14, output_10_733;
mixer gate_output_10_733(.a(output_11_733), .b(output_11_14), .y(output_10_733));
wire output_12_733, output_12_14, output_11_733;
mixer gate_output_11_733(.a(output_12_733), .b(output_12_14), .y(output_11_733));
wire output_13_733, output_13_14, output_12_733;
mixer gate_output_12_733(.a(output_13_733), .b(output_13_14), .y(output_12_733));
wire output_14_733, output_14_14, output_13_733;
mixer gate_output_13_733(.a(output_14_733), .b(output_14_14), .y(output_13_733));
wire output_15_733, output_15_14, output_14_733;
mixer gate_output_14_733(.a(output_15_733), .b(output_15_14), .y(output_14_733));
wire output_16_733, output_16_14, output_15_733;
mixer gate_output_15_733(.a(output_16_733), .b(output_16_14), .y(output_15_733));
wire output_1_734, output_1_15, output_0_734;
mixer gate_output_0_734(.a(output_1_734), .b(output_1_15), .y(output_0_734));
wire output_2_734, output_2_15, output_1_734;
mixer gate_output_1_734(.a(output_2_734), .b(output_2_15), .y(output_1_734));
wire output_3_734, output_3_15, output_2_734;
mixer gate_output_2_734(.a(output_3_734), .b(output_3_15), .y(output_2_734));
wire output_4_734, output_4_15, output_3_734;
mixer gate_output_3_734(.a(output_4_734), .b(output_4_15), .y(output_3_734));
wire output_5_734, output_5_15, output_4_734;
mixer gate_output_4_734(.a(output_5_734), .b(output_5_15), .y(output_4_734));
wire output_6_734, output_6_15, output_5_734;
mixer gate_output_5_734(.a(output_6_734), .b(output_6_15), .y(output_5_734));
wire output_7_734, output_7_15, output_6_734;
mixer gate_output_6_734(.a(output_7_734), .b(output_7_15), .y(output_6_734));
wire output_8_734, output_8_15, output_7_734;
mixer gate_output_7_734(.a(output_8_734), .b(output_8_15), .y(output_7_734));
wire output_9_734, output_9_15, output_8_734;
mixer gate_output_8_734(.a(output_9_734), .b(output_9_15), .y(output_8_734));
wire output_10_734, output_10_15, output_9_734;
mixer gate_output_9_734(.a(output_10_734), .b(output_10_15), .y(output_9_734));
wire output_11_734, output_11_15, output_10_734;
mixer gate_output_10_734(.a(output_11_734), .b(output_11_15), .y(output_10_734));
wire output_12_734, output_12_15, output_11_734;
mixer gate_output_11_734(.a(output_12_734), .b(output_12_15), .y(output_11_734));
wire output_13_734, output_13_15, output_12_734;
mixer gate_output_12_734(.a(output_13_734), .b(output_13_15), .y(output_12_734));
wire output_14_734, output_14_15, output_13_734;
mixer gate_output_13_734(.a(output_14_734), .b(output_14_15), .y(output_13_734));
wire output_15_734, output_15_15, output_14_734;
mixer gate_output_14_734(.a(output_15_734), .b(output_15_15), .y(output_14_734));
wire output_16_734, output_16_15, output_15_734;
mixer gate_output_15_734(.a(output_16_734), .b(output_16_15), .y(output_15_734));
wire output_1_735, output_1_0, output_0_735;
mixer gate_output_0_735(.a(output_1_735), .b(output_1_0), .y(output_0_735));
wire output_2_735, output_2_0, output_1_735;
mixer gate_output_1_735(.a(output_2_735), .b(output_2_0), .y(output_1_735));
wire output_3_735, output_3_0, output_2_735;
mixer gate_output_2_735(.a(output_3_735), .b(output_3_0), .y(output_2_735));
wire output_4_735, output_4_0, output_3_735;
mixer gate_output_3_735(.a(output_4_735), .b(output_4_0), .y(output_3_735));
wire output_5_735, output_5_0, output_4_735;
mixer gate_output_4_735(.a(output_5_735), .b(output_5_0), .y(output_4_735));
wire output_6_735, output_6_0, output_5_735;
mixer gate_output_5_735(.a(output_6_735), .b(output_6_0), .y(output_5_735));
wire output_7_735, output_7_0, output_6_735;
mixer gate_output_6_735(.a(output_7_735), .b(output_7_0), .y(output_6_735));
wire output_8_735, output_8_0, output_7_735;
mixer gate_output_7_735(.a(output_8_735), .b(output_8_0), .y(output_7_735));
wire output_9_735, output_9_0, output_8_735;
mixer gate_output_8_735(.a(output_9_735), .b(output_9_0), .y(output_8_735));
wire output_10_735, output_10_0, output_9_735;
mixer gate_output_9_735(.a(output_10_735), .b(output_10_0), .y(output_9_735));
wire output_11_735, output_11_0, output_10_735;
mixer gate_output_10_735(.a(output_11_735), .b(output_11_0), .y(output_10_735));
wire output_12_735, output_12_0, output_11_735;
mixer gate_output_11_735(.a(output_12_735), .b(output_12_0), .y(output_11_735));
wire output_13_735, output_13_0, output_12_735;
mixer gate_output_12_735(.a(output_13_735), .b(output_13_0), .y(output_12_735));
wire output_14_735, output_14_0, output_13_735;
mixer gate_output_13_735(.a(output_14_735), .b(output_14_0), .y(output_13_735));
wire output_15_735, output_15_0, output_14_735;
mixer gate_output_14_735(.a(output_15_735), .b(output_15_0), .y(output_14_735));
wire output_16_735, output_16_0, output_15_735;
mixer gate_output_15_735(.a(output_16_735), .b(output_16_0), .y(output_15_735));
wire output_1_736, output_1_1, output_0_736;
mixer gate_output_0_736(.a(output_1_736), .b(output_1_1), .y(output_0_736));
wire output_2_736, output_2_1, output_1_736;
mixer gate_output_1_736(.a(output_2_736), .b(output_2_1), .y(output_1_736));
wire output_3_736, output_3_1, output_2_736;
mixer gate_output_2_736(.a(output_3_736), .b(output_3_1), .y(output_2_736));
wire output_4_736, output_4_1, output_3_736;
mixer gate_output_3_736(.a(output_4_736), .b(output_4_1), .y(output_3_736));
wire output_5_736, output_5_1, output_4_736;
mixer gate_output_4_736(.a(output_5_736), .b(output_5_1), .y(output_4_736));
wire output_6_736, output_6_1, output_5_736;
mixer gate_output_5_736(.a(output_6_736), .b(output_6_1), .y(output_5_736));
wire output_7_736, output_7_1, output_6_736;
mixer gate_output_6_736(.a(output_7_736), .b(output_7_1), .y(output_6_736));
wire output_8_736, output_8_1, output_7_736;
mixer gate_output_7_736(.a(output_8_736), .b(output_8_1), .y(output_7_736));
wire output_9_736, output_9_1, output_8_736;
mixer gate_output_8_736(.a(output_9_736), .b(output_9_1), .y(output_8_736));
wire output_10_736, output_10_1, output_9_736;
mixer gate_output_9_736(.a(output_10_736), .b(output_10_1), .y(output_9_736));
wire output_11_736, output_11_1, output_10_736;
mixer gate_output_10_736(.a(output_11_736), .b(output_11_1), .y(output_10_736));
wire output_12_736, output_12_1, output_11_736;
mixer gate_output_11_736(.a(output_12_736), .b(output_12_1), .y(output_11_736));
wire output_13_736, output_13_1, output_12_736;
mixer gate_output_12_736(.a(output_13_736), .b(output_13_1), .y(output_12_736));
wire output_14_736, output_14_1, output_13_736;
mixer gate_output_13_736(.a(output_14_736), .b(output_14_1), .y(output_13_736));
wire output_15_736, output_15_1, output_14_736;
mixer gate_output_14_736(.a(output_15_736), .b(output_15_1), .y(output_14_736));
wire output_16_736, output_16_1, output_15_736;
mixer gate_output_15_736(.a(output_16_736), .b(output_16_1), .y(output_15_736));
wire output_1_737, output_1_2, output_0_737;
mixer gate_output_0_737(.a(output_1_737), .b(output_1_2), .y(output_0_737));
wire output_2_737, output_2_2, output_1_737;
mixer gate_output_1_737(.a(output_2_737), .b(output_2_2), .y(output_1_737));
wire output_3_737, output_3_2, output_2_737;
mixer gate_output_2_737(.a(output_3_737), .b(output_3_2), .y(output_2_737));
wire output_4_737, output_4_2, output_3_737;
mixer gate_output_3_737(.a(output_4_737), .b(output_4_2), .y(output_3_737));
wire output_5_737, output_5_2, output_4_737;
mixer gate_output_4_737(.a(output_5_737), .b(output_5_2), .y(output_4_737));
wire output_6_737, output_6_2, output_5_737;
mixer gate_output_5_737(.a(output_6_737), .b(output_6_2), .y(output_5_737));
wire output_7_737, output_7_2, output_6_737;
mixer gate_output_6_737(.a(output_7_737), .b(output_7_2), .y(output_6_737));
wire output_8_737, output_8_2, output_7_737;
mixer gate_output_7_737(.a(output_8_737), .b(output_8_2), .y(output_7_737));
wire output_9_737, output_9_2, output_8_737;
mixer gate_output_8_737(.a(output_9_737), .b(output_9_2), .y(output_8_737));
wire output_10_737, output_10_2, output_9_737;
mixer gate_output_9_737(.a(output_10_737), .b(output_10_2), .y(output_9_737));
wire output_11_737, output_11_2, output_10_737;
mixer gate_output_10_737(.a(output_11_737), .b(output_11_2), .y(output_10_737));
wire output_12_737, output_12_2, output_11_737;
mixer gate_output_11_737(.a(output_12_737), .b(output_12_2), .y(output_11_737));
wire output_13_737, output_13_2, output_12_737;
mixer gate_output_12_737(.a(output_13_737), .b(output_13_2), .y(output_12_737));
wire output_14_737, output_14_2, output_13_737;
mixer gate_output_13_737(.a(output_14_737), .b(output_14_2), .y(output_13_737));
wire output_15_737, output_15_2, output_14_737;
mixer gate_output_14_737(.a(output_15_737), .b(output_15_2), .y(output_14_737));
wire output_16_737, output_16_2, output_15_737;
mixer gate_output_15_737(.a(output_16_737), .b(output_16_2), .y(output_15_737));
wire output_1_738, output_1_3, output_0_738;
mixer gate_output_0_738(.a(output_1_738), .b(output_1_3), .y(output_0_738));
wire output_2_738, output_2_3, output_1_738;
mixer gate_output_1_738(.a(output_2_738), .b(output_2_3), .y(output_1_738));
wire output_3_738, output_3_3, output_2_738;
mixer gate_output_2_738(.a(output_3_738), .b(output_3_3), .y(output_2_738));
wire output_4_738, output_4_3, output_3_738;
mixer gate_output_3_738(.a(output_4_738), .b(output_4_3), .y(output_3_738));
wire output_5_738, output_5_3, output_4_738;
mixer gate_output_4_738(.a(output_5_738), .b(output_5_3), .y(output_4_738));
wire output_6_738, output_6_3, output_5_738;
mixer gate_output_5_738(.a(output_6_738), .b(output_6_3), .y(output_5_738));
wire output_7_738, output_7_3, output_6_738;
mixer gate_output_6_738(.a(output_7_738), .b(output_7_3), .y(output_6_738));
wire output_8_738, output_8_3, output_7_738;
mixer gate_output_7_738(.a(output_8_738), .b(output_8_3), .y(output_7_738));
wire output_9_738, output_9_3, output_8_738;
mixer gate_output_8_738(.a(output_9_738), .b(output_9_3), .y(output_8_738));
wire output_10_738, output_10_3, output_9_738;
mixer gate_output_9_738(.a(output_10_738), .b(output_10_3), .y(output_9_738));
wire output_11_738, output_11_3, output_10_738;
mixer gate_output_10_738(.a(output_11_738), .b(output_11_3), .y(output_10_738));
wire output_12_738, output_12_3, output_11_738;
mixer gate_output_11_738(.a(output_12_738), .b(output_12_3), .y(output_11_738));
wire output_13_738, output_13_3, output_12_738;
mixer gate_output_12_738(.a(output_13_738), .b(output_13_3), .y(output_12_738));
wire output_14_738, output_14_3, output_13_738;
mixer gate_output_13_738(.a(output_14_738), .b(output_14_3), .y(output_13_738));
wire output_15_738, output_15_3, output_14_738;
mixer gate_output_14_738(.a(output_15_738), .b(output_15_3), .y(output_14_738));
wire output_16_738, output_16_3, output_15_738;
mixer gate_output_15_738(.a(output_16_738), .b(output_16_3), .y(output_15_738));
wire output_1_739, output_1_4, output_0_739;
mixer gate_output_0_739(.a(output_1_739), .b(output_1_4), .y(output_0_739));
wire output_2_739, output_2_4, output_1_739;
mixer gate_output_1_739(.a(output_2_739), .b(output_2_4), .y(output_1_739));
wire output_3_739, output_3_4, output_2_739;
mixer gate_output_2_739(.a(output_3_739), .b(output_3_4), .y(output_2_739));
wire output_4_739, output_4_4, output_3_739;
mixer gate_output_3_739(.a(output_4_739), .b(output_4_4), .y(output_3_739));
wire output_5_739, output_5_4, output_4_739;
mixer gate_output_4_739(.a(output_5_739), .b(output_5_4), .y(output_4_739));
wire output_6_739, output_6_4, output_5_739;
mixer gate_output_5_739(.a(output_6_739), .b(output_6_4), .y(output_5_739));
wire output_7_739, output_7_4, output_6_739;
mixer gate_output_6_739(.a(output_7_739), .b(output_7_4), .y(output_6_739));
wire output_8_739, output_8_4, output_7_739;
mixer gate_output_7_739(.a(output_8_739), .b(output_8_4), .y(output_7_739));
wire output_9_739, output_9_4, output_8_739;
mixer gate_output_8_739(.a(output_9_739), .b(output_9_4), .y(output_8_739));
wire output_10_739, output_10_4, output_9_739;
mixer gate_output_9_739(.a(output_10_739), .b(output_10_4), .y(output_9_739));
wire output_11_739, output_11_4, output_10_739;
mixer gate_output_10_739(.a(output_11_739), .b(output_11_4), .y(output_10_739));
wire output_12_739, output_12_4, output_11_739;
mixer gate_output_11_739(.a(output_12_739), .b(output_12_4), .y(output_11_739));
wire output_13_739, output_13_4, output_12_739;
mixer gate_output_12_739(.a(output_13_739), .b(output_13_4), .y(output_12_739));
wire output_14_739, output_14_4, output_13_739;
mixer gate_output_13_739(.a(output_14_739), .b(output_14_4), .y(output_13_739));
wire output_15_739, output_15_4, output_14_739;
mixer gate_output_14_739(.a(output_15_739), .b(output_15_4), .y(output_14_739));
wire output_16_739, output_16_4, output_15_739;
mixer gate_output_15_739(.a(output_16_739), .b(output_16_4), .y(output_15_739));
wire output_1_740, output_1_5, output_0_740;
mixer gate_output_0_740(.a(output_1_740), .b(output_1_5), .y(output_0_740));
wire output_2_740, output_2_5, output_1_740;
mixer gate_output_1_740(.a(output_2_740), .b(output_2_5), .y(output_1_740));
wire output_3_740, output_3_5, output_2_740;
mixer gate_output_2_740(.a(output_3_740), .b(output_3_5), .y(output_2_740));
wire output_4_740, output_4_5, output_3_740;
mixer gate_output_3_740(.a(output_4_740), .b(output_4_5), .y(output_3_740));
wire output_5_740, output_5_5, output_4_740;
mixer gate_output_4_740(.a(output_5_740), .b(output_5_5), .y(output_4_740));
wire output_6_740, output_6_5, output_5_740;
mixer gate_output_5_740(.a(output_6_740), .b(output_6_5), .y(output_5_740));
wire output_7_740, output_7_5, output_6_740;
mixer gate_output_6_740(.a(output_7_740), .b(output_7_5), .y(output_6_740));
wire output_8_740, output_8_5, output_7_740;
mixer gate_output_7_740(.a(output_8_740), .b(output_8_5), .y(output_7_740));
wire output_9_740, output_9_5, output_8_740;
mixer gate_output_8_740(.a(output_9_740), .b(output_9_5), .y(output_8_740));
wire output_10_740, output_10_5, output_9_740;
mixer gate_output_9_740(.a(output_10_740), .b(output_10_5), .y(output_9_740));
wire output_11_740, output_11_5, output_10_740;
mixer gate_output_10_740(.a(output_11_740), .b(output_11_5), .y(output_10_740));
wire output_12_740, output_12_5, output_11_740;
mixer gate_output_11_740(.a(output_12_740), .b(output_12_5), .y(output_11_740));
wire output_13_740, output_13_5, output_12_740;
mixer gate_output_12_740(.a(output_13_740), .b(output_13_5), .y(output_12_740));
wire output_14_740, output_14_5, output_13_740;
mixer gate_output_13_740(.a(output_14_740), .b(output_14_5), .y(output_13_740));
wire output_15_740, output_15_5, output_14_740;
mixer gate_output_14_740(.a(output_15_740), .b(output_15_5), .y(output_14_740));
wire output_16_740, output_16_5, output_15_740;
mixer gate_output_15_740(.a(output_16_740), .b(output_16_5), .y(output_15_740));
wire output_1_741, output_1_6, output_0_741;
mixer gate_output_0_741(.a(output_1_741), .b(output_1_6), .y(output_0_741));
wire output_2_741, output_2_6, output_1_741;
mixer gate_output_1_741(.a(output_2_741), .b(output_2_6), .y(output_1_741));
wire output_3_741, output_3_6, output_2_741;
mixer gate_output_2_741(.a(output_3_741), .b(output_3_6), .y(output_2_741));
wire output_4_741, output_4_6, output_3_741;
mixer gate_output_3_741(.a(output_4_741), .b(output_4_6), .y(output_3_741));
wire output_5_741, output_5_6, output_4_741;
mixer gate_output_4_741(.a(output_5_741), .b(output_5_6), .y(output_4_741));
wire output_6_741, output_6_6, output_5_741;
mixer gate_output_5_741(.a(output_6_741), .b(output_6_6), .y(output_5_741));
wire output_7_741, output_7_6, output_6_741;
mixer gate_output_6_741(.a(output_7_741), .b(output_7_6), .y(output_6_741));
wire output_8_741, output_8_6, output_7_741;
mixer gate_output_7_741(.a(output_8_741), .b(output_8_6), .y(output_7_741));
wire output_9_741, output_9_6, output_8_741;
mixer gate_output_8_741(.a(output_9_741), .b(output_9_6), .y(output_8_741));
wire output_10_741, output_10_6, output_9_741;
mixer gate_output_9_741(.a(output_10_741), .b(output_10_6), .y(output_9_741));
wire output_11_741, output_11_6, output_10_741;
mixer gate_output_10_741(.a(output_11_741), .b(output_11_6), .y(output_10_741));
wire output_12_741, output_12_6, output_11_741;
mixer gate_output_11_741(.a(output_12_741), .b(output_12_6), .y(output_11_741));
wire output_13_741, output_13_6, output_12_741;
mixer gate_output_12_741(.a(output_13_741), .b(output_13_6), .y(output_12_741));
wire output_14_741, output_14_6, output_13_741;
mixer gate_output_13_741(.a(output_14_741), .b(output_14_6), .y(output_13_741));
wire output_15_741, output_15_6, output_14_741;
mixer gate_output_14_741(.a(output_15_741), .b(output_15_6), .y(output_14_741));
wire output_16_741, output_16_6, output_15_741;
mixer gate_output_15_741(.a(output_16_741), .b(output_16_6), .y(output_15_741));
wire output_1_742, output_1_7, output_0_742;
mixer gate_output_0_742(.a(output_1_742), .b(output_1_7), .y(output_0_742));
wire output_2_742, output_2_7, output_1_742;
mixer gate_output_1_742(.a(output_2_742), .b(output_2_7), .y(output_1_742));
wire output_3_742, output_3_7, output_2_742;
mixer gate_output_2_742(.a(output_3_742), .b(output_3_7), .y(output_2_742));
wire output_4_742, output_4_7, output_3_742;
mixer gate_output_3_742(.a(output_4_742), .b(output_4_7), .y(output_3_742));
wire output_5_742, output_5_7, output_4_742;
mixer gate_output_4_742(.a(output_5_742), .b(output_5_7), .y(output_4_742));
wire output_6_742, output_6_7, output_5_742;
mixer gate_output_5_742(.a(output_6_742), .b(output_6_7), .y(output_5_742));
wire output_7_742, output_7_7, output_6_742;
mixer gate_output_6_742(.a(output_7_742), .b(output_7_7), .y(output_6_742));
wire output_8_742, output_8_7, output_7_742;
mixer gate_output_7_742(.a(output_8_742), .b(output_8_7), .y(output_7_742));
wire output_9_742, output_9_7, output_8_742;
mixer gate_output_8_742(.a(output_9_742), .b(output_9_7), .y(output_8_742));
wire output_10_742, output_10_7, output_9_742;
mixer gate_output_9_742(.a(output_10_742), .b(output_10_7), .y(output_9_742));
wire output_11_742, output_11_7, output_10_742;
mixer gate_output_10_742(.a(output_11_742), .b(output_11_7), .y(output_10_742));
wire output_12_742, output_12_7, output_11_742;
mixer gate_output_11_742(.a(output_12_742), .b(output_12_7), .y(output_11_742));
wire output_13_742, output_13_7, output_12_742;
mixer gate_output_12_742(.a(output_13_742), .b(output_13_7), .y(output_12_742));
wire output_14_742, output_14_7, output_13_742;
mixer gate_output_13_742(.a(output_14_742), .b(output_14_7), .y(output_13_742));
wire output_15_742, output_15_7, output_14_742;
mixer gate_output_14_742(.a(output_15_742), .b(output_15_7), .y(output_14_742));
wire output_16_742, output_16_7, output_15_742;
mixer gate_output_15_742(.a(output_16_742), .b(output_16_7), .y(output_15_742));
wire output_1_743, output_1_8, output_0_743;
mixer gate_output_0_743(.a(output_1_743), .b(output_1_8), .y(output_0_743));
wire output_2_743, output_2_8, output_1_743;
mixer gate_output_1_743(.a(output_2_743), .b(output_2_8), .y(output_1_743));
wire output_3_743, output_3_8, output_2_743;
mixer gate_output_2_743(.a(output_3_743), .b(output_3_8), .y(output_2_743));
wire output_4_743, output_4_8, output_3_743;
mixer gate_output_3_743(.a(output_4_743), .b(output_4_8), .y(output_3_743));
wire output_5_743, output_5_8, output_4_743;
mixer gate_output_4_743(.a(output_5_743), .b(output_5_8), .y(output_4_743));
wire output_6_743, output_6_8, output_5_743;
mixer gate_output_5_743(.a(output_6_743), .b(output_6_8), .y(output_5_743));
wire output_7_743, output_7_8, output_6_743;
mixer gate_output_6_743(.a(output_7_743), .b(output_7_8), .y(output_6_743));
wire output_8_743, output_8_8, output_7_743;
mixer gate_output_7_743(.a(output_8_743), .b(output_8_8), .y(output_7_743));
wire output_9_743, output_9_8, output_8_743;
mixer gate_output_8_743(.a(output_9_743), .b(output_9_8), .y(output_8_743));
wire output_10_743, output_10_8, output_9_743;
mixer gate_output_9_743(.a(output_10_743), .b(output_10_8), .y(output_9_743));
wire output_11_743, output_11_8, output_10_743;
mixer gate_output_10_743(.a(output_11_743), .b(output_11_8), .y(output_10_743));
wire output_12_743, output_12_8, output_11_743;
mixer gate_output_11_743(.a(output_12_743), .b(output_12_8), .y(output_11_743));
wire output_13_743, output_13_8, output_12_743;
mixer gate_output_12_743(.a(output_13_743), .b(output_13_8), .y(output_12_743));
wire output_14_743, output_14_8, output_13_743;
mixer gate_output_13_743(.a(output_14_743), .b(output_14_8), .y(output_13_743));
wire output_15_743, output_15_8, output_14_743;
mixer gate_output_14_743(.a(output_15_743), .b(output_15_8), .y(output_14_743));
wire output_16_743, output_16_8, output_15_743;
mixer gate_output_15_743(.a(output_16_743), .b(output_16_8), .y(output_15_743));
wire output_1_744, output_1_9, output_0_744;
mixer gate_output_0_744(.a(output_1_744), .b(output_1_9), .y(output_0_744));
wire output_2_744, output_2_9, output_1_744;
mixer gate_output_1_744(.a(output_2_744), .b(output_2_9), .y(output_1_744));
wire output_3_744, output_3_9, output_2_744;
mixer gate_output_2_744(.a(output_3_744), .b(output_3_9), .y(output_2_744));
wire output_4_744, output_4_9, output_3_744;
mixer gate_output_3_744(.a(output_4_744), .b(output_4_9), .y(output_3_744));
wire output_5_744, output_5_9, output_4_744;
mixer gate_output_4_744(.a(output_5_744), .b(output_5_9), .y(output_4_744));
wire output_6_744, output_6_9, output_5_744;
mixer gate_output_5_744(.a(output_6_744), .b(output_6_9), .y(output_5_744));
wire output_7_744, output_7_9, output_6_744;
mixer gate_output_6_744(.a(output_7_744), .b(output_7_9), .y(output_6_744));
wire output_8_744, output_8_9, output_7_744;
mixer gate_output_7_744(.a(output_8_744), .b(output_8_9), .y(output_7_744));
wire output_9_744, output_9_9, output_8_744;
mixer gate_output_8_744(.a(output_9_744), .b(output_9_9), .y(output_8_744));
wire output_10_744, output_10_9, output_9_744;
mixer gate_output_9_744(.a(output_10_744), .b(output_10_9), .y(output_9_744));
wire output_11_744, output_11_9, output_10_744;
mixer gate_output_10_744(.a(output_11_744), .b(output_11_9), .y(output_10_744));
wire output_12_744, output_12_9, output_11_744;
mixer gate_output_11_744(.a(output_12_744), .b(output_12_9), .y(output_11_744));
wire output_13_744, output_13_9, output_12_744;
mixer gate_output_12_744(.a(output_13_744), .b(output_13_9), .y(output_12_744));
wire output_14_744, output_14_9, output_13_744;
mixer gate_output_13_744(.a(output_14_744), .b(output_14_9), .y(output_13_744));
wire output_15_744, output_15_9, output_14_744;
mixer gate_output_14_744(.a(output_15_744), .b(output_15_9), .y(output_14_744));
wire output_16_744, output_16_9, output_15_744;
mixer gate_output_15_744(.a(output_16_744), .b(output_16_9), .y(output_15_744));
wire output_1_745, output_1_10, output_0_745;
mixer gate_output_0_745(.a(output_1_745), .b(output_1_10), .y(output_0_745));
wire output_2_745, output_2_10, output_1_745;
mixer gate_output_1_745(.a(output_2_745), .b(output_2_10), .y(output_1_745));
wire output_3_745, output_3_10, output_2_745;
mixer gate_output_2_745(.a(output_3_745), .b(output_3_10), .y(output_2_745));
wire output_4_745, output_4_10, output_3_745;
mixer gate_output_3_745(.a(output_4_745), .b(output_4_10), .y(output_3_745));
wire output_5_745, output_5_10, output_4_745;
mixer gate_output_4_745(.a(output_5_745), .b(output_5_10), .y(output_4_745));
wire output_6_745, output_6_10, output_5_745;
mixer gate_output_5_745(.a(output_6_745), .b(output_6_10), .y(output_5_745));
wire output_7_745, output_7_10, output_6_745;
mixer gate_output_6_745(.a(output_7_745), .b(output_7_10), .y(output_6_745));
wire output_8_745, output_8_10, output_7_745;
mixer gate_output_7_745(.a(output_8_745), .b(output_8_10), .y(output_7_745));
wire output_9_745, output_9_10, output_8_745;
mixer gate_output_8_745(.a(output_9_745), .b(output_9_10), .y(output_8_745));
wire output_10_745, output_10_10, output_9_745;
mixer gate_output_9_745(.a(output_10_745), .b(output_10_10), .y(output_9_745));
wire output_11_745, output_11_10, output_10_745;
mixer gate_output_10_745(.a(output_11_745), .b(output_11_10), .y(output_10_745));
wire output_12_745, output_12_10, output_11_745;
mixer gate_output_11_745(.a(output_12_745), .b(output_12_10), .y(output_11_745));
wire output_13_745, output_13_10, output_12_745;
mixer gate_output_12_745(.a(output_13_745), .b(output_13_10), .y(output_12_745));
wire output_14_745, output_14_10, output_13_745;
mixer gate_output_13_745(.a(output_14_745), .b(output_14_10), .y(output_13_745));
wire output_15_745, output_15_10, output_14_745;
mixer gate_output_14_745(.a(output_15_745), .b(output_15_10), .y(output_14_745));
wire output_16_745, output_16_10, output_15_745;
mixer gate_output_15_745(.a(output_16_745), .b(output_16_10), .y(output_15_745));
wire output_1_746, output_1_11, output_0_746;
mixer gate_output_0_746(.a(output_1_746), .b(output_1_11), .y(output_0_746));
wire output_2_746, output_2_11, output_1_746;
mixer gate_output_1_746(.a(output_2_746), .b(output_2_11), .y(output_1_746));
wire output_3_746, output_3_11, output_2_746;
mixer gate_output_2_746(.a(output_3_746), .b(output_3_11), .y(output_2_746));
wire output_4_746, output_4_11, output_3_746;
mixer gate_output_3_746(.a(output_4_746), .b(output_4_11), .y(output_3_746));
wire output_5_746, output_5_11, output_4_746;
mixer gate_output_4_746(.a(output_5_746), .b(output_5_11), .y(output_4_746));
wire output_6_746, output_6_11, output_5_746;
mixer gate_output_5_746(.a(output_6_746), .b(output_6_11), .y(output_5_746));
wire output_7_746, output_7_11, output_6_746;
mixer gate_output_6_746(.a(output_7_746), .b(output_7_11), .y(output_6_746));
wire output_8_746, output_8_11, output_7_746;
mixer gate_output_7_746(.a(output_8_746), .b(output_8_11), .y(output_7_746));
wire output_9_746, output_9_11, output_8_746;
mixer gate_output_8_746(.a(output_9_746), .b(output_9_11), .y(output_8_746));
wire output_10_746, output_10_11, output_9_746;
mixer gate_output_9_746(.a(output_10_746), .b(output_10_11), .y(output_9_746));
wire output_11_746, output_11_11, output_10_746;
mixer gate_output_10_746(.a(output_11_746), .b(output_11_11), .y(output_10_746));
wire output_12_746, output_12_11, output_11_746;
mixer gate_output_11_746(.a(output_12_746), .b(output_12_11), .y(output_11_746));
wire output_13_746, output_13_11, output_12_746;
mixer gate_output_12_746(.a(output_13_746), .b(output_13_11), .y(output_12_746));
wire output_14_746, output_14_11, output_13_746;
mixer gate_output_13_746(.a(output_14_746), .b(output_14_11), .y(output_13_746));
wire output_15_746, output_15_11, output_14_746;
mixer gate_output_14_746(.a(output_15_746), .b(output_15_11), .y(output_14_746));
wire output_16_746, output_16_11, output_15_746;
mixer gate_output_15_746(.a(output_16_746), .b(output_16_11), .y(output_15_746));
wire output_1_747, output_1_12, output_0_747;
mixer gate_output_0_747(.a(output_1_747), .b(output_1_12), .y(output_0_747));
wire output_2_747, output_2_12, output_1_747;
mixer gate_output_1_747(.a(output_2_747), .b(output_2_12), .y(output_1_747));
wire output_3_747, output_3_12, output_2_747;
mixer gate_output_2_747(.a(output_3_747), .b(output_3_12), .y(output_2_747));
wire output_4_747, output_4_12, output_3_747;
mixer gate_output_3_747(.a(output_4_747), .b(output_4_12), .y(output_3_747));
wire output_5_747, output_5_12, output_4_747;
mixer gate_output_4_747(.a(output_5_747), .b(output_5_12), .y(output_4_747));
wire output_6_747, output_6_12, output_5_747;
mixer gate_output_5_747(.a(output_6_747), .b(output_6_12), .y(output_5_747));
wire output_7_747, output_7_12, output_6_747;
mixer gate_output_6_747(.a(output_7_747), .b(output_7_12), .y(output_6_747));
wire output_8_747, output_8_12, output_7_747;
mixer gate_output_7_747(.a(output_8_747), .b(output_8_12), .y(output_7_747));
wire output_9_747, output_9_12, output_8_747;
mixer gate_output_8_747(.a(output_9_747), .b(output_9_12), .y(output_8_747));
wire output_10_747, output_10_12, output_9_747;
mixer gate_output_9_747(.a(output_10_747), .b(output_10_12), .y(output_9_747));
wire output_11_747, output_11_12, output_10_747;
mixer gate_output_10_747(.a(output_11_747), .b(output_11_12), .y(output_10_747));
wire output_12_747, output_12_12, output_11_747;
mixer gate_output_11_747(.a(output_12_747), .b(output_12_12), .y(output_11_747));
wire output_13_747, output_13_12, output_12_747;
mixer gate_output_12_747(.a(output_13_747), .b(output_13_12), .y(output_12_747));
wire output_14_747, output_14_12, output_13_747;
mixer gate_output_13_747(.a(output_14_747), .b(output_14_12), .y(output_13_747));
wire output_15_747, output_15_12, output_14_747;
mixer gate_output_14_747(.a(output_15_747), .b(output_15_12), .y(output_14_747));
wire output_16_747, output_16_12, output_15_747;
mixer gate_output_15_747(.a(output_16_747), .b(output_16_12), .y(output_15_747));
wire output_1_748, output_1_13, output_0_748;
mixer gate_output_0_748(.a(output_1_748), .b(output_1_13), .y(output_0_748));
wire output_2_748, output_2_13, output_1_748;
mixer gate_output_1_748(.a(output_2_748), .b(output_2_13), .y(output_1_748));
wire output_3_748, output_3_13, output_2_748;
mixer gate_output_2_748(.a(output_3_748), .b(output_3_13), .y(output_2_748));
wire output_4_748, output_4_13, output_3_748;
mixer gate_output_3_748(.a(output_4_748), .b(output_4_13), .y(output_3_748));
wire output_5_748, output_5_13, output_4_748;
mixer gate_output_4_748(.a(output_5_748), .b(output_5_13), .y(output_4_748));
wire output_6_748, output_6_13, output_5_748;
mixer gate_output_5_748(.a(output_6_748), .b(output_6_13), .y(output_5_748));
wire output_7_748, output_7_13, output_6_748;
mixer gate_output_6_748(.a(output_7_748), .b(output_7_13), .y(output_6_748));
wire output_8_748, output_8_13, output_7_748;
mixer gate_output_7_748(.a(output_8_748), .b(output_8_13), .y(output_7_748));
wire output_9_748, output_9_13, output_8_748;
mixer gate_output_8_748(.a(output_9_748), .b(output_9_13), .y(output_8_748));
wire output_10_748, output_10_13, output_9_748;
mixer gate_output_9_748(.a(output_10_748), .b(output_10_13), .y(output_9_748));
wire output_11_748, output_11_13, output_10_748;
mixer gate_output_10_748(.a(output_11_748), .b(output_11_13), .y(output_10_748));
wire output_12_748, output_12_13, output_11_748;
mixer gate_output_11_748(.a(output_12_748), .b(output_12_13), .y(output_11_748));
wire output_13_748, output_13_13, output_12_748;
mixer gate_output_12_748(.a(output_13_748), .b(output_13_13), .y(output_12_748));
wire output_14_748, output_14_13, output_13_748;
mixer gate_output_13_748(.a(output_14_748), .b(output_14_13), .y(output_13_748));
wire output_15_748, output_15_13, output_14_748;
mixer gate_output_14_748(.a(output_15_748), .b(output_15_13), .y(output_14_748));
wire output_16_748, output_16_13, output_15_748;
mixer gate_output_15_748(.a(output_16_748), .b(output_16_13), .y(output_15_748));
wire output_1_749, output_1_14, output_0_749;
mixer gate_output_0_749(.a(output_1_749), .b(output_1_14), .y(output_0_749));
wire output_2_749, output_2_14, output_1_749;
mixer gate_output_1_749(.a(output_2_749), .b(output_2_14), .y(output_1_749));
wire output_3_749, output_3_14, output_2_749;
mixer gate_output_2_749(.a(output_3_749), .b(output_3_14), .y(output_2_749));
wire output_4_749, output_4_14, output_3_749;
mixer gate_output_3_749(.a(output_4_749), .b(output_4_14), .y(output_3_749));
wire output_5_749, output_5_14, output_4_749;
mixer gate_output_4_749(.a(output_5_749), .b(output_5_14), .y(output_4_749));
wire output_6_749, output_6_14, output_5_749;
mixer gate_output_5_749(.a(output_6_749), .b(output_6_14), .y(output_5_749));
wire output_7_749, output_7_14, output_6_749;
mixer gate_output_6_749(.a(output_7_749), .b(output_7_14), .y(output_6_749));
wire output_8_749, output_8_14, output_7_749;
mixer gate_output_7_749(.a(output_8_749), .b(output_8_14), .y(output_7_749));
wire output_9_749, output_9_14, output_8_749;
mixer gate_output_8_749(.a(output_9_749), .b(output_9_14), .y(output_8_749));
wire output_10_749, output_10_14, output_9_749;
mixer gate_output_9_749(.a(output_10_749), .b(output_10_14), .y(output_9_749));
wire output_11_749, output_11_14, output_10_749;
mixer gate_output_10_749(.a(output_11_749), .b(output_11_14), .y(output_10_749));
wire output_12_749, output_12_14, output_11_749;
mixer gate_output_11_749(.a(output_12_749), .b(output_12_14), .y(output_11_749));
wire output_13_749, output_13_14, output_12_749;
mixer gate_output_12_749(.a(output_13_749), .b(output_13_14), .y(output_12_749));
wire output_14_749, output_14_14, output_13_749;
mixer gate_output_13_749(.a(output_14_749), .b(output_14_14), .y(output_13_749));
wire output_15_749, output_15_14, output_14_749;
mixer gate_output_14_749(.a(output_15_749), .b(output_15_14), .y(output_14_749));
wire output_16_749, output_16_14, output_15_749;
mixer gate_output_15_749(.a(output_16_749), .b(output_16_14), .y(output_15_749));
wire output_1_750, output_1_15, output_0_750;
mixer gate_output_0_750(.a(output_1_750), .b(output_1_15), .y(output_0_750));
wire output_2_750, output_2_15, output_1_750;
mixer gate_output_1_750(.a(output_2_750), .b(output_2_15), .y(output_1_750));
wire output_3_750, output_3_15, output_2_750;
mixer gate_output_2_750(.a(output_3_750), .b(output_3_15), .y(output_2_750));
wire output_4_750, output_4_15, output_3_750;
mixer gate_output_3_750(.a(output_4_750), .b(output_4_15), .y(output_3_750));
wire output_5_750, output_5_15, output_4_750;
mixer gate_output_4_750(.a(output_5_750), .b(output_5_15), .y(output_4_750));
wire output_6_750, output_6_15, output_5_750;
mixer gate_output_5_750(.a(output_6_750), .b(output_6_15), .y(output_5_750));
wire output_7_750, output_7_15, output_6_750;
mixer gate_output_6_750(.a(output_7_750), .b(output_7_15), .y(output_6_750));
wire output_8_750, output_8_15, output_7_750;
mixer gate_output_7_750(.a(output_8_750), .b(output_8_15), .y(output_7_750));
wire output_9_750, output_9_15, output_8_750;
mixer gate_output_8_750(.a(output_9_750), .b(output_9_15), .y(output_8_750));
wire output_10_750, output_10_15, output_9_750;
mixer gate_output_9_750(.a(output_10_750), .b(output_10_15), .y(output_9_750));
wire output_11_750, output_11_15, output_10_750;
mixer gate_output_10_750(.a(output_11_750), .b(output_11_15), .y(output_10_750));
wire output_12_750, output_12_15, output_11_750;
mixer gate_output_11_750(.a(output_12_750), .b(output_12_15), .y(output_11_750));
wire output_13_750, output_13_15, output_12_750;
mixer gate_output_12_750(.a(output_13_750), .b(output_13_15), .y(output_12_750));
wire output_14_750, output_14_15, output_13_750;
mixer gate_output_13_750(.a(output_14_750), .b(output_14_15), .y(output_13_750));
wire output_15_750, output_15_15, output_14_750;
mixer gate_output_14_750(.a(output_15_750), .b(output_15_15), .y(output_14_750));
wire output_16_750, output_16_15, output_15_750;
mixer gate_output_15_750(.a(output_16_750), .b(output_16_15), .y(output_15_750));
wire output_1_751, output_1_0, output_0_751;
mixer gate_output_0_751(.a(output_1_751), .b(output_1_0), .y(output_0_751));
wire output_2_751, output_2_0, output_1_751;
mixer gate_output_1_751(.a(output_2_751), .b(output_2_0), .y(output_1_751));
wire output_3_751, output_3_0, output_2_751;
mixer gate_output_2_751(.a(output_3_751), .b(output_3_0), .y(output_2_751));
wire output_4_751, output_4_0, output_3_751;
mixer gate_output_3_751(.a(output_4_751), .b(output_4_0), .y(output_3_751));
wire output_5_751, output_5_0, output_4_751;
mixer gate_output_4_751(.a(output_5_751), .b(output_5_0), .y(output_4_751));
wire output_6_751, output_6_0, output_5_751;
mixer gate_output_5_751(.a(output_6_751), .b(output_6_0), .y(output_5_751));
wire output_7_751, output_7_0, output_6_751;
mixer gate_output_6_751(.a(output_7_751), .b(output_7_0), .y(output_6_751));
wire output_8_751, output_8_0, output_7_751;
mixer gate_output_7_751(.a(output_8_751), .b(output_8_0), .y(output_7_751));
wire output_9_751, output_9_0, output_8_751;
mixer gate_output_8_751(.a(output_9_751), .b(output_9_0), .y(output_8_751));
wire output_10_751, output_10_0, output_9_751;
mixer gate_output_9_751(.a(output_10_751), .b(output_10_0), .y(output_9_751));
wire output_11_751, output_11_0, output_10_751;
mixer gate_output_10_751(.a(output_11_751), .b(output_11_0), .y(output_10_751));
wire output_12_751, output_12_0, output_11_751;
mixer gate_output_11_751(.a(output_12_751), .b(output_12_0), .y(output_11_751));
wire output_13_751, output_13_0, output_12_751;
mixer gate_output_12_751(.a(output_13_751), .b(output_13_0), .y(output_12_751));
wire output_14_751, output_14_0, output_13_751;
mixer gate_output_13_751(.a(output_14_751), .b(output_14_0), .y(output_13_751));
wire output_15_751, output_15_0, output_14_751;
mixer gate_output_14_751(.a(output_15_751), .b(output_15_0), .y(output_14_751));
wire output_16_751, output_16_0, output_15_751;
mixer gate_output_15_751(.a(output_16_751), .b(output_16_0), .y(output_15_751));
wire output_1_752, output_1_1, output_0_752;
mixer gate_output_0_752(.a(output_1_752), .b(output_1_1), .y(output_0_752));
wire output_2_752, output_2_1, output_1_752;
mixer gate_output_1_752(.a(output_2_752), .b(output_2_1), .y(output_1_752));
wire output_3_752, output_3_1, output_2_752;
mixer gate_output_2_752(.a(output_3_752), .b(output_3_1), .y(output_2_752));
wire output_4_752, output_4_1, output_3_752;
mixer gate_output_3_752(.a(output_4_752), .b(output_4_1), .y(output_3_752));
wire output_5_752, output_5_1, output_4_752;
mixer gate_output_4_752(.a(output_5_752), .b(output_5_1), .y(output_4_752));
wire output_6_752, output_6_1, output_5_752;
mixer gate_output_5_752(.a(output_6_752), .b(output_6_1), .y(output_5_752));
wire output_7_752, output_7_1, output_6_752;
mixer gate_output_6_752(.a(output_7_752), .b(output_7_1), .y(output_6_752));
wire output_8_752, output_8_1, output_7_752;
mixer gate_output_7_752(.a(output_8_752), .b(output_8_1), .y(output_7_752));
wire output_9_752, output_9_1, output_8_752;
mixer gate_output_8_752(.a(output_9_752), .b(output_9_1), .y(output_8_752));
wire output_10_752, output_10_1, output_9_752;
mixer gate_output_9_752(.a(output_10_752), .b(output_10_1), .y(output_9_752));
wire output_11_752, output_11_1, output_10_752;
mixer gate_output_10_752(.a(output_11_752), .b(output_11_1), .y(output_10_752));
wire output_12_752, output_12_1, output_11_752;
mixer gate_output_11_752(.a(output_12_752), .b(output_12_1), .y(output_11_752));
wire output_13_752, output_13_1, output_12_752;
mixer gate_output_12_752(.a(output_13_752), .b(output_13_1), .y(output_12_752));
wire output_14_752, output_14_1, output_13_752;
mixer gate_output_13_752(.a(output_14_752), .b(output_14_1), .y(output_13_752));
wire output_15_752, output_15_1, output_14_752;
mixer gate_output_14_752(.a(output_15_752), .b(output_15_1), .y(output_14_752));
wire output_16_752, output_16_1, output_15_752;
mixer gate_output_15_752(.a(output_16_752), .b(output_16_1), .y(output_15_752));
wire output_1_753, output_1_2, output_0_753;
mixer gate_output_0_753(.a(output_1_753), .b(output_1_2), .y(output_0_753));
wire output_2_753, output_2_2, output_1_753;
mixer gate_output_1_753(.a(output_2_753), .b(output_2_2), .y(output_1_753));
wire output_3_753, output_3_2, output_2_753;
mixer gate_output_2_753(.a(output_3_753), .b(output_3_2), .y(output_2_753));
wire output_4_753, output_4_2, output_3_753;
mixer gate_output_3_753(.a(output_4_753), .b(output_4_2), .y(output_3_753));
wire output_5_753, output_5_2, output_4_753;
mixer gate_output_4_753(.a(output_5_753), .b(output_5_2), .y(output_4_753));
wire output_6_753, output_6_2, output_5_753;
mixer gate_output_5_753(.a(output_6_753), .b(output_6_2), .y(output_5_753));
wire output_7_753, output_7_2, output_6_753;
mixer gate_output_6_753(.a(output_7_753), .b(output_7_2), .y(output_6_753));
wire output_8_753, output_8_2, output_7_753;
mixer gate_output_7_753(.a(output_8_753), .b(output_8_2), .y(output_7_753));
wire output_9_753, output_9_2, output_8_753;
mixer gate_output_8_753(.a(output_9_753), .b(output_9_2), .y(output_8_753));
wire output_10_753, output_10_2, output_9_753;
mixer gate_output_9_753(.a(output_10_753), .b(output_10_2), .y(output_9_753));
wire output_11_753, output_11_2, output_10_753;
mixer gate_output_10_753(.a(output_11_753), .b(output_11_2), .y(output_10_753));
wire output_12_753, output_12_2, output_11_753;
mixer gate_output_11_753(.a(output_12_753), .b(output_12_2), .y(output_11_753));
wire output_13_753, output_13_2, output_12_753;
mixer gate_output_12_753(.a(output_13_753), .b(output_13_2), .y(output_12_753));
wire output_14_753, output_14_2, output_13_753;
mixer gate_output_13_753(.a(output_14_753), .b(output_14_2), .y(output_13_753));
wire output_15_753, output_15_2, output_14_753;
mixer gate_output_14_753(.a(output_15_753), .b(output_15_2), .y(output_14_753));
wire output_16_753, output_16_2, output_15_753;
mixer gate_output_15_753(.a(output_16_753), .b(output_16_2), .y(output_15_753));
wire output_1_754, output_1_3, output_0_754;
mixer gate_output_0_754(.a(output_1_754), .b(output_1_3), .y(output_0_754));
wire output_2_754, output_2_3, output_1_754;
mixer gate_output_1_754(.a(output_2_754), .b(output_2_3), .y(output_1_754));
wire output_3_754, output_3_3, output_2_754;
mixer gate_output_2_754(.a(output_3_754), .b(output_3_3), .y(output_2_754));
wire output_4_754, output_4_3, output_3_754;
mixer gate_output_3_754(.a(output_4_754), .b(output_4_3), .y(output_3_754));
wire output_5_754, output_5_3, output_4_754;
mixer gate_output_4_754(.a(output_5_754), .b(output_5_3), .y(output_4_754));
wire output_6_754, output_6_3, output_5_754;
mixer gate_output_5_754(.a(output_6_754), .b(output_6_3), .y(output_5_754));
wire output_7_754, output_7_3, output_6_754;
mixer gate_output_6_754(.a(output_7_754), .b(output_7_3), .y(output_6_754));
wire output_8_754, output_8_3, output_7_754;
mixer gate_output_7_754(.a(output_8_754), .b(output_8_3), .y(output_7_754));
wire output_9_754, output_9_3, output_8_754;
mixer gate_output_8_754(.a(output_9_754), .b(output_9_3), .y(output_8_754));
wire output_10_754, output_10_3, output_9_754;
mixer gate_output_9_754(.a(output_10_754), .b(output_10_3), .y(output_9_754));
wire output_11_754, output_11_3, output_10_754;
mixer gate_output_10_754(.a(output_11_754), .b(output_11_3), .y(output_10_754));
wire output_12_754, output_12_3, output_11_754;
mixer gate_output_11_754(.a(output_12_754), .b(output_12_3), .y(output_11_754));
wire output_13_754, output_13_3, output_12_754;
mixer gate_output_12_754(.a(output_13_754), .b(output_13_3), .y(output_12_754));
wire output_14_754, output_14_3, output_13_754;
mixer gate_output_13_754(.a(output_14_754), .b(output_14_3), .y(output_13_754));
wire output_15_754, output_15_3, output_14_754;
mixer gate_output_14_754(.a(output_15_754), .b(output_15_3), .y(output_14_754));
wire output_16_754, output_16_3, output_15_754;
mixer gate_output_15_754(.a(output_16_754), .b(output_16_3), .y(output_15_754));
wire output_1_755, output_1_4, output_0_755;
mixer gate_output_0_755(.a(output_1_755), .b(output_1_4), .y(output_0_755));
wire output_2_755, output_2_4, output_1_755;
mixer gate_output_1_755(.a(output_2_755), .b(output_2_4), .y(output_1_755));
wire output_3_755, output_3_4, output_2_755;
mixer gate_output_2_755(.a(output_3_755), .b(output_3_4), .y(output_2_755));
wire output_4_755, output_4_4, output_3_755;
mixer gate_output_3_755(.a(output_4_755), .b(output_4_4), .y(output_3_755));
wire output_5_755, output_5_4, output_4_755;
mixer gate_output_4_755(.a(output_5_755), .b(output_5_4), .y(output_4_755));
wire output_6_755, output_6_4, output_5_755;
mixer gate_output_5_755(.a(output_6_755), .b(output_6_4), .y(output_5_755));
wire output_7_755, output_7_4, output_6_755;
mixer gate_output_6_755(.a(output_7_755), .b(output_7_4), .y(output_6_755));
wire output_8_755, output_8_4, output_7_755;
mixer gate_output_7_755(.a(output_8_755), .b(output_8_4), .y(output_7_755));
wire output_9_755, output_9_4, output_8_755;
mixer gate_output_8_755(.a(output_9_755), .b(output_9_4), .y(output_8_755));
wire output_10_755, output_10_4, output_9_755;
mixer gate_output_9_755(.a(output_10_755), .b(output_10_4), .y(output_9_755));
wire output_11_755, output_11_4, output_10_755;
mixer gate_output_10_755(.a(output_11_755), .b(output_11_4), .y(output_10_755));
wire output_12_755, output_12_4, output_11_755;
mixer gate_output_11_755(.a(output_12_755), .b(output_12_4), .y(output_11_755));
wire output_13_755, output_13_4, output_12_755;
mixer gate_output_12_755(.a(output_13_755), .b(output_13_4), .y(output_12_755));
wire output_14_755, output_14_4, output_13_755;
mixer gate_output_13_755(.a(output_14_755), .b(output_14_4), .y(output_13_755));
wire output_15_755, output_15_4, output_14_755;
mixer gate_output_14_755(.a(output_15_755), .b(output_15_4), .y(output_14_755));
wire output_16_755, output_16_4, output_15_755;
mixer gate_output_15_755(.a(output_16_755), .b(output_16_4), .y(output_15_755));
wire output_1_756, output_1_5, output_0_756;
mixer gate_output_0_756(.a(output_1_756), .b(output_1_5), .y(output_0_756));
wire output_2_756, output_2_5, output_1_756;
mixer gate_output_1_756(.a(output_2_756), .b(output_2_5), .y(output_1_756));
wire output_3_756, output_3_5, output_2_756;
mixer gate_output_2_756(.a(output_3_756), .b(output_3_5), .y(output_2_756));
wire output_4_756, output_4_5, output_3_756;
mixer gate_output_3_756(.a(output_4_756), .b(output_4_5), .y(output_3_756));
wire output_5_756, output_5_5, output_4_756;
mixer gate_output_4_756(.a(output_5_756), .b(output_5_5), .y(output_4_756));
wire output_6_756, output_6_5, output_5_756;
mixer gate_output_5_756(.a(output_6_756), .b(output_6_5), .y(output_5_756));
wire output_7_756, output_7_5, output_6_756;
mixer gate_output_6_756(.a(output_7_756), .b(output_7_5), .y(output_6_756));
wire output_8_756, output_8_5, output_7_756;
mixer gate_output_7_756(.a(output_8_756), .b(output_8_5), .y(output_7_756));
wire output_9_756, output_9_5, output_8_756;
mixer gate_output_8_756(.a(output_9_756), .b(output_9_5), .y(output_8_756));
wire output_10_756, output_10_5, output_9_756;
mixer gate_output_9_756(.a(output_10_756), .b(output_10_5), .y(output_9_756));
wire output_11_756, output_11_5, output_10_756;
mixer gate_output_10_756(.a(output_11_756), .b(output_11_5), .y(output_10_756));
wire output_12_756, output_12_5, output_11_756;
mixer gate_output_11_756(.a(output_12_756), .b(output_12_5), .y(output_11_756));
wire output_13_756, output_13_5, output_12_756;
mixer gate_output_12_756(.a(output_13_756), .b(output_13_5), .y(output_12_756));
wire output_14_756, output_14_5, output_13_756;
mixer gate_output_13_756(.a(output_14_756), .b(output_14_5), .y(output_13_756));
wire output_15_756, output_15_5, output_14_756;
mixer gate_output_14_756(.a(output_15_756), .b(output_15_5), .y(output_14_756));
wire output_16_756, output_16_5, output_15_756;
mixer gate_output_15_756(.a(output_16_756), .b(output_16_5), .y(output_15_756));
wire output_1_757, output_1_6, output_0_757;
mixer gate_output_0_757(.a(output_1_757), .b(output_1_6), .y(output_0_757));
wire output_2_757, output_2_6, output_1_757;
mixer gate_output_1_757(.a(output_2_757), .b(output_2_6), .y(output_1_757));
wire output_3_757, output_3_6, output_2_757;
mixer gate_output_2_757(.a(output_3_757), .b(output_3_6), .y(output_2_757));
wire output_4_757, output_4_6, output_3_757;
mixer gate_output_3_757(.a(output_4_757), .b(output_4_6), .y(output_3_757));
wire output_5_757, output_5_6, output_4_757;
mixer gate_output_4_757(.a(output_5_757), .b(output_5_6), .y(output_4_757));
wire output_6_757, output_6_6, output_5_757;
mixer gate_output_5_757(.a(output_6_757), .b(output_6_6), .y(output_5_757));
wire output_7_757, output_7_6, output_6_757;
mixer gate_output_6_757(.a(output_7_757), .b(output_7_6), .y(output_6_757));
wire output_8_757, output_8_6, output_7_757;
mixer gate_output_7_757(.a(output_8_757), .b(output_8_6), .y(output_7_757));
wire output_9_757, output_9_6, output_8_757;
mixer gate_output_8_757(.a(output_9_757), .b(output_9_6), .y(output_8_757));
wire output_10_757, output_10_6, output_9_757;
mixer gate_output_9_757(.a(output_10_757), .b(output_10_6), .y(output_9_757));
wire output_11_757, output_11_6, output_10_757;
mixer gate_output_10_757(.a(output_11_757), .b(output_11_6), .y(output_10_757));
wire output_12_757, output_12_6, output_11_757;
mixer gate_output_11_757(.a(output_12_757), .b(output_12_6), .y(output_11_757));
wire output_13_757, output_13_6, output_12_757;
mixer gate_output_12_757(.a(output_13_757), .b(output_13_6), .y(output_12_757));
wire output_14_757, output_14_6, output_13_757;
mixer gate_output_13_757(.a(output_14_757), .b(output_14_6), .y(output_13_757));
wire output_15_757, output_15_6, output_14_757;
mixer gate_output_14_757(.a(output_15_757), .b(output_15_6), .y(output_14_757));
wire output_16_757, output_16_6, output_15_757;
mixer gate_output_15_757(.a(output_16_757), .b(output_16_6), .y(output_15_757));
wire output_1_758, output_1_7, output_0_758;
mixer gate_output_0_758(.a(output_1_758), .b(output_1_7), .y(output_0_758));
wire output_2_758, output_2_7, output_1_758;
mixer gate_output_1_758(.a(output_2_758), .b(output_2_7), .y(output_1_758));
wire output_3_758, output_3_7, output_2_758;
mixer gate_output_2_758(.a(output_3_758), .b(output_3_7), .y(output_2_758));
wire output_4_758, output_4_7, output_3_758;
mixer gate_output_3_758(.a(output_4_758), .b(output_4_7), .y(output_3_758));
wire output_5_758, output_5_7, output_4_758;
mixer gate_output_4_758(.a(output_5_758), .b(output_5_7), .y(output_4_758));
wire output_6_758, output_6_7, output_5_758;
mixer gate_output_5_758(.a(output_6_758), .b(output_6_7), .y(output_5_758));
wire output_7_758, output_7_7, output_6_758;
mixer gate_output_6_758(.a(output_7_758), .b(output_7_7), .y(output_6_758));
wire output_8_758, output_8_7, output_7_758;
mixer gate_output_7_758(.a(output_8_758), .b(output_8_7), .y(output_7_758));
wire output_9_758, output_9_7, output_8_758;
mixer gate_output_8_758(.a(output_9_758), .b(output_9_7), .y(output_8_758));
wire output_10_758, output_10_7, output_9_758;
mixer gate_output_9_758(.a(output_10_758), .b(output_10_7), .y(output_9_758));
wire output_11_758, output_11_7, output_10_758;
mixer gate_output_10_758(.a(output_11_758), .b(output_11_7), .y(output_10_758));
wire output_12_758, output_12_7, output_11_758;
mixer gate_output_11_758(.a(output_12_758), .b(output_12_7), .y(output_11_758));
wire output_13_758, output_13_7, output_12_758;
mixer gate_output_12_758(.a(output_13_758), .b(output_13_7), .y(output_12_758));
wire output_14_758, output_14_7, output_13_758;
mixer gate_output_13_758(.a(output_14_758), .b(output_14_7), .y(output_13_758));
wire output_15_758, output_15_7, output_14_758;
mixer gate_output_14_758(.a(output_15_758), .b(output_15_7), .y(output_14_758));
wire output_16_758, output_16_7, output_15_758;
mixer gate_output_15_758(.a(output_16_758), .b(output_16_7), .y(output_15_758));
wire output_1_759, output_1_8, output_0_759;
mixer gate_output_0_759(.a(output_1_759), .b(output_1_8), .y(output_0_759));
wire output_2_759, output_2_8, output_1_759;
mixer gate_output_1_759(.a(output_2_759), .b(output_2_8), .y(output_1_759));
wire output_3_759, output_3_8, output_2_759;
mixer gate_output_2_759(.a(output_3_759), .b(output_3_8), .y(output_2_759));
wire output_4_759, output_4_8, output_3_759;
mixer gate_output_3_759(.a(output_4_759), .b(output_4_8), .y(output_3_759));
wire output_5_759, output_5_8, output_4_759;
mixer gate_output_4_759(.a(output_5_759), .b(output_5_8), .y(output_4_759));
wire output_6_759, output_6_8, output_5_759;
mixer gate_output_5_759(.a(output_6_759), .b(output_6_8), .y(output_5_759));
wire output_7_759, output_7_8, output_6_759;
mixer gate_output_6_759(.a(output_7_759), .b(output_7_8), .y(output_6_759));
wire output_8_759, output_8_8, output_7_759;
mixer gate_output_7_759(.a(output_8_759), .b(output_8_8), .y(output_7_759));
wire output_9_759, output_9_8, output_8_759;
mixer gate_output_8_759(.a(output_9_759), .b(output_9_8), .y(output_8_759));
wire output_10_759, output_10_8, output_9_759;
mixer gate_output_9_759(.a(output_10_759), .b(output_10_8), .y(output_9_759));
wire output_11_759, output_11_8, output_10_759;
mixer gate_output_10_759(.a(output_11_759), .b(output_11_8), .y(output_10_759));
wire output_12_759, output_12_8, output_11_759;
mixer gate_output_11_759(.a(output_12_759), .b(output_12_8), .y(output_11_759));
wire output_13_759, output_13_8, output_12_759;
mixer gate_output_12_759(.a(output_13_759), .b(output_13_8), .y(output_12_759));
wire output_14_759, output_14_8, output_13_759;
mixer gate_output_13_759(.a(output_14_759), .b(output_14_8), .y(output_13_759));
wire output_15_759, output_15_8, output_14_759;
mixer gate_output_14_759(.a(output_15_759), .b(output_15_8), .y(output_14_759));
wire output_16_759, output_16_8, output_15_759;
mixer gate_output_15_759(.a(output_16_759), .b(output_16_8), .y(output_15_759));
wire output_1_760, output_1_9, output_0_760;
mixer gate_output_0_760(.a(output_1_760), .b(output_1_9), .y(output_0_760));
wire output_2_760, output_2_9, output_1_760;
mixer gate_output_1_760(.a(output_2_760), .b(output_2_9), .y(output_1_760));
wire output_3_760, output_3_9, output_2_760;
mixer gate_output_2_760(.a(output_3_760), .b(output_3_9), .y(output_2_760));
wire output_4_760, output_4_9, output_3_760;
mixer gate_output_3_760(.a(output_4_760), .b(output_4_9), .y(output_3_760));
wire output_5_760, output_5_9, output_4_760;
mixer gate_output_4_760(.a(output_5_760), .b(output_5_9), .y(output_4_760));
wire output_6_760, output_6_9, output_5_760;
mixer gate_output_5_760(.a(output_6_760), .b(output_6_9), .y(output_5_760));
wire output_7_760, output_7_9, output_6_760;
mixer gate_output_6_760(.a(output_7_760), .b(output_7_9), .y(output_6_760));
wire output_8_760, output_8_9, output_7_760;
mixer gate_output_7_760(.a(output_8_760), .b(output_8_9), .y(output_7_760));
wire output_9_760, output_9_9, output_8_760;
mixer gate_output_8_760(.a(output_9_760), .b(output_9_9), .y(output_8_760));
wire output_10_760, output_10_9, output_9_760;
mixer gate_output_9_760(.a(output_10_760), .b(output_10_9), .y(output_9_760));
wire output_11_760, output_11_9, output_10_760;
mixer gate_output_10_760(.a(output_11_760), .b(output_11_9), .y(output_10_760));
wire output_12_760, output_12_9, output_11_760;
mixer gate_output_11_760(.a(output_12_760), .b(output_12_9), .y(output_11_760));
wire output_13_760, output_13_9, output_12_760;
mixer gate_output_12_760(.a(output_13_760), .b(output_13_9), .y(output_12_760));
wire output_14_760, output_14_9, output_13_760;
mixer gate_output_13_760(.a(output_14_760), .b(output_14_9), .y(output_13_760));
wire output_15_760, output_15_9, output_14_760;
mixer gate_output_14_760(.a(output_15_760), .b(output_15_9), .y(output_14_760));
wire output_16_760, output_16_9, output_15_760;
mixer gate_output_15_760(.a(output_16_760), .b(output_16_9), .y(output_15_760));
wire output_1_761, output_1_10, output_0_761;
mixer gate_output_0_761(.a(output_1_761), .b(output_1_10), .y(output_0_761));
wire output_2_761, output_2_10, output_1_761;
mixer gate_output_1_761(.a(output_2_761), .b(output_2_10), .y(output_1_761));
wire output_3_761, output_3_10, output_2_761;
mixer gate_output_2_761(.a(output_3_761), .b(output_3_10), .y(output_2_761));
wire output_4_761, output_4_10, output_3_761;
mixer gate_output_3_761(.a(output_4_761), .b(output_4_10), .y(output_3_761));
wire output_5_761, output_5_10, output_4_761;
mixer gate_output_4_761(.a(output_5_761), .b(output_5_10), .y(output_4_761));
wire output_6_761, output_6_10, output_5_761;
mixer gate_output_5_761(.a(output_6_761), .b(output_6_10), .y(output_5_761));
wire output_7_761, output_7_10, output_6_761;
mixer gate_output_6_761(.a(output_7_761), .b(output_7_10), .y(output_6_761));
wire output_8_761, output_8_10, output_7_761;
mixer gate_output_7_761(.a(output_8_761), .b(output_8_10), .y(output_7_761));
wire output_9_761, output_9_10, output_8_761;
mixer gate_output_8_761(.a(output_9_761), .b(output_9_10), .y(output_8_761));
wire output_10_761, output_10_10, output_9_761;
mixer gate_output_9_761(.a(output_10_761), .b(output_10_10), .y(output_9_761));
wire output_11_761, output_11_10, output_10_761;
mixer gate_output_10_761(.a(output_11_761), .b(output_11_10), .y(output_10_761));
wire output_12_761, output_12_10, output_11_761;
mixer gate_output_11_761(.a(output_12_761), .b(output_12_10), .y(output_11_761));
wire output_13_761, output_13_10, output_12_761;
mixer gate_output_12_761(.a(output_13_761), .b(output_13_10), .y(output_12_761));
wire output_14_761, output_14_10, output_13_761;
mixer gate_output_13_761(.a(output_14_761), .b(output_14_10), .y(output_13_761));
wire output_15_761, output_15_10, output_14_761;
mixer gate_output_14_761(.a(output_15_761), .b(output_15_10), .y(output_14_761));
wire output_16_761, output_16_10, output_15_761;
mixer gate_output_15_761(.a(output_16_761), .b(output_16_10), .y(output_15_761));
wire output_1_762, output_1_11, output_0_762;
mixer gate_output_0_762(.a(output_1_762), .b(output_1_11), .y(output_0_762));
wire output_2_762, output_2_11, output_1_762;
mixer gate_output_1_762(.a(output_2_762), .b(output_2_11), .y(output_1_762));
wire output_3_762, output_3_11, output_2_762;
mixer gate_output_2_762(.a(output_3_762), .b(output_3_11), .y(output_2_762));
wire output_4_762, output_4_11, output_3_762;
mixer gate_output_3_762(.a(output_4_762), .b(output_4_11), .y(output_3_762));
wire output_5_762, output_5_11, output_4_762;
mixer gate_output_4_762(.a(output_5_762), .b(output_5_11), .y(output_4_762));
wire output_6_762, output_6_11, output_5_762;
mixer gate_output_5_762(.a(output_6_762), .b(output_6_11), .y(output_5_762));
wire output_7_762, output_7_11, output_6_762;
mixer gate_output_6_762(.a(output_7_762), .b(output_7_11), .y(output_6_762));
wire output_8_762, output_8_11, output_7_762;
mixer gate_output_7_762(.a(output_8_762), .b(output_8_11), .y(output_7_762));
wire output_9_762, output_9_11, output_8_762;
mixer gate_output_8_762(.a(output_9_762), .b(output_9_11), .y(output_8_762));
wire output_10_762, output_10_11, output_9_762;
mixer gate_output_9_762(.a(output_10_762), .b(output_10_11), .y(output_9_762));
wire output_11_762, output_11_11, output_10_762;
mixer gate_output_10_762(.a(output_11_762), .b(output_11_11), .y(output_10_762));
wire output_12_762, output_12_11, output_11_762;
mixer gate_output_11_762(.a(output_12_762), .b(output_12_11), .y(output_11_762));
wire output_13_762, output_13_11, output_12_762;
mixer gate_output_12_762(.a(output_13_762), .b(output_13_11), .y(output_12_762));
wire output_14_762, output_14_11, output_13_762;
mixer gate_output_13_762(.a(output_14_762), .b(output_14_11), .y(output_13_762));
wire output_15_762, output_15_11, output_14_762;
mixer gate_output_14_762(.a(output_15_762), .b(output_15_11), .y(output_14_762));
wire output_16_762, output_16_11, output_15_762;
mixer gate_output_15_762(.a(output_16_762), .b(output_16_11), .y(output_15_762));
wire output_1_763, output_1_12, output_0_763;
mixer gate_output_0_763(.a(output_1_763), .b(output_1_12), .y(output_0_763));
wire output_2_763, output_2_12, output_1_763;
mixer gate_output_1_763(.a(output_2_763), .b(output_2_12), .y(output_1_763));
wire output_3_763, output_3_12, output_2_763;
mixer gate_output_2_763(.a(output_3_763), .b(output_3_12), .y(output_2_763));
wire output_4_763, output_4_12, output_3_763;
mixer gate_output_3_763(.a(output_4_763), .b(output_4_12), .y(output_3_763));
wire output_5_763, output_5_12, output_4_763;
mixer gate_output_4_763(.a(output_5_763), .b(output_5_12), .y(output_4_763));
wire output_6_763, output_6_12, output_5_763;
mixer gate_output_5_763(.a(output_6_763), .b(output_6_12), .y(output_5_763));
wire output_7_763, output_7_12, output_6_763;
mixer gate_output_6_763(.a(output_7_763), .b(output_7_12), .y(output_6_763));
wire output_8_763, output_8_12, output_7_763;
mixer gate_output_7_763(.a(output_8_763), .b(output_8_12), .y(output_7_763));
wire output_9_763, output_9_12, output_8_763;
mixer gate_output_8_763(.a(output_9_763), .b(output_9_12), .y(output_8_763));
wire output_10_763, output_10_12, output_9_763;
mixer gate_output_9_763(.a(output_10_763), .b(output_10_12), .y(output_9_763));
wire output_11_763, output_11_12, output_10_763;
mixer gate_output_10_763(.a(output_11_763), .b(output_11_12), .y(output_10_763));
wire output_12_763, output_12_12, output_11_763;
mixer gate_output_11_763(.a(output_12_763), .b(output_12_12), .y(output_11_763));
wire output_13_763, output_13_12, output_12_763;
mixer gate_output_12_763(.a(output_13_763), .b(output_13_12), .y(output_12_763));
wire output_14_763, output_14_12, output_13_763;
mixer gate_output_13_763(.a(output_14_763), .b(output_14_12), .y(output_13_763));
wire output_15_763, output_15_12, output_14_763;
mixer gate_output_14_763(.a(output_15_763), .b(output_15_12), .y(output_14_763));
wire output_16_763, output_16_12, output_15_763;
mixer gate_output_15_763(.a(output_16_763), .b(output_16_12), .y(output_15_763));
wire output_1_764, output_1_13, output_0_764;
mixer gate_output_0_764(.a(output_1_764), .b(output_1_13), .y(output_0_764));
wire output_2_764, output_2_13, output_1_764;
mixer gate_output_1_764(.a(output_2_764), .b(output_2_13), .y(output_1_764));
wire output_3_764, output_3_13, output_2_764;
mixer gate_output_2_764(.a(output_3_764), .b(output_3_13), .y(output_2_764));
wire output_4_764, output_4_13, output_3_764;
mixer gate_output_3_764(.a(output_4_764), .b(output_4_13), .y(output_3_764));
wire output_5_764, output_5_13, output_4_764;
mixer gate_output_4_764(.a(output_5_764), .b(output_5_13), .y(output_4_764));
wire output_6_764, output_6_13, output_5_764;
mixer gate_output_5_764(.a(output_6_764), .b(output_6_13), .y(output_5_764));
wire output_7_764, output_7_13, output_6_764;
mixer gate_output_6_764(.a(output_7_764), .b(output_7_13), .y(output_6_764));
wire output_8_764, output_8_13, output_7_764;
mixer gate_output_7_764(.a(output_8_764), .b(output_8_13), .y(output_7_764));
wire output_9_764, output_9_13, output_8_764;
mixer gate_output_8_764(.a(output_9_764), .b(output_9_13), .y(output_8_764));
wire output_10_764, output_10_13, output_9_764;
mixer gate_output_9_764(.a(output_10_764), .b(output_10_13), .y(output_9_764));
wire output_11_764, output_11_13, output_10_764;
mixer gate_output_10_764(.a(output_11_764), .b(output_11_13), .y(output_10_764));
wire output_12_764, output_12_13, output_11_764;
mixer gate_output_11_764(.a(output_12_764), .b(output_12_13), .y(output_11_764));
wire output_13_764, output_13_13, output_12_764;
mixer gate_output_12_764(.a(output_13_764), .b(output_13_13), .y(output_12_764));
wire output_14_764, output_14_13, output_13_764;
mixer gate_output_13_764(.a(output_14_764), .b(output_14_13), .y(output_13_764));
wire output_15_764, output_15_13, output_14_764;
mixer gate_output_14_764(.a(output_15_764), .b(output_15_13), .y(output_14_764));
wire output_16_764, output_16_13, output_15_764;
mixer gate_output_15_764(.a(output_16_764), .b(output_16_13), .y(output_15_764));
wire output_1_765, output_1_14, output_0_765;
mixer gate_output_0_765(.a(output_1_765), .b(output_1_14), .y(output_0_765));
wire output_2_765, output_2_14, output_1_765;
mixer gate_output_1_765(.a(output_2_765), .b(output_2_14), .y(output_1_765));
wire output_3_765, output_3_14, output_2_765;
mixer gate_output_2_765(.a(output_3_765), .b(output_3_14), .y(output_2_765));
wire output_4_765, output_4_14, output_3_765;
mixer gate_output_3_765(.a(output_4_765), .b(output_4_14), .y(output_3_765));
wire output_5_765, output_5_14, output_4_765;
mixer gate_output_4_765(.a(output_5_765), .b(output_5_14), .y(output_4_765));
wire output_6_765, output_6_14, output_5_765;
mixer gate_output_5_765(.a(output_6_765), .b(output_6_14), .y(output_5_765));
wire output_7_765, output_7_14, output_6_765;
mixer gate_output_6_765(.a(output_7_765), .b(output_7_14), .y(output_6_765));
wire output_8_765, output_8_14, output_7_765;
mixer gate_output_7_765(.a(output_8_765), .b(output_8_14), .y(output_7_765));
wire output_9_765, output_9_14, output_8_765;
mixer gate_output_8_765(.a(output_9_765), .b(output_9_14), .y(output_8_765));
wire output_10_765, output_10_14, output_9_765;
mixer gate_output_9_765(.a(output_10_765), .b(output_10_14), .y(output_9_765));
wire output_11_765, output_11_14, output_10_765;
mixer gate_output_10_765(.a(output_11_765), .b(output_11_14), .y(output_10_765));
wire output_12_765, output_12_14, output_11_765;
mixer gate_output_11_765(.a(output_12_765), .b(output_12_14), .y(output_11_765));
wire output_13_765, output_13_14, output_12_765;
mixer gate_output_12_765(.a(output_13_765), .b(output_13_14), .y(output_12_765));
wire output_14_765, output_14_14, output_13_765;
mixer gate_output_13_765(.a(output_14_765), .b(output_14_14), .y(output_13_765));
wire output_15_765, output_15_14, output_14_765;
mixer gate_output_14_765(.a(output_15_765), .b(output_15_14), .y(output_14_765));
wire output_16_765, output_16_14, output_15_765;
mixer gate_output_15_765(.a(output_16_765), .b(output_16_14), .y(output_15_765));
wire output_1_766, output_1_15, output_0_766;
mixer gate_output_0_766(.a(output_1_766), .b(output_1_15), .y(output_0_766));
wire output_2_766, output_2_15, output_1_766;
mixer gate_output_1_766(.a(output_2_766), .b(output_2_15), .y(output_1_766));
wire output_3_766, output_3_15, output_2_766;
mixer gate_output_2_766(.a(output_3_766), .b(output_3_15), .y(output_2_766));
wire output_4_766, output_4_15, output_3_766;
mixer gate_output_3_766(.a(output_4_766), .b(output_4_15), .y(output_3_766));
wire output_5_766, output_5_15, output_4_766;
mixer gate_output_4_766(.a(output_5_766), .b(output_5_15), .y(output_4_766));
wire output_6_766, output_6_15, output_5_766;
mixer gate_output_5_766(.a(output_6_766), .b(output_6_15), .y(output_5_766));
wire output_7_766, output_7_15, output_6_766;
mixer gate_output_6_766(.a(output_7_766), .b(output_7_15), .y(output_6_766));
wire output_8_766, output_8_15, output_7_766;
mixer gate_output_7_766(.a(output_8_766), .b(output_8_15), .y(output_7_766));
wire output_9_766, output_9_15, output_8_766;
mixer gate_output_8_766(.a(output_9_766), .b(output_9_15), .y(output_8_766));
wire output_10_766, output_10_15, output_9_766;
mixer gate_output_9_766(.a(output_10_766), .b(output_10_15), .y(output_9_766));
wire output_11_766, output_11_15, output_10_766;
mixer gate_output_10_766(.a(output_11_766), .b(output_11_15), .y(output_10_766));
wire output_12_766, output_12_15, output_11_766;
mixer gate_output_11_766(.a(output_12_766), .b(output_12_15), .y(output_11_766));
wire output_13_766, output_13_15, output_12_766;
mixer gate_output_12_766(.a(output_13_766), .b(output_13_15), .y(output_12_766));
wire output_14_766, output_14_15, output_13_766;
mixer gate_output_13_766(.a(output_14_766), .b(output_14_15), .y(output_13_766));
wire output_15_766, output_15_15, output_14_766;
mixer gate_output_14_766(.a(output_15_766), .b(output_15_15), .y(output_14_766));
wire output_16_766, output_16_15, output_15_766;
mixer gate_output_15_766(.a(output_16_766), .b(output_16_15), .y(output_15_766));
wire output_1_767, output_1_0, output_0_767;
mixer gate_output_0_767(.a(output_1_767), .b(output_1_0), .y(output_0_767));
wire output_2_767, output_2_0, output_1_767;
mixer gate_output_1_767(.a(output_2_767), .b(output_2_0), .y(output_1_767));
wire output_3_767, output_3_0, output_2_767;
mixer gate_output_2_767(.a(output_3_767), .b(output_3_0), .y(output_2_767));
wire output_4_767, output_4_0, output_3_767;
mixer gate_output_3_767(.a(output_4_767), .b(output_4_0), .y(output_3_767));
wire output_5_767, output_5_0, output_4_767;
mixer gate_output_4_767(.a(output_5_767), .b(output_5_0), .y(output_4_767));
wire output_6_767, output_6_0, output_5_767;
mixer gate_output_5_767(.a(output_6_767), .b(output_6_0), .y(output_5_767));
wire output_7_767, output_7_0, output_6_767;
mixer gate_output_6_767(.a(output_7_767), .b(output_7_0), .y(output_6_767));
wire output_8_767, output_8_0, output_7_767;
mixer gate_output_7_767(.a(output_8_767), .b(output_8_0), .y(output_7_767));
wire output_9_767, output_9_0, output_8_767;
mixer gate_output_8_767(.a(output_9_767), .b(output_9_0), .y(output_8_767));
wire output_10_767, output_10_0, output_9_767;
mixer gate_output_9_767(.a(output_10_767), .b(output_10_0), .y(output_9_767));
wire output_11_767, output_11_0, output_10_767;
mixer gate_output_10_767(.a(output_11_767), .b(output_11_0), .y(output_10_767));
wire output_12_767, output_12_0, output_11_767;
mixer gate_output_11_767(.a(output_12_767), .b(output_12_0), .y(output_11_767));
wire output_13_767, output_13_0, output_12_767;
mixer gate_output_12_767(.a(output_13_767), .b(output_13_0), .y(output_12_767));
wire output_14_767, output_14_0, output_13_767;
mixer gate_output_13_767(.a(output_14_767), .b(output_14_0), .y(output_13_767));
wire output_15_767, output_15_0, output_14_767;
mixer gate_output_14_767(.a(output_15_767), .b(output_15_0), .y(output_14_767));
wire output_16_767, output_16_0, output_15_767;
mixer gate_output_15_767(.a(output_16_767), .b(output_16_0), .y(output_15_767));
wire output_1_768, output_1_1, output_0_768;
mixer gate_output_0_768(.a(output_1_768), .b(output_1_1), .y(output_0_768));
wire output_2_768, output_2_1, output_1_768;
mixer gate_output_1_768(.a(output_2_768), .b(output_2_1), .y(output_1_768));
wire output_3_768, output_3_1, output_2_768;
mixer gate_output_2_768(.a(output_3_768), .b(output_3_1), .y(output_2_768));
wire output_4_768, output_4_1, output_3_768;
mixer gate_output_3_768(.a(output_4_768), .b(output_4_1), .y(output_3_768));
wire output_5_768, output_5_1, output_4_768;
mixer gate_output_4_768(.a(output_5_768), .b(output_5_1), .y(output_4_768));
wire output_6_768, output_6_1, output_5_768;
mixer gate_output_5_768(.a(output_6_768), .b(output_6_1), .y(output_5_768));
wire output_7_768, output_7_1, output_6_768;
mixer gate_output_6_768(.a(output_7_768), .b(output_7_1), .y(output_6_768));
wire output_8_768, output_8_1, output_7_768;
mixer gate_output_7_768(.a(output_8_768), .b(output_8_1), .y(output_7_768));
wire output_9_768, output_9_1, output_8_768;
mixer gate_output_8_768(.a(output_9_768), .b(output_9_1), .y(output_8_768));
wire output_10_768, output_10_1, output_9_768;
mixer gate_output_9_768(.a(output_10_768), .b(output_10_1), .y(output_9_768));
wire output_11_768, output_11_1, output_10_768;
mixer gate_output_10_768(.a(output_11_768), .b(output_11_1), .y(output_10_768));
wire output_12_768, output_12_1, output_11_768;
mixer gate_output_11_768(.a(output_12_768), .b(output_12_1), .y(output_11_768));
wire output_13_768, output_13_1, output_12_768;
mixer gate_output_12_768(.a(output_13_768), .b(output_13_1), .y(output_12_768));
wire output_14_768, output_14_1, output_13_768;
mixer gate_output_13_768(.a(output_14_768), .b(output_14_1), .y(output_13_768));
wire output_15_768, output_15_1, output_14_768;
mixer gate_output_14_768(.a(output_15_768), .b(output_15_1), .y(output_14_768));
wire output_16_768, output_16_1, output_15_768;
mixer gate_output_15_768(.a(output_16_768), .b(output_16_1), .y(output_15_768));
wire output_1_769, output_1_2, output_0_769;
mixer gate_output_0_769(.a(output_1_769), .b(output_1_2), .y(output_0_769));
wire output_2_769, output_2_2, output_1_769;
mixer gate_output_1_769(.a(output_2_769), .b(output_2_2), .y(output_1_769));
wire output_3_769, output_3_2, output_2_769;
mixer gate_output_2_769(.a(output_3_769), .b(output_3_2), .y(output_2_769));
wire output_4_769, output_4_2, output_3_769;
mixer gate_output_3_769(.a(output_4_769), .b(output_4_2), .y(output_3_769));
wire output_5_769, output_5_2, output_4_769;
mixer gate_output_4_769(.a(output_5_769), .b(output_5_2), .y(output_4_769));
wire output_6_769, output_6_2, output_5_769;
mixer gate_output_5_769(.a(output_6_769), .b(output_6_2), .y(output_5_769));
wire output_7_769, output_7_2, output_6_769;
mixer gate_output_6_769(.a(output_7_769), .b(output_7_2), .y(output_6_769));
wire output_8_769, output_8_2, output_7_769;
mixer gate_output_7_769(.a(output_8_769), .b(output_8_2), .y(output_7_769));
wire output_9_769, output_9_2, output_8_769;
mixer gate_output_8_769(.a(output_9_769), .b(output_9_2), .y(output_8_769));
wire output_10_769, output_10_2, output_9_769;
mixer gate_output_9_769(.a(output_10_769), .b(output_10_2), .y(output_9_769));
wire output_11_769, output_11_2, output_10_769;
mixer gate_output_10_769(.a(output_11_769), .b(output_11_2), .y(output_10_769));
wire output_12_769, output_12_2, output_11_769;
mixer gate_output_11_769(.a(output_12_769), .b(output_12_2), .y(output_11_769));
wire output_13_769, output_13_2, output_12_769;
mixer gate_output_12_769(.a(output_13_769), .b(output_13_2), .y(output_12_769));
wire output_14_769, output_14_2, output_13_769;
mixer gate_output_13_769(.a(output_14_769), .b(output_14_2), .y(output_13_769));
wire output_15_769, output_15_2, output_14_769;
mixer gate_output_14_769(.a(output_15_769), .b(output_15_2), .y(output_14_769));
wire output_16_769, output_16_2, output_15_769;
mixer gate_output_15_769(.a(output_16_769), .b(output_16_2), .y(output_15_769));
wire output_1_770, output_1_3, output_0_770;
mixer gate_output_0_770(.a(output_1_770), .b(output_1_3), .y(output_0_770));
wire output_2_770, output_2_3, output_1_770;
mixer gate_output_1_770(.a(output_2_770), .b(output_2_3), .y(output_1_770));
wire output_3_770, output_3_3, output_2_770;
mixer gate_output_2_770(.a(output_3_770), .b(output_3_3), .y(output_2_770));
wire output_4_770, output_4_3, output_3_770;
mixer gate_output_3_770(.a(output_4_770), .b(output_4_3), .y(output_3_770));
wire output_5_770, output_5_3, output_4_770;
mixer gate_output_4_770(.a(output_5_770), .b(output_5_3), .y(output_4_770));
wire output_6_770, output_6_3, output_5_770;
mixer gate_output_5_770(.a(output_6_770), .b(output_6_3), .y(output_5_770));
wire output_7_770, output_7_3, output_6_770;
mixer gate_output_6_770(.a(output_7_770), .b(output_7_3), .y(output_6_770));
wire output_8_770, output_8_3, output_7_770;
mixer gate_output_7_770(.a(output_8_770), .b(output_8_3), .y(output_7_770));
wire output_9_770, output_9_3, output_8_770;
mixer gate_output_8_770(.a(output_9_770), .b(output_9_3), .y(output_8_770));
wire output_10_770, output_10_3, output_9_770;
mixer gate_output_9_770(.a(output_10_770), .b(output_10_3), .y(output_9_770));
wire output_11_770, output_11_3, output_10_770;
mixer gate_output_10_770(.a(output_11_770), .b(output_11_3), .y(output_10_770));
wire output_12_770, output_12_3, output_11_770;
mixer gate_output_11_770(.a(output_12_770), .b(output_12_3), .y(output_11_770));
wire output_13_770, output_13_3, output_12_770;
mixer gate_output_12_770(.a(output_13_770), .b(output_13_3), .y(output_12_770));
wire output_14_770, output_14_3, output_13_770;
mixer gate_output_13_770(.a(output_14_770), .b(output_14_3), .y(output_13_770));
wire output_15_770, output_15_3, output_14_770;
mixer gate_output_14_770(.a(output_15_770), .b(output_15_3), .y(output_14_770));
wire output_16_770, output_16_3, output_15_770;
mixer gate_output_15_770(.a(output_16_770), .b(output_16_3), .y(output_15_770));
wire output_1_771, output_1_4, output_0_771;
mixer gate_output_0_771(.a(output_1_771), .b(output_1_4), .y(output_0_771));
wire output_2_771, output_2_4, output_1_771;
mixer gate_output_1_771(.a(output_2_771), .b(output_2_4), .y(output_1_771));
wire output_3_771, output_3_4, output_2_771;
mixer gate_output_2_771(.a(output_3_771), .b(output_3_4), .y(output_2_771));
wire output_4_771, output_4_4, output_3_771;
mixer gate_output_3_771(.a(output_4_771), .b(output_4_4), .y(output_3_771));
wire output_5_771, output_5_4, output_4_771;
mixer gate_output_4_771(.a(output_5_771), .b(output_5_4), .y(output_4_771));
wire output_6_771, output_6_4, output_5_771;
mixer gate_output_5_771(.a(output_6_771), .b(output_6_4), .y(output_5_771));
wire output_7_771, output_7_4, output_6_771;
mixer gate_output_6_771(.a(output_7_771), .b(output_7_4), .y(output_6_771));
wire output_8_771, output_8_4, output_7_771;
mixer gate_output_7_771(.a(output_8_771), .b(output_8_4), .y(output_7_771));
wire output_9_771, output_9_4, output_8_771;
mixer gate_output_8_771(.a(output_9_771), .b(output_9_4), .y(output_8_771));
wire output_10_771, output_10_4, output_9_771;
mixer gate_output_9_771(.a(output_10_771), .b(output_10_4), .y(output_9_771));
wire output_11_771, output_11_4, output_10_771;
mixer gate_output_10_771(.a(output_11_771), .b(output_11_4), .y(output_10_771));
wire output_12_771, output_12_4, output_11_771;
mixer gate_output_11_771(.a(output_12_771), .b(output_12_4), .y(output_11_771));
wire output_13_771, output_13_4, output_12_771;
mixer gate_output_12_771(.a(output_13_771), .b(output_13_4), .y(output_12_771));
wire output_14_771, output_14_4, output_13_771;
mixer gate_output_13_771(.a(output_14_771), .b(output_14_4), .y(output_13_771));
wire output_15_771, output_15_4, output_14_771;
mixer gate_output_14_771(.a(output_15_771), .b(output_15_4), .y(output_14_771));
wire output_16_771, output_16_4, output_15_771;
mixer gate_output_15_771(.a(output_16_771), .b(output_16_4), .y(output_15_771));
wire output_1_772, output_1_5, output_0_772;
mixer gate_output_0_772(.a(output_1_772), .b(output_1_5), .y(output_0_772));
wire output_2_772, output_2_5, output_1_772;
mixer gate_output_1_772(.a(output_2_772), .b(output_2_5), .y(output_1_772));
wire output_3_772, output_3_5, output_2_772;
mixer gate_output_2_772(.a(output_3_772), .b(output_3_5), .y(output_2_772));
wire output_4_772, output_4_5, output_3_772;
mixer gate_output_3_772(.a(output_4_772), .b(output_4_5), .y(output_3_772));
wire output_5_772, output_5_5, output_4_772;
mixer gate_output_4_772(.a(output_5_772), .b(output_5_5), .y(output_4_772));
wire output_6_772, output_6_5, output_5_772;
mixer gate_output_5_772(.a(output_6_772), .b(output_6_5), .y(output_5_772));
wire output_7_772, output_7_5, output_6_772;
mixer gate_output_6_772(.a(output_7_772), .b(output_7_5), .y(output_6_772));
wire output_8_772, output_8_5, output_7_772;
mixer gate_output_7_772(.a(output_8_772), .b(output_8_5), .y(output_7_772));
wire output_9_772, output_9_5, output_8_772;
mixer gate_output_8_772(.a(output_9_772), .b(output_9_5), .y(output_8_772));
wire output_10_772, output_10_5, output_9_772;
mixer gate_output_9_772(.a(output_10_772), .b(output_10_5), .y(output_9_772));
wire output_11_772, output_11_5, output_10_772;
mixer gate_output_10_772(.a(output_11_772), .b(output_11_5), .y(output_10_772));
wire output_12_772, output_12_5, output_11_772;
mixer gate_output_11_772(.a(output_12_772), .b(output_12_5), .y(output_11_772));
wire output_13_772, output_13_5, output_12_772;
mixer gate_output_12_772(.a(output_13_772), .b(output_13_5), .y(output_12_772));
wire output_14_772, output_14_5, output_13_772;
mixer gate_output_13_772(.a(output_14_772), .b(output_14_5), .y(output_13_772));
wire output_15_772, output_15_5, output_14_772;
mixer gate_output_14_772(.a(output_15_772), .b(output_15_5), .y(output_14_772));
wire output_16_772, output_16_5, output_15_772;
mixer gate_output_15_772(.a(output_16_772), .b(output_16_5), .y(output_15_772));
wire output_1_773, output_1_6, output_0_773;
mixer gate_output_0_773(.a(output_1_773), .b(output_1_6), .y(output_0_773));
wire output_2_773, output_2_6, output_1_773;
mixer gate_output_1_773(.a(output_2_773), .b(output_2_6), .y(output_1_773));
wire output_3_773, output_3_6, output_2_773;
mixer gate_output_2_773(.a(output_3_773), .b(output_3_6), .y(output_2_773));
wire output_4_773, output_4_6, output_3_773;
mixer gate_output_3_773(.a(output_4_773), .b(output_4_6), .y(output_3_773));
wire output_5_773, output_5_6, output_4_773;
mixer gate_output_4_773(.a(output_5_773), .b(output_5_6), .y(output_4_773));
wire output_6_773, output_6_6, output_5_773;
mixer gate_output_5_773(.a(output_6_773), .b(output_6_6), .y(output_5_773));
wire output_7_773, output_7_6, output_6_773;
mixer gate_output_6_773(.a(output_7_773), .b(output_7_6), .y(output_6_773));
wire output_8_773, output_8_6, output_7_773;
mixer gate_output_7_773(.a(output_8_773), .b(output_8_6), .y(output_7_773));
wire output_9_773, output_9_6, output_8_773;
mixer gate_output_8_773(.a(output_9_773), .b(output_9_6), .y(output_8_773));
wire output_10_773, output_10_6, output_9_773;
mixer gate_output_9_773(.a(output_10_773), .b(output_10_6), .y(output_9_773));
wire output_11_773, output_11_6, output_10_773;
mixer gate_output_10_773(.a(output_11_773), .b(output_11_6), .y(output_10_773));
wire output_12_773, output_12_6, output_11_773;
mixer gate_output_11_773(.a(output_12_773), .b(output_12_6), .y(output_11_773));
wire output_13_773, output_13_6, output_12_773;
mixer gate_output_12_773(.a(output_13_773), .b(output_13_6), .y(output_12_773));
wire output_14_773, output_14_6, output_13_773;
mixer gate_output_13_773(.a(output_14_773), .b(output_14_6), .y(output_13_773));
wire output_15_773, output_15_6, output_14_773;
mixer gate_output_14_773(.a(output_15_773), .b(output_15_6), .y(output_14_773));
wire output_16_773, output_16_6, output_15_773;
mixer gate_output_15_773(.a(output_16_773), .b(output_16_6), .y(output_15_773));
wire output_1_774, output_1_7, output_0_774;
mixer gate_output_0_774(.a(output_1_774), .b(output_1_7), .y(output_0_774));
wire output_2_774, output_2_7, output_1_774;
mixer gate_output_1_774(.a(output_2_774), .b(output_2_7), .y(output_1_774));
wire output_3_774, output_3_7, output_2_774;
mixer gate_output_2_774(.a(output_3_774), .b(output_3_7), .y(output_2_774));
wire output_4_774, output_4_7, output_3_774;
mixer gate_output_3_774(.a(output_4_774), .b(output_4_7), .y(output_3_774));
wire output_5_774, output_5_7, output_4_774;
mixer gate_output_4_774(.a(output_5_774), .b(output_5_7), .y(output_4_774));
wire output_6_774, output_6_7, output_5_774;
mixer gate_output_5_774(.a(output_6_774), .b(output_6_7), .y(output_5_774));
wire output_7_774, output_7_7, output_6_774;
mixer gate_output_6_774(.a(output_7_774), .b(output_7_7), .y(output_6_774));
wire output_8_774, output_8_7, output_7_774;
mixer gate_output_7_774(.a(output_8_774), .b(output_8_7), .y(output_7_774));
wire output_9_774, output_9_7, output_8_774;
mixer gate_output_8_774(.a(output_9_774), .b(output_9_7), .y(output_8_774));
wire output_10_774, output_10_7, output_9_774;
mixer gate_output_9_774(.a(output_10_774), .b(output_10_7), .y(output_9_774));
wire output_11_774, output_11_7, output_10_774;
mixer gate_output_10_774(.a(output_11_774), .b(output_11_7), .y(output_10_774));
wire output_12_774, output_12_7, output_11_774;
mixer gate_output_11_774(.a(output_12_774), .b(output_12_7), .y(output_11_774));
wire output_13_774, output_13_7, output_12_774;
mixer gate_output_12_774(.a(output_13_774), .b(output_13_7), .y(output_12_774));
wire output_14_774, output_14_7, output_13_774;
mixer gate_output_13_774(.a(output_14_774), .b(output_14_7), .y(output_13_774));
wire output_15_774, output_15_7, output_14_774;
mixer gate_output_14_774(.a(output_15_774), .b(output_15_7), .y(output_14_774));
wire output_16_774, output_16_7, output_15_774;
mixer gate_output_15_774(.a(output_16_774), .b(output_16_7), .y(output_15_774));
wire output_1_775, output_1_8, output_0_775;
mixer gate_output_0_775(.a(output_1_775), .b(output_1_8), .y(output_0_775));
wire output_2_775, output_2_8, output_1_775;
mixer gate_output_1_775(.a(output_2_775), .b(output_2_8), .y(output_1_775));
wire output_3_775, output_3_8, output_2_775;
mixer gate_output_2_775(.a(output_3_775), .b(output_3_8), .y(output_2_775));
wire output_4_775, output_4_8, output_3_775;
mixer gate_output_3_775(.a(output_4_775), .b(output_4_8), .y(output_3_775));
wire output_5_775, output_5_8, output_4_775;
mixer gate_output_4_775(.a(output_5_775), .b(output_5_8), .y(output_4_775));
wire output_6_775, output_6_8, output_5_775;
mixer gate_output_5_775(.a(output_6_775), .b(output_6_8), .y(output_5_775));
wire output_7_775, output_7_8, output_6_775;
mixer gate_output_6_775(.a(output_7_775), .b(output_7_8), .y(output_6_775));
wire output_8_775, output_8_8, output_7_775;
mixer gate_output_7_775(.a(output_8_775), .b(output_8_8), .y(output_7_775));
wire output_9_775, output_9_8, output_8_775;
mixer gate_output_8_775(.a(output_9_775), .b(output_9_8), .y(output_8_775));
wire output_10_775, output_10_8, output_9_775;
mixer gate_output_9_775(.a(output_10_775), .b(output_10_8), .y(output_9_775));
wire output_11_775, output_11_8, output_10_775;
mixer gate_output_10_775(.a(output_11_775), .b(output_11_8), .y(output_10_775));
wire output_12_775, output_12_8, output_11_775;
mixer gate_output_11_775(.a(output_12_775), .b(output_12_8), .y(output_11_775));
wire output_13_775, output_13_8, output_12_775;
mixer gate_output_12_775(.a(output_13_775), .b(output_13_8), .y(output_12_775));
wire output_14_775, output_14_8, output_13_775;
mixer gate_output_13_775(.a(output_14_775), .b(output_14_8), .y(output_13_775));
wire output_15_775, output_15_8, output_14_775;
mixer gate_output_14_775(.a(output_15_775), .b(output_15_8), .y(output_14_775));
wire output_16_775, output_16_8, output_15_775;
mixer gate_output_15_775(.a(output_16_775), .b(output_16_8), .y(output_15_775));
wire output_1_776, output_1_9, output_0_776;
mixer gate_output_0_776(.a(output_1_776), .b(output_1_9), .y(output_0_776));
wire output_2_776, output_2_9, output_1_776;
mixer gate_output_1_776(.a(output_2_776), .b(output_2_9), .y(output_1_776));
wire output_3_776, output_3_9, output_2_776;
mixer gate_output_2_776(.a(output_3_776), .b(output_3_9), .y(output_2_776));
wire output_4_776, output_4_9, output_3_776;
mixer gate_output_3_776(.a(output_4_776), .b(output_4_9), .y(output_3_776));
wire output_5_776, output_5_9, output_4_776;
mixer gate_output_4_776(.a(output_5_776), .b(output_5_9), .y(output_4_776));
wire output_6_776, output_6_9, output_5_776;
mixer gate_output_5_776(.a(output_6_776), .b(output_6_9), .y(output_5_776));
wire output_7_776, output_7_9, output_6_776;
mixer gate_output_6_776(.a(output_7_776), .b(output_7_9), .y(output_6_776));
wire output_8_776, output_8_9, output_7_776;
mixer gate_output_7_776(.a(output_8_776), .b(output_8_9), .y(output_7_776));
wire output_9_776, output_9_9, output_8_776;
mixer gate_output_8_776(.a(output_9_776), .b(output_9_9), .y(output_8_776));
wire output_10_776, output_10_9, output_9_776;
mixer gate_output_9_776(.a(output_10_776), .b(output_10_9), .y(output_9_776));
wire output_11_776, output_11_9, output_10_776;
mixer gate_output_10_776(.a(output_11_776), .b(output_11_9), .y(output_10_776));
wire output_12_776, output_12_9, output_11_776;
mixer gate_output_11_776(.a(output_12_776), .b(output_12_9), .y(output_11_776));
wire output_13_776, output_13_9, output_12_776;
mixer gate_output_12_776(.a(output_13_776), .b(output_13_9), .y(output_12_776));
wire output_14_776, output_14_9, output_13_776;
mixer gate_output_13_776(.a(output_14_776), .b(output_14_9), .y(output_13_776));
wire output_15_776, output_15_9, output_14_776;
mixer gate_output_14_776(.a(output_15_776), .b(output_15_9), .y(output_14_776));
wire output_16_776, output_16_9, output_15_776;
mixer gate_output_15_776(.a(output_16_776), .b(output_16_9), .y(output_15_776));
wire output_1_777, output_1_10, output_0_777;
mixer gate_output_0_777(.a(output_1_777), .b(output_1_10), .y(output_0_777));
wire output_2_777, output_2_10, output_1_777;
mixer gate_output_1_777(.a(output_2_777), .b(output_2_10), .y(output_1_777));
wire output_3_777, output_3_10, output_2_777;
mixer gate_output_2_777(.a(output_3_777), .b(output_3_10), .y(output_2_777));
wire output_4_777, output_4_10, output_3_777;
mixer gate_output_3_777(.a(output_4_777), .b(output_4_10), .y(output_3_777));
wire output_5_777, output_5_10, output_4_777;
mixer gate_output_4_777(.a(output_5_777), .b(output_5_10), .y(output_4_777));
wire output_6_777, output_6_10, output_5_777;
mixer gate_output_5_777(.a(output_6_777), .b(output_6_10), .y(output_5_777));
wire output_7_777, output_7_10, output_6_777;
mixer gate_output_6_777(.a(output_7_777), .b(output_7_10), .y(output_6_777));
wire output_8_777, output_8_10, output_7_777;
mixer gate_output_7_777(.a(output_8_777), .b(output_8_10), .y(output_7_777));
wire output_9_777, output_9_10, output_8_777;
mixer gate_output_8_777(.a(output_9_777), .b(output_9_10), .y(output_8_777));
wire output_10_777, output_10_10, output_9_777;
mixer gate_output_9_777(.a(output_10_777), .b(output_10_10), .y(output_9_777));
wire output_11_777, output_11_10, output_10_777;
mixer gate_output_10_777(.a(output_11_777), .b(output_11_10), .y(output_10_777));
wire output_12_777, output_12_10, output_11_777;
mixer gate_output_11_777(.a(output_12_777), .b(output_12_10), .y(output_11_777));
wire output_13_777, output_13_10, output_12_777;
mixer gate_output_12_777(.a(output_13_777), .b(output_13_10), .y(output_12_777));
wire output_14_777, output_14_10, output_13_777;
mixer gate_output_13_777(.a(output_14_777), .b(output_14_10), .y(output_13_777));
wire output_15_777, output_15_10, output_14_777;
mixer gate_output_14_777(.a(output_15_777), .b(output_15_10), .y(output_14_777));
wire output_16_777, output_16_10, output_15_777;
mixer gate_output_15_777(.a(output_16_777), .b(output_16_10), .y(output_15_777));
wire output_1_778, output_1_11, output_0_778;
mixer gate_output_0_778(.a(output_1_778), .b(output_1_11), .y(output_0_778));
wire output_2_778, output_2_11, output_1_778;
mixer gate_output_1_778(.a(output_2_778), .b(output_2_11), .y(output_1_778));
wire output_3_778, output_3_11, output_2_778;
mixer gate_output_2_778(.a(output_3_778), .b(output_3_11), .y(output_2_778));
wire output_4_778, output_4_11, output_3_778;
mixer gate_output_3_778(.a(output_4_778), .b(output_4_11), .y(output_3_778));
wire output_5_778, output_5_11, output_4_778;
mixer gate_output_4_778(.a(output_5_778), .b(output_5_11), .y(output_4_778));
wire output_6_778, output_6_11, output_5_778;
mixer gate_output_5_778(.a(output_6_778), .b(output_6_11), .y(output_5_778));
wire output_7_778, output_7_11, output_6_778;
mixer gate_output_6_778(.a(output_7_778), .b(output_7_11), .y(output_6_778));
wire output_8_778, output_8_11, output_7_778;
mixer gate_output_7_778(.a(output_8_778), .b(output_8_11), .y(output_7_778));
wire output_9_778, output_9_11, output_8_778;
mixer gate_output_8_778(.a(output_9_778), .b(output_9_11), .y(output_8_778));
wire output_10_778, output_10_11, output_9_778;
mixer gate_output_9_778(.a(output_10_778), .b(output_10_11), .y(output_9_778));
wire output_11_778, output_11_11, output_10_778;
mixer gate_output_10_778(.a(output_11_778), .b(output_11_11), .y(output_10_778));
wire output_12_778, output_12_11, output_11_778;
mixer gate_output_11_778(.a(output_12_778), .b(output_12_11), .y(output_11_778));
wire output_13_778, output_13_11, output_12_778;
mixer gate_output_12_778(.a(output_13_778), .b(output_13_11), .y(output_12_778));
wire output_14_778, output_14_11, output_13_778;
mixer gate_output_13_778(.a(output_14_778), .b(output_14_11), .y(output_13_778));
wire output_15_778, output_15_11, output_14_778;
mixer gate_output_14_778(.a(output_15_778), .b(output_15_11), .y(output_14_778));
wire output_16_778, output_16_11, output_15_778;
mixer gate_output_15_778(.a(output_16_778), .b(output_16_11), .y(output_15_778));
wire output_1_779, output_1_12, output_0_779;
mixer gate_output_0_779(.a(output_1_779), .b(output_1_12), .y(output_0_779));
wire output_2_779, output_2_12, output_1_779;
mixer gate_output_1_779(.a(output_2_779), .b(output_2_12), .y(output_1_779));
wire output_3_779, output_3_12, output_2_779;
mixer gate_output_2_779(.a(output_3_779), .b(output_3_12), .y(output_2_779));
wire output_4_779, output_4_12, output_3_779;
mixer gate_output_3_779(.a(output_4_779), .b(output_4_12), .y(output_3_779));
wire output_5_779, output_5_12, output_4_779;
mixer gate_output_4_779(.a(output_5_779), .b(output_5_12), .y(output_4_779));
wire output_6_779, output_6_12, output_5_779;
mixer gate_output_5_779(.a(output_6_779), .b(output_6_12), .y(output_5_779));
wire output_7_779, output_7_12, output_6_779;
mixer gate_output_6_779(.a(output_7_779), .b(output_7_12), .y(output_6_779));
wire output_8_779, output_8_12, output_7_779;
mixer gate_output_7_779(.a(output_8_779), .b(output_8_12), .y(output_7_779));
wire output_9_779, output_9_12, output_8_779;
mixer gate_output_8_779(.a(output_9_779), .b(output_9_12), .y(output_8_779));
wire output_10_779, output_10_12, output_9_779;
mixer gate_output_9_779(.a(output_10_779), .b(output_10_12), .y(output_9_779));
wire output_11_779, output_11_12, output_10_779;
mixer gate_output_10_779(.a(output_11_779), .b(output_11_12), .y(output_10_779));
wire output_12_779, output_12_12, output_11_779;
mixer gate_output_11_779(.a(output_12_779), .b(output_12_12), .y(output_11_779));
wire output_13_779, output_13_12, output_12_779;
mixer gate_output_12_779(.a(output_13_779), .b(output_13_12), .y(output_12_779));
wire output_14_779, output_14_12, output_13_779;
mixer gate_output_13_779(.a(output_14_779), .b(output_14_12), .y(output_13_779));
wire output_15_779, output_15_12, output_14_779;
mixer gate_output_14_779(.a(output_15_779), .b(output_15_12), .y(output_14_779));
wire output_16_779, output_16_12, output_15_779;
mixer gate_output_15_779(.a(output_16_779), .b(output_16_12), .y(output_15_779));
wire output_1_780, output_1_13, output_0_780;
mixer gate_output_0_780(.a(output_1_780), .b(output_1_13), .y(output_0_780));
wire output_2_780, output_2_13, output_1_780;
mixer gate_output_1_780(.a(output_2_780), .b(output_2_13), .y(output_1_780));
wire output_3_780, output_3_13, output_2_780;
mixer gate_output_2_780(.a(output_3_780), .b(output_3_13), .y(output_2_780));
wire output_4_780, output_4_13, output_3_780;
mixer gate_output_3_780(.a(output_4_780), .b(output_4_13), .y(output_3_780));
wire output_5_780, output_5_13, output_4_780;
mixer gate_output_4_780(.a(output_5_780), .b(output_5_13), .y(output_4_780));
wire output_6_780, output_6_13, output_5_780;
mixer gate_output_5_780(.a(output_6_780), .b(output_6_13), .y(output_5_780));
wire output_7_780, output_7_13, output_6_780;
mixer gate_output_6_780(.a(output_7_780), .b(output_7_13), .y(output_6_780));
wire output_8_780, output_8_13, output_7_780;
mixer gate_output_7_780(.a(output_8_780), .b(output_8_13), .y(output_7_780));
wire output_9_780, output_9_13, output_8_780;
mixer gate_output_8_780(.a(output_9_780), .b(output_9_13), .y(output_8_780));
wire output_10_780, output_10_13, output_9_780;
mixer gate_output_9_780(.a(output_10_780), .b(output_10_13), .y(output_9_780));
wire output_11_780, output_11_13, output_10_780;
mixer gate_output_10_780(.a(output_11_780), .b(output_11_13), .y(output_10_780));
wire output_12_780, output_12_13, output_11_780;
mixer gate_output_11_780(.a(output_12_780), .b(output_12_13), .y(output_11_780));
wire output_13_780, output_13_13, output_12_780;
mixer gate_output_12_780(.a(output_13_780), .b(output_13_13), .y(output_12_780));
wire output_14_780, output_14_13, output_13_780;
mixer gate_output_13_780(.a(output_14_780), .b(output_14_13), .y(output_13_780));
wire output_15_780, output_15_13, output_14_780;
mixer gate_output_14_780(.a(output_15_780), .b(output_15_13), .y(output_14_780));
wire output_16_780, output_16_13, output_15_780;
mixer gate_output_15_780(.a(output_16_780), .b(output_16_13), .y(output_15_780));
wire output_1_781, output_1_14, output_0_781;
mixer gate_output_0_781(.a(output_1_781), .b(output_1_14), .y(output_0_781));
wire output_2_781, output_2_14, output_1_781;
mixer gate_output_1_781(.a(output_2_781), .b(output_2_14), .y(output_1_781));
wire output_3_781, output_3_14, output_2_781;
mixer gate_output_2_781(.a(output_3_781), .b(output_3_14), .y(output_2_781));
wire output_4_781, output_4_14, output_3_781;
mixer gate_output_3_781(.a(output_4_781), .b(output_4_14), .y(output_3_781));
wire output_5_781, output_5_14, output_4_781;
mixer gate_output_4_781(.a(output_5_781), .b(output_5_14), .y(output_4_781));
wire output_6_781, output_6_14, output_5_781;
mixer gate_output_5_781(.a(output_6_781), .b(output_6_14), .y(output_5_781));
wire output_7_781, output_7_14, output_6_781;
mixer gate_output_6_781(.a(output_7_781), .b(output_7_14), .y(output_6_781));
wire output_8_781, output_8_14, output_7_781;
mixer gate_output_7_781(.a(output_8_781), .b(output_8_14), .y(output_7_781));
wire output_9_781, output_9_14, output_8_781;
mixer gate_output_8_781(.a(output_9_781), .b(output_9_14), .y(output_8_781));
wire output_10_781, output_10_14, output_9_781;
mixer gate_output_9_781(.a(output_10_781), .b(output_10_14), .y(output_9_781));
wire output_11_781, output_11_14, output_10_781;
mixer gate_output_10_781(.a(output_11_781), .b(output_11_14), .y(output_10_781));
wire output_12_781, output_12_14, output_11_781;
mixer gate_output_11_781(.a(output_12_781), .b(output_12_14), .y(output_11_781));
wire output_13_781, output_13_14, output_12_781;
mixer gate_output_12_781(.a(output_13_781), .b(output_13_14), .y(output_12_781));
wire output_14_781, output_14_14, output_13_781;
mixer gate_output_13_781(.a(output_14_781), .b(output_14_14), .y(output_13_781));
wire output_15_781, output_15_14, output_14_781;
mixer gate_output_14_781(.a(output_15_781), .b(output_15_14), .y(output_14_781));
wire output_16_781, output_16_14, output_15_781;
mixer gate_output_15_781(.a(output_16_781), .b(output_16_14), .y(output_15_781));
wire output_1_782, output_1_15, output_0_782;
mixer gate_output_0_782(.a(output_1_782), .b(output_1_15), .y(output_0_782));
wire output_2_782, output_2_15, output_1_782;
mixer gate_output_1_782(.a(output_2_782), .b(output_2_15), .y(output_1_782));
wire output_3_782, output_3_15, output_2_782;
mixer gate_output_2_782(.a(output_3_782), .b(output_3_15), .y(output_2_782));
wire output_4_782, output_4_15, output_3_782;
mixer gate_output_3_782(.a(output_4_782), .b(output_4_15), .y(output_3_782));
wire output_5_782, output_5_15, output_4_782;
mixer gate_output_4_782(.a(output_5_782), .b(output_5_15), .y(output_4_782));
wire output_6_782, output_6_15, output_5_782;
mixer gate_output_5_782(.a(output_6_782), .b(output_6_15), .y(output_5_782));
wire output_7_782, output_7_15, output_6_782;
mixer gate_output_6_782(.a(output_7_782), .b(output_7_15), .y(output_6_782));
wire output_8_782, output_8_15, output_7_782;
mixer gate_output_7_782(.a(output_8_782), .b(output_8_15), .y(output_7_782));
wire output_9_782, output_9_15, output_8_782;
mixer gate_output_8_782(.a(output_9_782), .b(output_9_15), .y(output_8_782));
wire output_10_782, output_10_15, output_9_782;
mixer gate_output_9_782(.a(output_10_782), .b(output_10_15), .y(output_9_782));
wire output_11_782, output_11_15, output_10_782;
mixer gate_output_10_782(.a(output_11_782), .b(output_11_15), .y(output_10_782));
wire output_12_782, output_12_15, output_11_782;
mixer gate_output_11_782(.a(output_12_782), .b(output_12_15), .y(output_11_782));
wire output_13_782, output_13_15, output_12_782;
mixer gate_output_12_782(.a(output_13_782), .b(output_13_15), .y(output_12_782));
wire output_14_782, output_14_15, output_13_782;
mixer gate_output_13_782(.a(output_14_782), .b(output_14_15), .y(output_13_782));
wire output_15_782, output_15_15, output_14_782;
mixer gate_output_14_782(.a(output_15_782), .b(output_15_15), .y(output_14_782));
wire output_16_782, output_16_15, output_15_782;
mixer gate_output_15_782(.a(output_16_782), .b(output_16_15), .y(output_15_782));
wire output_1_783, output_1_0, output_0_783;
mixer gate_output_0_783(.a(output_1_783), .b(output_1_0), .y(output_0_783));
wire output_2_783, output_2_0, output_1_783;
mixer gate_output_1_783(.a(output_2_783), .b(output_2_0), .y(output_1_783));
wire output_3_783, output_3_0, output_2_783;
mixer gate_output_2_783(.a(output_3_783), .b(output_3_0), .y(output_2_783));
wire output_4_783, output_4_0, output_3_783;
mixer gate_output_3_783(.a(output_4_783), .b(output_4_0), .y(output_3_783));
wire output_5_783, output_5_0, output_4_783;
mixer gate_output_4_783(.a(output_5_783), .b(output_5_0), .y(output_4_783));
wire output_6_783, output_6_0, output_5_783;
mixer gate_output_5_783(.a(output_6_783), .b(output_6_0), .y(output_5_783));
wire output_7_783, output_7_0, output_6_783;
mixer gate_output_6_783(.a(output_7_783), .b(output_7_0), .y(output_6_783));
wire output_8_783, output_8_0, output_7_783;
mixer gate_output_7_783(.a(output_8_783), .b(output_8_0), .y(output_7_783));
wire output_9_783, output_9_0, output_8_783;
mixer gate_output_8_783(.a(output_9_783), .b(output_9_0), .y(output_8_783));
wire output_10_783, output_10_0, output_9_783;
mixer gate_output_9_783(.a(output_10_783), .b(output_10_0), .y(output_9_783));
wire output_11_783, output_11_0, output_10_783;
mixer gate_output_10_783(.a(output_11_783), .b(output_11_0), .y(output_10_783));
wire output_12_783, output_12_0, output_11_783;
mixer gate_output_11_783(.a(output_12_783), .b(output_12_0), .y(output_11_783));
wire output_13_783, output_13_0, output_12_783;
mixer gate_output_12_783(.a(output_13_783), .b(output_13_0), .y(output_12_783));
wire output_14_783, output_14_0, output_13_783;
mixer gate_output_13_783(.a(output_14_783), .b(output_14_0), .y(output_13_783));
wire output_15_783, output_15_0, output_14_783;
mixer gate_output_14_783(.a(output_15_783), .b(output_15_0), .y(output_14_783));
wire output_16_783, output_16_0, output_15_783;
mixer gate_output_15_783(.a(output_16_783), .b(output_16_0), .y(output_15_783));
wire output_1_784, output_1_1, output_0_784;
mixer gate_output_0_784(.a(output_1_784), .b(output_1_1), .y(output_0_784));
wire output_2_784, output_2_1, output_1_784;
mixer gate_output_1_784(.a(output_2_784), .b(output_2_1), .y(output_1_784));
wire output_3_784, output_3_1, output_2_784;
mixer gate_output_2_784(.a(output_3_784), .b(output_3_1), .y(output_2_784));
wire output_4_784, output_4_1, output_3_784;
mixer gate_output_3_784(.a(output_4_784), .b(output_4_1), .y(output_3_784));
wire output_5_784, output_5_1, output_4_784;
mixer gate_output_4_784(.a(output_5_784), .b(output_5_1), .y(output_4_784));
wire output_6_784, output_6_1, output_5_784;
mixer gate_output_5_784(.a(output_6_784), .b(output_6_1), .y(output_5_784));
wire output_7_784, output_7_1, output_6_784;
mixer gate_output_6_784(.a(output_7_784), .b(output_7_1), .y(output_6_784));
wire output_8_784, output_8_1, output_7_784;
mixer gate_output_7_784(.a(output_8_784), .b(output_8_1), .y(output_7_784));
wire output_9_784, output_9_1, output_8_784;
mixer gate_output_8_784(.a(output_9_784), .b(output_9_1), .y(output_8_784));
wire output_10_784, output_10_1, output_9_784;
mixer gate_output_9_784(.a(output_10_784), .b(output_10_1), .y(output_9_784));
wire output_11_784, output_11_1, output_10_784;
mixer gate_output_10_784(.a(output_11_784), .b(output_11_1), .y(output_10_784));
wire output_12_784, output_12_1, output_11_784;
mixer gate_output_11_784(.a(output_12_784), .b(output_12_1), .y(output_11_784));
wire output_13_784, output_13_1, output_12_784;
mixer gate_output_12_784(.a(output_13_784), .b(output_13_1), .y(output_12_784));
wire output_14_784, output_14_1, output_13_784;
mixer gate_output_13_784(.a(output_14_784), .b(output_14_1), .y(output_13_784));
wire output_15_784, output_15_1, output_14_784;
mixer gate_output_14_784(.a(output_15_784), .b(output_15_1), .y(output_14_784));
wire output_16_784, output_16_1, output_15_784;
mixer gate_output_15_784(.a(output_16_784), .b(output_16_1), .y(output_15_784));
wire output_1_785, output_1_2, output_0_785;
mixer gate_output_0_785(.a(output_1_785), .b(output_1_2), .y(output_0_785));
wire output_2_785, output_2_2, output_1_785;
mixer gate_output_1_785(.a(output_2_785), .b(output_2_2), .y(output_1_785));
wire output_3_785, output_3_2, output_2_785;
mixer gate_output_2_785(.a(output_3_785), .b(output_3_2), .y(output_2_785));
wire output_4_785, output_4_2, output_3_785;
mixer gate_output_3_785(.a(output_4_785), .b(output_4_2), .y(output_3_785));
wire output_5_785, output_5_2, output_4_785;
mixer gate_output_4_785(.a(output_5_785), .b(output_5_2), .y(output_4_785));
wire output_6_785, output_6_2, output_5_785;
mixer gate_output_5_785(.a(output_6_785), .b(output_6_2), .y(output_5_785));
wire output_7_785, output_7_2, output_6_785;
mixer gate_output_6_785(.a(output_7_785), .b(output_7_2), .y(output_6_785));
wire output_8_785, output_8_2, output_7_785;
mixer gate_output_7_785(.a(output_8_785), .b(output_8_2), .y(output_7_785));
wire output_9_785, output_9_2, output_8_785;
mixer gate_output_8_785(.a(output_9_785), .b(output_9_2), .y(output_8_785));
wire output_10_785, output_10_2, output_9_785;
mixer gate_output_9_785(.a(output_10_785), .b(output_10_2), .y(output_9_785));
wire output_11_785, output_11_2, output_10_785;
mixer gate_output_10_785(.a(output_11_785), .b(output_11_2), .y(output_10_785));
wire output_12_785, output_12_2, output_11_785;
mixer gate_output_11_785(.a(output_12_785), .b(output_12_2), .y(output_11_785));
wire output_13_785, output_13_2, output_12_785;
mixer gate_output_12_785(.a(output_13_785), .b(output_13_2), .y(output_12_785));
wire output_14_785, output_14_2, output_13_785;
mixer gate_output_13_785(.a(output_14_785), .b(output_14_2), .y(output_13_785));
wire output_15_785, output_15_2, output_14_785;
mixer gate_output_14_785(.a(output_15_785), .b(output_15_2), .y(output_14_785));
wire output_16_785, output_16_2, output_15_785;
mixer gate_output_15_785(.a(output_16_785), .b(output_16_2), .y(output_15_785));
wire output_1_786, output_1_3, output_0_786;
mixer gate_output_0_786(.a(output_1_786), .b(output_1_3), .y(output_0_786));
wire output_2_786, output_2_3, output_1_786;
mixer gate_output_1_786(.a(output_2_786), .b(output_2_3), .y(output_1_786));
wire output_3_786, output_3_3, output_2_786;
mixer gate_output_2_786(.a(output_3_786), .b(output_3_3), .y(output_2_786));
wire output_4_786, output_4_3, output_3_786;
mixer gate_output_3_786(.a(output_4_786), .b(output_4_3), .y(output_3_786));
wire output_5_786, output_5_3, output_4_786;
mixer gate_output_4_786(.a(output_5_786), .b(output_5_3), .y(output_4_786));
wire output_6_786, output_6_3, output_5_786;
mixer gate_output_5_786(.a(output_6_786), .b(output_6_3), .y(output_5_786));
wire output_7_786, output_7_3, output_6_786;
mixer gate_output_6_786(.a(output_7_786), .b(output_7_3), .y(output_6_786));
wire output_8_786, output_8_3, output_7_786;
mixer gate_output_7_786(.a(output_8_786), .b(output_8_3), .y(output_7_786));
wire output_9_786, output_9_3, output_8_786;
mixer gate_output_8_786(.a(output_9_786), .b(output_9_3), .y(output_8_786));
wire output_10_786, output_10_3, output_9_786;
mixer gate_output_9_786(.a(output_10_786), .b(output_10_3), .y(output_9_786));
wire output_11_786, output_11_3, output_10_786;
mixer gate_output_10_786(.a(output_11_786), .b(output_11_3), .y(output_10_786));
wire output_12_786, output_12_3, output_11_786;
mixer gate_output_11_786(.a(output_12_786), .b(output_12_3), .y(output_11_786));
wire output_13_786, output_13_3, output_12_786;
mixer gate_output_12_786(.a(output_13_786), .b(output_13_3), .y(output_12_786));
wire output_14_786, output_14_3, output_13_786;
mixer gate_output_13_786(.a(output_14_786), .b(output_14_3), .y(output_13_786));
wire output_15_786, output_15_3, output_14_786;
mixer gate_output_14_786(.a(output_15_786), .b(output_15_3), .y(output_14_786));
wire output_16_786, output_16_3, output_15_786;
mixer gate_output_15_786(.a(output_16_786), .b(output_16_3), .y(output_15_786));
wire output_1_787, output_1_4, output_0_787;
mixer gate_output_0_787(.a(output_1_787), .b(output_1_4), .y(output_0_787));
wire output_2_787, output_2_4, output_1_787;
mixer gate_output_1_787(.a(output_2_787), .b(output_2_4), .y(output_1_787));
wire output_3_787, output_3_4, output_2_787;
mixer gate_output_2_787(.a(output_3_787), .b(output_3_4), .y(output_2_787));
wire output_4_787, output_4_4, output_3_787;
mixer gate_output_3_787(.a(output_4_787), .b(output_4_4), .y(output_3_787));
wire output_5_787, output_5_4, output_4_787;
mixer gate_output_4_787(.a(output_5_787), .b(output_5_4), .y(output_4_787));
wire output_6_787, output_6_4, output_5_787;
mixer gate_output_5_787(.a(output_6_787), .b(output_6_4), .y(output_5_787));
wire output_7_787, output_7_4, output_6_787;
mixer gate_output_6_787(.a(output_7_787), .b(output_7_4), .y(output_6_787));
wire output_8_787, output_8_4, output_7_787;
mixer gate_output_7_787(.a(output_8_787), .b(output_8_4), .y(output_7_787));
wire output_9_787, output_9_4, output_8_787;
mixer gate_output_8_787(.a(output_9_787), .b(output_9_4), .y(output_8_787));
wire output_10_787, output_10_4, output_9_787;
mixer gate_output_9_787(.a(output_10_787), .b(output_10_4), .y(output_9_787));
wire output_11_787, output_11_4, output_10_787;
mixer gate_output_10_787(.a(output_11_787), .b(output_11_4), .y(output_10_787));
wire output_12_787, output_12_4, output_11_787;
mixer gate_output_11_787(.a(output_12_787), .b(output_12_4), .y(output_11_787));
wire output_13_787, output_13_4, output_12_787;
mixer gate_output_12_787(.a(output_13_787), .b(output_13_4), .y(output_12_787));
wire output_14_787, output_14_4, output_13_787;
mixer gate_output_13_787(.a(output_14_787), .b(output_14_4), .y(output_13_787));
wire output_15_787, output_15_4, output_14_787;
mixer gate_output_14_787(.a(output_15_787), .b(output_15_4), .y(output_14_787));
wire output_16_787, output_16_4, output_15_787;
mixer gate_output_15_787(.a(output_16_787), .b(output_16_4), .y(output_15_787));
wire output_1_788, output_1_5, output_0_788;
mixer gate_output_0_788(.a(output_1_788), .b(output_1_5), .y(output_0_788));
wire output_2_788, output_2_5, output_1_788;
mixer gate_output_1_788(.a(output_2_788), .b(output_2_5), .y(output_1_788));
wire output_3_788, output_3_5, output_2_788;
mixer gate_output_2_788(.a(output_3_788), .b(output_3_5), .y(output_2_788));
wire output_4_788, output_4_5, output_3_788;
mixer gate_output_3_788(.a(output_4_788), .b(output_4_5), .y(output_3_788));
wire output_5_788, output_5_5, output_4_788;
mixer gate_output_4_788(.a(output_5_788), .b(output_5_5), .y(output_4_788));
wire output_6_788, output_6_5, output_5_788;
mixer gate_output_5_788(.a(output_6_788), .b(output_6_5), .y(output_5_788));
wire output_7_788, output_7_5, output_6_788;
mixer gate_output_6_788(.a(output_7_788), .b(output_7_5), .y(output_6_788));
wire output_8_788, output_8_5, output_7_788;
mixer gate_output_7_788(.a(output_8_788), .b(output_8_5), .y(output_7_788));
wire output_9_788, output_9_5, output_8_788;
mixer gate_output_8_788(.a(output_9_788), .b(output_9_5), .y(output_8_788));
wire output_10_788, output_10_5, output_9_788;
mixer gate_output_9_788(.a(output_10_788), .b(output_10_5), .y(output_9_788));
wire output_11_788, output_11_5, output_10_788;
mixer gate_output_10_788(.a(output_11_788), .b(output_11_5), .y(output_10_788));
wire output_12_788, output_12_5, output_11_788;
mixer gate_output_11_788(.a(output_12_788), .b(output_12_5), .y(output_11_788));
wire output_13_788, output_13_5, output_12_788;
mixer gate_output_12_788(.a(output_13_788), .b(output_13_5), .y(output_12_788));
wire output_14_788, output_14_5, output_13_788;
mixer gate_output_13_788(.a(output_14_788), .b(output_14_5), .y(output_13_788));
wire output_15_788, output_15_5, output_14_788;
mixer gate_output_14_788(.a(output_15_788), .b(output_15_5), .y(output_14_788));
wire output_16_788, output_16_5, output_15_788;
mixer gate_output_15_788(.a(output_16_788), .b(output_16_5), .y(output_15_788));
wire output_1_789, output_1_6, output_0_789;
mixer gate_output_0_789(.a(output_1_789), .b(output_1_6), .y(output_0_789));
wire output_2_789, output_2_6, output_1_789;
mixer gate_output_1_789(.a(output_2_789), .b(output_2_6), .y(output_1_789));
wire output_3_789, output_3_6, output_2_789;
mixer gate_output_2_789(.a(output_3_789), .b(output_3_6), .y(output_2_789));
wire output_4_789, output_4_6, output_3_789;
mixer gate_output_3_789(.a(output_4_789), .b(output_4_6), .y(output_3_789));
wire output_5_789, output_5_6, output_4_789;
mixer gate_output_4_789(.a(output_5_789), .b(output_5_6), .y(output_4_789));
wire output_6_789, output_6_6, output_5_789;
mixer gate_output_5_789(.a(output_6_789), .b(output_6_6), .y(output_5_789));
wire output_7_789, output_7_6, output_6_789;
mixer gate_output_6_789(.a(output_7_789), .b(output_7_6), .y(output_6_789));
wire output_8_789, output_8_6, output_7_789;
mixer gate_output_7_789(.a(output_8_789), .b(output_8_6), .y(output_7_789));
wire output_9_789, output_9_6, output_8_789;
mixer gate_output_8_789(.a(output_9_789), .b(output_9_6), .y(output_8_789));
wire output_10_789, output_10_6, output_9_789;
mixer gate_output_9_789(.a(output_10_789), .b(output_10_6), .y(output_9_789));
wire output_11_789, output_11_6, output_10_789;
mixer gate_output_10_789(.a(output_11_789), .b(output_11_6), .y(output_10_789));
wire output_12_789, output_12_6, output_11_789;
mixer gate_output_11_789(.a(output_12_789), .b(output_12_6), .y(output_11_789));
wire output_13_789, output_13_6, output_12_789;
mixer gate_output_12_789(.a(output_13_789), .b(output_13_6), .y(output_12_789));
wire output_14_789, output_14_6, output_13_789;
mixer gate_output_13_789(.a(output_14_789), .b(output_14_6), .y(output_13_789));
wire output_15_789, output_15_6, output_14_789;
mixer gate_output_14_789(.a(output_15_789), .b(output_15_6), .y(output_14_789));
wire output_16_789, output_16_6, output_15_789;
mixer gate_output_15_789(.a(output_16_789), .b(output_16_6), .y(output_15_789));
wire output_1_790, output_1_7, output_0_790;
mixer gate_output_0_790(.a(output_1_790), .b(output_1_7), .y(output_0_790));
wire output_2_790, output_2_7, output_1_790;
mixer gate_output_1_790(.a(output_2_790), .b(output_2_7), .y(output_1_790));
wire output_3_790, output_3_7, output_2_790;
mixer gate_output_2_790(.a(output_3_790), .b(output_3_7), .y(output_2_790));
wire output_4_790, output_4_7, output_3_790;
mixer gate_output_3_790(.a(output_4_790), .b(output_4_7), .y(output_3_790));
wire output_5_790, output_5_7, output_4_790;
mixer gate_output_4_790(.a(output_5_790), .b(output_5_7), .y(output_4_790));
wire output_6_790, output_6_7, output_5_790;
mixer gate_output_5_790(.a(output_6_790), .b(output_6_7), .y(output_5_790));
wire output_7_790, output_7_7, output_6_790;
mixer gate_output_6_790(.a(output_7_790), .b(output_7_7), .y(output_6_790));
wire output_8_790, output_8_7, output_7_790;
mixer gate_output_7_790(.a(output_8_790), .b(output_8_7), .y(output_7_790));
wire output_9_790, output_9_7, output_8_790;
mixer gate_output_8_790(.a(output_9_790), .b(output_9_7), .y(output_8_790));
wire output_10_790, output_10_7, output_9_790;
mixer gate_output_9_790(.a(output_10_790), .b(output_10_7), .y(output_9_790));
wire output_11_790, output_11_7, output_10_790;
mixer gate_output_10_790(.a(output_11_790), .b(output_11_7), .y(output_10_790));
wire output_12_790, output_12_7, output_11_790;
mixer gate_output_11_790(.a(output_12_790), .b(output_12_7), .y(output_11_790));
wire output_13_790, output_13_7, output_12_790;
mixer gate_output_12_790(.a(output_13_790), .b(output_13_7), .y(output_12_790));
wire output_14_790, output_14_7, output_13_790;
mixer gate_output_13_790(.a(output_14_790), .b(output_14_7), .y(output_13_790));
wire output_15_790, output_15_7, output_14_790;
mixer gate_output_14_790(.a(output_15_790), .b(output_15_7), .y(output_14_790));
wire output_16_790, output_16_7, output_15_790;
mixer gate_output_15_790(.a(output_16_790), .b(output_16_7), .y(output_15_790));
wire output_1_791, output_1_8, output_0_791;
mixer gate_output_0_791(.a(output_1_791), .b(output_1_8), .y(output_0_791));
wire output_2_791, output_2_8, output_1_791;
mixer gate_output_1_791(.a(output_2_791), .b(output_2_8), .y(output_1_791));
wire output_3_791, output_3_8, output_2_791;
mixer gate_output_2_791(.a(output_3_791), .b(output_3_8), .y(output_2_791));
wire output_4_791, output_4_8, output_3_791;
mixer gate_output_3_791(.a(output_4_791), .b(output_4_8), .y(output_3_791));
wire output_5_791, output_5_8, output_4_791;
mixer gate_output_4_791(.a(output_5_791), .b(output_5_8), .y(output_4_791));
wire output_6_791, output_6_8, output_5_791;
mixer gate_output_5_791(.a(output_6_791), .b(output_6_8), .y(output_5_791));
wire output_7_791, output_7_8, output_6_791;
mixer gate_output_6_791(.a(output_7_791), .b(output_7_8), .y(output_6_791));
wire output_8_791, output_8_8, output_7_791;
mixer gate_output_7_791(.a(output_8_791), .b(output_8_8), .y(output_7_791));
wire output_9_791, output_9_8, output_8_791;
mixer gate_output_8_791(.a(output_9_791), .b(output_9_8), .y(output_8_791));
wire output_10_791, output_10_8, output_9_791;
mixer gate_output_9_791(.a(output_10_791), .b(output_10_8), .y(output_9_791));
wire output_11_791, output_11_8, output_10_791;
mixer gate_output_10_791(.a(output_11_791), .b(output_11_8), .y(output_10_791));
wire output_12_791, output_12_8, output_11_791;
mixer gate_output_11_791(.a(output_12_791), .b(output_12_8), .y(output_11_791));
wire output_13_791, output_13_8, output_12_791;
mixer gate_output_12_791(.a(output_13_791), .b(output_13_8), .y(output_12_791));
wire output_14_791, output_14_8, output_13_791;
mixer gate_output_13_791(.a(output_14_791), .b(output_14_8), .y(output_13_791));
wire output_15_791, output_15_8, output_14_791;
mixer gate_output_14_791(.a(output_15_791), .b(output_15_8), .y(output_14_791));
wire output_16_791, output_16_8, output_15_791;
mixer gate_output_15_791(.a(output_16_791), .b(output_16_8), .y(output_15_791));
wire output_1_792, output_1_9, output_0_792;
mixer gate_output_0_792(.a(output_1_792), .b(output_1_9), .y(output_0_792));
wire output_2_792, output_2_9, output_1_792;
mixer gate_output_1_792(.a(output_2_792), .b(output_2_9), .y(output_1_792));
wire output_3_792, output_3_9, output_2_792;
mixer gate_output_2_792(.a(output_3_792), .b(output_3_9), .y(output_2_792));
wire output_4_792, output_4_9, output_3_792;
mixer gate_output_3_792(.a(output_4_792), .b(output_4_9), .y(output_3_792));
wire output_5_792, output_5_9, output_4_792;
mixer gate_output_4_792(.a(output_5_792), .b(output_5_9), .y(output_4_792));
wire output_6_792, output_6_9, output_5_792;
mixer gate_output_5_792(.a(output_6_792), .b(output_6_9), .y(output_5_792));
wire output_7_792, output_7_9, output_6_792;
mixer gate_output_6_792(.a(output_7_792), .b(output_7_9), .y(output_6_792));
wire output_8_792, output_8_9, output_7_792;
mixer gate_output_7_792(.a(output_8_792), .b(output_8_9), .y(output_7_792));
wire output_9_792, output_9_9, output_8_792;
mixer gate_output_8_792(.a(output_9_792), .b(output_9_9), .y(output_8_792));
wire output_10_792, output_10_9, output_9_792;
mixer gate_output_9_792(.a(output_10_792), .b(output_10_9), .y(output_9_792));
wire output_11_792, output_11_9, output_10_792;
mixer gate_output_10_792(.a(output_11_792), .b(output_11_9), .y(output_10_792));
wire output_12_792, output_12_9, output_11_792;
mixer gate_output_11_792(.a(output_12_792), .b(output_12_9), .y(output_11_792));
wire output_13_792, output_13_9, output_12_792;
mixer gate_output_12_792(.a(output_13_792), .b(output_13_9), .y(output_12_792));
wire output_14_792, output_14_9, output_13_792;
mixer gate_output_13_792(.a(output_14_792), .b(output_14_9), .y(output_13_792));
wire output_15_792, output_15_9, output_14_792;
mixer gate_output_14_792(.a(output_15_792), .b(output_15_9), .y(output_14_792));
wire output_16_792, output_16_9, output_15_792;
mixer gate_output_15_792(.a(output_16_792), .b(output_16_9), .y(output_15_792));
wire output_1_793, output_1_10, output_0_793;
mixer gate_output_0_793(.a(output_1_793), .b(output_1_10), .y(output_0_793));
wire output_2_793, output_2_10, output_1_793;
mixer gate_output_1_793(.a(output_2_793), .b(output_2_10), .y(output_1_793));
wire output_3_793, output_3_10, output_2_793;
mixer gate_output_2_793(.a(output_3_793), .b(output_3_10), .y(output_2_793));
wire output_4_793, output_4_10, output_3_793;
mixer gate_output_3_793(.a(output_4_793), .b(output_4_10), .y(output_3_793));
wire output_5_793, output_5_10, output_4_793;
mixer gate_output_4_793(.a(output_5_793), .b(output_5_10), .y(output_4_793));
wire output_6_793, output_6_10, output_5_793;
mixer gate_output_5_793(.a(output_6_793), .b(output_6_10), .y(output_5_793));
wire output_7_793, output_7_10, output_6_793;
mixer gate_output_6_793(.a(output_7_793), .b(output_7_10), .y(output_6_793));
wire output_8_793, output_8_10, output_7_793;
mixer gate_output_7_793(.a(output_8_793), .b(output_8_10), .y(output_7_793));
wire output_9_793, output_9_10, output_8_793;
mixer gate_output_8_793(.a(output_9_793), .b(output_9_10), .y(output_8_793));
wire output_10_793, output_10_10, output_9_793;
mixer gate_output_9_793(.a(output_10_793), .b(output_10_10), .y(output_9_793));
wire output_11_793, output_11_10, output_10_793;
mixer gate_output_10_793(.a(output_11_793), .b(output_11_10), .y(output_10_793));
wire output_12_793, output_12_10, output_11_793;
mixer gate_output_11_793(.a(output_12_793), .b(output_12_10), .y(output_11_793));
wire output_13_793, output_13_10, output_12_793;
mixer gate_output_12_793(.a(output_13_793), .b(output_13_10), .y(output_12_793));
wire output_14_793, output_14_10, output_13_793;
mixer gate_output_13_793(.a(output_14_793), .b(output_14_10), .y(output_13_793));
wire output_15_793, output_15_10, output_14_793;
mixer gate_output_14_793(.a(output_15_793), .b(output_15_10), .y(output_14_793));
wire output_16_793, output_16_10, output_15_793;
mixer gate_output_15_793(.a(output_16_793), .b(output_16_10), .y(output_15_793));
wire output_1_794, output_1_11, output_0_794;
mixer gate_output_0_794(.a(output_1_794), .b(output_1_11), .y(output_0_794));
wire output_2_794, output_2_11, output_1_794;
mixer gate_output_1_794(.a(output_2_794), .b(output_2_11), .y(output_1_794));
wire output_3_794, output_3_11, output_2_794;
mixer gate_output_2_794(.a(output_3_794), .b(output_3_11), .y(output_2_794));
wire output_4_794, output_4_11, output_3_794;
mixer gate_output_3_794(.a(output_4_794), .b(output_4_11), .y(output_3_794));
wire output_5_794, output_5_11, output_4_794;
mixer gate_output_4_794(.a(output_5_794), .b(output_5_11), .y(output_4_794));
wire output_6_794, output_6_11, output_5_794;
mixer gate_output_5_794(.a(output_6_794), .b(output_6_11), .y(output_5_794));
wire output_7_794, output_7_11, output_6_794;
mixer gate_output_6_794(.a(output_7_794), .b(output_7_11), .y(output_6_794));
wire output_8_794, output_8_11, output_7_794;
mixer gate_output_7_794(.a(output_8_794), .b(output_8_11), .y(output_7_794));
wire output_9_794, output_9_11, output_8_794;
mixer gate_output_8_794(.a(output_9_794), .b(output_9_11), .y(output_8_794));
wire output_10_794, output_10_11, output_9_794;
mixer gate_output_9_794(.a(output_10_794), .b(output_10_11), .y(output_9_794));
wire output_11_794, output_11_11, output_10_794;
mixer gate_output_10_794(.a(output_11_794), .b(output_11_11), .y(output_10_794));
wire output_12_794, output_12_11, output_11_794;
mixer gate_output_11_794(.a(output_12_794), .b(output_12_11), .y(output_11_794));
wire output_13_794, output_13_11, output_12_794;
mixer gate_output_12_794(.a(output_13_794), .b(output_13_11), .y(output_12_794));
wire output_14_794, output_14_11, output_13_794;
mixer gate_output_13_794(.a(output_14_794), .b(output_14_11), .y(output_13_794));
wire output_15_794, output_15_11, output_14_794;
mixer gate_output_14_794(.a(output_15_794), .b(output_15_11), .y(output_14_794));
wire output_16_794, output_16_11, output_15_794;
mixer gate_output_15_794(.a(output_16_794), .b(output_16_11), .y(output_15_794));
wire output_1_795, output_1_12, output_0_795;
mixer gate_output_0_795(.a(output_1_795), .b(output_1_12), .y(output_0_795));
wire output_2_795, output_2_12, output_1_795;
mixer gate_output_1_795(.a(output_2_795), .b(output_2_12), .y(output_1_795));
wire output_3_795, output_3_12, output_2_795;
mixer gate_output_2_795(.a(output_3_795), .b(output_3_12), .y(output_2_795));
wire output_4_795, output_4_12, output_3_795;
mixer gate_output_3_795(.a(output_4_795), .b(output_4_12), .y(output_3_795));
wire output_5_795, output_5_12, output_4_795;
mixer gate_output_4_795(.a(output_5_795), .b(output_5_12), .y(output_4_795));
wire output_6_795, output_6_12, output_5_795;
mixer gate_output_5_795(.a(output_6_795), .b(output_6_12), .y(output_5_795));
wire output_7_795, output_7_12, output_6_795;
mixer gate_output_6_795(.a(output_7_795), .b(output_7_12), .y(output_6_795));
wire output_8_795, output_8_12, output_7_795;
mixer gate_output_7_795(.a(output_8_795), .b(output_8_12), .y(output_7_795));
wire output_9_795, output_9_12, output_8_795;
mixer gate_output_8_795(.a(output_9_795), .b(output_9_12), .y(output_8_795));
wire output_10_795, output_10_12, output_9_795;
mixer gate_output_9_795(.a(output_10_795), .b(output_10_12), .y(output_9_795));
wire output_11_795, output_11_12, output_10_795;
mixer gate_output_10_795(.a(output_11_795), .b(output_11_12), .y(output_10_795));
wire output_12_795, output_12_12, output_11_795;
mixer gate_output_11_795(.a(output_12_795), .b(output_12_12), .y(output_11_795));
wire output_13_795, output_13_12, output_12_795;
mixer gate_output_12_795(.a(output_13_795), .b(output_13_12), .y(output_12_795));
wire output_14_795, output_14_12, output_13_795;
mixer gate_output_13_795(.a(output_14_795), .b(output_14_12), .y(output_13_795));
wire output_15_795, output_15_12, output_14_795;
mixer gate_output_14_795(.a(output_15_795), .b(output_15_12), .y(output_14_795));
wire output_16_795, output_16_12, output_15_795;
mixer gate_output_15_795(.a(output_16_795), .b(output_16_12), .y(output_15_795));
wire output_1_796, output_1_13, output_0_796;
mixer gate_output_0_796(.a(output_1_796), .b(output_1_13), .y(output_0_796));
wire output_2_796, output_2_13, output_1_796;
mixer gate_output_1_796(.a(output_2_796), .b(output_2_13), .y(output_1_796));
wire output_3_796, output_3_13, output_2_796;
mixer gate_output_2_796(.a(output_3_796), .b(output_3_13), .y(output_2_796));
wire output_4_796, output_4_13, output_3_796;
mixer gate_output_3_796(.a(output_4_796), .b(output_4_13), .y(output_3_796));
wire output_5_796, output_5_13, output_4_796;
mixer gate_output_4_796(.a(output_5_796), .b(output_5_13), .y(output_4_796));
wire output_6_796, output_6_13, output_5_796;
mixer gate_output_5_796(.a(output_6_796), .b(output_6_13), .y(output_5_796));
wire output_7_796, output_7_13, output_6_796;
mixer gate_output_6_796(.a(output_7_796), .b(output_7_13), .y(output_6_796));
wire output_8_796, output_8_13, output_7_796;
mixer gate_output_7_796(.a(output_8_796), .b(output_8_13), .y(output_7_796));
wire output_9_796, output_9_13, output_8_796;
mixer gate_output_8_796(.a(output_9_796), .b(output_9_13), .y(output_8_796));
wire output_10_796, output_10_13, output_9_796;
mixer gate_output_9_796(.a(output_10_796), .b(output_10_13), .y(output_9_796));
wire output_11_796, output_11_13, output_10_796;
mixer gate_output_10_796(.a(output_11_796), .b(output_11_13), .y(output_10_796));
wire output_12_796, output_12_13, output_11_796;
mixer gate_output_11_796(.a(output_12_796), .b(output_12_13), .y(output_11_796));
wire output_13_796, output_13_13, output_12_796;
mixer gate_output_12_796(.a(output_13_796), .b(output_13_13), .y(output_12_796));
wire output_14_796, output_14_13, output_13_796;
mixer gate_output_13_796(.a(output_14_796), .b(output_14_13), .y(output_13_796));
wire output_15_796, output_15_13, output_14_796;
mixer gate_output_14_796(.a(output_15_796), .b(output_15_13), .y(output_14_796));
wire output_16_796, output_16_13, output_15_796;
mixer gate_output_15_796(.a(output_16_796), .b(output_16_13), .y(output_15_796));
wire output_1_797, output_1_14, output_0_797;
mixer gate_output_0_797(.a(output_1_797), .b(output_1_14), .y(output_0_797));
wire output_2_797, output_2_14, output_1_797;
mixer gate_output_1_797(.a(output_2_797), .b(output_2_14), .y(output_1_797));
wire output_3_797, output_3_14, output_2_797;
mixer gate_output_2_797(.a(output_3_797), .b(output_3_14), .y(output_2_797));
wire output_4_797, output_4_14, output_3_797;
mixer gate_output_3_797(.a(output_4_797), .b(output_4_14), .y(output_3_797));
wire output_5_797, output_5_14, output_4_797;
mixer gate_output_4_797(.a(output_5_797), .b(output_5_14), .y(output_4_797));
wire output_6_797, output_6_14, output_5_797;
mixer gate_output_5_797(.a(output_6_797), .b(output_6_14), .y(output_5_797));
wire output_7_797, output_7_14, output_6_797;
mixer gate_output_6_797(.a(output_7_797), .b(output_7_14), .y(output_6_797));
wire output_8_797, output_8_14, output_7_797;
mixer gate_output_7_797(.a(output_8_797), .b(output_8_14), .y(output_7_797));
wire output_9_797, output_9_14, output_8_797;
mixer gate_output_8_797(.a(output_9_797), .b(output_9_14), .y(output_8_797));
wire output_10_797, output_10_14, output_9_797;
mixer gate_output_9_797(.a(output_10_797), .b(output_10_14), .y(output_9_797));
wire output_11_797, output_11_14, output_10_797;
mixer gate_output_10_797(.a(output_11_797), .b(output_11_14), .y(output_10_797));
wire output_12_797, output_12_14, output_11_797;
mixer gate_output_11_797(.a(output_12_797), .b(output_12_14), .y(output_11_797));
wire output_13_797, output_13_14, output_12_797;
mixer gate_output_12_797(.a(output_13_797), .b(output_13_14), .y(output_12_797));
wire output_14_797, output_14_14, output_13_797;
mixer gate_output_13_797(.a(output_14_797), .b(output_14_14), .y(output_13_797));
wire output_15_797, output_15_14, output_14_797;
mixer gate_output_14_797(.a(output_15_797), .b(output_15_14), .y(output_14_797));
wire output_16_797, output_16_14, output_15_797;
mixer gate_output_15_797(.a(output_16_797), .b(output_16_14), .y(output_15_797));
wire output_1_798, output_1_15, output_0_798;
mixer gate_output_0_798(.a(output_1_798), .b(output_1_15), .y(output_0_798));
wire output_2_798, output_2_15, output_1_798;
mixer gate_output_1_798(.a(output_2_798), .b(output_2_15), .y(output_1_798));
wire output_3_798, output_3_15, output_2_798;
mixer gate_output_2_798(.a(output_3_798), .b(output_3_15), .y(output_2_798));
wire output_4_798, output_4_15, output_3_798;
mixer gate_output_3_798(.a(output_4_798), .b(output_4_15), .y(output_3_798));
wire output_5_798, output_5_15, output_4_798;
mixer gate_output_4_798(.a(output_5_798), .b(output_5_15), .y(output_4_798));
wire output_6_798, output_6_15, output_5_798;
mixer gate_output_5_798(.a(output_6_798), .b(output_6_15), .y(output_5_798));
wire output_7_798, output_7_15, output_6_798;
mixer gate_output_6_798(.a(output_7_798), .b(output_7_15), .y(output_6_798));
wire output_8_798, output_8_15, output_7_798;
mixer gate_output_7_798(.a(output_8_798), .b(output_8_15), .y(output_7_798));
wire output_9_798, output_9_15, output_8_798;
mixer gate_output_8_798(.a(output_9_798), .b(output_9_15), .y(output_8_798));
wire output_10_798, output_10_15, output_9_798;
mixer gate_output_9_798(.a(output_10_798), .b(output_10_15), .y(output_9_798));
wire output_11_798, output_11_15, output_10_798;
mixer gate_output_10_798(.a(output_11_798), .b(output_11_15), .y(output_10_798));
wire output_12_798, output_12_15, output_11_798;
mixer gate_output_11_798(.a(output_12_798), .b(output_12_15), .y(output_11_798));
wire output_13_798, output_13_15, output_12_798;
mixer gate_output_12_798(.a(output_13_798), .b(output_13_15), .y(output_12_798));
wire output_14_798, output_14_15, output_13_798;
mixer gate_output_13_798(.a(output_14_798), .b(output_14_15), .y(output_13_798));
wire output_15_798, output_15_15, output_14_798;
mixer gate_output_14_798(.a(output_15_798), .b(output_15_15), .y(output_14_798));
wire output_16_798, output_16_15, output_15_798;
mixer gate_output_15_798(.a(output_16_798), .b(output_16_15), .y(output_15_798));
wire output_1_799, output_1_0, output_0_799;
mixer gate_output_0_799(.a(output_1_799), .b(output_1_0), .y(output_0_799));
wire output_2_799, output_2_0, output_1_799;
mixer gate_output_1_799(.a(output_2_799), .b(output_2_0), .y(output_1_799));
wire output_3_799, output_3_0, output_2_799;
mixer gate_output_2_799(.a(output_3_799), .b(output_3_0), .y(output_2_799));
wire output_4_799, output_4_0, output_3_799;
mixer gate_output_3_799(.a(output_4_799), .b(output_4_0), .y(output_3_799));
wire output_5_799, output_5_0, output_4_799;
mixer gate_output_4_799(.a(output_5_799), .b(output_5_0), .y(output_4_799));
wire output_6_799, output_6_0, output_5_799;
mixer gate_output_5_799(.a(output_6_799), .b(output_6_0), .y(output_5_799));
wire output_7_799, output_7_0, output_6_799;
mixer gate_output_6_799(.a(output_7_799), .b(output_7_0), .y(output_6_799));
wire output_8_799, output_8_0, output_7_799;
mixer gate_output_7_799(.a(output_8_799), .b(output_8_0), .y(output_7_799));
wire output_9_799, output_9_0, output_8_799;
mixer gate_output_8_799(.a(output_9_799), .b(output_9_0), .y(output_8_799));
wire output_10_799, output_10_0, output_9_799;
mixer gate_output_9_799(.a(output_10_799), .b(output_10_0), .y(output_9_799));
wire output_11_799, output_11_0, output_10_799;
mixer gate_output_10_799(.a(output_11_799), .b(output_11_0), .y(output_10_799));
wire output_12_799, output_12_0, output_11_799;
mixer gate_output_11_799(.a(output_12_799), .b(output_12_0), .y(output_11_799));
wire output_13_799, output_13_0, output_12_799;
mixer gate_output_12_799(.a(output_13_799), .b(output_13_0), .y(output_12_799));
wire output_14_799, output_14_0, output_13_799;
mixer gate_output_13_799(.a(output_14_799), .b(output_14_0), .y(output_13_799));
wire output_15_799, output_15_0, output_14_799;
mixer gate_output_14_799(.a(output_15_799), .b(output_15_0), .y(output_14_799));
wire output_16_799, output_16_0, output_15_799;
mixer gate_output_15_799(.a(output_16_799), .b(output_16_0), .y(output_15_799));
wire output_1_800, output_1_1, output_0_800;
mixer gate_output_0_800(.a(output_1_800), .b(output_1_1), .y(output_0_800));
wire output_2_800, output_2_1, output_1_800;
mixer gate_output_1_800(.a(output_2_800), .b(output_2_1), .y(output_1_800));
wire output_3_800, output_3_1, output_2_800;
mixer gate_output_2_800(.a(output_3_800), .b(output_3_1), .y(output_2_800));
wire output_4_800, output_4_1, output_3_800;
mixer gate_output_3_800(.a(output_4_800), .b(output_4_1), .y(output_3_800));
wire output_5_800, output_5_1, output_4_800;
mixer gate_output_4_800(.a(output_5_800), .b(output_5_1), .y(output_4_800));
wire output_6_800, output_6_1, output_5_800;
mixer gate_output_5_800(.a(output_6_800), .b(output_6_1), .y(output_5_800));
wire output_7_800, output_7_1, output_6_800;
mixer gate_output_6_800(.a(output_7_800), .b(output_7_1), .y(output_6_800));
wire output_8_800, output_8_1, output_7_800;
mixer gate_output_7_800(.a(output_8_800), .b(output_8_1), .y(output_7_800));
wire output_9_800, output_9_1, output_8_800;
mixer gate_output_8_800(.a(output_9_800), .b(output_9_1), .y(output_8_800));
wire output_10_800, output_10_1, output_9_800;
mixer gate_output_9_800(.a(output_10_800), .b(output_10_1), .y(output_9_800));
wire output_11_800, output_11_1, output_10_800;
mixer gate_output_10_800(.a(output_11_800), .b(output_11_1), .y(output_10_800));
wire output_12_800, output_12_1, output_11_800;
mixer gate_output_11_800(.a(output_12_800), .b(output_12_1), .y(output_11_800));
wire output_13_800, output_13_1, output_12_800;
mixer gate_output_12_800(.a(output_13_800), .b(output_13_1), .y(output_12_800));
wire output_14_800, output_14_1, output_13_800;
mixer gate_output_13_800(.a(output_14_800), .b(output_14_1), .y(output_13_800));
wire output_15_800, output_15_1, output_14_800;
mixer gate_output_14_800(.a(output_15_800), .b(output_15_1), .y(output_14_800));
wire output_16_800, output_16_1, output_15_800;
mixer gate_output_15_800(.a(output_16_800), .b(output_16_1), .y(output_15_800));
wire output_1_801, output_1_2, output_0_801;
mixer gate_output_0_801(.a(output_1_801), .b(output_1_2), .y(output_0_801));
wire output_2_801, output_2_2, output_1_801;
mixer gate_output_1_801(.a(output_2_801), .b(output_2_2), .y(output_1_801));
wire output_3_801, output_3_2, output_2_801;
mixer gate_output_2_801(.a(output_3_801), .b(output_3_2), .y(output_2_801));
wire output_4_801, output_4_2, output_3_801;
mixer gate_output_3_801(.a(output_4_801), .b(output_4_2), .y(output_3_801));
wire output_5_801, output_5_2, output_4_801;
mixer gate_output_4_801(.a(output_5_801), .b(output_5_2), .y(output_4_801));
wire output_6_801, output_6_2, output_5_801;
mixer gate_output_5_801(.a(output_6_801), .b(output_6_2), .y(output_5_801));
wire output_7_801, output_7_2, output_6_801;
mixer gate_output_6_801(.a(output_7_801), .b(output_7_2), .y(output_6_801));
wire output_8_801, output_8_2, output_7_801;
mixer gate_output_7_801(.a(output_8_801), .b(output_8_2), .y(output_7_801));
wire output_9_801, output_9_2, output_8_801;
mixer gate_output_8_801(.a(output_9_801), .b(output_9_2), .y(output_8_801));
wire output_10_801, output_10_2, output_9_801;
mixer gate_output_9_801(.a(output_10_801), .b(output_10_2), .y(output_9_801));
wire output_11_801, output_11_2, output_10_801;
mixer gate_output_10_801(.a(output_11_801), .b(output_11_2), .y(output_10_801));
wire output_12_801, output_12_2, output_11_801;
mixer gate_output_11_801(.a(output_12_801), .b(output_12_2), .y(output_11_801));
wire output_13_801, output_13_2, output_12_801;
mixer gate_output_12_801(.a(output_13_801), .b(output_13_2), .y(output_12_801));
wire output_14_801, output_14_2, output_13_801;
mixer gate_output_13_801(.a(output_14_801), .b(output_14_2), .y(output_13_801));
wire output_15_801, output_15_2, output_14_801;
mixer gate_output_14_801(.a(output_15_801), .b(output_15_2), .y(output_14_801));
wire output_16_801, output_16_2, output_15_801;
mixer gate_output_15_801(.a(output_16_801), .b(output_16_2), .y(output_15_801));
wire output_1_802, output_1_3, output_0_802;
mixer gate_output_0_802(.a(output_1_802), .b(output_1_3), .y(output_0_802));
wire output_2_802, output_2_3, output_1_802;
mixer gate_output_1_802(.a(output_2_802), .b(output_2_3), .y(output_1_802));
wire output_3_802, output_3_3, output_2_802;
mixer gate_output_2_802(.a(output_3_802), .b(output_3_3), .y(output_2_802));
wire output_4_802, output_4_3, output_3_802;
mixer gate_output_3_802(.a(output_4_802), .b(output_4_3), .y(output_3_802));
wire output_5_802, output_5_3, output_4_802;
mixer gate_output_4_802(.a(output_5_802), .b(output_5_3), .y(output_4_802));
wire output_6_802, output_6_3, output_5_802;
mixer gate_output_5_802(.a(output_6_802), .b(output_6_3), .y(output_5_802));
wire output_7_802, output_7_3, output_6_802;
mixer gate_output_6_802(.a(output_7_802), .b(output_7_3), .y(output_6_802));
wire output_8_802, output_8_3, output_7_802;
mixer gate_output_7_802(.a(output_8_802), .b(output_8_3), .y(output_7_802));
wire output_9_802, output_9_3, output_8_802;
mixer gate_output_8_802(.a(output_9_802), .b(output_9_3), .y(output_8_802));
wire output_10_802, output_10_3, output_9_802;
mixer gate_output_9_802(.a(output_10_802), .b(output_10_3), .y(output_9_802));
wire output_11_802, output_11_3, output_10_802;
mixer gate_output_10_802(.a(output_11_802), .b(output_11_3), .y(output_10_802));
wire output_12_802, output_12_3, output_11_802;
mixer gate_output_11_802(.a(output_12_802), .b(output_12_3), .y(output_11_802));
wire output_13_802, output_13_3, output_12_802;
mixer gate_output_12_802(.a(output_13_802), .b(output_13_3), .y(output_12_802));
wire output_14_802, output_14_3, output_13_802;
mixer gate_output_13_802(.a(output_14_802), .b(output_14_3), .y(output_13_802));
wire output_15_802, output_15_3, output_14_802;
mixer gate_output_14_802(.a(output_15_802), .b(output_15_3), .y(output_14_802));
wire output_16_802, output_16_3, output_15_802;
mixer gate_output_15_802(.a(output_16_802), .b(output_16_3), .y(output_15_802));
wire output_1_803, output_1_4, output_0_803;
mixer gate_output_0_803(.a(output_1_803), .b(output_1_4), .y(output_0_803));
wire output_2_803, output_2_4, output_1_803;
mixer gate_output_1_803(.a(output_2_803), .b(output_2_4), .y(output_1_803));
wire output_3_803, output_3_4, output_2_803;
mixer gate_output_2_803(.a(output_3_803), .b(output_3_4), .y(output_2_803));
wire output_4_803, output_4_4, output_3_803;
mixer gate_output_3_803(.a(output_4_803), .b(output_4_4), .y(output_3_803));
wire output_5_803, output_5_4, output_4_803;
mixer gate_output_4_803(.a(output_5_803), .b(output_5_4), .y(output_4_803));
wire output_6_803, output_6_4, output_5_803;
mixer gate_output_5_803(.a(output_6_803), .b(output_6_4), .y(output_5_803));
wire output_7_803, output_7_4, output_6_803;
mixer gate_output_6_803(.a(output_7_803), .b(output_7_4), .y(output_6_803));
wire output_8_803, output_8_4, output_7_803;
mixer gate_output_7_803(.a(output_8_803), .b(output_8_4), .y(output_7_803));
wire output_9_803, output_9_4, output_8_803;
mixer gate_output_8_803(.a(output_9_803), .b(output_9_4), .y(output_8_803));
wire output_10_803, output_10_4, output_9_803;
mixer gate_output_9_803(.a(output_10_803), .b(output_10_4), .y(output_9_803));
wire output_11_803, output_11_4, output_10_803;
mixer gate_output_10_803(.a(output_11_803), .b(output_11_4), .y(output_10_803));
wire output_12_803, output_12_4, output_11_803;
mixer gate_output_11_803(.a(output_12_803), .b(output_12_4), .y(output_11_803));
wire output_13_803, output_13_4, output_12_803;
mixer gate_output_12_803(.a(output_13_803), .b(output_13_4), .y(output_12_803));
wire output_14_803, output_14_4, output_13_803;
mixer gate_output_13_803(.a(output_14_803), .b(output_14_4), .y(output_13_803));
wire output_15_803, output_15_4, output_14_803;
mixer gate_output_14_803(.a(output_15_803), .b(output_15_4), .y(output_14_803));
wire output_16_803, output_16_4, output_15_803;
mixer gate_output_15_803(.a(output_16_803), .b(output_16_4), .y(output_15_803));
wire output_1_804, output_1_5, output_0_804;
mixer gate_output_0_804(.a(output_1_804), .b(output_1_5), .y(output_0_804));
wire output_2_804, output_2_5, output_1_804;
mixer gate_output_1_804(.a(output_2_804), .b(output_2_5), .y(output_1_804));
wire output_3_804, output_3_5, output_2_804;
mixer gate_output_2_804(.a(output_3_804), .b(output_3_5), .y(output_2_804));
wire output_4_804, output_4_5, output_3_804;
mixer gate_output_3_804(.a(output_4_804), .b(output_4_5), .y(output_3_804));
wire output_5_804, output_5_5, output_4_804;
mixer gate_output_4_804(.a(output_5_804), .b(output_5_5), .y(output_4_804));
wire output_6_804, output_6_5, output_5_804;
mixer gate_output_5_804(.a(output_6_804), .b(output_6_5), .y(output_5_804));
wire output_7_804, output_7_5, output_6_804;
mixer gate_output_6_804(.a(output_7_804), .b(output_7_5), .y(output_6_804));
wire output_8_804, output_8_5, output_7_804;
mixer gate_output_7_804(.a(output_8_804), .b(output_8_5), .y(output_7_804));
wire output_9_804, output_9_5, output_8_804;
mixer gate_output_8_804(.a(output_9_804), .b(output_9_5), .y(output_8_804));
wire output_10_804, output_10_5, output_9_804;
mixer gate_output_9_804(.a(output_10_804), .b(output_10_5), .y(output_9_804));
wire output_11_804, output_11_5, output_10_804;
mixer gate_output_10_804(.a(output_11_804), .b(output_11_5), .y(output_10_804));
wire output_12_804, output_12_5, output_11_804;
mixer gate_output_11_804(.a(output_12_804), .b(output_12_5), .y(output_11_804));
wire output_13_804, output_13_5, output_12_804;
mixer gate_output_12_804(.a(output_13_804), .b(output_13_5), .y(output_12_804));
wire output_14_804, output_14_5, output_13_804;
mixer gate_output_13_804(.a(output_14_804), .b(output_14_5), .y(output_13_804));
wire output_15_804, output_15_5, output_14_804;
mixer gate_output_14_804(.a(output_15_804), .b(output_15_5), .y(output_14_804));
wire output_16_804, output_16_5, output_15_804;
mixer gate_output_15_804(.a(output_16_804), .b(output_16_5), .y(output_15_804));
wire output_1_805, output_1_6, output_0_805;
mixer gate_output_0_805(.a(output_1_805), .b(output_1_6), .y(output_0_805));
wire output_2_805, output_2_6, output_1_805;
mixer gate_output_1_805(.a(output_2_805), .b(output_2_6), .y(output_1_805));
wire output_3_805, output_3_6, output_2_805;
mixer gate_output_2_805(.a(output_3_805), .b(output_3_6), .y(output_2_805));
wire output_4_805, output_4_6, output_3_805;
mixer gate_output_3_805(.a(output_4_805), .b(output_4_6), .y(output_3_805));
wire output_5_805, output_5_6, output_4_805;
mixer gate_output_4_805(.a(output_5_805), .b(output_5_6), .y(output_4_805));
wire output_6_805, output_6_6, output_5_805;
mixer gate_output_5_805(.a(output_6_805), .b(output_6_6), .y(output_5_805));
wire output_7_805, output_7_6, output_6_805;
mixer gate_output_6_805(.a(output_7_805), .b(output_7_6), .y(output_6_805));
wire output_8_805, output_8_6, output_7_805;
mixer gate_output_7_805(.a(output_8_805), .b(output_8_6), .y(output_7_805));
wire output_9_805, output_9_6, output_8_805;
mixer gate_output_8_805(.a(output_9_805), .b(output_9_6), .y(output_8_805));
wire output_10_805, output_10_6, output_9_805;
mixer gate_output_9_805(.a(output_10_805), .b(output_10_6), .y(output_9_805));
wire output_11_805, output_11_6, output_10_805;
mixer gate_output_10_805(.a(output_11_805), .b(output_11_6), .y(output_10_805));
wire output_12_805, output_12_6, output_11_805;
mixer gate_output_11_805(.a(output_12_805), .b(output_12_6), .y(output_11_805));
wire output_13_805, output_13_6, output_12_805;
mixer gate_output_12_805(.a(output_13_805), .b(output_13_6), .y(output_12_805));
wire output_14_805, output_14_6, output_13_805;
mixer gate_output_13_805(.a(output_14_805), .b(output_14_6), .y(output_13_805));
wire output_15_805, output_15_6, output_14_805;
mixer gate_output_14_805(.a(output_15_805), .b(output_15_6), .y(output_14_805));
wire output_16_805, output_16_6, output_15_805;
mixer gate_output_15_805(.a(output_16_805), .b(output_16_6), .y(output_15_805));
wire output_1_806, output_1_7, output_0_806;
mixer gate_output_0_806(.a(output_1_806), .b(output_1_7), .y(output_0_806));
wire output_2_806, output_2_7, output_1_806;
mixer gate_output_1_806(.a(output_2_806), .b(output_2_7), .y(output_1_806));
wire output_3_806, output_3_7, output_2_806;
mixer gate_output_2_806(.a(output_3_806), .b(output_3_7), .y(output_2_806));
wire output_4_806, output_4_7, output_3_806;
mixer gate_output_3_806(.a(output_4_806), .b(output_4_7), .y(output_3_806));
wire output_5_806, output_5_7, output_4_806;
mixer gate_output_4_806(.a(output_5_806), .b(output_5_7), .y(output_4_806));
wire output_6_806, output_6_7, output_5_806;
mixer gate_output_5_806(.a(output_6_806), .b(output_6_7), .y(output_5_806));
wire output_7_806, output_7_7, output_6_806;
mixer gate_output_6_806(.a(output_7_806), .b(output_7_7), .y(output_6_806));
wire output_8_806, output_8_7, output_7_806;
mixer gate_output_7_806(.a(output_8_806), .b(output_8_7), .y(output_7_806));
wire output_9_806, output_9_7, output_8_806;
mixer gate_output_8_806(.a(output_9_806), .b(output_9_7), .y(output_8_806));
wire output_10_806, output_10_7, output_9_806;
mixer gate_output_9_806(.a(output_10_806), .b(output_10_7), .y(output_9_806));
wire output_11_806, output_11_7, output_10_806;
mixer gate_output_10_806(.a(output_11_806), .b(output_11_7), .y(output_10_806));
wire output_12_806, output_12_7, output_11_806;
mixer gate_output_11_806(.a(output_12_806), .b(output_12_7), .y(output_11_806));
wire output_13_806, output_13_7, output_12_806;
mixer gate_output_12_806(.a(output_13_806), .b(output_13_7), .y(output_12_806));
wire output_14_806, output_14_7, output_13_806;
mixer gate_output_13_806(.a(output_14_806), .b(output_14_7), .y(output_13_806));
wire output_15_806, output_15_7, output_14_806;
mixer gate_output_14_806(.a(output_15_806), .b(output_15_7), .y(output_14_806));
wire output_16_806, output_16_7, output_15_806;
mixer gate_output_15_806(.a(output_16_806), .b(output_16_7), .y(output_15_806));
wire output_1_807, output_1_8, output_0_807;
mixer gate_output_0_807(.a(output_1_807), .b(output_1_8), .y(output_0_807));
wire output_2_807, output_2_8, output_1_807;
mixer gate_output_1_807(.a(output_2_807), .b(output_2_8), .y(output_1_807));
wire output_3_807, output_3_8, output_2_807;
mixer gate_output_2_807(.a(output_3_807), .b(output_3_8), .y(output_2_807));
wire output_4_807, output_4_8, output_3_807;
mixer gate_output_3_807(.a(output_4_807), .b(output_4_8), .y(output_3_807));
wire output_5_807, output_5_8, output_4_807;
mixer gate_output_4_807(.a(output_5_807), .b(output_5_8), .y(output_4_807));
wire output_6_807, output_6_8, output_5_807;
mixer gate_output_5_807(.a(output_6_807), .b(output_6_8), .y(output_5_807));
wire output_7_807, output_7_8, output_6_807;
mixer gate_output_6_807(.a(output_7_807), .b(output_7_8), .y(output_6_807));
wire output_8_807, output_8_8, output_7_807;
mixer gate_output_7_807(.a(output_8_807), .b(output_8_8), .y(output_7_807));
wire output_9_807, output_9_8, output_8_807;
mixer gate_output_8_807(.a(output_9_807), .b(output_9_8), .y(output_8_807));
wire output_10_807, output_10_8, output_9_807;
mixer gate_output_9_807(.a(output_10_807), .b(output_10_8), .y(output_9_807));
wire output_11_807, output_11_8, output_10_807;
mixer gate_output_10_807(.a(output_11_807), .b(output_11_8), .y(output_10_807));
wire output_12_807, output_12_8, output_11_807;
mixer gate_output_11_807(.a(output_12_807), .b(output_12_8), .y(output_11_807));
wire output_13_807, output_13_8, output_12_807;
mixer gate_output_12_807(.a(output_13_807), .b(output_13_8), .y(output_12_807));
wire output_14_807, output_14_8, output_13_807;
mixer gate_output_13_807(.a(output_14_807), .b(output_14_8), .y(output_13_807));
wire output_15_807, output_15_8, output_14_807;
mixer gate_output_14_807(.a(output_15_807), .b(output_15_8), .y(output_14_807));
wire output_16_807, output_16_8, output_15_807;
mixer gate_output_15_807(.a(output_16_807), .b(output_16_8), .y(output_15_807));
wire output_1_808, output_1_9, output_0_808;
mixer gate_output_0_808(.a(output_1_808), .b(output_1_9), .y(output_0_808));
wire output_2_808, output_2_9, output_1_808;
mixer gate_output_1_808(.a(output_2_808), .b(output_2_9), .y(output_1_808));
wire output_3_808, output_3_9, output_2_808;
mixer gate_output_2_808(.a(output_3_808), .b(output_3_9), .y(output_2_808));
wire output_4_808, output_4_9, output_3_808;
mixer gate_output_3_808(.a(output_4_808), .b(output_4_9), .y(output_3_808));
wire output_5_808, output_5_9, output_4_808;
mixer gate_output_4_808(.a(output_5_808), .b(output_5_9), .y(output_4_808));
wire output_6_808, output_6_9, output_5_808;
mixer gate_output_5_808(.a(output_6_808), .b(output_6_9), .y(output_5_808));
wire output_7_808, output_7_9, output_6_808;
mixer gate_output_6_808(.a(output_7_808), .b(output_7_9), .y(output_6_808));
wire output_8_808, output_8_9, output_7_808;
mixer gate_output_7_808(.a(output_8_808), .b(output_8_9), .y(output_7_808));
wire output_9_808, output_9_9, output_8_808;
mixer gate_output_8_808(.a(output_9_808), .b(output_9_9), .y(output_8_808));
wire output_10_808, output_10_9, output_9_808;
mixer gate_output_9_808(.a(output_10_808), .b(output_10_9), .y(output_9_808));
wire output_11_808, output_11_9, output_10_808;
mixer gate_output_10_808(.a(output_11_808), .b(output_11_9), .y(output_10_808));
wire output_12_808, output_12_9, output_11_808;
mixer gate_output_11_808(.a(output_12_808), .b(output_12_9), .y(output_11_808));
wire output_13_808, output_13_9, output_12_808;
mixer gate_output_12_808(.a(output_13_808), .b(output_13_9), .y(output_12_808));
wire output_14_808, output_14_9, output_13_808;
mixer gate_output_13_808(.a(output_14_808), .b(output_14_9), .y(output_13_808));
wire output_15_808, output_15_9, output_14_808;
mixer gate_output_14_808(.a(output_15_808), .b(output_15_9), .y(output_14_808));
wire output_16_808, output_16_9, output_15_808;
mixer gate_output_15_808(.a(output_16_808), .b(output_16_9), .y(output_15_808));
wire output_1_809, output_1_10, output_0_809;
mixer gate_output_0_809(.a(output_1_809), .b(output_1_10), .y(output_0_809));
wire output_2_809, output_2_10, output_1_809;
mixer gate_output_1_809(.a(output_2_809), .b(output_2_10), .y(output_1_809));
wire output_3_809, output_3_10, output_2_809;
mixer gate_output_2_809(.a(output_3_809), .b(output_3_10), .y(output_2_809));
wire output_4_809, output_4_10, output_3_809;
mixer gate_output_3_809(.a(output_4_809), .b(output_4_10), .y(output_3_809));
wire output_5_809, output_5_10, output_4_809;
mixer gate_output_4_809(.a(output_5_809), .b(output_5_10), .y(output_4_809));
wire output_6_809, output_6_10, output_5_809;
mixer gate_output_5_809(.a(output_6_809), .b(output_6_10), .y(output_5_809));
wire output_7_809, output_7_10, output_6_809;
mixer gate_output_6_809(.a(output_7_809), .b(output_7_10), .y(output_6_809));
wire output_8_809, output_8_10, output_7_809;
mixer gate_output_7_809(.a(output_8_809), .b(output_8_10), .y(output_7_809));
wire output_9_809, output_9_10, output_8_809;
mixer gate_output_8_809(.a(output_9_809), .b(output_9_10), .y(output_8_809));
wire output_10_809, output_10_10, output_9_809;
mixer gate_output_9_809(.a(output_10_809), .b(output_10_10), .y(output_9_809));
wire output_11_809, output_11_10, output_10_809;
mixer gate_output_10_809(.a(output_11_809), .b(output_11_10), .y(output_10_809));
wire output_12_809, output_12_10, output_11_809;
mixer gate_output_11_809(.a(output_12_809), .b(output_12_10), .y(output_11_809));
wire output_13_809, output_13_10, output_12_809;
mixer gate_output_12_809(.a(output_13_809), .b(output_13_10), .y(output_12_809));
wire output_14_809, output_14_10, output_13_809;
mixer gate_output_13_809(.a(output_14_809), .b(output_14_10), .y(output_13_809));
wire output_15_809, output_15_10, output_14_809;
mixer gate_output_14_809(.a(output_15_809), .b(output_15_10), .y(output_14_809));
wire output_16_809, output_16_10, output_15_809;
mixer gate_output_15_809(.a(output_16_809), .b(output_16_10), .y(output_15_809));
wire output_1_810, output_1_11, output_0_810;
mixer gate_output_0_810(.a(output_1_810), .b(output_1_11), .y(output_0_810));
wire output_2_810, output_2_11, output_1_810;
mixer gate_output_1_810(.a(output_2_810), .b(output_2_11), .y(output_1_810));
wire output_3_810, output_3_11, output_2_810;
mixer gate_output_2_810(.a(output_3_810), .b(output_3_11), .y(output_2_810));
wire output_4_810, output_4_11, output_3_810;
mixer gate_output_3_810(.a(output_4_810), .b(output_4_11), .y(output_3_810));
wire output_5_810, output_5_11, output_4_810;
mixer gate_output_4_810(.a(output_5_810), .b(output_5_11), .y(output_4_810));
wire output_6_810, output_6_11, output_5_810;
mixer gate_output_5_810(.a(output_6_810), .b(output_6_11), .y(output_5_810));
wire output_7_810, output_7_11, output_6_810;
mixer gate_output_6_810(.a(output_7_810), .b(output_7_11), .y(output_6_810));
wire output_8_810, output_8_11, output_7_810;
mixer gate_output_7_810(.a(output_8_810), .b(output_8_11), .y(output_7_810));
wire output_9_810, output_9_11, output_8_810;
mixer gate_output_8_810(.a(output_9_810), .b(output_9_11), .y(output_8_810));
wire output_10_810, output_10_11, output_9_810;
mixer gate_output_9_810(.a(output_10_810), .b(output_10_11), .y(output_9_810));
wire output_11_810, output_11_11, output_10_810;
mixer gate_output_10_810(.a(output_11_810), .b(output_11_11), .y(output_10_810));
wire output_12_810, output_12_11, output_11_810;
mixer gate_output_11_810(.a(output_12_810), .b(output_12_11), .y(output_11_810));
wire output_13_810, output_13_11, output_12_810;
mixer gate_output_12_810(.a(output_13_810), .b(output_13_11), .y(output_12_810));
wire output_14_810, output_14_11, output_13_810;
mixer gate_output_13_810(.a(output_14_810), .b(output_14_11), .y(output_13_810));
wire output_15_810, output_15_11, output_14_810;
mixer gate_output_14_810(.a(output_15_810), .b(output_15_11), .y(output_14_810));
wire output_16_810, output_16_11, output_15_810;
mixer gate_output_15_810(.a(output_16_810), .b(output_16_11), .y(output_15_810));
wire output_1_811, output_1_12, output_0_811;
mixer gate_output_0_811(.a(output_1_811), .b(output_1_12), .y(output_0_811));
wire output_2_811, output_2_12, output_1_811;
mixer gate_output_1_811(.a(output_2_811), .b(output_2_12), .y(output_1_811));
wire output_3_811, output_3_12, output_2_811;
mixer gate_output_2_811(.a(output_3_811), .b(output_3_12), .y(output_2_811));
wire output_4_811, output_4_12, output_3_811;
mixer gate_output_3_811(.a(output_4_811), .b(output_4_12), .y(output_3_811));
wire output_5_811, output_5_12, output_4_811;
mixer gate_output_4_811(.a(output_5_811), .b(output_5_12), .y(output_4_811));
wire output_6_811, output_6_12, output_5_811;
mixer gate_output_5_811(.a(output_6_811), .b(output_6_12), .y(output_5_811));
wire output_7_811, output_7_12, output_6_811;
mixer gate_output_6_811(.a(output_7_811), .b(output_7_12), .y(output_6_811));
wire output_8_811, output_8_12, output_7_811;
mixer gate_output_7_811(.a(output_8_811), .b(output_8_12), .y(output_7_811));
wire output_9_811, output_9_12, output_8_811;
mixer gate_output_8_811(.a(output_9_811), .b(output_9_12), .y(output_8_811));
wire output_10_811, output_10_12, output_9_811;
mixer gate_output_9_811(.a(output_10_811), .b(output_10_12), .y(output_9_811));
wire output_11_811, output_11_12, output_10_811;
mixer gate_output_10_811(.a(output_11_811), .b(output_11_12), .y(output_10_811));
wire output_12_811, output_12_12, output_11_811;
mixer gate_output_11_811(.a(output_12_811), .b(output_12_12), .y(output_11_811));
wire output_13_811, output_13_12, output_12_811;
mixer gate_output_12_811(.a(output_13_811), .b(output_13_12), .y(output_12_811));
wire output_14_811, output_14_12, output_13_811;
mixer gate_output_13_811(.a(output_14_811), .b(output_14_12), .y(output_13_811));
wire output_15_811, output_15_12, output_14_811;
mixer gate_output_14_811(.a(output_15_811), .b(output_15_12), .y(output_14_811));
wire output_16_811, output_16_12, output_15_811;
mixer gate_output_15_811(.a(output_16_811), .b(output_16_12), .y(output_15_811));
wire output_1_812, output_1_13, output_0_812;
mixer gate_output_0_812(.a(output_1_812), .b(output_1_13), .y(output_0_812));
wire output_2_812, output_2_13, output_1_812;
mixer gate_output_1_812(.a(output_2_812), .b(output_2_13), .y(output_1_812));
wire output_3_812, output_3_13, output_2_812;
mixer gate_output_2_812(.a(output_3_812), .b(output_3_13), .y(output_2_812));
wire output_4_812, output_4_13, output_3_812;
mixer gate_output_3_812(.a(output_4_812), .b(output_4_13), .y(output_3_812));
wire output_5_812, output_5_13, output_4_812;
mixer gate_output_4_812(.a(output_5_812), .b(output_5_13), .y(output_4_812));
wire output_6_812, output_6_13, output_5_812;
mixer gate_output_5_812(.a(output_6_812), .b(output_6_13), .y(output_5_812));
wire output_7_812, output_7_13, output_6_812;
mixer gate_output_6_812(.a(output_7_812), .b(output_7_13), .y(output_6_812));
wire output_8_812, output_8_13, output_7_812;
mixer gate_output_7_812(.a(output_8_812), .b(output_8_13), .y(output_7_812));
wire output_9_812, output_9_13, output_8_812;
mixer gate_output_8_812(.a(output_9_812), .b(output_9_13), .y(output_8_812));
wire output_10_812, output_10_13, output_9_812;
mixer gate_output_9_812(.a(output_10_812), .b(output_10_13), .y(output_9_812));
wire output_11_812, output_11_13, output_10_812;
mixer gate_output_10_812(.a(output_11_812), .b(output_11_13), .y(output_10_812));
wire output_12_812, output_12_13, output_11_812;
mixer gate_output_11_812(.a(output_12_812), .b(output_12_13), .y(output_11_812));
wire output_13_812, output_13_13, output_12_812;
mixer gate_output_12_812(.a(output_13_812), .b(output_13_13), .y(output_12_812));
wire output_14_812, output_14_13, output_13_812;
mixer gate_output_13_812(.a(output_14_812), .b(output_14_13), .y(output_13_812));
wire output_15_812, output_15_13, output_14_812;
mixer gate_output_14_812(.a(output_15_812), .b(output_15_13), .y(output_14_812));
wire output_16_812, output_16_13, output_15_812;
mixer gate_output_15_812(.a(output_16_812), .b(output_16_13), .y(output_15_812));
wire output_1_813, output_1_14, output_0_813;
mixer gate_output_0_813(.a(output_1_813), .b(output_1_14), .y(output_0_813));
wire output_2_813, output_2_14, output_1_813;
mixer gate_output_1_813(.a(output_2_813), .b(output_2_14), .y(output_1_813));
wire output_3_813, output_3_14, output_2_813;
mixer gate_output_2_813(.a(output_3_813), .b(output_3_14), .y(output_2_813));
wire output_4_813, output_4_14, output_3_813;
mixer gate_output_3_813(.a(output_4_813), .b(output_4_14), .y(output_3_813));
wire output_5_813, output_5_14, output_4_813;
mixer gate_output_4_813(.a(output_5_813), .b(output_5_14), .y(output_4_813));
wire output_6_813, output_6_14, output_5_813;
mixer gate_output_5_813(.a(output_6_813), .b(output_6_14), .y(output_5_813));
wire output_7_813, output_7_14, output_6_813;
mixer gate_output_6_813(.a(output_7_813), .b(output_7_14), .y(output_6_813));
wire output_8_813, output_8_14, output_7_813;
mixer gate_output_7_813(.a(output_8_813), .b(output_8_14), .y(output_7_813));
wire output_9_813, output_9_14, output_8_813;
mixer gate_output_8_813(.a(output_9_813), .b(output_9_14), .y(output_8_813));
wire output_10_813, output_10_14, output_9_813;
mixer gate_output_9_813(.a(output_10_813), .b(output_10_14), .y(output_9_813));
wire output_11_813, output_11_14, output_10_813;
mixer gate_output_10_813(.a(output_11_813), .b(output_11_14), .y(output_10_813));
wire output_12_813, output_12_14, output_11_813;
mixer gate_output_11_813(.a(output_12_813), .b(output_12_14), .y(output_11_813));
wire output_13_813, output_13_14, output_12_813;
mixer gate_output_12_813(.a(output_13_813), .b(output_13_14), .y(output_12_813));
wire output_14_813, output_14_14, output_13_813;
mixer gate_output_13_813(.a(output_14_813), .b(output_14_14), .y(output_13_813));
wire output_15_813, output_15_14, output_14_813;
mixer gate_output_14_813(.a(output_15_813), .b(output_15_14), .y(output_14_813));
wire output_16_813, output_16_14, output_15_813;
mixer gate_output_15_813(.a(output_16_813), .b(output_16_14), .y(output_15_813));
wire output_1_814, output_1_15, output_0_814;
mixer gate_output_0_814(.a(output_1_814), .b(output_1_15), .y(output_0_814));
wire output_2_814, output_2_15, output_1_814;
mixer gate_output_1_814(.a(output_2_814), .b(output_2_15), .y(output_1_814));
wire output_3_814, output_3_15, output_2_814;
mixer gate_output_2_814(.a(output_3_814), .b(output_3_15), .y(output_2_814));
wire output_4_814, output_4_15, output_3_814;
mixer gate_output_3_814(.a(output_4_814), .b(output_4_15), .y(output_3_814));
wire output_5_814, output_5_15, output_4_814;
mixer gate_output_4_814(.a(output_5_814), .b(output_5_15), .y(output_4_814));
wire output_6_814, output_6_15, output_5_814;
mixer gate_output_5_814(.a(output_6_814), .b(output_6_15), .y(output_5_814));
wire output_7_814, output_7_15, output_6_814;
mixer gate_output_6_814(.a(output_7_814), .b(output_7_15), .y(output_6_814));
wire output_8_814, output_8_15, output_7_814;
mixer gate_output_7_814(.a(output_8_814), .b(output_8_15), .y(output_7_814));
wire output_9_814, output_9_15, output_8_814;
mixer gate_output_8_814(.a(output_9_814), .b(output_9_15), .y(output_8_814));
wire output_10_814, output_10_15, output_9_814;
mixer gate_output_9_814(.a(output_10_814), .b(output_10_15), .y(output_9_814));
wire output_11_814, output_11_15, output_10_814;
mixer gate_output_10_814(.a(output_11_814), .b(output_11_15), .y(output_10_814));
wire output_12_814, output_12_15, output_11_814;
mixer gate_output_11_814(.a(output_12_814), .b(output_12_15), .y(output_11_814));
wire output_13_814, output_13_15, output_12_814;
mixer gate_output_12_814(.a(output_13_814), .b(output_13_15), .y(output_12_814));
wire output_14_814, output_14_15, output_13_814;
mixer gate_output_13_814(.a(output_14_814), .b(output_14_15), .y(output_13_814));
wire output_15_814, output_15_15, output_14_814;
mixer gate_output_14_814(.a(output_15_814), .b(output_15_15), .y(output_14_814));
wire output_16_814, output_16_15, output_15_814;
mixer gate_output_15_814(.a(output_16_814), .b(output_16_15), .y(output_15_814));
wire output_1_815, output_1_0, output_0_815;
mixer gate_output_0_815(.a(output_1_815), .b(output_1_0), .y(output_0_815));
wire output_2_815, output_2_0, output_1_815;
mixer gate_output_1_815(.a(output_2_815), .b(output_2_0), .y(output_1_815));
wire output_3_815, output_3_0, output_2_815;
mixer gate_output_2_815(.a(output_3_815), .b(output_3_0), .y(output_2_815));
wire output_4_815, output_4_0, output_3_815;
mixer gate_output_3_815(.a(output_4_815), .b(output_4_0), .y(output_3_815));
wire output_5_815, output_5_0, output_4_815;
mixer gate_output_4_815(.a(output_5_815), .b(output_5_0), .y(output_4_815));
wire output_6_815, output_6_0, output_5_815;
mixer gate_output_5_815(.a(output_6_815), .b(output_6_0), .y(output_5_815));
wire output_7_815, output_7_0, output_6_815;
mixer gate_output_6_815(.a(output_7_815), .b(output_7_0), .y(output_6_815));
wire output_8_815, output_8_0, output_7_815;
mixer gate_output_7_815(.a(output_8_815), .b(output_8_0), .y(output_7_815));
wire output_9_815, output_9_0, output_8_815;
mixer gate_output_8_815(.a(output_9_815), .b(output_9_0), .y(output_8_815));
wire output_10_815, output_10_0, output_9_815;
mixer gate_output_9_815(.a(output_10_815), .b(output_10_0), .y(output_9_815));
wire output_11_815, output_11_0, output_10_815;
mixer gate_output_10_815(.a(output_11_815), .b(output_11_0), .y(output_10_815));
wire output_12_815, output_12_0, output_11_815;
mixer gate_output_11_815(.a(output_12_815), .b(output_12_0), .y(output_11_815));
wire output_13_815, output_13_0, output_12_815;
mixer gate_output_12_815(.a(output_13_815), .b(output_13_0), .y(output_12_815));
wire output_14_815, output_14_0, output_13_815;
mixer gate_output_13_815(.a(output_14_815), .b(output_14_0), .y(output_13_815));
wire output_15_815, output_15_0, output_14_815;
mixer gate_output_14_815(.a(output_15_815), .b(output_15_0), .y(output_14_815));
wire output_16_815, output_16_0, output_15_815;
mixer gate_output_15_815(.a(output_16_815), .b(output_16_0), .y(output_15_815));
wire output_1_816, output_1_1, output_0_816;
mixer gate_output_0_816(.a(output_1_816), .b(output_1_1), .y(output_0_816));
wire output_2_816, output_2_1, output_1_816;
mixer gate_output_1_816(.a(output_2_816), .b(output_2_1), .y(output_1_816));
wire output_3_816, output_3_1, output_2_816;
mixer gate_output_2_816(.a(output_3_816), .b(output_3_1), .y(output_2_816));
wire output_4_816, output_4_1, output_3_816;
mixer gate_output_3_816(.a(output_4_816), .b(output_4_1), .y(output_3_816));
wire output_5_816, output_5_1, output_4_816;
mixer gate_output_4_816(.a(output_5_816), .b(output_5_1), .y(output_4_816));
wire output_6_816, output_6_1, output_5_816;
mixer gate_output_5_816(.a(output_6_816), .b(output_6_1), .y(output_5_816));
wire output_7_816, output_7_1, output_6_816;
mixer gate_output_6_816(.a(output_7_816), .b(output_7_1), .y(output_6_816));
wire output_8_816, output_8_1, output_7_816;
mixer gate_output_7_816(.a(output_8_816), .b(output_8_1), .y(output_7_816));
wire output_9_816, output_9_1, output_8_816;
mixer gate_output_8_816(.a(output_9_816), .b(output_9_1), .y(output_8_816));
wire output_10_816, output_10_1, output_9_816;
mixer gate_output_9_816(.a(output_10_816), .b(output_10_1), .y(output_9_816));
wire output_11_816, output_11_1, output_10_816;
mixer gate_output_10_816(.a(output_11_816), .b(output_11_1), .y(output_10_816));
wire output_12_816, output_12_1, output_11_816;
mixer gate_output_11_816(.a(output_12_816), .b(output_12_1), .y(output_11_816));
wire output_13_816, output_13_1, output_12_816;
mixer gate_output_12_816(.a(output_13_816), .b(output_13_1), .y(output_12_816));
wire output_14_816, output_14_1, output_13_816;
mixer gate_output_13_816(.a(output_14_816), .b(output_14_1), .y(output_13_816));
wire output_15_816, output_15_1, output_14_816;
mixer gate_output_14_816(.a(output_15_816), .b(output_15_1), .y(output_14_816));
wire output_16_816, output_16_1, output_15_816;
mixer gate_output_15_816(.a(output_16_816), .b(output_16_1), .y(output_15_816));
wire output_1_817, output_1_2, output_0_817;
mixer gate_output_0_817(.a(output_1_817), .b(output_1_2), .y(output_0_817));
wire output_2_817, output_2_2, output_1_817;
mixer gate_output_1_817(.a(output_2_817), .b(output_2_2), .y(output_1_817));
wire output_3_817, output_3_2, output_2_817;
mixer gate_output_2_817(.a(output_3_817), .b(output_3_2), .y(output_2_817));
wire output_4_817, output_4_2, output_3_817;
mixer gate_output_3_817(.a(output_4_817), .b(output_4_2), .y(output_3_817));
wire output_5_817, output_5_2, output_4_817;
mixer gate_output_4_817(.a(output_5_817), .b(output_5_2), .y(output_4_817));
wire output_6_817, output_6_2, output_5_817;
mixer gate_output_5_817(.a(output_6_817), .b(output_6_2), .y(output_5_817));
wire output_7_817, output_7_2, output_6_817;
mixer gate_output_6_817(.a(output_7_817), .b(output_7_2), .y(output_6_817));
wire output_8_817, output_8_2, output_7_817;
mixer gate_output_7_817(.a(output_8_817), .b(output_8_2), .y(output_7_817));
wire output_9_817, output_9_2, output_8_817;
mixer gate_output_8_817(.a(output_9_817), .b(output_9_2), .y(output_8_817));
wire output_10_817, output_10_2, output_9_817;
mixer gate_output_9_817(.a(output_10_817), .b(output_10_2), .y(output_9_817));
wire output_11_817, output_11_2, output_10_817;
mixer gate_output_10_817(.a(output_11_817), .b(output_11_2), .y(output_10_817));
wire output_12_817, output_12_2, output_11_817;
mixer gate_output_11_817(.a(output_12_817), .b(output_12_2), .y(output_11_817));
wire output_13_817, output_13_2, output_12_817;
mixer gate_output_12_817(.a(output_13_817), .b(output_13_2), .y(output_12_817));
wire output_14_817, output_14_2, output_13_817;
mixer gate_output_13_817(.a(output_14_817), .b(output_14_2), .y(output_13_817));
wire output_15_817, output_15_2, output_14_817;
mixer gate_output_14_817(.a(output_15_817), .b(output_15_2), .y(output_14_817));
wire output_16_817, output_16_2, output_15_817;
mixer gate_output_15_817(.a(output_16_817), .b(output_16_2), .y(output_15_817));
wire output_1_818, output_1_3, output_0_818;
mixer gate_output_0_818(.a(output_1_818), .b(output_1_3), .y(output_0_818));
wire output_2_818, output_2_3, output_1_818;
mixer gate_output_1_818(.a(output_2_818), .b(output_2_3), .y(output_1_818));
wire output_3_818, output_3_3, output_2_818;
mixer gate_output_2_818(.a(output_3_818), .b(output_3_3), .y(output_2_818));
wire output_4_818, output_4_3, output_3_818;
mixer gate_output_3_818(.a(output_4_818), .b(output_4_3), .y(output_3_818));
wire output_5_818, output_5_3, output_4_818;
mixer gate_output_4_818(.a(output_5_818), .b(output_5_3), .y(output_4_818));
wire output_6_818, output_6_3, output_5_818;
mixer gate_output_5_818(.a(output_6_818), .b(output_6_3), .y(output_5_818));
wire output_7_818, output_7_3, output_6_818;
mixer gate_output_6_818(.a(output_7_818), .b(output_7_3), .y(output_6_818));
wire output_8_818, output_8_3, output_7_818;
mixer gate_output_7_818(.a(output_8_818), .b(output_8_3), .y(output_7_818));
wire output_9_818, output_9_3, output_8_818;
mixer gate_output_8_818(.a(output_9_818), .b(output_9_3), .y(output_8_818));
wire output_10_818, output_10_3, output_9_818;
mixer gate_output_9_818(.a(output_10_818), .b(output_10_3), .y(output_9_818));
wire output_11_818, output_11_3, output_10_818;
mixer gate_output_10_818(.a(output_11_818), .b(output_11_3), .y(output_10_818));
wire output_12_818, output_12_3, output_11_818;
mixer gate_output_11_818(.a(output_12_818), .b(output_12_3), .y(output_11_818));
wire output_13_818, output_13_3, output_12_818;
mixer gate_output_12_818(.a(output_13_818), .b(output_13_3), .y(output_12_818));
wire output_14_818, output_14_3, output_13_818;
mixer gate_output_13_818(.a(output_14_818), .b(output_14_3), .y(output_13_818));
wire output_15_818, output_15_3, output_14_818;
mixer gate_output_14_818(.a(output_15_818), .b(output_15_3), .y(output_14_818));
wire output_16_818, output_16_3, output_15_818;
mixer gate_output_15_818(.a(output_16_818), .b(output_16_3), .y(output_15_818));
wire output_1_819, output_1_4, output_0_819;
mixer gate_output_0_819(.a(output_1_819), .b(output_1_4), .y(output_0_819));
wire output_2_819, output_2_4, output_1_819;
mixer gate_output_1_819(.a(output_2_819), .b(output_2_4), .y(output_1_819));
wire output_3_819, output_3_4, output_2_819;
mixer gate_output_2_819(.a(output_3_819), .b(output_3_4), .y(output_2_819));
wire output_4_819, output_4_4, output_3_819;
mixer gate_output_3_819(.a(output_4_819), .b(output_4_4), .y(output_3_819));
wire output_5_819, output_5_4, output_4_819;
mixer gate_output_4_819(.a(output_5_819), .b(output_5_4), .y(output_4_819));
wire output_6_819, output_6_4, output_5_819;
mixer gate_output_5_819(.a(output_6_819), .b(output_6_4), .y(output_5_819));
wire output_7_819, output_7_4, output_6_819;
mixer gate_output_6_819(.a(output_7_819), .b(output_7_4), .y(output_6_819));
wire output_8_819, output_8_4, output_7_819;
mixer gate_output_7_819(.a(output_8_819), .b(output_8_4), .y(output_7_819));
wire output_9_819, output_9_4, output_8_819;
mixer gate_output_8_819(.a(output_9_819), .b(output_9_4), .y(output_8_819));
wire output_10_819, output_10_4, output_9_819;
mixer gate_output_9_819(.a(output_10_819), .b(output_10_4), .y(output_9_819));
wire output_11_819, output_11_4, output_10_819;
mixer gate_output_10_819(.a(output_11_819), .b(output_11_4), .y(output_10_819));
wire output_12_819, output_12_4, output_11_819;
mixer gate_output_11_819(.a(output_12_819), .b(output_12_4), .y(output_11_819));
wire output_13_819, output_13_4, output_12_819;
mixer gate_output_12_819(.a(output_13_819), .b(output_13_4), .y(output_12_819));
wire output_14_819, output_14_4, output_13_819;
mixer gate_output_13_819(.a(output_14_819), .b(output_14_4), .y(output_13_819));
wire output_15_819, output_15_4, output_14_819;
mixer gate_output_14_819(.a(output_15_819), .b(output_15_4), .y(output_14_819));
wire output_16_819, output_16_4, output_15_819;
mixer gate_output_15_819(.a(output_16_819), .b(output_16_4), .y(output_15_819));
wire output_1_820, output_1_5, output_0_820;
mixer gate_output_0_820(.a(output_1_820), .b(output_1_5), .y(output_0_820));
wire output_2_820, output_2_5, output_1_820;
mixer gate_output_1_820(.a(output_2_820), .b(output_2_5), .y(output_1_820));
wire output_3_820, output_3_5, output_2_820;
mixer gate_output_2_820(.a(output_3_820), .b(output_3_5), .y(output_2_820));
wire output_4_820, output_4_5, output_3_820;
mixer gate_output_3_820(.a(output_4_820), .b(output_4_5), .y(output_3_820));
wire output_5_820, output_5_5, output_4_820;
mixer gate_output_4_820(.a(output_5_820), .b(output_5_5), .y(output_4_820));
wire output_6_820, output_6_5, output_5_820;
mixer gate_output_5_820(.a(output_6_820), .b(output_6_5), .y(output_5_820));
wire output_7_820, output_7_5, output_6_820;
mixer gate_output_6_820(.a(output_7_820), .b(output_7_5), .y(output_6_820));
wire output_8_820, output_8_5, output_7_820;
mixer gate_output_7_820(.a(output_8_820), .b(output_8_5), .y(output_7_820));
wire output_9_820, output_9_5, output_8_820;
mixer gate_output_8_820(.a(output_9_820), .b(output_9_5), .y(output_8_820));
wire output_10_820, output_10_5, output_9_820;
mixer gate_output_9_820(.a(output_10_820), .b(output_10_5), .y(output_9_820));
wire output_11_820, output_11_5, output_10_820;
mixer gate_output_10_820(.a(output_11_820), .b(output_11_5), .y(output_10_820));
wire output_12_820, output_12_5, output_11_820;
mixer gate_output_11_820(.a(output_12_820), .b(output_12_5), .y(output_11_820));
wire output_13_820, output_13_5, output_12_820;
mixer gate_output_12_820(.a(output_13_820), .b(output_13_5), .y(output_12_820));
wire output_14_820, output_14_5, output_13_820;
mixer gate_output_13_820(.a(output_14_820), .b(output_14_5), .y(output_13_820));
wire output_15_820, output_15_5, output_14_820;
mixer gate_output_14_820(.a(output_15_820), .b(output_15_5), .y(output_14_820));
wire output_16_820, output_16_5, output_15_820;
mixer gate_output_15_820(.a(output_16_820), .b(output_16_5), .y(output_15_820));
wire output_1_821, output_1_6, output_0_821;
mixer gate_output_0_821(.a(output_1_821), .b(output_1_6), .y(output_0_821));
wire output_2_821, output_2_6, output_1_821;
mixer gate_output_1_821(.a(output_2_821), .b(output_2_6), .y(output_1_821));
wire output_3_821, output_3_6, output_2_821;
mixer gate_output_2_821(.a(output_3_821), .b(output_3_6), .y(output_2_821));
wire output_4_821, output_4_6, output_3_821;
mixer gate_output_3_821(.a(output_4_821), .b(output_4_6), .y(output_3_821));
wire output_5_821, output_5_6, output_4_821;
mixer gate_output_4_821(.a(output_5_821), .b(output_5_6), .y(output_4_821));
wire output_6_821, output_6_6, output_5_821;
mixer gate_output_5_821(.a(output_6_821), .b(output_6_6), .y(output_5_821));
wire output_7_821, output_7_6, output_6_821;
mixer gate_output_6_821(.a(output_7_821), .b(output_7_6), .y(output_6_821));
wire output_8_821, output_8_6, output_7_821;
mixer gate_output_7_821(.a(output_8_821), .b(output_8_6), .y(output_7_821));
wire output_9_821, output_9_6, output_8_821;
mixer gate_output_8_821(.a(output_9_821), .b(output_9_6), .y(output_8_821));
wire output_10_821, output_10_6, output_9_821;
mixer gate_output_9_821(.a(output_10_821), .b(output_10_6), .y(output_9_821));
wire output_11_821, output_11_6, output_10_821;
mixer gate_output_10_821(.a(output_11_821), .b(output_11_6), .y(output_10_821));
wire output_12_821, output_12_6, output_11_821;
mixer gate_output_11_821(.a(output_12_821), .b(output_12_6), .y(output_11_821));
wire output_13_821, output_13_6, output_12_821;
mixer gate_output_12_821(.a(output_13_821), .b(output_13_6), .y(output_12_821));
wire output_14_821, output_14_6, output_13_821;
mixer gate_output_13_821(.a(output_14_821), .b(output_14_6), .y(output_13_821));
wire output_15_821, output_15_6, output_14_821;
mixer gate_output_14_821(.a(output_15_821), .b(output_15_6), .y(output_14_821));
wire output_16_821, output_16_6, output_15_821;
mixer gate_output_15_821(.a(output_16_821), .b(output_16_6), .y(output_15_821));
wire output_1_822, output_1_7, output_0_822;
mixer gate_output_0_822(.a(output_1_822), .b(output_1_7), .y(output_0_822));
wire output_2_822, output_2_7, output_1_822;
mixer gate_output_1_822(.a(output_2_822), .b(output_2_7), .y(output_1_822));
wire output_3_822, output_3_7, output_2_822;
mixer gate_output_2_822(.a(output_3_822), .b(output_3_7), .y(output_2_822));
wire output_4_822, output_4_7, output_3_822;
mixer gate_output_3_822(.a(output_4_822), .b(output_4_7), .y(output_3_822));
wire output_5_822, output_5_7, output_4_822;
mixer gate_output_4_822(.a(output_5_822), .b(output_5_7), .y(output_4_822));
wire output_6_822, output_6_7, output_5_822;
mixer gate_output_5_822(.a(output_6_822), .b(output_6_7), .y(output_5_822));
wire output_7_822, output_7_7, output_6_822;
mixer gate_output_6_822(.a(output_7_822), .b(output_7_7), .y(output_6_822));
wire output_8_822, output_8_7, output_7_822;
mixer gate_output_7_822(.a(output_8_822), .b(output_8_7), .y(output_7_822));
wire output_9_822, output_9_7, output_8_822;
mixer gate_output_8_822(.a(output_9_822), .b(output_9_7), .y(output_8_822));
wire output_10_822, output_10_7, output_9_822;
mixer gate_output_9_822(.a(output_10_822), .b(output_10_7), .y(output_9_822));
wire output_11_822, output_11_7, output_10_822;
mixer gate_output_10_822(.a(output_11_822), .b(output_11_7), .y(output_10_822));
wire output_12_822, output_12_7, output_11_822;
mixer gate_output_11_822(.a(output_12_822), .b(output_12_7), .y(output_11_822));
wire output_13_822, output_13_7, output_12_822;
mixer gate_output_12_822(.a(output_13_822), .b(output_13_7), .y(output_12_822));
wire output_14_822, output_14_7, output_13_822;
mixer gate_output_13_822(.a(output_14_822), .b(output_14_7), .y(output_13_822));
wire output_15_822, output_15_7, output_14_822;
mixer gate_output_14_822(.a(output_15_822), .b(output_15_7), .y(output_14_822));
wire output_16_822, output_16_7, output_15_822;
mixer gate_output_15_822(.a(output_16_822), .b(output_16_7), .y(output_15_822));
wire output_1_823, output_1_8, output_0_823;
mixer gate_output_0_823(.a(output_1_823), .b(output_1_8), .y(output_0_823));
wire output_2_823, output_2_8, output_1_823;
mixer gate_output_1_823(.a(output_2_823), .b(output_2_8), .y(output_1_823));
wire output_3_823, output_3_8, output_2_823;
mixer gate_output_2_823(.a(output_3_823), .b(output_3_8), .y(output_2_823));
wire output_4_823, output_4_8, output_3_823;
mixer gate_output_3_823(.a(output_4_823), .b(output_4_8), .y(output_3_823));
wire output_5_823, output_5_8, output_4_823;
mixer gate_output_4_823(.a(output_5_823), .b(output_5_8), .y(output_4_823));
wire output_6_823, output_6_8, output_5_823;
mixer gate_output_5_823(.a(output_6_823), .b(output_6_8), .y(output_5_823));
wire output_7_823, output_7_8, output_6_823;
mixer gate_output_6_823(.a(output_7_823), .b(output_7_8), .y(output_6_823));
wire output_8_823, output_8_8, output_7_823;
mixer gate_output_7_823(.a(output_8_823), .b(output_8_8), .y(output_7_823));
wire output_9_823, output_9_8, output_8_823;
mixer gate_output_8_823(.a(output_9_823), .b(output_9_8), .y(output_8_823));
wire output_10_823, output_10_8, output_9_823;
mixer gate_output_9_823(.a(output_10_823), .b(output_10_8), .y(output_9_823));
wire output_11_823, output_11_8, output_10_823;
mixer gate_output_10_823(.a(output_11_823), .b(output_11_8), .y(output_10_823));
wire output_12_823, output_12_8, output_11_823;
mixer gate_output_11_823(.a(output_12_823), .b(output_12_8), .y(output_11_823));
wire output_13_823, output_13_8, output_12_823;
mixer gate_output_12_823(.a(output_13_823), .b(output_13_8), .y(output_12_823));
wire output_14_823, output_14_8, output_13_823;
mixer gate_output_13_823(.a(output_14_823), .b(output_14_8), .y(output_13_823));
wire output_15_823, output_15_8, output_14_823;
mixer gate_output_14_823(.a(output_15_823), .b(output_15_8), .y(output_14_823));
wire output_16_823, output_16_8, output_15_823;
mixer gate_output_15_823(.a(output_16_823), .b(output_16_8), .y(output_15_823));
wire output_1_824, output_1_9, output_0_824;
mixer gate_output_0_824(.a(output_1_824), .b(output_1_9), .y(output_0_824));
wire output_2_824, output_2_9, output_1_824;
mixer gate_output_1_824(.a(output_2_824), .b(output_2_9), .y(output_1_824));
wire output_3_824, output_3_9, output_2_824;
mixer gate_output_2_824(.a(output_3_824), .b(output_3_9), .y(output_2_824));
wire output_4_824, output_4_9, output_3_824;
mixer gate_output_3_824(.a(output_4_824), .b(output_4_9), .y(output_3_824));
wire output_5_824, output_5_9, output_4_824;
mixer gate_output_4_824(.a(output_5_824), .b(output_5_9), .y(output_4_824));
wire output_6_824, output_6_9, output_5_824;
mixer gate_output_5_824(.a(output_6_824), .b(output_6_9), .y(output_5_824));
wire output_7_824, output_7_9, output_6_824;
mixer gate_output_6_824(.a(output_7_824), .b(output_7_9), .y(output_6_824));
wire output_8_824, output_8_9, output_7_824;
mixer gate_output_7_824(.a(output_8_824), .b(output_8_9), .y(output_7_824));
wire output_9_824, output_9_9, output_8_824;
mixer gate_output_8_824(.a(output_9_824), .b(output_9_9), .y(output_8_824));
wire output_10_824, output_10_9, output_9_824;
mixer gate_output_9_824(.a(output_10_824), .b(output_10_9), .y(output_9_824));
wire output_11_824, output_11_9, output_10_824;
mixer gate_output_10_824(.a(output_11_824), .b(output_11_9), .y(output_10_824));
wire output_12_824, output_12_9, output_11_824;
mixer gate_output_11_824(.a(output_12_824), .b(output_12_9), .y(output_11_824));
wire output_13_824, output_13_9, output_12_824;
mixer gate_output_12_824(.a(output_13_824), .b(output_13_9), .y(output_12_824));
wire output_14_824, output_14_9, output_13_824;
mixer gate_output_13_824(.a(output_14_824), .b(output_14_9), .y(output_13_824));
wire output_15_824, output_15_9, output_14_824;
mixer gate_output_14_824(.a(output_15_824), .b(output_15_9), .y(output_14_824));
wire output_16_824, output_16_9, output_15_824;
mixer gate_output_15_824(.a(output_16_824), .b(output_16_9), .y(output_15_824));
wire output_1_825, output_1_10, output_0_825;
mixer gate_output_0_825(.a(output_1_825), .b(output_1_10), .y(output_0_825));
wire output_2_825, output_2_10, output_1_825;
mixer gate_output_1_825(.a(output_2_825), .b(output_2_10), .y(output_1_825));
wire output_3_825, output_3_10, output_2_825;
mixer gate_output_2_825(.a(output_3_825), .b(output_3_10), .y(output_2_825));
wire output_4_825, output_4_10, output_3_825;
mixer gate_output_3_825(.a(output_4_825), .b(output_4_10), .y(output_3_825));
wire output_5_825, output_5_10, output_4_825;
mixer gate_output_4_825(.a(output_5_825), .b(output_5_10), .y(output_4_825));
wire output_6_825, output_6_10, output_5_825;
mixer gate_output_5_825(.a(output_6_825), .b(output_6_10), .y(output_5_825));
wire output_7_825, output_7_10, output_6_825;
mixer gate_output_6_825(.a(output_7_825), .b(output_7_10), .y(output_6_825));
wire output_8_825, output_8_10, output_7_825;
mixer gate_output_7_825(.a(output_8_825), .b(output_8_10), .y(output_7_825));
wire output_9_825, output_9_10, output_8_825;
mixer gate_output_8_825(.a(output_9_825), .b(output_9_10), .y(output_8_825));
wire output_10_825, output_10_10, output_9_825;
mixer gate_output_9_825(.a(output_10_825), .b(output_10_10), .y(output_9_825));
wire output_11_825, output_11_10, output_10_825;
mixer gate_output_10_825(.a(output_11_825), .b(output_11_10), .y(output_10_825));
wire output_12_825, output_12_10, output_11_825;
mixer gate_output_11_825(.a(output_12_825), .b(output_12_10), .y(output_11_825));
wire output_13_825, output_13_10, output_12_825;
mixer gate_output_12_825(.a(output_13_825), .b(output_13_10), .y(output_12_825));
wire output_14_825, output_14_10, output_13_825;
mixer gate_output_13_825(.a(output_14_825), .b(output_14_10), .y(output_13_825));
wire output_15_825, output_15_10, output_14_825;
mixer gate_output_14_825(.a(output_15_825), .b(output_15_10), .y(output_14_825));
wire output_16_825, output_16_10, output_15_825;
mixer gate_output_15_825(.a(output_16_825), .b(output_16_10), .y(output_15_825));
wire output_1_826, output_1_11, output_0_826;
mixer gate_output_0_826(.a(output_1_826), .b(output_1_11), .y(output_0_826));
wire output_2_826, output_2_11, output_1_826;
mixer gate_output_1_826(.a(output_2_826), .b(output_2_11), .y(output_1_826));
wire output_3_826, output_3_11, output_2_826;
mixer gate_output_2_826(.a(output_3_826), .b(output_3_11), .y(output_2_826));
wire output_4_826, output_4_11, output_3_826;
mixer gate_output_3_826(.a(output_4_826), .b(output_4_11), .y(output_3_826));
wire output_5_826, output_5_11, output_4_826;
mixer gate_output_4_826(.a(output_5_826), .b(output_5_11), .y(output_4_826));
wire output_6_826, output_6_11, output_5_826;
mixer gate_output_5_826(.a(output_6_826), .b(output_6_11), .y(output_5_826));
wire output_7_826, output_7_11, output_6_826;
mixer gate_output_6_826(.a(output_7_826), .b(output_7_11), .y(output_6_826));
wire output_8_826, output_8_11, output_7_826;
mixer gate_output_7_826(.a(output_8_826), .b(output_8_11), .y(output_7_826));
wire output_9_826, output_9_11, output_8_826;
mixer gate_output_8_826(.a(output_9_826), .b(output_9_11), .y(output_8_826));
wire output_10_826, output_10_11, output_9_826;
mixer gate_output_9_826(.a(output_10_826), .b(output_10_11), .y(output_9_826));
wire output_11_826, output_11_11, output_10_826;
mixer gate_output_10_826(.a(output_11_826), .b(output_11_11), .y(output_10_826));
wire output_12_826, output_12_11, output_11_826;
mixer gate_output_11_826(.a(output_12_826), .b(output_12_11), .y(output_11_826));
wire output_13_826, output_13_11, output_12_826;
mixer gate_output_12_826(.a(output_13_826), .b(output_13_11), .y(output_12_826));
wire output_14_826, output_14_11, output_13_826;
mixer gate_output_13_826(.a(output_14_826), .b(output_14_11), .y(output_13_826));
wire output_15_826, output_15_11, output_14_826;
mixer gate_output_14_826(.a(output_15_826), .b(output_15_11), .y(output_14_826));
wire output_16_826, output_16_11, output_15_826;
mixer gate_output_15_826(.a(output_16_826), .b(output_16_11), .y(output_15_826));
wire output_1_827, output_1_12, output_0_827;
mixer gate_output_0_827(.a(output_1_827), .b(output_1_12), .y(output_0_827));
wire output_2_827, output_2_12, output_1_827;
mixer gate_output_1_827(.a(output_2_827), .b(output_2_12), .y(output_1_827));
wire output_3_827, output_3_12, output_2_827;
mixer gate_output_2_827(.a(output_3_827), .b(output_3_12), .y(output_2_827));
wire output_4_827, output_4_12, output_3_827;
mixer gate_output_3_827(.a(output_4_827), .b(output_4_12), .y(output_3_827));
wire output_5_827, output_5_12, output_4_827;
mixer gate_output_4_827(.a(output_5_827), .b(output_5_12), .y(output_4_827));
wire output_6_827, output_6_12, output_5_827;
mixer gate_output_5_827(.a(output_6_827), .b(output_6_12), .y(output_5_827));
wire output_7_827, output_7_12, output_6_827;
mixer gate_output_6_827(.a(output_7_827), .b(output_7_12), .y(output_6_827));
wire output_8_827, output_8_12, output_7_827;
mixer gate_output_7_827(.a(output_8_827), .b(output_8_12), .y(output_7_827));
wire output_9_827, output_9_12, output_8_827;
mixer gate_output_8_827(.a(output_9_827), .b(output_9_12), .y(output_8_827));
wire output_10_827, output_10_12, output_9_827;
mixer gate_output_9_827(.a(output_10_827), .b(output_10_12), .y(output_9_827));
wire output_11_827, output_11_12, output_10_827;
mixer gate_output_10_827(.a(output_11_827), .b(output_11_12), .y(output_10_827));
wire output_12_827, output_12_12, output_11_827;
mixer gate_output_11_827(.a(output_12_827), .b(output_12_12), .y(output_11_827));
wire output_13_827, output_13_12, output_12_827;
mixer gate_output_12_827(.a(output_13_827), .b(output_13_12), .y(output_12_827));
wire output_14_827, output_14_12, output_13_827;
mixer gate_output_13_827(.a(output_14_827), .b(output_14_12), .y(output_13_827));
wire output_15_827, output_15_12, output_14_827;
mixer gate_output_14_827(.a(output_15_827), .b(output_15_12), .y(output_14_827));
wire output_16_827, output_16_12, output_15_827;
mixer gate_output_15_827(.a(output_16_827), .b(output_16_12), .y(output_15_827));
wire output_1_828, output_1_13, output_0_828;
mixer gate_output_0_828(.a(output_1_828), .b(output_1_13), .y(output_0_828));
wire output_2_828, output_2_13, output_1_828;
mixer gate_output_1_828(.a(output_2_828), .b(output_2_13), .y(output_1_828));
wire output_3_828, output_3_13, output_2_828;
mixer gate_output_2_828(.a(output_3_828), .b(output_3_13), .y(output_2_828));
wire output_4_828, output_4_13, output_3_828;
mixer gate_output_3_828(.a(output_4_828), .b(output_4_13), .y(output_3_828));
wire output_5_828, output_5_13, output_4_828;
mixer gate_output_4_828(.a(output_5_828), .b(output_5_13), .y(output_4_828));
wire output_6_828, output_6_13, output_5_828;
mixer gate_output_5_828(.a(output_6_828), .b(output_6_13), .y(output_5_828));
wire output_7_828, output_7_13, output_6_828;
mixer gate_output_6_828(.a(output_7_828), .b(output_7_13), .y(output_6_828));
wire output_8_828, output_8_13, output_7_828;
mixer gate_output_7_828(.a(output_8_828), .b(output_8_13), .y(output_7_828));
wire output_9_828, output_9_13, output_8_828;
mixer gate_output_8_828(.a(output_9_828), .b(output_9_13), .y(output_8_828));
wire output_10_828, output_10_13, output_9_828;
mixer gate_output_9_828(.a(output_10_828), .b(output_10_13), .y(output_9_828));
wire output_11_828, output_11_13, output_10_828;
mixer gate_output_10_828(.a(output_11_828), .b(output_11_13), .y(output_10_828));
wire output_12_828, output_12_13, output_11_828;
mixer gate_output_11_828(.a(output_12_828), .b(output_12_13), .y(output_11_828));
wire output_13_828, output_13_13, output_12_828;
mixer gate_output_12_828(.a(output_13_828), .b(output_13_13), .y(output_12_828));
wire output_14_828, output_14_13, output_13_828;
mixer gate_output_13_828(.a(output_14_828), .b(output_14_13), .y(output_13_828));
wire output_15_828, output_15_13, output_14_828;
mixer gate_output_14_828(.a(output_15_828), .b(output_15_13), .y(output_14_828));
wire output_16_828, output_16_13, output_15_828;
mixer gate_output_15_828(.a(output_16_828), .b(output_16_13), .y(output_15_828));
wire output_1_829, output_1_14, output_0_829;
mixer gate_output_0_829(.a(output_1_829), .b(output_1_14), .y(output_0_829));
wire output_2_829, output_2_14, output_1_829;
mixer gate_output_1_829(.a(output_2_829), .b(output_2_14), .y(output_1_829));
wire output_3_829, output_3_14, output_2_829;
mixer gate_output_2_829(.a(output_3_829), .b(output_3_14), .y(output_2_829));
wire output_4_829, output_4_14, output_3_829;
mixer gate_output_3_829(.a(output_4_829), .b(output_4_14), .y(output_3_829));
wire output_5_829, output_5_14, output_4_829;
mixer gate_output_4_829(.a(output_5_829), .b(output_5_14), .y(output_4_829));
wire output_6_829, output_6_14, output_5_829;
mixer gate_output_5_829(.a(output_6_829), .b(output_6_14), .y(output_5_829));
wire output_7_829, output_7_14, output_6_829;
mixer gate_output_6_829(.a(output_7_829), .b(output_7_14), .y(output_6_829));
wire output_8_829, output_8_14, output_7_829;
mixer gate_output_7_829(.a(output_8_829), .b(output_8_14), .y(output_7_829));
wire output_9_829, output_9_14, output_8_829;
mixer gate_output_8_829(.a(output_9_829), .b(output_9_14), .y(output_8_829));
wire output_10_829, output_10_14, output_9_829;
mixer gate_output_9_829(.a(output_10_829), .b(output_10_14), .y(output_9_829));
wire output_11_829, output_11_14, output_10_829;
mixer gate_output_10_829(.a(output_11_829), .b(output_11_14), .y(output_10_829));
wire output_12_829, output_12_14, output_11_829;
mixer gate_output_11_829(.a(output_12_829), .b(output_12_14), .y(output_11_829));
wire output_13_829, output_13_14, output_12_829;
mixer gate_output_12_829(.a(output_13_829), .b(output_13_14), .y(output_12_829));
wire output_14_829, output_14_14, output_13_829;
mixer gate_output_13_829(.a(output_14_829), .b(output_14_14), .y(output_13_829));
wire output_15_829, output_15_14, output_14_829;
mixer gate_output_14_829(.a(output_15_829), .b(output_15_14), .y(output_14_829));
wire output_16_829, output_16_14, output_15_829;
mixer gate_output_15_829(.a(output_16_829), .b(output_16_14), .y(output_15_829));
wire output_1_830, output_1_15, output_0_830;
mixer gate_output_0_830(.a(output_1_830), .b(output_1_15), .y(output_0_830));
wire output_2_830, output_2_15, output_1_830;
mixer gate_output_1_830(.a(output_2_830), .b(output_2_15), .y(output_1_830));
wire output_3_830, output_3_15, output_2_830;
mixer gate_output_2_830(.a(output_3_830), .b(output_3_15), .y(output_2_830));
wire output_4_830, output_4_15, output_3_830;
mixer gate_output_3_830(.a(output_4_830), .b(output_4_15), .y(output_3_830));
wire output_5_830, output_5_15, output_4_830;
mixer gate_output_4_830(.a(output_5_830), .b(output_5_15), .y(output_4_830));
wire output_6_830, output_6_15, output_5_830;
mixer gate_output_5_830(.a(output_6_830), .b(output_6_15), .y(output_5_830));
wire output_7_830, output_7_15, output_6_830;
mixer gate_output_6_830(.a(output_7_830), .b(output_7_15), .y(output_6_830));
wire output_8_830, output_8_15, output_7_830;
mixer gate_output_7_830(.a(output_8_830), .b(output_8_15), .y(output_7_830));
wire output_9_830, output_9_15, output_8_830;
mixer gate_output_8_830(.a(output_9_830), .b(output_9_15), .y(output_8_830));
wire output_10_830, output_10_15, output_9_830;
mixer gate_output_9_830(.a(output_10_830), .b(output_10_15), .y(output_9_830));
wire output_11_830, output_11_15, output_10_830;
mixer gate_output_10_830(.a(output_11_830), .b(output_11_15), .y(output_10_830));
wire output_12_830, output_12_15, output_11_830;
mixer gate_output_11_830(.a(output_12_830), .b(output_12_15), .y(output_11_830));
wire output_13_830, output_13_15, output_12_830;
mixer gate_output_12_830(.a(output_13_830), .b(output_13_15), .y(output_12_830));
wire output_14_830, output_14_15, output_13_830;
mixer gate_output_13_830(.a(output_14_830), .b(output_14_15), .y(output_13_830));
wire output_15_830, output_15_15, output_14_830;
mixer gate_output_14_830(.a(output_15_830), .b(output_15_15), .y(output_14_830));
wire output_16_830, output_16_15, output_15_830;
mixer gate_output_15_830(.a(output_16_830), .b(output_16_15), .y(output_15_830));
wire output_1_831, output_1_0, output_0_831;
mixer gate_output_0_831(.a(output_1_831), .b(output_1_0), .y(output_0_831));
wire output_2_831, output_2_0, output_1_831;
mixer gate_output_1_831(.a(output_2_831), .b(output_2_0), .y(output_1_831));
wire output_3_831, output_3_0, output_2_831;
mixer gate_output_2_831(.a(output_3_831), .b(output_3_0), .y(output_2_831));
wire output_4_831, output_4_0, output_3_831;
mixer gate_output_3_831(.a(output_4_831), .b(output_4_0), .y(output_3_831));
wire output_5_831, output_5_0, output_4_831;
mixer gate_output_4_831(.a(output_5_831), .b(output_5_0), .y(output_4_831));
wire output_6_831, output_6_0, output_5_831;
mixer gate_output_5_831(.a(output_6_831), .b(output_6_0), .y(output_5_831));
wire output_7_831, output_7_0, output_6_831;
mixer gate_output_6_831(.a(output_7_831), .b(output_7_0), .y(output_6_831));
wire output_8_831, output_8_0, output_7_831;
mixer gate_output_7_831(.a(output_8_831), .b(output_8_0), .y(output_7_831));
wire output_9_831, output_9_0, output_8_831;
mixer gate_output_8_831(.a(output_9_831), .b(output_9_0), .y(output_8_831));
wire output_10_831, output_10_0, output_9_831;
mixer gate_output_9_831(.a(output_10_831), .b(output_10_0), .y(output_9_831));
wire output_11_831, output_11_0, output_10_831;
mixer gate_output_10_831(.a(output_11_831), .b(output_11_0), .y(output_10_831));
wire output_12_831, output_12_0, output_11_831;
mixer gate_output_11_831(.a(output_12_831), .b(output_12_0), .y(output_11_831));
wire output_13_831, output_13_0, output_12_831;
mixer gate_output_12_831(.a(output_13_831), .b(output_13_0), .y(output_12_831));
wire output_14_831, output_14_0, output_13_831;
mixer gate_output_13_831(.a(output_14_831), .b(output_14_0), .y(output_13_831));
wire output_15_831, output_15_0, output_14_831;
mixer gate_output_14_831(.a(output_15_831), .b(output_15_0), .y(output_14_831));
wire output_16_831, output_16_0, output_15_831;
mixer gate_output_15_831(.a(output_16_831), .b(output_16_0), .y(output_15_831));
wire output_1_832, output_1_1, output_0_832;
mixer gate_output_0_832(.a(output_1_832), .b(output_1_1), .y(output_0_832));
wire output_2_832, output_2_1, output_1_832;
mixer gate_output_1_832(.a(output_2_832), .b(output_2_1), .y(output_1_832));
wire output_3_832, output_3_1, output_2_832;
mixer gate_output_2_832(.a(output_3_832), .b(output_3_1), .y(output_2_832));
wire output_4_832, output_4_1, output_3_832;
mixer gate_output_3_832(.a(output_4_832), .b(output_4_1), .y(output_3_832));
wire output_5_832, output_5_1, output_4_832;
mixer gate_output_4_832(.a(output_5_832), .b(output_5_1), .y(output_4_832));
wire output_6_832, output_6_1, output_5_832;
mixer gate_output_5_832(.a(output_6_832), .b(output_6_1), .y(output_5_832));
wire output_7_832, output_7_1, output_6_832;
mixer gate_output_6_832(.a(output_7_832), .b(output_7_1), .y(output_6_832));
wire output_8_832, output_8_1, output_7_832;
mixer gate_output_7_832(.a(output_8_832), .b(output_8_1), .y(output_7_832));
wire output_9_832, output_9_1, output_8_832;
mixer gate_output_8_832(.a(output_9_832), .b(output_9_1), .y(output_8_832));
wire output_10_832, output_10_1, output_9_832;
mixer gate_output_9_832(.a(output_10_832), .b(output_10_1), .y(output_9_832));
wire output_11_832, output_11_1, output_10_832;
mixer gate_output_10_832(.a(output_11_832), .b(output_11_1), .y(output_10_832));
wire output_12_832, output_12_1, output_11_832;
mixer gate_output_11_832(.a(output_12_832), .b(output_12_1), .y(output_11_832));
wire output_13_832, output_13_1, output_12_832;
mixer gate_output_12_832(.a(output_13_832), .b(output_13_1), .y(output_12_832));
wire output_14_832, output_14_1, output_13_832;
mixer gate_output_13_832(.a(output_14_832), .b(output_14_1), .y(output_13_832));
wire output_15_832, output_15_1, output_14_832;
mixer gate_output_14_832(.a(output_15_832), .b(output_15_1), .y(output_14_832));
wire output_16_832, output_16_1, output_15_832;
mixer gate_output_15_832(.a(output_16_832), .b(output_16_1), .y(output_15_832));
wire output_1_833, output_1_2, output_0_833;
mixer gate_output_0_833(.a(output_1_833), .b(output_1_2), .y(output_0_833));
wire output_2_833, output_2_2, output_1_833;
mixer gate_output_1_833(.a(output_2_833), .b(output_2_2), .y(output_1_833));
wire output_3_833, output_3_2, output_2_833;
mixer gate_output_2_833(.a(output_3_833), .b(output_3_2), .y(output_2_833));
wire output_4_833, output_4_2, output_3_833;
mixer gate_output_3_833(.a(output_4_833), .b(output_4_2), .y(output_3_833));
wire output_5_833, output_5_2, output_4_833;
mixer gate_output_4_833(.a(output_5_833), .b(output_5_2), .y(output_4_833));
wire output_6_833, output_6_2, output_5_833;
mixer gate_output_5_833(.a(output_6_833), .b(output_6_2), .y(output_5_833));
wire output_7_833, output_7_2, output_6_833;
mixer gate_output_6_833(.a(output_7_833), .b(output_7_2), .y(output_6_833));
wire output_8_833, output_8_2, output_7_833;
mixer gate_output_7_833(.a(output_8_833), .b(output_8_2), .y(output_7_833));
wire output_9_833, output_9_2, output_8_833;
mixer gate_output_8_833(.a(output_9_833), .b(output_9_2), .y(output_8_833));
wire output_10_833, output_10_2, output_9_833;
mixer gate_output_9_833(.a(output_10_833), .b(output_10_2), .y(output_9_833));
wire output_11_833, output_11_2, output_10_833;
mixer gate_output_10_833(.a(output_11_833), .b(output_11_2), .y(output_10_833));
wire output_12_833, output_12_2, output_11_833;
mixer gate_output_11_833(.a(output_12_833), .b(output_12_2), .y(output_11_833));
wire output_13_833, output_13_2, output_12_833;
mixer gate_output_12_833(.a(output_13_833), .b(output_13_2), .y(output_12_833));
wire output_14_833, output_14_2, output_13_833;
mixer gate_output_13_833(.a(output_14_833), .b(output_14_2), .y(output_13_833));
wire output_15_833, output_15_2, output_14_833;
mixer gate_output_14_833(.a(output_15_833), .b(output_15_2), .y(output_14_833));
wire output_16_833, output_16_2, output_15_833;
mixer gate_output_15_833(.a(output_16_833), .b(output_16_2), .y(output_15_833));
wire output_1_834, output_1_3, output_0_834;
mixer gate_output_0_834(.a(output_1_834), .b(output_1_3), .y(output_0_834));
wire output_2_834, output_2_3, output_1_834;
mixer gate_output_1_834(.a(output_2_834), .b(output_2_3), .y(output_1_834));
wire output_3_834, output_3_3, output_2_834;
mixer gate_output_2_834(.a(output_3_834), .b(output_3_3), .y(output_2_834));
wire output_4_834, output_4_3, output_3_834;
mixer gate_output_3_834(.a(output_4_834), .b(output_4_3), .y(output_3_834));
wire output_5_834, output_5_3, output_4_834;
mixer gate_output_4_834(.a(output_5_834), .b(output_5_3), .y(output_4_834));
wire output_6_834, output_6_3, output_5_834;
mixer gate_output_5_834(.a(output_6_834), .b(output_6_3), .y(output_5_834));
wire output_7_834, output_7_3, output_6_834;
mixer gate_output_6_834(.a(output_7_834), .b(output_7_3), .y(output_6_834));
wire output_8_834, output_8_3, output_7_834;
mixer gate_output_7_834(.a(output_8_834), .b(output_8_3), .y(output_7_834));
wire output_9_834, output_9_3, output_8_834;
mixer gate_output_8_834(.a(output_9_834), .b(output_9_3), .y(output_8_834));
wire output_10_834, output_10_3, output_9_834;
mixer gate_output_9_834(.a(output_10_834), .b(output_10_3), .y(output_9_834));
wire output_11_834, output_11_3, output_10_834;
mixer gate_output_10_834(.a(output_11_834), .b(output_11_3), .y(output_10_834));
wire output_12_834, output_12_3, output_11_834;
mixer gate_output_11_834(.a(output_12_834), .b(output_12_3), .y(output_11_834));
wire output_13_834, output_13_3, output_12_834;
mixer gate_output_12_834(.a(output_13_834), .b(output_13_3), .y(output_12_834));
wire output_14_834, output_14_3, output_13_834;
mixer gate_output_13_834(.a(output_14_834), .b(output_14_3), .y(output_13_834));
wire output_15_834, output_15_3, output_14_834;
mixer gate_output_14_834(.a(output_15_834), .b(output_15_3), .y(output_14_834));
wire output_16_834, output_16_3, output_15_834;
mixer gate_output_15_834(.a(output_16_834), .b(output_16_3), .y(output_15_834));
wire output_1_835, output_1_4, output_0_835;
mixer gate_output_0_835(.a(output_1_835), .b(output_1_4), .y(output_0_835));
wire output_2_835, output_2_4, output_1_835;
mixer gate_output_1_835(.a(output_2_835), .b(output_2_4), .y(output_1_835));
wire output_3_835, output_3_4, output_2_835;
mixer gate_output_2_835(.a(output_3_835), .b(output_3_4), .y(output_2_835));
wire output_4_835, output_4_4, output_3_835;
mixer gate_output_3_835(.a(output_4_835), .b(output_4_4), .y(output_3_835));
wire output_5_835, output_5_4, output_4_835;
mixer gate_output_4_835(.a(output_5_835), .b(output_5_4), .y(output_4_835));
wire output_6_835, output_6_4, output_5_835;
mixer gate_output_5_835(.a(output_6_835), .b(output_6_4), .y(output_5_835));
wire output_7_835, output_7_4, output_6_835;
mixer gate_output_6_835(.a(output_7_835), .b(output_7_4), .y(output_6_835));
wire output_8_835, output_8_4, output_7_835;
mixer gate_output_7_835(.a(output_8_835), .b(output_8_4), .y(output_7_835));
wire output_9_835, output_9_4, output_8_835;
mixer gate_output_8_835(.a(output_9_835), .b(output_9_4), .y(output_8_835));
wire output_10_835, output_10_4, output_9_835;
mixer gate_output_9_835(.a(output_10_835), .b(output_10_4), .y(output_9_835));
wire output_11_835, output_11_4, output_10_835;
mixer gate_output_10_835(.a(output_11_835), .b(output_11_4), .y(output_10_835));
wire output_12_835, output_12_4, output_11_835;
mixer gate_output_11_835(.a(output_12_835), .b(output_12_4), .y(output_11_835));
wire output_13_835, output_13_4, output_12_835;
mixer gate_output_12_835(.a(output_13_835), .b(output_13_4), .y(output_12_835));
wire output_14_835, output_14_4, output_13_835;
mixer gate_output_13_835(.a(output_14_835), .b(output_14_4), .y(output_13_835));
wire output_15_835, output_15_4, output_14_835;
mixer gate_output_14_835(.a(output_15_835), .b(output_15_4), .y(output_14_835));
wire output_16_835, output_16_4, output_15_835;
mixer gate_output_15_835(.a(output_16_835), .b(output_16_4), .y(output_15_835));
wire output_1_836, output_1_5, output_0_836;
mixer gate_output_0_836(.a(output_1_836), .b(output_1_5), .y(output_0_836));
wire output_2_836, output_2_5, output_1_836;
mixer gate_output_1_836(.a(output_2_836), .b(output_2_5), .y(output_1_836));
wire output_3_836, output_3_5, output_2_836;
mixer gate_output_2_836(.a(output_3_836), .b(output_3_5), .y(output_2_836));
wire output_4_836, output_4_5, output_3_836;
mixer gate_output_3_836(.a(output_4_836), .b(output_4_5), .y(output_3_836));
wire output_5_836, output_5_5, output_4_836;
mixer gate_output_4_836(.a(output_5_836), .b(output_5_5), .y(output_4_836));
wire output_6_836, output_6_5, output_5_836;
mixer gate_output_5_836(.a(output_6_836), .b(output_6_5), .y(output_5_836));
wire output_7_836, output_7_5, output_6_836;
mixer gate_output_6_836(.a(output_7_836), .b(output_7_5), .y(output_6_836));
wire output_8_836, output_8_5, output_7_836;
mixer gate_output_7_836(.a(output_8_836), .b(output_8_5), .y(output_7_836));
wire output_9_836, output_9_5, output_8_836;
mixer gate_output_8_836(.a(output_9_836), .b(output_9_5), .y(output_8_836));
wire output_10_836, output_10_5, output_9_836;
mixer gate_output_9_836(.a(output_10_836), .b(output_10_5), .y(output_9_836));
wire output_11_836, output_11_5, output_10_836;
mixer gate_output_10_836(.a(output_11_836), .b(output_11_5), .y(output_10_836));
wire output_12_836, output_12_5, output_11_836;
mixer gate_output_11_836(.a(output_12_836), .b(output_12_5), .y(output_11_836));
wire output_13_836, output_13_5, output_12_836;
mixer gate_output_12_836(.a(output_13_836), .b(output_13_5), .y(output_12_836));
wire output_14_836, output_14_5, output_13_836;
mixer gate_output_13_836(.a(output_14_836), .b(output_14_5), .y(output_13_836));
wire output_15_836, output_15_5, output_14_836;
mixer gate_output_14_836(.a(output_15_836), .b(output_15_5), .y(output_14_836));
wire output_16_836, output_16_5, output_15_836;
mixer gate_output_15_836(.a(output_16_836), .b(output_16_5), .y(output_15_836));
wire output_1_837, output_1_6, output_0_837;
mixer gate_output_0_837(.a(output_1_837), .b(output_1_6), .y(output_0_837));
wire output_2_837, output_2_6, output_1_837;
mixer gate_output_1_837(.a(output_2_837), .b(output_2_6), .y(output_1_837));
wire output_3_837, output_3_6, output_2_837;
mixer gate_output_2_837(.a(output_3_837), .b(output_3_6), .y(output_2_837));
wire output_4_837, output_4_6, output_3_837;
mixer gate_output_3_837(.a(output_4_837), .b(output_4_6), .y(output_3_837));
wire output_5_837, output_5_6, output_4_837;
mixer gate_output_4_837(.a(output_5_837), .b(output_5_6), .y(output_4_837));
wire output_6_837, output_6_6, output_5_837;
mixer gate_output_5_837(.a(output_6_837), .b(output_6_6), .y(output_5_837));
wire output_7_837, output_7_6, output_6_837;
mixer gate_output_6_837(.a(output_7_837), .b(output_7_6), .y(output_6_837));
wire output_8_837, output_8_6, output_7_837;
mixer gate_output_7_837(.a(output_8_837), .b(output_8_6), .y(output_7_837));
wire output_9_837, output_9_6, output_8_837;
mixer gate_output_8_837(.a(output_9_837), .b(output_9_6), .y(output_8_837));
wire output_10_837, output_10_6, output_9_837;
mixer gate_output_9_837(.a(output_10_837), .b(output_10_6), .y(output_9_837));
wire output_11_837, output_11_6, output_10_837;
mixer gate_output_10_837(.a(output_11_837), .b(output_11_6), .y(output_10_837));
wire output_12_837, output_12_6, output_11_837;
mixer gate_output_11_837(.a(output_12_837), .b(output_12_6), .y(output_11_837));
wire output_13_837, output_13_6, output_12_837;
mixer gate_output_12_837(.a(output_13_837), .b(output_13_6), .y(output_12_837));
wire output_14_837, output_14_6, output_13_837;
mixer gate_output_13_837(.a(output_14_837), .b(output_14_6), .y(output_13_837));
wire output_15_837, output_15_6, output_14_837;
mixer gate_output_14_837(.a(output_15_837), .b(output_15_6), .y(output_14_837));
wire output_16_837, output_16_6, output_15_837;
mixer gate_output_15_837(.a(output_16_837), .b(output_16_6), .y(output_15_837));
wire output_1_838, output_1_7, output_0_838;
mixer gate_output_0_838(.a(output_1_838), .b(output_1_7), .y(output_0_838));
wire output_2_838, output_2_7, output_1_838;
mixer gate_output_1_838(.a(output_2_838), .b(output_2_7), .y(output_1_838));
wire output_3_838, output_3_7, output_2_838;
mixer gate_output_2_838(.a(output_3_838), .b(output_3_7), .y(output_2_838));
wire output_4_838, output_4_7, output_3_838;
mixer gate_output_3_838(.a(output_4_838), .b(output_4_7), .y(output_3_838));
wire output_5_838, output_5_7, output_4_838;
mixer gate_output_4_838(.a(output_5_838), .b(output_5_7), .y(output_4_838));
wire output_6_838, output_6_7, output_5_838;
mixer gate_output_5_838(.a(output_6_838), .b(output_6_7), .y(output_5_838));
wire output_7_838, output_7_7, output_6_838;
mixer gate_output_6_838(.a(output_7_838), .b(output_7_7), .y(output_6_838));
wire output_8_838, output_8_7, output_7_838;
mixer gate_output_7_838(.a(output_8_838), .b(output_8_7), .y(output_7_838));
wire output_9_838, output_9_7, output_8_838;
mixer gate_output_8_838(.a(output_9_838), .b(output_9_7), .y(output_8_838));
wire output_10_838, output_10_7, output_9_838;
mixer gate_output_9_838(.a(output_10_838), .b(output_10_7), .y(output_9_838));
wire output_11_838, output_11_7, output_10_838;
mixer gate_output_10_838(.a(output_11_838), .b(output_11_7), .y(output_10_838));
wire output_12_838, output_12_7, output_11_838;
mixer gate_output_11_838(.a(output_12_838), .b(output_12_7), .y(output_11_838));
wire output_13_838, output_13_7, output_12_838;
mixer gate_output_12_838(.a(output_13_838), .b(output_13_7), .y(output_12_838));
wire output_14_838, output_14_7, output_13_838;
mixer gate_output_13_838(.a(output_14_838), .b(output_14_7), .y(output_13_838));
wire output_15_838, output_15_7, output_14_838;
mixer gate_output_14_838(.a(output_15_838), .b(output_15_7), .y(output_14_838));
wire output_16_838, output_16_7, output_15_838;
mixer gate_output_15_838(.a(output_16_838), .b(output_16_7), .y(output_15_838));
wire output_1_839, output_1_8, output_0_839;
mixer gate_output_0_839(.a(output_1_839), .b(output_1_8), .y(output_0_839));
wire output_2_839, output_2_8, output_1_839;
mixer gate_output_1_839(.a(output_2_839), .b(output_2_8), .y(output_1_839));
wire output_3_839, output_3_8, output_2_839;
mixer gate_output_2_839(.a(output_3_839), .b(output_3_8), .y(output_2_839));
wire output_4_839, output_4_8, output_3_839;
mixer gate_output_3_839(.a(output_4_839), .b(output_4_8), .y(output_3_839));
wire output_5_839, output_5_8, output_4_839;
mixer gate_output_4_839(.a(output_5_839), .b(output_5_8), .y(output_4_839));
wire output_6_839, output_6_8, output_5_839;
mixer gate_output_5_839(.a(output_6_839), .b(output_6_8), .y(output_5_839));
wire output_7_839, output_7_8, output_6_839;
mixer gate_output_6_839(.a(output_7_839), .b(output_7_8), .y(output_6_839));
wire output_8_839, output_8_8, output_7_839;
mixer gate_output_7_839(.a(output_8_839), .b(output_8_8), .y(output_7_839));
wire output_9_839, output_9_8, output_8_839;
mixer gate_output_8_839(.a(output_9_839), .b(output_9_8), .y(output_8_839));
wire output_10_839, output_10_8, output_9_839;
mixer gate_output_9_839(.a(output_10_839), .b(output_10_8), .y(output_9_839));
wire output_11_839, output_11_8, output_10_839;
mixer gate_output_10_839(.a(output_11_839), .b(output_11_8), .y(output_10_839));
wire output_12_839, output_12_8, output_11_839;
mixer gate_output_11_839(.a(output_12_839), .b(output_12_8), .y(output_11_839));
wire output_13_839, output_13_8, output_12_839;
mixer gate_output_12_839(.a(output_13_839), .b(output_13_8), .y(output_12_839));
wire output_14_839, output_14_8, output_13_839;
mixer gate_output_13_839(.a(output_14_839), .b(output_14_8), .y(output_13_839));
wire output_15_839, output_15_8, output_14_839;
mixer gate_output_14_839(.a(output_15_839), .b(output_15_8), .y(output_14_839));
wire output_16_839, output_16_8, output_15_839;
mixer gate_output_15_839(.a(output_16_839), .b(output_16_8), .y(output_15_839));
wire output_1_840, output_1_9, output_0_840;
mixer gate_output_0_840(.a(output_1_840), .b(output_1_9), .y(output_0_840));
wire output_2_840, output_2_9, output_1_840;
mixer gate_output_1_840(.a(output_2_840), .b(output_2_9), .y(output_1_840));
wire output_3_840, output_3_9, output_2_840;
mixer gate_output_2_840(.a(output_3_840), .b(output_3_9), .y(output_2_840));
wire output_4_840, output_4_9, output_3_840;
mixer gate_output_3_840(.a(output_4_840), .b(output_4_9), .y(output_3_840));
wire output_5_840, output_5_9, output_4_840;
mixer gate_output_4_840(.a(output_5_840), .b(output_5_9), .y(output_4_840));
wire output_6_840, output_6_9, output_5_840;
mixer gate_output_5_840(.a(output_6_840), .b(output_6_9), .y(output_5_840));
wire output_7_840, output_7_9, output_6_840;
mixer gate_output_6_840(.a(output_7_840), .b(output_7_9), .y(output_6_840));
wire output_8_840, output_8_9, output_7_840;
mixer gate_output_7_840(.a(output_8_840), .b(output_8_9), .y(output_7_840));
wire output_9_840, output_9_9, output_8_840;
mixer gate_output_8_840(.a(output_9_840), .b(output_9_9), .y(output_8_840));
wire output_10_840, output_10_9, output_9_840;
mixer gate_output_9_840(.a(output_10_840), .b(output_10_9), .y(output_9_840));
wire output_11_840, output_11_9, output_10_840;
mixer gate_output_10_840(.a(output_11_840), .b(output_11_9), .y(output_10_840));
wire output_12_840, output_12_9, output_11_840;
mixer gate_output_11_840(.a(output_12_840), .b(output_12_9), .y(output_11_840));
wire output_13_840, output_13_9, output_12_840;
mixer gate_output_12_840(.a(output_13_840), .b(output_13_9), .y(output_12_840));
wire output_14_840, output_14_9, output_13_840;
mixer gate_output_13_840(.a(output_14_840), .b(output_14_9), .y(output_13_840));
wire output_15_840, output_15_9, output_14_840;
mixer gate_output_14_840(.a(output_15_840), .b(output_15_9), .y(output_14_840));
wire output_16_840, output_16_9, output_15_840;
mixer gate_output_15_840(.a(output_16_840), .b(output_16_9), .y(output_15_840));
wire output_1_841, output_1_10, output_0_841;
mixer gate_output_0_841(.a(output_1_841), .b(output_1_10), .y(output_0_841));
wire output_2_841, output_2_10, output_1_841;
mixer gate_output_1_841(.a(output_2_841), .b(output_2_10), .y(output_1_841));
wire output_3_841, output_3_10, output_2_841;
mixer gate_output_2_841(.a(output_3_841), .b(output_3_10), .y(output_2_841));
wire output_4_841, output_4_10, output_3_841;
mixer gate_output_3_841(.a(output_4_841), .b(output_4_10), .y(output_3_841));
wire output_5_841, output_5_10, output_4_841;
mixer gate_output_4_841(.a(output_5_841), .b(output_5_10), .y(output_4_841));
wire output_6_841, output_6_10, output_5_841;
mixer gate_output_5_841(.a(output_6_841), .b(output_6_10), .y(output_5_841));
wire output_7_841, output_7_10, output_6_841;
mixer gate_output_6_841(.a(output_7_841), .b(output_7_10), .y(output_6_841));
wire output_8_841, output_8_10, output_7_841;
mixer gate_output_7_841(.a(output_8_841), .b(output_8_10), .y(output_7_841));
wire output_9_841, output_9_10, output_8_841;
mixer gate_output_8_841(.a(output_9_841), .b(output_9_10), .y(output_8_841));
wire output_10_841, output_10_10, output_9_841;
mixer gate_output_9_841(.a(output_10_841), .b(output_10_10), .y(output_9_841));
wire output_11_841, output_11_10, output_10_841;
mixer gate_output_10_841(.a(output_11_841), .b(output_11_10), .y(output_10_841));
wire output_12_841, output_12_10, output_11_841;
mixer gate_output_11_841(.a(output_12_841), .b(output_12_10), .y(output_11_841));
wire output_13_841, output_13_10, output_12_841;
mixer gate_output_12_841(.a(output_13_841), .b(output_13_10), .y(output_12_841));
wire output_14_841, output_14_10, output_13_841;
mixer gate_output_13_841(.a(output_14_841), .b(output_14_10), .y(output_13_841));
wire output_15_841, output_15_10, output_14_841;
mixer gate_output_14_841(.a(output_15_841), .b(output_15_10), .y(output_14_841));
wire output_16_841, output_16_10, output_15_841;
mixer gate_output_15_841(.a(output_16_841), .b(output_16_10), .y(output_15_841));
wire output_1_842, output_1_11, output_0_842;
mixer gate_output_0_842(.a(output_1_842), .b(output_1_11), .y(output_0_842));
wire output_2_842, output_2_11, output_1_842;
mixer gate_output_1_842(.a(output_2_842), .b(output_2_11), .y(output_1_842));
wire output_3_842, output_3_11, output_2_842;
mixer gate_output_2_842(.a(output_3_842), .b(output_3_11), .y(output_2_842));
wire output_4_842, output_4_11, output_3_842;
mixer gate_output_3_842(.a(output_4_842), .b(output_4_11), .y(output_3_842));
wire output_5_842, output_5_11, output_4_842;
mixer gate_output_4_842(.a(output_5_842), .b(output_5_11), .y(output_4_842));
wire output_6_842, output_6_11, output_5_842;
mixer gate_output_5_842(.a(output_6_842), .b(output_6_11), .y(output_5_842));
wire output_7_842, output_7_11, output_6_842;
mixer gate_output_6_842(.a(output_7_842), .b(output_7_11), .y(output_6_842));
wire output_8_842, output_8_11, output_7_842;
mixer gate_output_7_842(.a(output_8_842), .b(output_8_11), .y(output_7_842));
wire output_9_842, output_9_11, output_8_842;
mixer gate_output_8_842(.a(output_9_842), .b(output_9_11), .y(output_8_842));
wire output_10_842, output_10_11, output_9_842;
mixer gate_output_9_842(.a(output_10_842), .b(output_10_11), .y(output_9_842));
wire output_11_842, output_11_11, output_10_842;
mixer gate_output_10_842(.a(output_11_842), .b(output_11_11), .y(output_10_842));
wire output_12_842, output_12_11, output_11_842;
mixer gate_output_11_842(.a(output_12_842), .b(output_12_11), .y(output_11_842));
wire output_13_842, output_13_11, output_12_842;
mixer gate_output_12_842(.a(output_13_842), .b(output_13_11), .y(output_12_842));
wire output_14_842, output_14_11, output_13_842;
mixer gate_output_13_842(.a(output_14_842), .b(output_14_11), .y(output_13_842));
wire output_15_842, output_15_11, output_14_842;
mixer gate_output_14_842(.a(output_15_842), .b(output_15_11), .y(output_14_842));
wire output_16_842, output_16_11, output_15_842;
mixer gate_output_15_842(.a(output_16_842), .b(output_16_11), .y(output_15_842));
wire output_1_843, output_1_12, output_0_843;
mixer gate_output_0_843(.a(output_1_843), .b(output_1_12), .y(output_0_843));
wire output_2_843, output_2_12, output_1_843;
mixer gate_output_1_843(.a(output_2_843), .b(output_2_12), .y(output_1_843));
wire output_3_843, output_3_12, output_2_843;
mixer gate_output_2_843(.a(output_3_843), .b(output_3_12), .y(output_2_843));
wire output_4_843, output_4_12, output_3_843;
mixer gate_output_3_843(.a(output_4_843), .b(output_4_12), .y(output_3_843));
wire output_5_843, output_5_12, output_4_843;
mixer gate_output_4_843(.a(output_5_843), .b(output_5_12), .y(output_4_843));
wire output_6_843, output_6_12, output_5_843;
mixer gate_output_5_843(.a(output_6_843), .b(output_6_12), .y(output_5_843));
wire output_7_843, output_7_12, output_6_843;
mixer gate_output_6_843(.a(output_7_843), .b(output_7_12), .y(output_6_843));
wire output_8_843, output_8_12, output_7_843;
mixer gate_output_7_843(.a(output_8_843), .b(output_8_12), .y(output_7_843));
wire output_9_843, output_9_12, output_8_843;
mixer gate_output_8_843(.a(output_9_843), .b(output_9_12), .y(output_8_843));
wire output_10_843, output_10_12, output_9_843;
mixer gate_output_9_843(.a(output_10_843), .b(output_10_12), .y(output_9_843));
wire output_11_843, output_11_12, output_10_843;
mixer gate_output_10_843(.a(output_11_843), .b(output_11_12), .y(output_10_843));
wire output_12_843, output_12_12, output_11_843;
mixer gate_output_11_843(.a(output_12_843), .b(output_12_12), .y(output_11_843));
wire output_13_843, output_13_12, output_12_843;
mixer gate_output_12_843(.a(output_13_843), .b(output_13_12), .y(output_12_843));
wire output_14_843, output_14_12, output_13_843;
mixer gate_output_13_843(.a(output_14_843), .b(output_14_12), .y(output_13_843));
wire output_15_843, output_15_12, output_14_843;
mixer gate_output_14_843(.a(output_15_843), .b(output_15_12), .y(output_14_843));
wire output_16_843, output_16_12, output_15_843;
mixer gate_output_15_843(.a(output_16_843), .b(output_16_12), .y(output_15_843));
wire output_1_844, output_1_13, output_0_844;
mixer gate_output_0_844(.a(output_1_844), .b(output_1_13), .y(output_0_844));
wire output_2_844, output_2_13, output_1_844;
mixer gate_output_1_844(.a(output_2_844), .b(output_2_13), .y(output_1_844));
wire output_3_844, output_3_13, output_2_844;
mixer gate_output_2_844(.a(output_3_844), .b(output_3_13), .y(output_2_844));
wire output_4_844, output_4_13, output_3_844;
mixer gate_output_3_844(.a(output_4_844), .b(output_4_13), .y(output_3_844));
wire output_5_844, output_5_13, output_4_844;
mixer gate_output_4_844(.a(output_5_844), .b(output_5_13), .y(output_4_844));
wire output_6_844, output_6_13, output_5_844;
mixer gate_output_5_844(.a(output_6_844), .b(output_6_13), .y(output_5_844));
wire output_7_844, output_7_13, output_6_844;
mixer gate_output_6_844(.a(output_7_844), .b(output_7_13), .y(output_6_844));
wire output_8_844, output_8_13, output_7_844;
mixer gate_output_7_844(.a(output_8_844), .b(output_8_13), .y(output_7_844));
wire output_9_844, output_9_13, output_8_844;
mixer gate_output_8_844(.a(output_9_844), .b(output_9_13), .y(output_8_844));
wire output_10_844, output_10_13, output_9_844;
mixer gate_output_9_844(.a(output_10_844), .b(output_10_13), .y(output_9_844));
wire output_11_844, output_11_13, output_10_844;
mixer gate_output_10_844(.a(output_11_844), .b(output_11_13), .y(output_10_844));
wire output_12_844, output_12_13, output_11_844;
mixer gate_output_11_844(.a(output_12_844), .b(output_12_13), .y(output_11_844));
wire output_13_844, output_13_13, output_12_844;
mixer gate_output_12_844(.a(output_13_844), .b(output_13_13), .y(output_12_844));
wire output_14_844, output_14_13, output_13_844;
mixer gate_output_13_844(.a(output_14_844), .b(output_14_13), .y(output_13_844));
wire output_15_844, output_15_13, output_14_844;
mixer gate_output_14_844(.a(output_15_844), .b(output_15_13), .y(output_14_844));
wire output_16_844, output_16_13, output_15_844;
mixer gate_output_15_844(.a(output_16_844), .b(output_16_13), .y(output_15_844));
wire output_1_845, output_1_14, output_0_845;
mixer gate_output_0_845(.a(output_1_845), .b(output_1_14), .y(output_0_845));
wire output_2_845, output_2_14, output_1_845;
mixer gate_output_1_845(.a(output_2_845), .b(output_2_14), .y(output_1_845));
wire output_3_845, output_3_14, output_2_845;
mixer gate_output_2_845(.a(output_3_845), .b(output_3_14), .y(output_2_845));
wire output_4_845, output_4_14, output_3_845;
mixer gate_output_3_845(.a(output_4_845), .b(output_4_14), .y(output_3_845));
wire output_5_845, output_5_14, output_4_845;
mixer gate_output_4_845(.a(output_5_845), .b(output_5_14), .y(output_4_845));
wire output_6_845, output_6_14, output_5_845;
mixer gate_output_5_845(.a(output_6_845), .b(output_6_14), .y(output_5_845));
wire output_7_845, output_7_14, output_6_845;
mixer gate_output_6_845(.a(output_7_845), .b(output_7_14), .y(output_6_845));
wire output_8_845, output_8_14, output_7_845;
mixer gate_output_7_845(.a(output_8_845), .b(output_8_14), .y(output_7_845));
wire output_9_845, output_9_14, output_8_845;
mixer gate_output_8_845(.a(output_9_845), .b(output_9_14), .y(output_8_845));
wire output_10_845, output_10_14, output_9_845;
mixer gate_output_9_845(.a(output_10_845), .b(output_10_14), .y(output_9_845));
wire output_11_845, output_11_14, output_10_845;
mixer gate_output_10_845(.a(output_11_845), .b(output_11_14), .y(output_10_845));
wire output_12_845, output_12_14, output_11_845;
mixer gate_output_11_845(.a(output_12_845), .b(output_12_14), .y(output_11_845));
wire output_13_845, output_13_14, output_12_845;
mixer gate_output_12_845(.a(output_13_845), .b(output_13_14), .y(output_12_845));
wire output_14_845, output_14_14, output_13_845;
mixer gate_output_13_845(.a(output_14_845), .b(output_14_14), .y(output_13_845));
wire output_15_845, output_15_14, output_14_845;
mixer gate_output_14_845(.a(output_15_845), .b(output_15_14), .y(output_14_845));
wire output_16_845, output_16_14, output_15_845;
mixer gate_output_15_845(.a(output_16_845), .b(output_16_14), .y(output_15_845));
wire output_1_846, output_1_15, output_0_846;
mixer gate_output_0_846(.a(output_1_846), .b(output_1_15), .y(output_0_846));
wire output_2_846, output_2_15, output_1_846;
mixer gate_output_1_846(.a(output_2_846), .b(output_2_15), .y(output_1_846));
wire output_3_846, output_3_15, output_2_846;
mixer gate_output_2_846(.a(output_3_846), .b(output_3_15), .y(output_2_846));
wire output_4_846, output_4_15, output_3_846;
mixer gate_output_3_846(.a(output_4_846), .b(output_4_15), .y(output_3_846));
wire output_5_846, output_5_15, output_4_846;
mixer gate_output_4_846(.a(output_5_846), .b(output_5_15), .y(output_4_846));
wire output_6_846, output_6_15, output_5_846;
mixer gate_output_5_846(.a(output_6_846), .b(output_6_15), .y(output_5_846));
wire output_7_846, output_7_15, output_6_846;
mixer gate_output_6_846(.a(output_7_846), .b(output_7_15), .y(output_6_846));
wire output_8_846, output_8_15, output_7_846;
mixer gate_output_7_846(.a(output_8_846), .b(output_8_15), .y(output_7_846));
wire output_9_846, output_9_15, output_8_846;
mixer gate_output_8_846(.a(output_9_846), .b(output_9_15), .y(output_8_846));
wire output_10_846, output_10_15, output_9_846;
mixer gate_output_9_846(.a(output_10_846), .b(output_10_15), .y(output_9_846));
wire output_11_846, output_11_15, output_10_846;
mixer gate_output_10_846(.a(output_11_846), .b(output_11_15), .y(output_10_846));
wire output_12_846, output_12_15, output_11_846;
mixer gate_output_11_846(.a(output_12_846), .b(output_12_15), .y(output_11_846));
wire output_13_846, output_13_15, output_12_846;
mixer gate_output_12_846(.a(output_13_846), .b(output_13_15), .y(output_12_846));
wire output_14_846, output_14_15, output_13_846;
mixer gate_output_13_846(.a(output_14_846), .b(output_14_15), .y(output_13_846));
wire output_15_846, output_15_15, output_14_846;
mixer gate_output_14_846(.a(output_15_846), .b(output_15_15), .y(output_14_846));
wire output_16_846, output_16_15, output_15_846;
mixer gate_output_15_846(.a(output_16_846), .b(output_16_15), .y(output_15_846));
wire output_1_847, output_1_0, output_0_847;
mixer gate_output_0_847(.a(output_1_847), .b(output_1_0), .y(output_0_847));
wire output_2_847, output_2_0, output_1_847;
mixer gate_output_1_847(.a(output_2_847), .b(output_2_0), .y(output_1_847));
wire output_3_847, output_3_0, output_2_847;
mixer gate_output_2_847(.a(output_3_847), .b(output_3_0), .y(output_2_847));
wire output_4_847, output_4_0, output_3_847;
mixer gate_output_3_847(.a(output_4_847), .b(output_4_0), .y(output_3_847));
wire output_5_847, output_5_0, output_4_847;
mixer gate_output_4_847(.a(output_5_847), .b(output_5_0), .y(output_4_847));
wire output_6_847, output_6_0, output_5_847;
mixer gate_output_5_847(.a(output_6_847), .b(output_6_0), .y(output_5_847));
wire output_7_847, output_7_0, output_6_847;
mixer gate_output_6_847(.a(output_7_847), .b(output_7_0), .y(output_6_847));
wire output_8_847, output_8_0, output_7_847;
mixer gate_output_7_847(.a(output_8_847), .b(output_8_0), .y(output_7_847));
wire output_9_847, output_9_0, output_8_847;
mixer gate_output_8_847(.a(output_9_847), .b(output_9_0), .y(output_8_847));
wire output_10_847, output_10_0, output_9_847;
mixer gate_output_9_847(.a(output_10_847), .b(output_10_0), .y(output_9_847));
wire output_11_847, output_11_0, output_10_847;
mixer gate_output_10_847(.a(output_11_847), .b(output_11_0), .y(output_10_847));
wire output_12_847, output_12_0, output_11_847;
mixer gate_output_11_847(.a(output_12_847), .b(output_12_0), .y(output_11_847));
wire output_13_847, output_13_0, output_12_847;
mixer gate_output_12_847(.a(output_13_847), .b(output_13_0), .y(output_12_847));
wire output_14_847, output_14_0, output_13_847;
mixer gate_output_13_847(.a(output_14_847), .b(output_14_0), .y(output_13_847));
wire output_15_847, output_15_0, output_14_847;
mixer gate_output_14_847(.a(output_15_847), .b(output_15_0), .y(output_14_847));
wire output_16_847, output_16_0, output_15_847;
mixer gate_output_15_847(.a(output_16_847), .b(output_16_0), .y(output_15_847));
wire output_1_848, output_1_1, output_0_848;
mixer gate_output_0_848(.a(output_1_848), .b(output_1_1), .y(output_0_848));
wire output_2_848, output_2_1, output_1_848;
mixer gate_output_1_848(.a(output_2_848), .b(output_2_1), .y(output_1_848));
wire output_3_848, output_3_1, output_2_848;
mixer gate_output_2_848(.a(output_3_848), .b(output_3_1), .y(output_2_848));
wire output_4_848, output_4_1, output_3_848;
mixer gate_output_3_848(.a(output_4_848), .b(output_4_1), .y(output_3_848));
wire output_5_848, output_5_1, output_4_848;
mixer gate_output_4_848(.a(output_5_848), .b(output_5_1), .y(output_4_848));
wire output_6_848, output_6_1, output_5_848;
mixer gate_output_5_848(.a(output_6_848), .b(output_6_1), .y(output_5_848));
wire output_7_848, output_7_1, output_6_848;
mixer gate_output_6_848(.a(output_7_848), .b(output_7_1), .y(output_6_848));
wire output_8_848, output_8_1, output_7_848;
mixer gate_output_7_848(.a(output_8_848), .b(output_8_1), .y(output_7_848));
wire output_9_848, output_9_1, output_8_848;
mixer gate_output_8_848(.a(output_9_848), .b(output_9_1), .y(output_8_848));
wire output_10_848, output_10_1, output_9_848;
mixer gate_output_9_848(.a(output_10_848), .b(output_10_1), .y(output_9_848));
wire output_11_848, output_11_1, output_10_848;
mixer gate_output_10_848(.a(output_11_848), .b(output_11_1), .y(output_10_848));
wire output_12_848, output_12_1, output_11_848;
mixer gate_output_11_848(.a(output_12_848), .b(output_12_1), .y(output_11_848));
wire output_13_848, output_13_1, output_12_848;
mixer gate_output_12_848(.a(output_13_848), .b(output_13_1), .y(output_12_848));
wire output_14_848, output_14_1, output_13_848;
mixer gate_output_13_848(.a(output_14_848), .b(output_14_1), .y(output_13_848));
wire output_15_848, output_15_1, output_14_848;
mixer gate_output_14_848(.a(output_15_848), .b(output_15_1), .y(output_14_848));
wire output_16_848, output_16_1, output_15_848;
mixer gate_output_15_848(.a(output_16_848), .b(output_16_1), .y(output_15_848));
wire output_1_849, output_1_2, output_0_849;
mixer gate_output_0_849(.a(output_1_849), .b(output_1_2), .y(output_0_849));
wire output_2_849, output_2_2, output_1_849;
mixer gate_output_1_849(.a(output_2_849), .b(output_2_2), .y(output_1_849));
wire output_3_849, output_3_2, output_2_849;
mixer gate_output_2_849(.a(output_3_849), .b(output_3_2), .y(output_2_849));
wire output_4_849, output_4_2, output_3_849;
mixer gate_output_3_849(.a(output_4_849), .b(output_4_2), .y(output_3_849));
wire output_5_849, output_5_2, output_4_849;
mixer gate_output_4_849(.a(output_5_849), .b(output_5_2), .y(output_4_849));
wire output_6_849, output_6_2, output_5_849;
mixer gate_output_5_849(.a(output_6_849), .b(output_6_2), .y(output_5_849));
wire output_7_849, output_7_2, output_6_849;
mixer gate_output_6_849(.a(output_7_849), .b(output_7_2), .y(output_6_849));
wire output_8_849, output_8_2, output_7_849;
mixer gate_output_7_849(.a(output_8_849), .b(output_8_2), .y(output_7_849));
wire output_9_849, output_9_2, output_8_849;
mixer gate_output_8_849(.a(output_9_849), .b(output_9_2), .y(output_8_849));
wire output_10_849, output_10_2, output_9_849;
mixer gate_output_9_849(.a(output_10_849), .b(output_10_2), .y(output_9_849));
wire output_11_849, output_11_2, output_10_849;
mixer gate_output_10_849(.a(output_11_849), .b(output_11_2), .y(output_10_849));
wire output_12_849, output_12_2, output_11_849;
mixer gate_output_11_849(.a(output_12_849), .b(output_12_2), .y(output_11_849));
wire output_13_849, output_13_2, output_12_849;
mixer gate_output_12_849(.a(output_13_849), .b(output_13_2), .y(output_12_849));
wire output_14_849, output_14_2, output_13_849;
mixer gate_output_13_849(.a(output_14_849), .b(output_14_2), .y(output_13_849));
wire output_15_849, output_15_2, output_14_849;
mixer gate_output_14_849(.a(output_15_849), .b(output_15_2), .y(output_14_849));
wire output_16_849, output_16_2, output_15_849;
mixer gate_output_15_849(.a(output_16_849), .b(output_16_2), .y(output_15_849));
wire output_1_850, output_1_3, output_0_850;
mixer gate_output_0_850(.a(output_1_850), .b(output_1_3), .y(output_0_850));
wire output_2_850, output_2_3, output_1_850;
mixer gate_output_1_850(.a(output_2_850), .b(output_2_3), .y(output_1_850));
wire output_3_850, output_3_3, output_2_850;
mixer gate_output_2_850(.a(output_3_850), .b(output_3_3), .y(output_2_850));
wire output_4_850, output_4_3, output_3_850;
mixer gate_output_3_850(.a(output_4_850), .b(output_4_3), .y(output_3_850));
wire output_5_850, output_5_3, output_4_850;
mixer gate_output_4_850(.a(output_5_850), .b(output_5_3), .y(output_4_850));
wire output_6_850, output_6_3, output_5_850;
mixer gate_output_5_850(.a(output_6_850), .b(output_6_3), .y(output_5_850));
wire output_7_850, output_7_3, output_6_850;
mixer gate_output_6_850(.a(output_7_850), .b(output_7_3), .y(output_6_850));
wire output_8_850, output_8_3, output_7_850;
mixer gate_output_7_850(.a(output_8_850), .b(output_8_3), .y(output_7_850));
wire output_9_850, output_9_3, output_8_850;
mixer gate_output_8_850(.a(output_9_850), .b(output_9_3), .y(output_8_850));
wire output_10_850, output_10_3, output_9_850;
mixer gate_output_9_850(.a(output_10_850), .b(output_10_3), .y(output_9_850));
wire output_11_850, output_11_3, output_10_850;
mixer gate_output_10_850(.a(output_11_850), .b(output_11_3), .y(output_10_850));
wire output_12_850, output_12_3, output_11_850;
mixer gate_output_11_850(.a(output_12_850), .b(output_12_3), .y(output_11_850));
wire output_13_850, output_13_3, output_12_850;
mixer gate_output_12_850(.a(output_13_850), .b(output_13_3), .y(output_12_850));
wire output_14_850, output_14_3, output_13_850;
mixer gate_output_13_850(.a(output_14_850), .b(output_14_3), .y(output_13_850));
wire output_15_850, output_15_3, output_14_850;
mixer gate_output_14_850(.a(output_15_850), .b(output_15_3), .y(output_14_850));
wire output_16_850, output_16_3, output_15_850;
mixer gate_output_15_850(.a(output_16_850), .b(output_16_3), .y(output_15_850));
wire output_1_851, output_1_4, output_0_851;
mixer gate_output_0_851(.a(output_1_851), .b(output_1_4), .y(output_0_851));
wire output_2_851, output_2_4, output_1_851;
mixer gate_output_1_851(.a(output_2_851), .b(output_2_4), .y(output_1_851));
wire output_3_851, output_3_4, output_2_851;
mixer gate_output_2_851(.a(output_3_851), .b(output_3_4), .y(output_2_851));
wire output_4_851, output_4_4, output_3_851;
mixer gate_output_3_851(.a(output_4_851), .b(output_4_4), .y(output_3_851));
wire output_5_851, output_5_4, output_4_851;
mixer gate_output_4_851(.a(output_5_851), .b(output_5_4), .y(output_4_851));
wire output_6_851, output_6_4, output_5_851;
mixer gate_output_5_851(.a(output_6_851), .b(output_6_4), .y(output_5_851));
wire output_7_851, output_7_4, output_6_851;
mixer gate_output_6_851(.a(output_7_851), .b(output_7_4), .y(output_6_851));
wire output_8_851, output_8_4, output_7_851;
mixer gate_output_7_851(.a(output_8_851), .b(output_8_4), .y(output_7_851));
wire output_9_851, output_9_4, output_8_851;
mixer gate_output_8_851(.a(output_9_851), .b(output_9_4), .y(output_8_851));
wire output_10_851, output_10_4, output_9_851;
mixer gate_output_9_851(.a(output_10_851), .b(output_10_4), .y(output_9_851));
wire output_11_851, output_11_4, output_10_851;
mixer gate_output_10_851(.a(output_11_851), .b(output_11_4), .y(output_10_851));
wire output_12_851, output_12_4, output_11_851;
mixer gate_output_11_851(.a(output_12_851), .b(output_12_4), .y(output_11_851));
wire output_13_851, output_13_4, output_12_851;
mixer gate_output_12_851(.a(output_13_851), .b(output_13_4), .y(output_12_851));
wire output_14_851, output_14_4, output_13_851;
mixer gate_output_13_851(.a(output_14_851), .b(output_14_4), .y(output_13_851));
wire output_15_851, output_15_4, output_14_851;
mixer gate_output_14_851(.a(output_15_851), .b(output_15_4), .y(output_14_851));
wire output_16_851, output_16_4, output_15_851;
mixer gate_output_15_851(.a(output_16_851), .b(output_16_4), .y(output_15_851));
wire output_1_852, output_1_5, output_0_852;
mixer gate_output_0_852(.a(output_1_852), .b(output_1_5), .y(output_0_852));
wire output_2_852, output_2_5, output_1_852;
mixer gate_output_1_852(.a(output_2_852), .b(output_2_5), .y(output_1_852));
wire output_3_852, output_3_5, output_2_852;
mixer gate_output_2_852(.a(output_3_852), .b(output_3_5), .y(output_2_852));
wire output_4_852, output_4_5, output_3_852;
mixer gate_output_3_852(.a(output_4_852), .b(output_4_5), .y(output_3_852));
wire output_5_852, output_5_5, output_4_852;
mixer gate_output_4_852(.a(output_5_852), .b(output_5_5), .y(output_4_852));
wire output_6_852, output_6_5, output_5_852;
mixer gate_output_5_852(.a(output_6_852), .b(output_6_5), .y(output_5_852));
wire output_7_852, output_7_5, output_6_852;
mixer gate_output_6_852(.a(output_7_852), .b(output_7_5), .y(output_6_852));
wire output_8_852, output_8_5, output_7_852;
mixer gate_output_7_852(.a(output_8_852), .b(output_8_5), .y(output_7_852));
wire output_9_852, output_9_5, output_8_852;
mixer gate_output_8_852(.a(output_9_852), .b(output_9_5), .y(output_8_852));
wire output_10_852, output_10_5, output_9_852;
mixer gate_output_9_852(.a(output_10_852), .b(output_10_5), .y(output_9_852));
wire output_11_852, output_11_5, output_10_852;
mixer gate_output_10_852(.a(output_11_852), .b(output_11_5), .y(output_10_852));
wire output_12_852, output_12_5, output_11_852;
mixer gate_output_11_852(.a(output_12_852), .b(output_12_5), .y(output_11_852));
wire output_13_852, output_13_5, output_12_852;
mixer gate_output_12_852(.a(output_13_852), .b(output_13_5), .y(output_12_852));
wire output_14_852, output_14_5, output_13_852;
mixer gate_output_13_852(.a(output_14_852), .b(output_14_5), .y(output_13_852));
wire output_15_852, output_15_5, output_14_852;
mixer gate_output_14_852(.a(output_15_852), .b(output_15_5), .y(output_14_852));
wire output_16_852, output_16_5, output_15_852;
mixer gate_output_15_852(.a(output_16_852), .b(output_16_5), .y(output_15_852));
wire output_1_853, output_1_6, output_0_853;
mixer gate_output_0_853(.a(output_1_853), .b(output_1_6), .y(output_0_853));
wire output_2_853, output_2_6, output_1_853;
mixer gate_output_1_853(.a(output_2_853), .b(output_2_6), .y(output_1_853));
wire output_3_853, output_3_6, output_2_853;
mixer gate_output_2_853(.a(output_3_853), .b(output_3_6), .y(output_2_853));
wire output_4_853, output_4_6, output_3_853;
mixer gate_output_3_853(.a(output_4_853), .b(output_4_6), .y(output_3_853));
wire output_5_853, output_5_6, output_4_853;
mixer gate_output_4_853(.a(output_5_853), .b(output_5_6), .y(output_4_853));
wire output_6_853, output_6_6, output_5_853;
mixer gate_output_5_853(.a(output_6_853), .b(output_6_6), .y(output_5_853));
wire output_7_853, output_7_6, output_6_853;
mixer gate_output_6_853(.a(output_7_853), .b(output_7_6), .y(output_6_853));
wire output_8_853, output_8_6, output_7_853;
mixer gate_output_7_853(.a(output_8_853), .b(output_8_6), .y(output_7_853));
wire output_9_853, output_9_6, output_8_853;
mixer gate_output_8_853(.a(output_9_853), .b(output_9_6), .y(output_8_853));
wire output_10_853, output_10_6, output_9_853;
mixer gate_output_9_853(.a(output_10_853), .b(output_10_6), .y(output_9_853));
wire output_11_853, output_11_6, output_10_853;
mixer gate_output_10_853(.a(output_11_853), .b(output_11_6), .y(output_10_853));
wire output_12_853, output_12_6, output_11_853;
mixer gate_output_11_853(.a(output_12_853), .b(output_12_6), .y(output_11_853));
wire output_13_853, output_13_6, output_12_853;
mixer gate_output_12_853(.a(output_13_853), .b(output_13_6), .y(output_12_853));
wire output_14_853, output_14_6, output_13_853;
mixer gate_output_13_853(.a(output_14_853), .b(output_14_6), .y(output_13_853));
wire output_15_853, output_15_6, output_14_853;
mixer gate_output_14_853(.a(output_15_853), .b(output_15_6), .y(output_14_853));
wire output_16_853, output_16_6, output_15_853;
mixer gate_output_15_853(.a(output_16_853), .b(output_16_6), .y(output_15_853));
wire output_1_854, output_1_7, output_0_854;
mixer gate_output_0_854(.a(output_1_854), .b(output_1_7), .y(output_0_854));
wire output_2_854, output_2_7, output_1_854;
mixer gate_output_1_854(.a(output_2_854), .b(output_2_7), .y(output_1_854));
wire output_3_854, output_3_7, output_2_854;
mixer gate_output_2_854(.a(output_3_854), .b(output_3_7), .y(output_2_854));
wire output_4_854, output_4_7, output_3_854;
mixer gate_output_3_854(.a(output_4_854), .b(output_4_7), .y(output_3_854));
wire output_5_854, output_5_7, output_4_854;
mixer gate_output_4_854(.a(output_5_854), .b(output_5_7), .y(output_4_854));
wire output_6_854, output_6_7, output_5_854;
mixer gate_output_5_854(.a(output_6_854), .b(output_6_7), .y(output_5_854));
wire output_7_854, output_7_7, output_6_854;
mixer gate_output_6_854(.a(output_7_854), .b(output_7_7), .y(output_6_854));
wire output_8_854, output_8_7, output_7_854;
mixer gate_output_7_854(.a(output_8_854), .b(output_8_7), .y(output_7_854));
wire output_9_854, output_9_7, output_8_854;
mixer gate_output_8_854(.a(output_9_854), .b(output_9_7), .y(output_8_854));
wire output_10_854, output_10_7, output_9_854;
mixer gate_output_9_854(.a(output_10_854), .b(output_10_7), .y(output_9_854));
wire output_11_854, output_11_7, output_10_854;
mixer gate_output_10_854(.a(output_11_854), .b(output_11_7), .y(output_10_854));
wire output_12_854, output_12_7, output_11_854;
mixer gate_output_11_854(.a(output_12_854), .b(output_12_7), .y(output_11_854));
wire output_13_854, output_13_7, output_12_854;
mixer gate_output_12_854(.a(output_13_854), .b(output_13_7), .y(output_12_854));
wire output_14_854, output_14_7, output_13_854;
mixer gate_output_13_854(.a(output_14_854), .b(output_14_7), .y(output_13_854));
wire output_15_854, output_15_7, output_14_854;
mixer gate_output_14_854(.a(output_15_854), .b(output_15_7), .y(output_14_854));
wire output_16_854, output_16_7, output_15_854;
mixer gate_output_15_854(.a(output_16_854), .b(output_16_7), .y(output_15_854));
wire output_1_855, output_1_8, output_0_855;
mixer gate_output_0_855(.a(output_1_855), .b(output_1_8), .y(output_0_855));
wire output_2_855, output_2_8, output_1_855;
mixer gate_output_1_855(.a(output_2_855), .b(output_2_8), .y(output_1_855));
wire output_3_855, output_3_8, output_2_855;
mixer gate_output_2_855(.a(output_3_855), .b(output_3_8), .y(output_2_855));
wire output_4_855, output_4_8, output_3_855;
mixer gate_output_3_855(.a(output_4_855), .b(output_4_8), .y(output_3_855));
wire output_5_855, output_5_8, output_4_855;
mixer gate_output_4_855(.a(output_5_855), .b(output_5_8), .y(output_4_855));
wire output_6_855, output_6_8, output_5_855;
mixer gate_output_5_855(.a(output_6_855), .b(output_6_8), .y(output_5_855));
wire output_7_855, output_7_8, output_6_855;
mixer gate_output_6_855(.a(output_7_855), .b(output_7_8), .y(output_6_855));
wire output_8_855, output_8_8, output_7_855;
mixer gate_output_7_855(.a(output_8_855), .b(output_8_8), .y(output_7_855));
wire output_9_855, output_9_8, output_8_855;
mixer gate_output_8_855(.a(output_9_855), .b(output_9_8), .y(output_8_855));
wire output_10_855, output_10_8, output_9_855;
mixer gate_output_9_855(.a(output_10_855), .b(output_10_8), .y(output_9_855));
wire output_11_855, output_11_8, output_10_855;
mixer gate_output_10_855(.a(output_11_855), .b(output_11_8), .y(output_10_855));
wire output_12_855, output_12_8, output_11_855;
mixer gate_output_11_855(.a(output_12_855), .b(output_12_8), .y(output_11_855));
wire output_13_855, output_13_8, output_12_855;
mixer gate_output_12_855(.a(output_13_855), .b(output_13_8), .y(output_12_855));
wire output_14_855, output_14_8, output_13_855;
mixer gate_output_13_855(.a(output_14_855), .b(output_14_8), .y(output_13_855));
wire output_15_855, output_15_8, output_14_855;
mixer gate_output_14_855(.a(output_15_855), .b(output_15_8), .y(output_14_855));
wire output_16_855, output_16_8, output_15_855;
mixer gate_output_15_855(.a(output_16_855), .b(output_16_8), .y(output_15_855));
wire output_1_856, output_1_9, output_0_856;
mixer gate_output_0_856(.a(output_1_856), .b(output_1_9), .y(output_0_856));
wire output_2_856, output_2_9, output_1_856;
mixer gate_output_1_856(.a(output_2_856), .b(output_2_9), .y(output_1_856));
wire output_3_856, output_3_9, output_2_856;
mixer gate_output_2_856(.a(output_3_856), .b(output_3_9), .y(output_2_856));
wire output_4_856, output_4_9, output_3_856;
mixer gate_output_3_856(.a(output_4_856), .b(output_4_9), .y(output_3_856));
wire output_5_856, output_5_9, output_4_856;
mixer gate_output_4_856(.a(output_5_856), .b(output_5_9), .y(output_4_856));
wire output_6_856, output_6_9, output_5_856;
mixer gate_output_5_856(.a(output_6_856), .b(output_6_9), .y(output_5_856));
wire output_7_856, output_7_9, output_6_856;
mixer gate_output_6_856(.a(output_7_856), .b(output_7_9), .y(output_6_856));
wire output_8_856, output_8_9, output_7_856;
mixer gate_output_7_856(.a(output_8_856), .b(output_8_9), .y(output_7_856));
wire output_9_856, output_9_9, output_8_856;
mixer gate_output_8_856(.a(output_9_856), .b(output_9_9), .y(output_8_856));
wire output_10_856, output_10_9, output_9_856;
mixer gate_output_9_856(.a(output_10_856), .b(output_10_9), .y(output_9_856));
wire output_11_856, output_11_9, output_10_856;
mixer gate_output_10_856(.a(output_11_856), .b(output_11_9), .y(output_10_856));
wire output_12_856, output_12_9, output_11_856;
mixer gate_output_11_856(.a(output_12_856), .b(output_12_9), .y(output_11_856));
wire output_13_856, output_13_9, output_12_856;
mixer gate_output_12_856(.a(output_13_856), .b(output_13_9), .y(output_12_856));
wire output_14_856, output_14_9, output_13_856;
mixer gate_output_13_856(.a(output_14_856), .b(output_14_9), .y(output_13_856));
wire output_15_856, output_15_9, output_14_856;
mixer gate_output_14_856(.a(output_15_856), .b(output_15_9), .y(output_14_856));
wire output_16_856, output_16_9, output_15_856;
mixer gate_output_15_856(.a(output_16_856), .b(output_16_9), .y(output_15_856));
wire output_1_857, output_1_10, output_0_857;
mixer gate_output_0_857(.a(output_1_857), .b(output_1_10), .y(output_0_857));
wire output_2_857, output_2_10, output_1_857;
mixer gate_output_1_857(.a(output_2_857), .b(output_2_10), .y(output_1_857));
wire output_3_857, output_3_10, output_2_857;
mixer gate_output_2_857(.a(output_3_857), .b(output_3_10), .y(output_2_857));
wire output_4_857, output_4_10, output_3_857;
mixer gate_output_3_857(.a(output_4_857), .b(output_4_10), .y(output_3_857));
wire output_5_857, output_5_10, output_4_857;
mixer gate_output_4_857(.a(output_5_857), .b(output_5_10), .y(output_4_857));
wire output_6_857, output_6_10, output_5_857;
mixer gate_output_5_857(.a(output_6_857), .b(output_6_10), .y(output_5_857));
wire output_7_857, output_7_10, output_6_857;
mixer gate_output_6_857(.a(output_7_857), .b(output_7_10), .y(output_6_857));
wire output_8_857, output_8_10, output_7_857;
mixer gate_output_7_857(.a(output_8_857), .b(output_8_10), .y(output_7_857));
wire output_9_857, output_9_10, output_8_857;
mixer gate_output_8_857(.a(output_9_857), .b(output_9_10), .y(output_8_857));
wire output_10_857, output_10_10, output_9_857;
mixer gate_output_9_857(.a(output_10_857), .b(output_10_10), .y(output_9_857));
wire output_11_857, output_11_10, output_10_857;
mixer gate_output_10_857(.a(output_11_857), .b(output_11_10), .y(output_10_857));
wire output_12_857, output_12_10, output_11_857;
mixer gate_output_11_857(.a(output_12_857), .b(output_12_10), .y(output_11_857));
wire output_13_857, output_13_10, output_12_857;
mixer gate_output_12_857(.a(output_13_857), .b(output_13_10), .y(output_12_857));
wire output_14_857, output_14_10, output_13_857;
mixer gate_output_13_857(.a(output_14_857), .b(output_14_10), .y(output_13_857));
wire output_15_857, output_15_10, output_14_857;
mixer gate_output_14_857(.a(output_15_857), .b(output_15_10), .y(output_14_857));
wire output_16_857, output_16_10, output_15_857;
mixer gate_output_15_857(.a(output_16_857), .b(output_16_10), .y(output_15_857));
wire output_1_858, output_1_11, output_0_858;
mixer gate_output_0_858(.a(output_1_858), .b(output_1_11), .y(output_0_858));
wire output_2_858, output_2_11, output_1_858;
mixer gate_output_1_858(.a(output_2_858), .b(output_2_11), .y(output_1_858));
wire output_3_858, output_3_11, output_2_858;
mixer gate_output_2_858(.a(output_3_858), .b(output_3_11), .y(output_2_858));
wire output_4_858, output_4_11, output_3_858;
mixer gate_output_3_858(.a(output_4_858), .b(output_4_11), .y(output_3_858));
wire output_5_858, output_5_11, output_4_858;
mixer gate_output_4_858(.a(output_5_858), .b(output_5_11), .y(output_4_858));
wire output_6_858, output_6_11, output_5_858;
mixer gate_output_5_858(.a(output_6_858), .b(output_6_11), .y(output_5_858));
wire output_7_858, output_7_11, output_6_858;
mixer gate_output_6_858(.a(output_7_858), .b(output_7_11), .y(output_6_858));
wire output_8_858, output_8_11, output_7_858;
mixer gate_output_7_858(.a(output_8_858), .b(output_8_11), .y(output_7_858));
wire output_9_858, output_9_11, output_8_858;
mixer gate_output_8_858(.a(output_9_858), .b(output_9_11), .y(output_8_858));
wire output_10_858, output_10_11, output_9_858;
mixer gate_output_9_858(.a(output_10_858), .b(output_10_11), .y(output_9_858));
wire output_11_858, output_11_11, output_10_858;
mixer gate_output_10_858(.a(output_11_858), .b(output_11_11), .y(output_10_858));
wire output_12_858, output_12_11, output_11_858;
mixer gate_output_11_858(.a(output_12_858), .b(output_12_11), .y(output_11_858));
wire output_13_858, output_13_11, output_12_858;
mixer gate_output_12_858(.a(output_13_858), .b(output_13_11), .y(output_12_858));
wire output_14_858, output_14_11, output_13_858;
mixer gate_output_13_858(.a(output_14_858), .b(output_14_11), .y(output_13_858));
wire output_15_858, output_15_11, output_14_858;
mixer gate_output_14_858(.a(output_15_858), .b(output_15_11), .y(output_14_858));
wire output_16_858, output_16_11, output_15_858;
mixer gate_output_15_858(.a(output_16_858), .b(output_16_11), .y(output_15_858));
wire output_1_859, output_1_12, output_0_859;
mixer gate_output_0_859(.a(output_1_859), .b(output_1_12), .y(output_0_859));
wire output_2_859, output_2_12, output_1_859;
mixer gate_output_1_859(.a(output_2_859), .b(output_2_12), .y(output_1_859));
wire output_3_859, output_3_12, output_2_859;
mixer gate_output_2_859(.a(output_3_859), .b(output_3_12), .y(output_2_859));
wire output_4_859, output_4_12, output_3_859;
mixer gate_output_3_859(.a(output_4_859), .b(output_4_12), .y(output_3_859));
wire output_5_859, output_5_12, output_4_859;
mixer gate_output_4_859(.a(output_5_859), .b(output_5_12), .y(output_4_859));
wire output_6_859, output_6_12, output_5_859;
mixer gate_output_5_859(.a(output_6_859), .b(output_6_12), .y(output_5_859));
wire output_7_859, output_7_12, output_6_859;
mixer gate_output_6_859(.a(output_7_859), .b(output_7_12), .y(output_6_859));
wire output_8_859, output_8_12, output_7_859;
mixer gate_output_7_859(.a(output_8_859), .b(output_8_12), .y(output_7_859));
wire output_9_859, output_9_12, output_8_859;
mixer gate_output_8_859(.a(output_9_859), .b(output_9_12), .y(output_8_859));
wire output_10_859, output_10_12, output_9_859;
mixer gate_output_9_859(.a(output_10_859), .b(output_10_12), .y(output_9_859));
wire output_11_859, output_11_12, output_10_859;
mixer gate_output_10_859(.a(output_11_859), .b(output_11_12), .y(output_10_859));
wire output_12_859, output_12_12, output_11_859;
mixer gate_output_11_859(.a(output_12_859), .b(output_12_12), .y(output_11_859));
wire output_13_859, output_13_12, output_12_859;
mixer gate_output_12_859(.a(output_13_859), .b(output_13_12), .y(output_12_859));
wire output_14_859, output_14_12, output_13_859;
mixer gate_output_13_859(.a(output_14_859), .b(output_14_12), .y(output_13_859));
wire output_15_859, output_15_12, output_14_859;
mixer gate_output_14_859(.a(output_15_859), .b(output_15_12), .y(output_14_859));
wire output_16_859, output_16_12, output_15_859;
mixer gate_output_15_859(.a(output_16_859), .b(output_16_12), .y(output_15_859));
wire output_1_860, output_1_13, output_0_860;
mixer gate_output_0_860(.a(output_1_860), .b(output_1_13), .y(output_0_860));
wire output_2_860, output_2_13, output_1_860;
mixer gate_output_1_860(.a(output_2_860), .b(output_2_13), .y(output_1_860));
wire output_3_860, output_3_13, output_2_860;
mixer gate_output_2_860(.a(output_3_860), .b(output_3_13), .y(output_2_860));
wire output_4_860, output_4_13, output_3_860;
mixer gate_output_3_860(.a(output_4_860), .b(output_4_13), .y(output_3_860));
wire output_5_860, output_5_13, output_4_860;
mixer gate_output_4_860(.a(output_5_860), .b(output_5_13), .y(output_4_860));
wire output_6_860, output_6_13, output_5_860;
mixer gate_output_5_860(.a(output_6_860), .b(output_6_13), .y(output_5_860));
wire output_7_860, output_7_13, output_6_860;
mixer gate_output_6_860(.a(output_7_860), .b(output_7_13), .y(output_6_860));
wire output_8_860, output_8_13, output_7_860;
mixer gate_output_7_860(.a(output_8_860), .b(output_8_13), .y(output_7_860));
wire output_9_860, output_9_13, output_8_860;
mixer gate_output_8_860(.a(output_9_860), .b(output_9_13), .y(output_8_860));
wire output_10_860, output_10_13, output_9_860;
mixer gate_output_9_860(.a(output_10_860), .b(output_10_13), .y(output_9_860));
wire output_11_860, output_11_13, output_10_860;
mixer gate_output_10_860(.a(output_11_860), .b(output_11_13), .y(output_10_860));
wire output_12_860, output_12_13, output_11_860;
mixer gate_output_11_860(.a(output_12_860), .b(output_12_13), .y(output_11_860));
wire output_13_860, output_13_13, output_12_860;
mixer gate_output_12_860(.a(output_13_860), .b(output_13_13), .y(output_12_860));
wire output_14_860, output_14_13, output_13_860;
mixer gate_output_13_860(.a(output_14_860), .b(output_14_13), .y(output_13_860));
wire output_15_860, output_15_13, output_14_860;
mixer gate_output_14_860(.a(output_15_860), .b(output_15_13), .y(output_14_860));
wire output_16_860, output_16_13, output_15_860;
mixer gate_output_15_860(.a(output_16_860), .b(output_16_13), .y(output_15_860));
wire output_1_861, output_1_14, output_0_861;
mixer gate_output_0_861(.a(output_1_861), .b(output_1_14), .y(output_0_861));
wire output_2_861, output_2_14, output_1_861;
mixer gate_output_1_861(.a(output_2_861), .b(output_2_14), .y(output_1_861));
wire output_3_861, output_3_14, output_2_861;
mixer gate_output_2_861(.a(output_3_861), .b(output_3_14), .y(output_2_861));
wire output_4_861, output_4_14, output_3_861;
mixer gate_output_3_861(.a(output_4_861), .b(output_4_14), .y(output_3_861));
wire output_5_861, output_5_14, output_4_861;
mixer gate_output_4_861(.a(output_5_861), .b(output_5_14), .y(output_4_861));
wire output_6_861, output_6_14, output_5_861;
mixer gate_output_5_861(.a(output_6_861), .b(output_6_14), .y(output_5_861));
wire output_7_861, output_7_14, output_6_861;
mixer gate_output_6_861(.a(output_7_861), .b(output_7_14), .y(output_6_861));
wire output_8_861, output_8_14, output_7_861;
mixer gate_output_7_861(.a(output_8_861), .b(output_8_14), .y(output_7_861));
wire output_9_861, output_9_14, output_8_861;
mixer gate_output_8_861(.a(output_9_861), .b(output_9_14), .y(output_8_861));
wire output_10_861, output_10_14, output_9_861;
mixer gate_output_9_861(.a(output_10_861), .b(output_10_14), .y(output_9_861));
wire output_11_861, output_11_14, output_10_861;
mixer gate_output_10_861(.a(output_11_861), .b(output_11_14), .y(output_10_861));
wire output_12_861, output_12_14, output_11_861;
mixer gate_output_11_861(.a(output_12_861), .b(output_12_14), .y(output_11_861));
wire output_13_861, output_13_14, output_12_861;
mixer gate_output_12_861(.a(output_13_861), .b(output_13_14), .y(output_12_861));
wire output_14_861, output_14_14, output_13_861;
mixer gate_output_13_861(.a(output_14_861), .b(output_14_14), .y(output_13_861));
wire output_15_861, output_15_14, output_14_861;
mixer gate_output_14_861(.a(output_15_861), .b(output_15_14), .y(output_14_861));
wire output_16_861, output_16_14, output_15_861;
mixer gate_output_15_861(.a(output_16_861), .b(output_16_14), .y(output_15_861));
wire output_1_862, output_1_15, output_0_862;
mixer gate_output_0_862(.a(output_1_862), .b(output_1_15), .y(output_0_862));
wire output_2_862, output_2_15, output_1_862;
mixer gate_output_1_862(.a(output_2_862), .b(output_2_15), .y(output_1_862));
wire output_3_862, output_3_15, output_2_862;
mixer gate_output_2_862(.a(output_3_862), .b(output_3_15), .y(output_2_862));
wire output_4_862, output_4_15, output_3_862;
mixer gate_output_3_862(.a(output_4_862), .b(output_4_15), .y(output_3_862));
wire output_5_862, output_5_15, output_4_862;
mixer gate_output_4_862(.a(output_5_862), .b(output_5_15), .y(output_4_862));
wire output_6_862, output_6_15, output_5_862;
mixer gate_output_5_862(.a(output_6_862), .b(output_6_15), .y(output_5_862));
wire output_7_862, output_7_15, output_6_862;
mixer gate_output_6_862(.a(output_7_862), .b(output_7_15), .y(output_6_862));
wire output_8_862, output_8_15, output_7_862;
mixer gate_output_7_862(.a(output_8_862), .b(output_8_15), .y(output_7_862));
wire output_9_862, output_9_15, output_8_862;
mixer gate_output_8_862(.a(output_9_862), .b(output_9_15), .y(output_8_862));
wire output_10_862, output_10_15, output_9_862;
mixer gate_output_9_862(.a(output_10_862), .b(output_10_15), .y(output_9_862));
wire output_11_862, output_11_15, output_10_862;
mixer gate_output_10_862(.a(output_11_862), .b(output_11_15), .y(output_10_862));
wire output_12_862, output_12_15, output_11_862;
mixer gate_output_11_862(.a(output_12_862), .b(output_12_15), .y(output_11_862));
wire output_13_862, output_13_15, output_12_862;
mixer gate_output_12_862(.a(output_13_862), .b(output_13_15), .y(output_12_862));
wire output_14_862, output_14_15, output_13_862;
mixer gate_output_13_862(.a(output_14_862), .b(output_14_15), .y(output_13_862));
wire output_15_862, output_15_15, output_14_862;
mixer gate_output_14_862(.a(output_15_862), .b(output_15_15), .y(output_14_862));
wire output_16_862, output_16_15, output_15_862;
mixer gate_output_15_862(.a(output_16_862), .b(output_16_15), .y(output_15_862));
wire output_1_863, output_1_0, output_0_863;
mixer gate_output_0_863(.a(output_1_863), .b(output_1_0), .y(output_0_863));
wire output_2_863, output_2_0, output_1_863;
mixer gate_output_1_863(.a(output_2_863), .b(output_2_0), .y(output_1_863));
wire output_3_863, output_3_0, output_2_863;
mixer gate_output_2_863(.a(output_3_863), .b(output_3_0), .y(output_2_863));
wire output_4_863, output_4_0, output_3_863;
mixer gate_output_3_863(.a(output_4_863), .b(output_4_0), .y(output_3_863));
wire output_5_863, output_5_0, output_4_863;
mixer gate_output_4_863(.a(output_5_863), .b(output_5_0), .y(output_4_863));
wire output_6_863, output_6_0, output_5_863;
mixer gate_output_5_863(.a(output_6_863), .b(output_6_0), .y(output_5_863));
wire output_7_863, output_7_0, output_6_863;
mixer gate_output_6_863(.a(output_7_863), .b(output_7_0), .y(output_6_863));
wire output_8_863, output_8_0, output_7_863;
mixer gate_output_7_863(.a(output_8_863), .b(output_8_0), .y(output_7_863));
wire output_9_863, output_9_0, output_8_863;
mixer gate_output_8_863(.a(output_9_863), .b(output_9_0), .y(output_8_863));
wire output_10_863, output_10_0, output_9_863;
mixer gate_output_9_863(.a(output_10_863), .b(output_10_0), .y(output_9_863));
wire output_11_863, output_11_0, output_10_863;
mixer gate_output_10_863(.a(output_11_863), .b(output_11_0), .y(output_10_863));
wire output_12_863, output_12_0, output_11_863;
mixer gate_output_11_863(.a(output_12_863), .b(output_12_0), .y(output_11_863));
wire output_13_863, output_13_0, output_12_863;
mixer gate_output_12_863(.a(output_13_863), .b(output_13_0), .y(output_12_863));
wire output_14_863, output_14_0, output_13_863;
mixer gate_output_13_863(.a(output_14_863), .b(output_14_0), .y(output_13_863));
wire output_15_863, output_15_0, output_14_863;
mixer gate_output_14_863(.a(output_15_863), .b(output_15_0), .y(output_14_863));
wire output_16_863, output_16_0, output_15_863;
mixer gate_output_15_863(.a(output_16_863), .b(output_16_0), .y(output_15_863));
wire output_1_864, output_1_1, output_0_864;
mixer gate_output_0_864(.a(output_1_864), .b(output_1_1), .y(output_0_864));
wire output_2_864, output_2_1, output_1_864;
mixer gate_output_1_864(.a(output_2_864), .b(output_2_1), .y(output_1_864));
wire output_3_864, output_3_1, output_2_864;
mixer gate_output_2_864(.a(output_3_864), .b(output_3_1), .y(output_2_864));
wire output_4_864, output_4_1, output_3_864;
mixer gate_output_3_864(.a(output_4_864), .b(output_4_1), .y(output_3_864));
wire output_5_864, output_5_1, output_4_864;
mixer gate_output_4_864(.a(output_5_864), .b(output_5_1), .y(output_4_864));
wire output_6_864, output_6_1, output_5_864;
mixer gate_output_5_864(.a(output_6_864), .b(output_6_1), .y(output_5_864));
wire output_7_864, output_7_1, output_6_864;
mixer gate_output_6_864(.a(output_7_864), .b(output_7_1), .y(output_6_864));
wire output_8_864, output_8_1, output_7_864;
mixer gate_output_7_864(.a(output_8_864), .b(output_8_1), .y(output_7_864));
wire output_9_864, output_9_1, output_8_864;
mixer gate_output_8_864(.a(output_9_864), .b(output_9_1), .y(output_8_864));
wire output_10_864, output_10_1, output_9_864;
mixer gate_output_9_864(.a(output_10_864), .b(output_10_1), .y(output_9_864));
wire output_11_864, output_11_1, output_10_864;
mixer gate_output_10_864(.a(output_11_864), .b(output_11_1), .y(output_10_864));
wire output_12_864, output_12_1, output_11_864;
mixer gate_output_11_864(.a(output_12_864), .b(output_12_1), .y(output_11_864));
wire output_13_864, output_13_1, output_12_864;
mixer gate_output_12_864(.a(output_13_864), .b(output_13_1), .y(output_12_864));
wire output_14_864, output_14_1, output_13_864;
mixer gate_output_13_864(.a(output_14_864), .b(output_14_1), .y(output_13_864));
wire output_15_864, output_15_1, output_14_864;
mixer gate_output_14_864(.a(output_15_864), .b(output_15_1), .y(output_14_864));
wire output_16_864, output_16_1, output_15_864;
mixer gate_output_15_864(.a(output_16_864), .b(output_16_1), .y(output_15_864));
wire output_1_865, output_1_2, output_0_865;
mixer gate_output_0_865(.a(output_1_865), .b(output_1_2), .y(output_0_865));
wire output_2_865, output_2_2, output_1_865;
mixer gate_output_1_865(.a(output_2_865), .b(output_2_2), .y(output_1_865));
wire output_3_865, output_3_2, output_2_865;
mixer gate_output_2_865(.a(output_3_865), .b(output_3_2), .y(output_2_865));
wire output_4_865, output_4_2, output_3_865;
mixer gate_output_3_865(.a(output_4_865), .b(output_4_2), .y(output_3_865));
wire output_5_865, output_5_2, output_4_865;
mixer gate_output_4_865(.a(output_5_865), .b(output_5_2), .y(output_4_865));
wire output_6_865, output_6_2, output_5_865;
mixer gate_output_5_865(.a(output_6_865), .b(output_6_2), .y(output_5_865));
wire output_7_865, output_7_2, output_6_865;
mixer gate_output_6_865(.a(output_7_865), .b(output_7_2), .y(output_6_865));
wire output_8_865, output_8_2, output_7_865;
mixer gate_output_7_865(.a(output_8_865), .b(output_8_2), .y(output_7_865));
wire output_9_865, output_9_2, output_8_865;
mixer gate_output_8_865(.a(output_9_865), .b(output_9_2), .y(output_8_865));
wire output_10_865, output_10_2, output_9_865;
mixer gate_output_9_865(.a(output_10_865), .b(output_10_2), .y(output_9_865));
wire output_11_865, output_11_2, output_10_865;
mixer gate_output_10_865(.a(output_11_865), .b(output_11_2), .y(output_10_865));
wire output_12_865, output_12_2, output_11_865;
mixer gate_output_11_865(.a(output_12_865), .b(output_12_2), .y(output_11_865));
wire output_13_865, output_13_2, output_12_865;
mixer gate_output_12_865(.a(output_13_865), .b(output_13_2), .y(output_12_865));
wire output_14_865, output_14_2, output_13_865;
mixer gate_output_13_865(.a(output_14_865), .b(output_14_2), .y(output_13_865));
wire output_15_865, output_15_2, output_14_865;
mixer gate_output_14_865(.a(output_15_865), .b(output_15_2), .y(output_14_865));
wire output_16_865, output_16_2, output_15_865;
mixer gate_output_15_865(.a(output_16_865), .b(output_16_2), .y(output_15_865));
wire output_1_866, output_1_3, output_0_866;
mixer gate_output_0_866(.a(output_1_866), .b(output_1_3), .y(output_0_866));
wire output_2_866, output_2_3, output_1_866;
mixer gate_output_1_866(.a(output_2_866), .b(output_2_3), .y(output_1_866));
wire output_3_866, output_3_3, output_2_866;
mixer gate_output_2_866(.a(output_3_866), .b(output_3_3), .y(output_2_866));
wire output_4_866, output_4_3, output_3_866;
mixer gate_output_3_866(.a(output_4_866), .b(output_4_3), .y(output_3_866));
wire output_5_866, output_5_3, output_4_866;
mixer gate_output_4_866(.a(output_5_866), .b(output_5_3), .y(output_4_866));
wire output_6_866, output_6_3, output_5_866;
mixer gate_output_5_866(.a(output_6_866), .b(output_6_3), .y(output_5_866));
wire output_7_866, output_7_3, output_6_866;
mixer gate_output_6_866(.a(output_7_866), .b(output_7_3), .y(output_6_866));
wire output_8_866, output_8_3, output_7_866;
mixer gate_output_7_866(.a(output_8_866), .b(output_8_3), .y(output_7_866));
wire output_9_866, output_9_3, output_8_866;
mixer gate_output_8_866(.a(output_9_866), .b(output_9_3), .y(output_8_866));
wire output_10_866, output_10_3, output_9_866;
mixer gate_output_9_866(.a(output_10_866), .b(output_10_3), .y(output_9_866));
wire output_11_866, output_11_3, output_10_866;
mixer gate_output_10_866(.a(output_11_866), .b(output_11_3), .y(output_10_866));
wire output_12_866, output_12_3, output_11_866;
mixer gate_output_11_866(.a(output_12_866), .b(output_12_3), .y(output_11_866));
wire output_13_866, output_13_3, output_12_866;
mixer gate_output_12_866(.a(output_13_866), .b(output_13_3), .y(output_12_866));
wire output_14_866, output_14_3, output_13_866;
mixer gate_output_13_866(.a(output_14_866), .b(output_14_3), .y(output_13_866));
wire output_15_866, output_15_3, output_14_866;
mixer gate_output_14_866(.a(output_15_866), .b(output_15_3), .y(output_14_866));
wire output_16_866, output_16_3, output_15_866;
mixer gate_output_15_866(.a(output_16_866), .b(output_16_3), .y(output_15_866));
wire output_1_867, output_1_4, output_0_867;
mixer gate_output_0_867(.a(output_1_867), .b(output_1_4), .y(output_0_867));
wire output_2_867, output_2_4, output_1_867;
mixer gate_output_1_867(.a(output_2_867), .b(output_2_4), .y(output_1_867));
wire output_3_867, output_3_4, output_2_867;
mixer gate_output_2_867(.a(output_3_867), .b(output_3_4), .y(output_2_867));
wire output_4_867, output_4_4, output_3_867;
mixer gate_output_3_867(.a(output_4_867), .b(output_4_4), .y(output_3_867));
wire output_5_867, output_5_4, output_4_867;
mixer gate_output_4_867(.a(output_5_867), .b(output_5_4), .y(output_4_867));
wire output_6_867, output_6_4, output_5_867;
mixer gate_output_5_867(.a(output_6_867), .b(output_6_4), .y(output_5_867));
wire output_7_867, output_7_4, output_6_867;
mixer gate_output_6_867(.a(output_7_867), .b(output_7_4), .y(output_6_867));
wire output_8_867, output_8_4, output_7_867;
mixer gate_output_7_867(.a(output_8_867), .b(output_8_4), .y(output_7_867));
wire output_9_867, output_9_4, output_8_867;
mixer gate_output_8_867(.a(output_9_867), .b(output_9_4), .y(output_8_867));
wire output_10_867, output_10_4, output_9_867;
mixer gate_output_9_867(.a(output_10_867), .b(output_10_4), .y(output_9_867));
wire output_11_867, output_11_4, output_10_867;
mixer gate_output_10_867(.a(output_11_867), .b(output_11_4), .y(output_10_867));
wire output_12_867, output_12_4, output_11_867;
mixer gate_output_11_867(.a(output_12_867), .b(output_12_4), .y(output_11_867));
wire output_13_867, output_13_4, output_12_867;
mixer gate_output_12_867(.a(output_13_867), .b(output_13_4), .y(output_12_867));
wire output_14_867, output_14_4, output_13_867;
mixer gate_output_13_867(.a(output_14_867), .b(output_14_4), .y(output_13_867));
wire output_15_867, output_15_4, output_14_867;
mixer gate_output_14_867(.a(output_15_867), .b(output_15_4), .y(output_14_867));
wire output_16_867, output_16_4, output_15_867;
mixer gate_output_15_867(.a(output_16_867), .b(output_16_4), .y(output_15_867));
wire output_1_868, output_1_5, output_0_868;
mixer gate_output_0_868(.a(output_1_868), .b(output_1_5), .y(output_0_868));
wire output_2_868, output_2_5, output_1_868;
mixer gate_output_1_868(.a(output_2_868), .b(output_2_5), .y(output_1_868));
wire output_3_868, output_3_5, output_2_868;
mixer gate_output_2_868(.a(output_3_868), .b(output_3_5), .y(output_2_868));
wire output_4_868, output_4_5, output_3_868;
mixer gate_output_3_868(.a(output_4_868), .b(output_4_5), .y(output_3_868));
wire output_5_868, output_5_5, output_4_868;
mixer gate_output_4_868(.a(output_5_868), .b(output_5_5), .y(output_4_868));
wire output_6_868, output_6_5, output_5_868;
mixer gate_output_5_868(.a(output_6_868), .b(output_6_5), .y(output_5_868));
wire output_7_868, output_7_5, output_6_868;
mixer gate_output_6_868(.a(output_7_868), .b(output_7_5), .y(output_6_868));
wire output_8_868, output_8_5, output_7_868;
mixer gate_output_7_868(.a(output_8_868), .b(output_8_5), .y(output_7_868));
wire output_9_868, output_9_5, output_8_868;
mixer gate_output_8_868(.a(output_9_868), .b(output_9_5), .y(output_8_868));
wire output_10_868, output_10_5, output_9_868;
mixer gate_output_9_868(.a(output_10_868), .b(output_10_5), .y(output_9_868));
wire output_11_868, output_11_5, output_10_868;
mixer gate_output_10_868(.a(output_11_868), .b(output_11_5), .y(output_10_868));
wire output_12_868, output_12_5, output_11_868;
mixer gate_output_11_868(.a(output_12_868), .b(output_12_5), .y(output_11_868));
wire output_13_868, output_13_5, output_12_868;
mixer gate_output_12_868(.a(output_13_868), .b(output_13_5), .y(output_12_868));
wire output_14_868, output_14_5, output_13_868;
mixer gate_output_13_868(.a(output_14_868), .b(output_14_5), .y(output_13_868));
wire output_15_868, output_15_5, output_14_868;
mixer gate_output_14_868(.a(output_15_868), .b(output_15_5), .y(output_14_868));
wire output_16_868, output_16_5, output_15_868;
mixer gate_output_15_868(.a(output_16_868), .b(output_16_5), .y(output_15_868));
wire output_1_869, output_1_6, output_0_869;
mixer gate_output_0_869(.a(output_1_869), .b(output_1_6), .y(output_0_869));
wire output_2_869, output_2_6, output_1_869;
mixer gate_output_1_869(.a(output_2_869), .b(output_2_6), .y(output_1_869));
wire output_3_869, output_3_6, output_2_869;
mixer gate_output_2_869(.a(output_3_869), .b(output_3_6), .y(output_2_869));
wire output_4_869, output_4_6, output_3_869;
mixer gate_output_3_869(.a(output_4_869), .b(output_4_6), .y(output_3_869));
wire output_5_869, output_5_6, output_4_869;
mixer gate_output_4_869(.a(output_5_869), .b(output_5_6), .y(output_4_869));
wire output_6_869, output_6_6, output_5_869;
mixer gate_output_5_869(.a(output_6_869), .b(output_6_6), .y(output_5_869));
wire output_7_869, output_7_6, output_6_869;
mixer gate_output_6_869(.a(output_7_869), .b(output_7_6), .y(output_6_869));
wire output_8_869, output_8_6, output_7_869;
mixer gate_output_7_869(.a(output_8_869), .b(output_8_6), .y(output_7_869));
wire output_9_869, output_9_6, output_8_869;
mixer gate_output_8_869(.a(output_9_869), .b(output_9_6), .y(output_8_869));
wire output_10_869, output_10_6, output_9_869;
mixer gate_output_9_869(.a(output_10_869), .b(output_10_6), .y(output_9_869));
wire output_11_869, output_11_6, output_10_869;
mixer gate_output_10_869(.a(output_11_869), .b(output_11_6), .y(output_10_869));
wire output_12_869, output_12_6, output_11_869;
mixer gate_output_11_869(.a(output_12_869), .b(output_12_6), .y(output_11_869));
wire output_13_869, output_13_6, output_12_869;
mixer gate_output_12_869(.a(output_13_869), .b(output_13_6), .y(output_12_869));
wire output_14_869, output_14_6, output_13_869;
mixer gate_output_13_869(.a(output_14_869), .b(output_14_6), .y(output_13_869));
wire output_15_869, output_15_6, output_14_869;
mixer gate_output_14_869(.a(output_15_869), .b(output_15_6), .y(output_14_869));
wire output_16_869, output_16_6, output_15_869;
mixer gate_output_15_869(.a(output_16_869), .b(output_16_6), .y(output_15_869));
wire output_1_870, output_1_7, output_0_870;
mixer gate_output_0_870(.a(output_1_870), .b(output_1_7), .y(output_0_870));
wire output_2_870, output_2_7, output_1_870;
mixer gate_output_1_870(.a(output_2_870), .b(output_2_7), .y(output_1_870));
wire output_3_870, output_3_7, output_2_870;
mixer gate_output_2_870(.a(output_3_870), .b(output_3_7), .y(output_2_870));
wire output_4_870, output_4_7, output_3_870;
mixer gate_output_3_870(.a(output_4_870), .b(output_4_7), .y(output_3_870));
wire output_5_870, output_5_7, output_4_870;
mixer gate_output_4_870(.a(output_5_870), .b(output_5_7), .y(output_4_870));
wire output_6_870, output_6_7, output_5_870;
mixer gate_output_5_870(.a(output_6_870), .b(output_6_7), .y(output_5_870));
wire output_7_870, output_7_7, output_6_870;
mixer gate_output_6_870(.a(output_7_870), .b(output_7_7), .y(output_6_870));
wire output_8_870, output_8_7, output_7_870;
mixer gate_output_7_870(.a(output_8_870), .b(output_8_7), .y(output_7_870));
wire output_9_870, output_9_7, output_8_870;
mixer gate_output_8_870(.a(output_9_870), .b(output_9_7), .y(output_8_870));
wire output_10_870, output_10_7, output_9_870;
mixer gate_output_9_870(.a(output_10_870), .b(output_10_7), .y(output_9_870));
wire output_11_870, output_11_7, output_10_870;
mixer gate_output_10_870(.a(output_11_870), .b(output_11_7), .y(output_10_870));
wire output_12_870, output_12_7, output_11_870;
mixer gate_output_11_870(.a(output_12_870), .b(output_12_7), .y(output_11_870));
wire output_13_870, output_13_7, output_12_870;
mixer gate_output_12_870(.a(output_13_870), .b(output_13_7), .y(output_12_870));
wire output_14_870, output_14_7, output_13_870;
mixer gate_output_13_870(.a(output_14_870), .b(output_14_7), .y(output_13_870));
wire output_15_870, output_15_7, output_14_870;
mixer gate_output_14_870(.a(output_15_870), .b(output_15_7), .y(output_14_870));
wire output_16_870, output_16_7, output_15_870;
mixer gate_output_15_870(.a(output_16_870), .b(output_16_7), .y(output_15_870));
wire output_1_871, output_1_8, output_0_871;
mixer gate_output_0_871(.a(output_1_871), .b(output_1_8), .y(output_0_871));
wire output_2_871, output_2_8, output_1_871;
mixer gate_output_1_871(.a(output_2_871), .b(output_2_8), .y(output_1_871));
wire output_3_871, output_3_8, output_2_871;
mixer gate_output_2_871(.a(output_3_871), .b(output_3_8), .y(output_2_871));
wire output_4_871, output_4_8, output_3_871;
mixer gate_output_3_871(.a(output_4_871), .b(output_4_8), .y(output_3_871));
wire output_5_871, output_5_8, output_4_871;
mixer gate_output_4_871(.a(output_5_871), .b(output_5_8), .y(output_4_871));
wire output_6_871, output_6_8, output_5_871;
mixer gate_output_5_871(.a(output_6_871), .b(output_6_8), .y(output_5_871));
wire output_7_871, output_7_8, output_6_871;
mixer gate_output_6_871(.a(output_7_871), .b(output_7_8), .y(output_6_871));
wire output_8_871, output_8_8, output_7_871;
mixer gate_output_7_871(.a(output_8_871), .b(output_8_8), .y(output_7_871));
wire output_9_871, output_9_8, output_8_871;
mixer gate_output_8_871(.a(output_9_871), .b(output_9_8), .y(output_8_871));
wire output_10_871, output_10_8, output_9_871;
mixer gate_output_9_871(.a(output_10_871), .b(output_10_8), .y(output_9_871));
wire output_11_871, output_11_8, output_10_871;
mixer gate_output_10_871(.a(output_11_871), .b(output_11_8), .y(output_10_871));
wire output_12_871, output_12_8, output_11_871;
mixer gate_output_11_871(.a(output_12_871), .b(output_12_8), .y(output_11_871));
wire output_13_871, output_13_8, output_12_871;
mixer gate_output_12_871(.a(output_13_871), .b(output_13_8), .y(output_12_871));
wire output_14_871, output_14_8, output_13_871;
mixer gate_output_13_871(.a(output_14_871), .b(output_14_8), .y(output_13_871));
wire output_15_871, output_15_8, output_14_871;
mixer gate_output_14_871(.a(output_15_871), .b(output_15_8), .y(output_14_871));
wire output_16_871, output_16_8, output_15_871;
mixer gate_output_15_871(.a(output_16_871), .b(output_16_8), .y(output_15_871));
wire output_1_872, output_1_9, output_0_872;
mixer gate_output_0_872(.a(output_1_872), .b(output_1_9), .y(output_0_872));
wire output_2_872, output_2_9, output_1_872;
mixer gate_output_1_872(.a(output_2_872), .b(output_2_9), .y(output_1_872));
wire output_3_872, output_3_9, output_2_872;
mixer gate_output_2_872(.a(output_3_872), .b(output_3_9), .y(output_2_872));
wire output_4_872, output_4_9, output_3_872;
mixer gate_output_3_872(.a(output_4_872), .b(output_4_9), .y(output_3_872));
wire output_5_872, output_5_9, output_4_872;
mixer gate_output_4_872(.a(output_5_872), .b(output_5_9), .y(output_4_872));
wire output_6_872, output_6_9, output_5_872;
mixer gate_output_5_872(.a(output_6_872), .b(output_6_9), .y(output_5_872));
wire output_7_872, output_7_9, output_6_872;
mixer gate_output_6_872(.a(output_7_872), .b(output_7_9), .y(output_6_872));
wire output_8_872, output_8_9, output_7_872;
mixer gate_output_7_872(.a(output_8_872), .b(output_8_9), .y(output_7_872));
wire output_9_872, output_9_9, output_8_872;
mixer gate_output_8_872(.a(output_9_872), .b(output_9_9), .y(output_8_872));
wire output_10_872, output_10_9, output_9_872;
mixer gate_output_9_872(.a(output_10_872), .b(output_10_9), .y(output_9_872));
wire output_11_872, output_11_9, output_10_872;
mixer gate_output_10_872(.a(output_11_872), .b(output_11_9), .y(output_10_872));
wire output_12_872, output_12_9, output_11_872;
mixer gate_output_11_872(.a(output_12_872), .b(output_12_9), .y(output_11_872));
wire output_13_872, output_13_9, output_12_872;
mixer gate_output_12_872(.a(output_13_872), .b(output_13_9), .y(output_12_872));
wire output_14_872, output_14_9, output_13_872;
mixer gate_output_13_872(.a(output_14_872), .b(output_14_9), .y(output_13_872));
wire output_15_872, output_15_9, output_14_872;
mixer gate_output_14_872(.a(output_15_872), .b(output_15_9), .y(output_14_872));
wire output_16_872, output_16_9, output_15_872;
mixer gate_output_15_872(.a(output_16_872), .b(output_16_9), .y(output_15_872));
wire output_1_873, output_1_10, output_0_873;
mixer gate_output_0_873(.a(output_1_873), .b(output_1_10), .y(output_0_873));
wire output_2_873, output_2_10, output_1_873;
mixer gate_output_1_873(.a(output_2_873), .b(output_2_10), .y(output_1_873));
wire output_3_873, output_3_10, output_2_873;
mixer gate_output_2_873(.a(output_3_873), .b(output_3_10), .y(output_2_873));
wire output_4_873, output_4_10, output_3_873;
mixer gate_output_3_873(.a(output_4_873), .b(output_4_10), .y(output_3_873));
wire output_5_873, output_5_10, output_4_873;
mixer gate_output_4_873(.a(output_5_873), .b(output_5_10), .y(output_4_873));
wire output_6_873, output_6_10, output_5_873;
mixer gate_output_5_873(.a(output_6_873), .b(output_6_10), .y(output_5_873));
wire output_7_873, output_7_10, output_6_873;
mixer gate_output_6_873(.a(output_7_873), .b(output_7_10), .y(output_6_873));
wire output_8_873, output_8_10, output_7_873;
mixer gate_output_7_873(.a(output_8_873), .b(output_8_10), .y(output_7_873));
wire output_9_873, output_9_10, output_8_873;
mixer gate_output_8_873(.a(output_9_873), .b(output_9_10), .y(output_8_873));
wire output_10_873, output_10_10, output_9_873;
mixer gate_output_9_873(.a(output_10_873), .b(output_10_10), .y(output_9_873));
wire output_11_873, output_11_10, output_10_873;
mixer gate_output_10_873(.a(output_11_873), .b(output_11_10), .y(output_10_873));
wire output_12_873, output_12_10, output_11_873;
mixer gate_output_11_873(.a(output_12_873), .b(output_12_10), .y(output_11_873));
wire output_13_873, output_13_10, output_12_873;
mixer gate_output_12_873(.a(output_13_873), .b(output_13_10), .y(output_12_873));
wire output_14_873, output_14_10, output_13_873;
mixer gate_output_13_873(.a(output_14_873), .b(output_14_10), .y(output_13_873));
wire output_15_873, output_15_10, output_14_873;
mixer gate_output_14_873(.a(output_15_873), .b(output_15_10), .y(output_14_873));
wire output_16_873, output_16_10, output_15_873;
mixer gate_output_15_873(.a(output_16_873), .b(output_16_10), .y(output_15_873));
wire output_1_874, output_1_11, output_0_874;
mixer gate_output_0_874(.a(output_1_874), .b(output_1_11), .y(output_0_874));
wire output_2_874, output_2_11, output_1_874;
mixer gate_output_1_874(.a(output_2_874), .b(output_2_11), .y(output_1_874));
wire output_3_874, output_3_11, output_2_874;
mixer gate_output_2_874(.a(output_3_874), .b(output_3_11), .y(output_2_874));
wire output_4_874, output_4_11, output_3_874;
mixer gate_output_3_874(.a(output_4_874), .b(output_4_11), .y(output_3_874));
wire output_5_874, output_5_11, output_4_874;
mixer gate_output_4_874(.a(output_5_874), .b(output_5_11), .y(output_4_874));
wire output_6_874, output_6_11, output_5_874;
mixer gate_output_5_874(.a(output_6_874), .b(output_6_11), .y(output_5_874));
wire output_7_874, output_7_11, output_6_874;
mixer gate_output_6_874(.a(output_7_874), .b(output_7_11), .y(output_6_874));
wire output_8_874, output_8_11, output_7_874;
mixer gate_output_7_874(.a(output_8_874), .b(output_8_11), .y(output_7_874));
wire output_9_874, output_9_11, output_8_874;
mixer gate_output_8_874(.a(output_9_874), .b(output_9_11), .y(output_8_874));
wire output_10_874, output_10_11, output_9_874;
mixer gate_output_9_874(.a(output_10_874), .b(output_10_11), .y(output_9_874));
wire output_11_874, output_11_11, output_10_874;
mixer gate_output_10_874(.a(output_11_874), .b(output_11_11), .y(output_10_874));
wire output_12_874, output_12_11, output_11_874;
mixer gate_output_11_874(.a(output_12_874), .b(output_12_11), .y(output_11_874));
wire output_13_874, output_13_11, output_12_874;
mixer gate_output_12_874(.a(output_13_874), .b(output_13_11), .y(output_12_874));
wire output_14_874, output_14_11, output_13_874;
mixer gate_output_13_874(.a(output_14_874), .b(output_14_11), .y(output_13_874));
wire output_15_874, output_15_11, output_14_874;
mixer gate_output_14_874(.a(output_15_874), .b(output_15_11), .y(output_14_874));
wire output_16_874, output_16_11, output_15_874;
mixer gate_output_15_874(.a(output_16_874), .b(output_16_11), .y(output_15_874));
wire output_1_875, output_1_12, output_0_875;
mixer gate_output_0_875(.a(output_1_875), .b(output_1_12), .y(output_0_875));
wire output_2_875, output_2_12, output_1_875;
mixer gate_output_1_875(.a(output_2_875), .b(output_2_12), .y(output_1_875));
wire output_3_875, output_3_12, output_2_875;
mixer gate_output_2_875(.a(output_3_875), .b(output_3_12), .y(output_2_875));
wire output_4_875, output_4_12, output_3_875;
mixer gate_output_3_875(.a(output_4_875), .b(output_4_12), .y(output_3_875));
wire output_5_875, output_5_12, output_4_875;
mixer gate_output_4_875(.a(output_5_875), .b(output_5_12), .y(output_4_875));
wire output_6_875, output_6_12, output_5_875;
mixer gate_output_5_875(.a(output_6_875), .b(output_6_12), .y(output_5_875));
wire output_7_875, output_7_12, output_6_875;
mixer gate_output_6_875(.a(output_7_875), .b(output_7_12), .y(output_6_875));
wire output_8_875, output_8_12, output_7_875;
mixer gate_output_7_875(.a(output_8_875), .b(output_8_12), .y(output_7_875));
wire output_9_875, output_9_12, output_8_875;
mixer gate_output_8_875(.a(output_9_875), .b(output_9_12), .y(output_8_875));
wire output_10_875, output_10_12, output_9_875;
mixer gate_output_9_875(.a(output_10_875), .b(output_10_12), .y(output_9_875));
wire output_11_875, output_11_12, output_10_875;
mixer gate_output_10_875(.a(output_11_875), .b(output_11_12), .y(output_10_875));
wire output_12_875, output_12_12, output_11_875;
mixer gate_output_11_875(.a(output_12_875), .b(output_12_12), .y(output_11_875));
wire output_13_875, output_13_12, output_12_875;
mixer gate_output_12_875(.a(output_13_875), .b(output_13_12), .y(output_12_875));
wire output_14_875, output_14_12, output_13_875;
mixer gate_output_13_875(.a(output_14_875), .b(output_14_12), .y(output_13_875));
wire output_15_875, output_15_12, output_14_875;
mixer gate_output_14_875(.a(output_15_875), .b(output_15_12), .y(output_14_875));
wire output_16_875, output_16_12, output_15_875;
mixer gate_output_15_875(.a(output_16_875), .b(output_16_12), .y(output_15_875));
wire output_1_876, output_1_13, output_0_876;
mixer gate_output_0_876(.a(output_1_876), .b(output_1_13), .y(output_0_876));
wire output_2_876, output_2_13, output_1_876;
mixer gate_output_1_876(.a(output_2_876), .b(output_2_13), .y(output_1_876));
wire output_3_876, output_3_13, output_2_876;
mixer gate_output_2_876(.a(output_3_876), .b(output_3_13), .y(output_2_876));
wire output_4_876, output_4_13, output_3_876;
mixer gate_output_3_876(.a(output_4_876), .b(output_4_13), .y(output_3_876));
wire output_5_876, output_5_13, output_4_876;
mixer gate_output_4_876(.a(output_5_876), .b(output_5_13), .y(output_4_876));
wire output_6_876, output_6_13, output_5_876;
mixer gate_output_5_876(.a(output_6_876), .b(output_6_13), .y(output_5_876));
wire output_7_876, output_7_13, output_6_876;
mixer gate_output_6_876(.a(output_7_876), .b(output_7_13), .y(output_6_876));
wire output_8_876, output_8_13, output_7_876;
mixer gate_output_7_876(.a(output_8_876), .b(output_8_13), .y(output_7_876));
wire output_9_876, output_9_13, output_8_876;
mixer gate_output_8_876(.a(output_9_876), .b(output_9_13), .y(output_8_876));
wire output_10_876, output_10_13, output_9_876;
mixer gate_output_9_876(.a(output_10_876), .b(output_10_13), .y(output_9_876));
wire output_11_876, output_11_13, output_10_876;
mixer gate_output_10_876(.a(output_11_876), .b(output_11_13), .y(output_10_876));
wire output_12_876, output_12_13, output_11_876;
mixer gate_output_11_876(.a(output_12_876), .b(output_12_13), .y(output_11_876));
wire output_13_876, output_13_13, output_12_876;
mixer gate_output_12_876(.a(output_13_876), .b(output_13_13), .y(output_12_876));
wire output_14_876, output_14_13, output_13_876;
mixer gate_output_13_876(.a(output_14_876), .b(output_14_13), .y(output_13_876));
wire output_15_876, output_15_13, output_14_876;
mixer gate_output_14_876(.a(output_15_876), .b(output_15_13), .y(output_14_876));
wire output_16_876, output_16_13, output_15_876;
mixer gate_output_15_876(.a(output_16_876), .b(output_16_13), .y(output_15_876));
wire output_1_877, output_1_14, output_0_877;
mixer gate_output_0_877(.a(output_1_877), .b(output_1_14), .y(output_0_877));
wire output_2_877, output_2_14, output_1_877;
mixer gate_output_1_877(.a(output_2_877), .b(output_2_14), .y(output_1_877));
wire output_3_877, output_3_14, output_2_877;
mixer gate_output_2_877(.a(output_3_877), .b(output_3_14), .y(output_2_877));
wire output_4_877, output_4_14, output_3_877;
mixer gate_output_3_877(.a(output_4_877), .b(output_4_14), .y(output_3_877));
wire output_5_877, output_5_14, output_4_877;
mixer gate_output_4_877(.a(output_5_877), .b(output_5_14), .y(output_4_877));
wire output_6_877, output_6_14, output_5_877;
mixer gate_output_5_877(.a(output_6_877), .b(output_6_14), .y(output_5_877));
wire output_7_877, output_7_14, output_6_877;
mixer gate_output_6_877(.a(output_7_877), .b(output_7_14), .y(output_6_877));
wire output_8_877, output_8_14, output_7_877;
mixer gate_output_7_877(.a(output_8_877), .b(output_8_14), .y(output_7_877));
wire output_9_877, output_9_14, output_8_877;
mixer gate_output_8_877(.a(output_9_877), .b(output_9_14), .y(output_8_877));
wire output_10_877, output_10_14, output_9_877;
mixer gate_output_9_877(.a(output_10_877), .b(output_10_14), .y(output_9_877));
wire output_11_877, output_11_14, output_10_877;
mixer gate_output_10_877(.a(output_11_877), .b(output_11_14), .y(output_10_877));
wire output_12_877, output_12_14, output_11_877;
mixer gate_output_11_877(.a(output_12_877), .b(output_12_14), .y(output_11_877));
wire output_13_877, output_13_14, output_12_877;
mixer gate_output_12_877(.a(output_13_877), .b(output_13_14), .y(output_12_877));
wire output_14_877, output_14_14, output_13_877;
mixer gate_output_13_877(.a(output_14_877), .b(output_14_14), .y(output_13_877));
wire output_15_877, output_15_14, output_14_877;
mixer gate_output_14_877(.a(output_15_877), .b(output_15_14), .y(output_14_877));
wire output_16_877, output_16_14, output_15_877;
mixer gate_output_15_877(.a(output_16_877), .b(output_16_14), .y(output_15_877));
wire output_1_878, output_1_15, output_0_878;
mixer gate_output_0_878(.a(output_1_878), .b(output_1_15), .y(output_0_878));
wire output_2_878, output_2_15, output_1_878;
mixer gate_output_1_878(.a(output_2_878), .b(output_2_15), .y(output_1_878));
wire output_3_878, output_3_15, output_2_878;
mixer gate_output_2_878(.a(output_3_878), .b(output_3_15), .y(output_2_878));
wire output_4_878, output_4_15, output_3_878;
mixer gate_output_3_878(.a(output_4_878), .b(output_4_15), .y(output_3_878));
wire output_5_878, output_5_15, output_4_878;
mixer gate_output_4_878(.a(output_5_878), .b(output_5_15), .y(output_4_878));
wire output_6_878, output_6_15, output_5_878;
mixer gate_output_5_878(.a(output_6_878), .b(output_6_15), .y(output_5_878));
wire output_7_878, output_7_15, output_6_878;
mixer gate_output_6_878(.a(output_7_878), .b(output_7_15), .y(output_6_878));
wire output_8_878, output_8_15, output_7_878;
mixer gate_output_7_878(.a(output_8_878), .b(output_8_15), .y(output_7_878));
wire output_9_878, output_9_15, output_8_878;
mixer gate_output_8_878(.a(output_9_878), .b(output_9_15), .y(output_8_878));
wire output_10_878, output_10_15, output_9_878;
mixer gate_output_9_878(.a(output_10_878), .b(output_10_15), .y(output_9_878));
wire output_11_878, output_11_15, output_10_878;
mixer gate_output_10_878(.a(output_11_878), .b(output_11_15), .y(output_10_878));
wire output_12_878, output_12_15, output_11_878;
mixer gate_output_11_878(.a(output_12_878), .b(output_12_15), .y(output_11_878));
wire output_13_878, output_13_15, output_12_878;
mixer gate_output_12_878(.a(output_13_878), .b(output_13_15), .y(output_12_878));
wire output_14_878, output_14_15, output_13_878;
mixer gate_output_13_878(.a(output_14_878), .b(output_14_15), .y(output_13_878));
wire output_15_878, output_15_15, output_14_878;
mixer gate_output_14_878(.a(output_15_878), .b(output_15_15), .y(output_14_878));
wire output_16_878, output_16_15, output_15_878;
mixer gate_output_15_878(.a(output_16_878), .b(output_16_15), .y(output_15_878));
wire output_1_879, output_1_0, output_0_879;
mixer gate_output_0_879(.a(output_1_879), .b(output_1_0), .y(output_0_879));
wire output_2_879, output_2_0, output_1_879;
mixer gate_output_1_879(.a(output_2_879), .b(output_2_0), .y(output_1_879));
wire output_3_879, output_3_0, output_2_879;
mixer gate_output_2_879(.a(output_3_879), .b(output_3_0), .y(output_2_879));
wire output_4_879, output_4_0, output_3_879;
mixer gate_output_3_879(.a(output_4_879), .b(output_4_0), .y(output_3_879));
wire output_5_879, output_5_0, output_4_879;
mixer gate_output_4_879(.a(output_5_879), .b(output_5_0), .y(output_4_879));
wire output_6_879, output_6_0, output_5_879;
mixer gate_output_5_879(.a(output_6_879), .b(output_6_0), .y(output_5_879));
wire output_7_879, output_7_0, output_6_879;
mixer gate_output_6_879(.a(output_7_879), .b(output_7_0), .y(output_6_879));
wire output_8_879, output_8_0, output_7_879;
mixer gate_output_7_879(.a(output_8_879), .b(output_8_0), .y(output_7_879));
wire output_9_879, output_9_0, output_8_879;
mixer gate_output_8_879(.a(output_9_879), .b(output_9_0), .y(output_8_879));
wire output_10_879, output_10_0, output_9_879;
mixer gate_output_9_879(.a(output_10_879), .b(output_10_0), .y(output_9_879));
wire output_11_879, output_11_0, output_10_879;
mixer gate_output_10_879(.a(output_11_879), .b(output_11_0), .y(output_10_879));
wire output_12_879, output_12_0, output_11_879;
mixer gate_output_11_879(.a(output_12_879), .b(output_12_0), .y(output_11_879));
wire output_13_879, output_13_0, output_12_879;
mixer gate_output_12_879(.a(output_13_879), .b(output_13_0), .y(output_12_879));
wire output_14_879, output_14_0, output_13_879;
mixer gate_output_13_879(.a(output_14_879), .b(output_14_0), .y(output_13_879));
wire output_15_879, output_15_0, output_14_879;
mixer gate_output_14_879(.a(output_15_879), .b(output_15_0), .y(output_14_879));
wire output_16_879, output_16_0, output_15_879;
mixer gate_output_15_879(.a(output_16_879), .b(output_16_0), .y(output_15_879));
wire output_1_880, output_1_1, output_0_880;
mixer gate_output_0_880(.a(output_1_880), .b(output_1_1), .y(output_0_880));
wire output_2_880, output_2_1, output_1_880;
mixer gate_output_1_880(.a(output_2_880), .b(output_2_1), .y(output_1_880));
wire output_3_880, output_3_1, output_2_880;
mixer gate_output_2_880(.a(output_3_880), .b(output_3_1), .y(output_2_880));
wire output_4_880, output_4_1, output_3_880;
mixer gate_output_3_880(.a(output_4_880), .b(output_4_1), .y(output_3_880));
wire output_5_880, output_5_1, output_4_880;
mixer gate_output_4_880(.a(output_5_880), .b(output_5_1), .y(output_4_880));
wire output_6_880, output_6_1, output_5_880;
mixer gate_output_5_880(.a(output_6_880), .b(output_6_1), .y(output_5_880));
wire output_7_880, output_7_1, output_6_880;
mixer gate_output_6_880(.a(output_7_880), .b(output_7_1), .y(output_6_880));
wire output_8_880, output_8_1, output_7_880;
mixer gate_output_7_880(.a(output_8_880), .b(output_8_1), .y(output_7_880));
wire output_9_880, output_9_1, output_8_880;
mixer gate_output_8_880(.a(output_9_880), .b(output_9_1), .y(output_8_880));
wire output_10_880, output_10_1, output_9_880;
mixer gate_output_9_880(.a(output_10_880), .b(output_10_1), .y(output_9_880));
wire output_11_880, output_11_1, output_10_880;
mixer gate_output_10_880(.a(output_11_880), .b(output_11_1), .y(output_10_880));
wire output_12_880, output_12_1, output_11_880;
mixer gate_output_11_880(.a(output_12_880), .b(output_12_1), .y(output_11_880));
wire output_13_880, output_13_1, output_12_880;
mixer gate_output_12_880(.a(output_13_880), .b(output_13_1), .y(output_12_880));
wire output_14_880, output_14_1, output_13_880;
mixer gate_output_13_880(.a(output_14_880), .b(output_14_1), .y(output_13_880));
wire output_15_880, output_15_1, output_14_880;
mixer gate_output_14_880(.a(output_15_880), .b(output_15_1), .y(output_14_880));
wire output_16_880, output_16_1, output_15_880;
mixer gate_output_15_880(.a(output_16_880), .b(output_16_1), .y(output_15_880));
wire output_1_881, output_1_2, output_0_881;
mixer gate_output_0_881(.a(output_1_881), .b(output_1_2), .y(output_0_881));
wire output_2_881, output_2_2, output_1_881;
mixer gate_output_1_881(.a(output_2_881), .b(output_2_2), .y(output_1_881));
wire output_3_881, output_3_2, output_2_881;
mixer gate_output_2_881(.a(output_3_881), .b(output_3_2), .y(output_2_881));
wire output_4_881, output_4_2, output_3_881;
mixer gate_output_3_881(.a(output_4_881), .b(output_4_2), .y(output_3_881));
wire output_5_881, output_5_2, output_4_881;
mixer gate_output_4_881(.a(output_5_881), .b(output_5_2), .y(output_4_881));
wire output_6_881, output_6_2, output_5_881;
mixer gate_output_5_881(.a(output_6_881), .b(output_6_2), .y(output_5_881));
wire output_7_881, output_7_2, output_6_881;
mixer gate_output_6_881(.a(output_7_881), .b(output_7_2), .y(output_6_881));
wire output_8_881, output_8_2, output_7_881;
mixer gate_output_7_881(.a(output_8_881), .b(output_8_2), .y(output_7_881));
wire output_9_881, output_9_2, output_8_881;
mixer gate_output_8_881(.a(output_9_881), .b(output_9_2), .y(output_8_881));
wire output_10_881, output_10_2, output_9_881;
mixer gate_output_9_881(.a(output_10_881), .b(output_10_2), .y(output_9_881));
wire output_11_881, output_11_2, output_10_881;
mixer gate_output_10_881(.a(output_11_881), .b(output_11_2), .y(output_10_881));
wire output_12_881, output_12_2, output_11_881;
mixer gate_output_11_881(.a(output_12_881), .b(output_12_2), .y(output_11_881));
wire output_13_881, output_13_2, output_12_881;
mixer gate_output_12_881(.a(output_13_881), .b(output_13_2), .y(output_12_881));
wire output_14_881, output_14_2, output_13_881;
mixer gate_output_13_881(.a(output_14_881), .b(output_14_2), .y(output_13_881));
wire output_15_881, output_15_2, output_14_881;
mixer gate_output_14_881(.a(output_15_881), .b(output_15_2), .y(output_14_881));
wire output_16_881, output_16_2, output_15_881;
mixer gate_output_15_881(.a(output_16_881), .b(output_16_2), .y(output_15_881));
wire output_1_882, output_1_3, output_0_882;
mixer gate_output_0_882(.a(output_1_882), .b(output_1_3), .y(output_0_882));
wire output_2_882, output_2_3, output_1_882;
mixer gate_output_1_882(.a(output_2_882), .b(output_2_3), .y(output_1_882));
wire output_3_882, output_3_3, output_2_882;
mixer gate_output_2_882(.a(output_3_882), .b(output_3_3), .y(output_2_882));
wire output_4_882, output_4_3, output_3_882;
mixer gate_output_3_882(.a(output_4_882), .b(output_4_3), .y(output_3_882));
wire output_5_882, output_5_3, output_4_882;
mixer gate_output_4_882(.a(output_5_882), .b(output_5_3), .y(output_4_882));
wire output_6_882, output_6_3, output_5_882;
mixer gate_output_5_882(.a(output_6_882), .b(output_6_3), .y(output_5_882));
wire output_7_882, output_7_3, output_6_882;
mixer gate_output_6_882(.a(output_7_882), .b(output_7_3), .y(output_6_882));
wire output_8_882, output_8_3, output_7_882;
mixer gate_output_7_882(.a(output_8_882), .b(output_8_3), .y(output_7_882));
wire output_9_882, output_9_3, output_8_882;
mixer gate_output_8_882(.a(output_9_882), .b(output_9_3), .y(output_8_882));
wire output_10_882, output_10_3, output_9_882;
mixer gate_output_9_882(.a(output_10_882), .b(output_10_3), .y(output_9_882));
wire output_11_882, output_11_3, output_10_882;
mixer gate_output_10_882(.a(output_11_882), .b(output_11_3), .y(output_10_882));
wire output_12_882, output_12_3, output_11_882;
mixer gate_output_11_882(.a(output_12_882), .b(output_12_3), .y(output_11_882));
wire output_13_882, output_13_3, output_12_882;
mixer gate_output_12_882(.a(output_13_882), .b(output_13_3), .y(output_12_882));
wire output_14_882, output_14_3, output_13_882;
mixer gate_output_13_882(.a(output_14_882), .b(output_14_3), .y(output_13_882));
wire output_15_882, output_15_3, output_14_882;
mixer gate_output_14_882(.a(output_15_882), .b(output_15_3), .y(output_14_882));
wire output_16_882, output_16_3, output_15_882;
mixer gate_output_15_882(.a(output_16_882), .b(output_16_3), .y(output_15_882));
wire output_1_883, output_1_4, output_0_883;
mixer gate_output_0_883(.a(output_1_883), .b(output_1_4), .y(output_0_883));
wire output_2_883, output_2_4, output_1_883;
mixer gate_output_1_883(.a(output_2_883), .b(output_2_4), .y(output_1_883));
wire output_3_883, output_3_4, output_2_883;
mixer gate_output_2_883(.a(output_3_883), .b(output_3_4), .y(output_2_883));
wire output_4_883, output_4_4, output_3_883;
mixer gate_output_3_883(.a(output_4_883), .b(output_4_4), .y(output_3_883));
wire output_5_883, output_5_4, output_4_883;
mixer gate_output_4_883(.a(output_5_883), .b(output_5_4), .y(output_4_883));
wire output_6_883, output_6_4, output_5_883;
mixer gate_output_5_883(.a(output_6_883), .b(output_6_4), .y(output_5_883));
wire output_7_883, output_7_4, output_6_883;
mixer gate_output_6_883(.a(output_7_883), .b(output_7_4), .y(output_6_883));
wire output_8_883, output_8_4, output_7_883;
mixer gate_output_7_883(.a(output_8_883), .b(output_8_4), .y(output_7_883));
wire output_9_883, output_9_4, output_8_883;
mixer gate_output_8_883(.a(output_9_883), .b(output_9_4), .y(output_8_883));
wire output_10_883, output_10_4, output_9_883;
mixer gate_output_9_883(.a(output_10_883), .b(output_10_4), .y(output_9_883));
wire output_11_883, output_11_4, output_10_883;
mixer gate_output_10_883(.a(output_11_883), .b(output_11_4), .y(output_10_883));
wire output_12_883, output_12_4, output_11_883;
mixer gate_output_11_883(.a(output_12_883), .b(output_12_4), .y(output_11_883));
wire output_13_883, output_13_4, output_12_883;
mixer gate_output_12_883(.a(output_13_883), .b(output_13_4), .y(output_12_883));
wire output_14_883, output_14_4, output_13_883;
mixer gate_output_13_883(.a(output_14_883), .b(output_14_4), .y(output_13_883));
wire output_15_883, output_15_4, output_14_883;
mixer gate_output_14_883(.a(output_15_883), .b(output_15_4), .y(output_14_883));
wire output_16_883, output_16_4, output_15_883;
mixer gate_output_15_883(.a(output_16_883), .b(output_16_4), .y(output_15_883));
wire output_1_884, output_1_5, output_0_884;
mixer gate_output_0_884(.a(output_1_884), .b(output_1_5), .y(output_0_884));
wire output_2_884, output_2_5, output_1_884;
mixer gate_output_1_884(.a(output_2_884), .b(output_2_5), .y(output_1_884));
wire output_3_884, output_3_5, output_2_884;
mixer gate_output_2_884(.a(output_3_884), .b(output_3_5), .y(output_2_884));
wire output_4_884, output_4_5, output_3_884;
mixer gate_output_3_884(.a(output_4_884), .b(output_4_5), .y(output_3_884));
wire output_5_884, output_5_5, output_4_884;
mixer gate_output_4_884(.a(output_5_884), .b(output_5_5), .y(output_4_884));
wire output_6_884, output_6_5, output_5_884;
mixer gate_output_5_884(.a(output_6_884), .b(output_6_5), .y(output_5_884));
wire output_7_884, output_7_5, output_6_884;
mixer gate_output_6_884(.a(output_7_884), .b(output_7_5), .y(output_6_884));
wire output_8_884, output_8_5, output_7_884;
mixer gate_output_7_884(.a(output_8_884), .b(output_8_5), .y(output_7_884));
wire output_9_884, output_9_5, output_8_884;
mixer gate_output_8_884(.a(output_9_884), .b(output_9_5), .y(output_8_884));
wire output_10_884, output_10_5, output_9_884;
mixer gate_output_9_884(.a(output_10_884), .b(output_10_5), .y(output_9_884));
wire output_11_884, output_11_5, output_10_884;
mixer gate_output_10_884(.a(output_11_884), .b(output_11_5), .y(output_10_884));
wire output_12_884, output_12_5, output_11_884;
mixer gate_output_11_884(.a(output_12_884), .b(output_12_5), .y(output_11_884));
wire output_13_884, output_13_5, output_12_884;
mixer gate_output_12_884(.a(output_13_884), .b(output_13_5), .y(output_12_884));
wire output_14_884, output_14_5, output_13_884;
mixer gate_output_13_884(.a(output_14_884), .b(output_14_5), .y(output_13_884));
wire output_15_884, output_15_5, output_14_884;
mixer gate_output_14_884(.a(output_15_884), .b(output_15_5), .y(output_14_884));
wire output_16_884, output_16_5, output_15_884;
mixer gate_output_15_884(.a(output_16_884), .b(output_16_5), .y(output_15_884));
wire output_1_885, output_1_6, output_0_885;
mixer gate_output_0_885(.a(output_1_885), .b(output_1_6), .y(output_0_885));
wire output_2_885, output_2_6, output_1_885;
mixer gate_output_1_885(.a(output_2_885), .b(output_2_6), .y(output_1_885));
wire output_3_885, output_3_6, output_2_885;
mixer gate_output_2_885(.a(output_3_885), .b(output_3_6), .y(output_2_885));
wire output_4_885, output_4_6, output_3_885;
mixer gate_output_3_885(.a(output_4_885), .b(output_4_6), .y(output_3_885));
wire output_5_885, output_5_6, output_4_885;
mixer gate_output_4_885(.a(output_5_885), .b(output_5_6), .y(output_4_885));
wire output_6_885, output_6_6, output_5_885;
mixer gate_output_5_885(.a(output_6_885), .b(output_6_6), .y(output_5_885));
wire output_7_885, output_7_6, output_6_885;
mixer gate_output_6_885(.a(output_7_885), .b(output_7_6), .y(output_6_885));
wire output_8_885, output_8_6, output_7_885;
mixer gate_output_7_885(.a(output_8_885), .b(output_8_6), .y(output_7_885));
wire output_9_885, output_9_6, output_8_885;
mixer gate_output_8_885(.a(output_9_885), .b(output_9_6), .y(output_8_885));
wire output_10_885, output_10_6, output_9_885;
mixer gate_output_9_885(.a(output_10_885), .b(output_10_6), .y(output_9_885));
wire output_11_885, output_11_6, output_10_885;
mixer gate_output_10_885(.a(output_11_885), .b(output_11_6), .y(output_10_885));
wire output_12_885, output_12_6, output_11_885;
mixer gate_output_11_885(.a(output_12_885), .b(output_12_6), .y(output_11_885));
wire output_13_885, output_13_6, output_12_885;
mixer gate_output_12_885(.a(output_13_885), .b(output_13_6), .y(output_12_885));
wire output_14_885, output_14_6, output_13_885;
mixer gate_output_13_885(.a(output_14_885), .b(output_14_6), .y(output_13_885));
wire output_15_885, output_15_6, output_14_885;
mixer gate_output_14_885(.a(output_15_885), .b(output_15_6), .y(output_14_885));
wire output_16_885, output_16_6, output_15_885;
mixer gate_output_15_885(.a(output_16_885), .b(output_16_6), .y(output_15_885));
wire output_1_886, output_1_7, output_0_886;
mixer gate_output_0_886(.a(output_1_886), .b(output_1_7), .y(output_0_886));
wire output_2_886, output_2_7, output_1_886;
mixer gate_output_1_886(.a(output_2_886), .b(output_2_7), .y(output_1_886));
wire output_3_886, output_3_7, output_2_886;
mixer gate_output_2_886(.a(output_3_886), .b(output_3_7), .y(output_2_886));
wire output_4_886, output_4_7, output_3_886;
mixer gate_output_3_886(.a(output_4_886), .b(output_4_7), .y(output_3_886));
wire output_5_886, output_5_7, output_4_886;
mixer gate_output_4_886(.a(output_5_886), .b(output_5_7), .y(output_4_886));
wire output_6_886, output_6_7, output_5_886;
mixer gate_output_5_886(.a(output_6_886), .b(output_6_7), .y(output_5_886));
wire output_7_886, output_7_7, output_6_886;
mixer gate_output_6_886(.a(output_7_886), .b(output_7_7), .y(output_6_886));
wire output_8_886, output_8_7, output_7_886;
mixer gate_output_7_886(.a(output_8_886), .b(output_8_7), .y(output_7_886));
wire output_9_886, output_9_7, output_8_886;
mixer gate_output_8_886(.a(output_9_886), .b(output_9_7), .y(output_8_886));
wire output_10_886, output_10_7, output_9_886;
mixer gate_output_9_886(.a(output_10_886), .b(output_10_7), .y(output_9_886));
wire output_11_886, output_11_7, output_10_886;
mixer gate_output_10_886(.a(output_11_886), .b(output_11_7), .y(output_10_886));
wire output_12_886, output_12_7, output_11_886;
mixer gate_output_11_886(.a(output_12_886), .b(output_12_7), .y(output_11_886));
wire output_13_886, output_13_7, output_12_886;
mixer gate_output_12_886(.a(output_13_886), .b(output_13_7), .y(output_12_886));
wire output_14_886, output_14_7, output_13_886;
mixer gate_output_13_886(.a(output_14_886), .b(output_14_7), .y(output_13_886));
wire output_15_886, output_15_7, output_14_886;
mixer gate_output_14_886(.a(output_15_886), .b(output_15_7), .y(output_14_886));
wire output_16_886, output_16_7, output_15_886;
mixer gate_output_15_886(.a(output_16_886), .b(output_16_7), .y(output_15_886));
wire output_1_887, output_1_8, output_0_887;
mixer gate_output_0_887(.a(output_1_887), .b(output_1_8), .y(output_0_887));
wire output_2_887, output_2_8, output_1_887;
mixer gate_output_1_887(.a(output_2_887), .b(output_2_8), .y(output_1_887));
wire output_3_887, output_3_8, output_2_887;
mixer gate_output_2_887(.a(output_3_887), .b(output_3_8), .y(output_2_887));
wire output_4_887, output_4_8, output_3_887;
mixer gate_output_3_887(.a(output_4_887), .b(output_4_8), .y(output_3_887));
wire output_5_887, output_5_8, output_4_887;
mixer gate_output_4_887(.a(output_5_887), .b(output_5_8), .y(output_4_887));
wire output_6_887, output_6_8, output_5_887;
mixer gate_output_5_887(.a(output_6_887), .b(output_6_8), .y(output_5_887));
wire output_7_887, output_7_8, output_6_887;
mixer gate_output_6_887(.a(output_7_887), .b(output_7_8), .y(output_6_887));
wire output_8_887, output_8_8, output_7_887;
mixer gate_output_7_887(.a(output_8_887), .b(output_8_8), .y(output_7_887));
wire output_9_887, output_9_8, output_8_887;
mixer gate_output_8_887(.a(output_9_887), .b(output_9_8), .y(output_8_887));
wire output_10_887, output_10_8, output_9_887;
mixer gate_output_9_887(.a(output_10_887), .b(output_10_8), .y(output_9_887));
wire output_11_887, output_11_8, output_10_887;
mixer gate_output_10_887(.a(output_11_887), .b(output_11_8), .y(output_10_887));
wire output_12_887, output_12_8, output_11_887;
mixer gate_output_11_887(.a(output_12_887), .b(output_12_8), .y(output_11_887));
wire output_13_887, output_13_8, output_12_887;
mixer gate_output_12_887(.a(output_13_887), .b(output_13_8), .y(output_12_887));
wire output_14_887, output_14_8, output_13_887;
mixer gate_output_13_887(.a(output_14_887), .b(output_14_8), .y(output_13_887));
wire output_15_887, output_15_8, output_14_887;
mixer gate_output_14_887(.a(output_15_887), .b(output_15_8), .y(output_14_887));
wire output_16_887, output_16_8, output_15_887;
mixer gate_output_15_887(.a(output_16_887), .b(output_16_8), .y(output_15_887));
wire output_1_888, output_1_9, output_0_888;
mixer gate_output_0_888(.a(output_1_888), .b(output_1_9), .y(output_0_888));
wire output_2_888, output_2_9, output_1_888;
mixer gate_output_1_888(.a(output_2_888), .b(output_2_9), .y(output_1_888));
wire output_3_888, output_3_9, output_2_888;
mixer gate_output_2_888(.a(output_3_888), .b(output_3_9), .y(output_2_888));
wire output_4_888, output_4_9, output_3_888;
mixer gate_output_3_888(.a(output_4_888), .b(output_4_9), .y(output_3_888));
wire output_5_888, output_5_9, output_4_888;
mixer gate_output_4_888(.a(output_5_888), .b(output_5_9), .y(output_4_888));
wire output_6_888, output_6_9, output_5_888;
mixer gate_output_5_888(.a(output_6_888), .b(output_6_9), .y(output_5_888));
wire output_7_888, output_7_9, output_6_888;
mixer gate_output_6_888(.a(output_7_888), .b(output_7_9), .y(output_6_888));
wire output_8_888, output_8_9, output_7_888;
mixer gate_output_7_888(.a(output_8_888), .b(output_8_9), .y(output_7_888));
wire output_9_888, output_9_9, output_8_888;
mixer gate_output_8_888(.a(output_9_888), .b(output_9_9), .y(output_8_888));
wire output_10_888, output_10_9, output_9_888;
mixer gate_output_9_888(.a(output_10_888), .b(output_10_9), .y(output_9_888));
wire output_11_888, output_11_9, output_10_888;
mixer gate_output_10_888(.a(output_11_888), .b(output_11_9), .y(output_10_888));
wire output_12_888, output_12_9, output_11_888;
mixer gate_output_11_888(.a(output_12_888), .b(output_12_9), .y(output_11_888));
wire output_13_888, output_13_9, output_12_888;
mixer gate_output_12_888(.a(output_13_888), .b(output_13_9), .y(output_12_888));
wire output_14_888, output_14_9, output_13_888;
mixer gate_output_13_888(.a(output_14_888), .b(output_14_9), .y(output_13_888));
wire output_15_888, output_15_9, output_14_888;
mixer gate_output_14_888(.a(output_15_888), .b(output_15_9), .y(output_14_888));
wire output_16_888, output_16_9, output_15_888;
mixer gate_output_15_888(.a(output_16_888), .b(output_16_9), .y(output_15_888));
wire output_1_889, output_1_10, output_0_889;
mixer gate_output_0_889(.a(output_1_889), .b(output_1_10), .y(output_0_889));
wire output_2_889, output_2_10, output_1_889;
mixer gate_output_1_889(.a(output_2_889), .b(output_2_10), .y(output_1_889));
wire output_3_889, output_3_10, output_2_889;
mixer gate_output_2_889(.a(output_3_889), .b(output_3_10), .y(output_2_889));
wire output_4_889, output_4_10, output_3_889;
mixer gate_output_3_889(.a(output_4_889), .b(output_4_10), .y(output_3_889));
wire output_5_889, output_5_10, output_4_889;
mixer gate_output_4_889(.a(output_5_889), .b(output_5_10), .y(output_4_889));
wire output_6_889, output_6_10, output_5_889;
mixer gate_output_5_889(.a(output_6_889), .b(output_6_10), .y(output_5_889));
wire output_7_889, output_7_10, output_6_889;
mixer gate_output_6_889(.a(output_7_889), .b(output_7_10), .y(output_6_889));
wire output_8_889, output_8_10, output_7_889;
mixer gate_output_7_889(.a(output_8_889), .b(output_8_10), .y(output_7_889));
wire output_9_889, output_9_10, output_8_889;
mixer gate_output_8_889(.a(output_9_889), .b(output_9_10), .y(output_8_889));
wire output_10_889, output_10_10, output_9_889;
mixer gate_output_9_889(.a(output_10_889), .b(output_10_10), .y(output_9_889));
wire output_11_889, output_11_10, output_10_889;
mixer gate_output_10_889(.a(output_11_889), .b(output_11_10), .y(output_10_889));
wire output_12_889, output_12_10, output_11_889;
mixer gate_output_11_889(.a(output_12_889), .b(output_12_10), .y(output_11_889));
wire output_13_889, output_13_10, output_12_889;
mixer gate_output_12_889(.a(output_13_889), .b(output_13_10), .y(output_12_889));
wire output_14_889, output_14_10, output_13_889;
mixer gate_output_13_889(.a(output_14_889), .b(output_14_10), .y(output_13_889));
wire output_15_889, output_15_10, output_14_889;
mixer gate_output_14_889(.a(output_15_889), .b(output_15_10), .y(output_14_889));
wire output_16_889, output_16_10, output_15_889;
mixer gate_output_15_889(.a(output_16_889), .b(output_16_10), .y(output_15_889));
wire output_1_890, output_1_11, output_0_890;
mixer gate_output_0_890(.a(output_1_890), .b(output_1_11), .y(output_0_890));
wire output_2_890, output_2_11, output_1_890;
mixer gate_output_1_890(.a(output_2_890), .b(output_2_11), .y(output_1_890));
wire output_3_890, output_3_11, output_2_890;
mixer gate_output_2_890(.a(output_3_890), .b(output_3_11), .y(output_2_890));
wire output_4_890, output_4_11, output_3_890;
mixer gate_output_3_890(.a(output_4_890), .b(output_4_11), .y(output_3_890));
wire output_5_890, output_5_11, output_4_890;
mixer gate_output_4_890(.a(output_5_890), .b(output_5_11), .y(output_4_890));
wire output_6_890, output_6_11, output_5_890;
mixer gate_output_5_890(.a(output_6_890), .b(output_6_11), .y(output_5_890));
wire output_7_890, output_7_11, output_6_890;
mixer gate_output_6_890(.a(output_7_890), .b(output_7_11), .y(output_6_890));
wire output_8_890, output_8_11, output_7_890;
mixer gate_output_7_890(.a(output_8_890), .b(output_8_11), .y(output_7_890));
wire output_9_890, output_9_11, output_8_890;
mixer gate_output_8_890(.a(output_9_890), .b(output_9_11), .y(output_8_890));
wire output_10_890, output_10_11, output_9_890;
mixer gate_output_9_890(.a(output_10_890), .b(output_10_11), .y(output_9_890));
wire output_11_890, output_11_11, output_10_890;
mixer gate_output_10_890(.a(output_11_890), .b(output_11_11), .y(output_10_890));
wire output_12_890, output_12_11, output_11_890;
mixer gate_output_11_890(.a(output_12_890), .b(output_12_11), .y(output_11_890));
wire output_13_890, output_13_11, output_12_890;
mixer gate_output_12_890(.a(output_13_890), .b(output_13_11), .y(output_12_890));
wire output_14_890, output_14_11, output_13_890;
mixer gate_output_13_890(.a(output_14_890), .b(output_14_11), .y(output_13_890));
wire output_15_890, output_15_11, output_14_890;
mixer gate_output_14_890(.a(output_15_890), .b(output_15_11), .y(output_14_890));
wire output_16_890, output_16_11, output_15_890;
mixer gate_output_15_890(.a(output_16_890), .b(output_16_11), .y(output_15_890));
wire output_1_891, output_1_12, output_0_891;
mixer gate_output_0_891(.a(output_1_891), .b(output_1_12), .y(output_0_891));
wire output_2_891, output_2_12, output_1_891;
mixer gate_output_1_891(.a(output_2_891), .b(output_2_12), .y(output_1_891));
wire output_3_891, output_3_12, output_2_891;
mixer gate_output_2_891(.a(output_3_891), .b(output_3_12), .y(output_2_891));
wire output_4_891, output_4_12, output_3_891;
mixer gate_output_3_891(.a(output_4_891), .b(output_4_12), .y(output_3_891));
wire output_5_891, output_5_12, output_4_891;
mixer gate_output_4_891(.a(output_5_891), .b(output_5_12), .y(output_4_891));
wire output_6_891, output_6_12, output_5_891;
mixer gate_output_5_891(.a(output_6_891), .b(output_6_12), .y(output_5_891));
wire output_7_891, output_7_12, output_6_891;
mixer gate_output_6_891(.a(output_7_891), .b(output_7_12), .y(output_6_891));
wire output_8_891, output_8_12, output_7_891;
mixer gate_output_7_891(.a(output_8_891), .b(output_8_12), .y(output_7_891));
wire output_9_891, output_9_12, output_8_891;
mixer gate_output_8_891(.a(output_9_891), .b(output_9_12), .y(output_8_891));
wire output_10_891, output_10_12, output_9_891;
mixer gate_output_9_891(.a(output_10_891), .b(output_10_12), .y(output_9_891));
wire output_11_891, output_11_12, output_10_891;
mixer gate_output_10_891(.a(output_11_891), .b(output_11_12), .y(output_10_891));
wire output_12_891, output_12_12, output_11_891;
mixer gate_output_11_891(.a(output_12_891), .b(output_12_12), .y(output_11_891));
wire output_13_891, output_13_12, output_12_891;
mixer gate_output_12_891(.a(output_13_891), .b(output_13_12), .y(output_12_891));
wire output_14_891, output_14_12, output_13_891;
mixer gate_output_13_891(.a(output_14_891), .b(output_14_12), .y(output_13_891));
wire output_15_891, output_15_12, output_14_891;
mixer gate_output_14_891(.a(output_15_891), .b(output_15_12), .y(output_14_891));
wire output_16_891, output_16_12, output_15_891;
mixer gate_output_15_891(.a(output_16_891), .b(output_16_12), .y(output_15_891));
wire output_1_892, output_1_13, output_0_892;
mixer gate_output_0_892(.a(output_1_892), .b(output_1_13), .y(output_0_892));
wire output_2_892, output_2_13, output_1_892;
mixer gate_output_1_892(.a(output_2_892), .b(output_2_13), .y(output_1_892));
wire output_3_892, output_3_13, output_2_892;
mixer gate_output_2_892(.a(output_3_892), .b(output_3_13), .y(output_2_892));
wire output_4_892, output_4_13, output_3_892;
mixer gate_output_3_892(.a(output_4_892), .b(output_4_13), .y(output_3_892));
wire output_5_892, output_5_13, output_4_892;
mixer gate_output_4_892(.a(output_5_892), .b(output_5_13), .y(output_4_892));
wire output_6_892, output_6_13, output_5_892;
mixer gate_output_5_892(.a(output_6_892), .b(output_6_13), .y(output_5_892));
wire output_7_892, output_7_13, output_6_892;
mixer gate_output_6_892(.a(output_7_892), .b(output_7_13), .y(output_6_892));
wire output_8_892, output_8_13, output_7_892;
mixer gate_output_7_892(.a(output_8_892), .b(output_8_13), .y(output_7_892));
wire output_9_892, output_9_13, output_8_892;
mixer gate_output_8_892(.a(output_9_892), .b(output_9_13), .y(output_8_892));
wire output_10_892, output_10_13, output_9_892;
mixer gate_output_9_892(.a(output_10_892), .b(output_10_13), .y(output_9_892));
wire output_11_892, output_11_13, output_10_892;
mixer gate_output_10_892(.a(output_11_892), .b(output_11_13), .y(output_10_892));
wire output_12_892, output_12_13, output_11_892;
mixer gate_output_11_892(.a(output_12_892), .b(output_12_13), .y(output_11_892));
wire output_13_892, output_13_13, output_12_892;
mixer gate_output_12_892(.a(output_13_892), .b(output_13_13), .y(output_12_892));
wire output_14_892, output_14_13, output_13_892;
mixer gate_output_13_892(.a(output_14_892), .b(output_14_13), .y(output_13_892));
wire output_15_892, output_15_13, output_14_892;
mixer gate_output_14_892(.a(output_15_892), .b(output_15_13), .y(output_14_892));
wire output_16_892, output_16_13, output_15_892;
mixer gate_output_15_892(.a(output_16_892), .b(output_16_13), .y(output_15_892));
wire output_1_893, output_1_14, output_0_893;
mixer gate_output_0_893(.a(output_1_893), .b(output_1_14), .y(output_0_893));
wire output_2_893, output_2_14, output_1_893;
mixer gate_output_1_893(.a(output_2_893), .b(output_2_14), .y(output_1_893));
wire output_3_893, output_3_14, output_2_893;
mixer gate_output_2_893(.a(output_3_893), .b(output_3_14), .y(output_2_893));
wire output_4_893, output_4_14, output_3_893;
mixer gate_output_3_893(.a(output_4_893), .b(output_4_14), .y(output_3_893));
wire output_5_893, output_5_14, output_4_893;
mixer gate_output_4_893(.a(output_5_893), .b(output_5_14), .y(output_4_893));
wire output_6_893, output_6_14, output_5_893;
mixer gate_output_5_893(.a(output_6_893), .b(output_6_14), .y(output_5_893));
wire output_7_893, output_7_14, output_6_893;
mixer gate_output_6_893(.a(output_7_893), .b(output_7_14), .y(output_6_893));
wire output_8_893, output_8_14, output_7_893;
mixer gate_output_7_893(.a(output_8_893), .b(output_8_14), .y(output_7_893));
wire output_9_893, output_9_14, output_8_893;
mixer gate_output_8_893(.a(output_9_893), .b(output_9_14), .y(output_8_893));
wire output_10_893, output_10_14, output_9_893;
mixer gate_output_9_893(.a(output_10_893), .b(output_10_14), .y(output_9_893));
wire output_11_893, output_11_14, output_10_893;
mixer gate_output_10_893(.a(output_11_893), .b(output_11_14), .y(output_10_893));
wire output_12_893, output_12_14, output_11_893;
mixer gate_output_11_893(.a(output_12_893), .b(output_12_14), .y(output_11_893));
wire output_13_893, output_13_14, output_12_893;
mixer gate_output_12_893(.a(output_13_893), .b(output_13_14), .y(output_12_893));
wire output_14_893, output_14_14, output_13_893;
mixer gate_output_13_893(.a(output_14_893), .b(output_14_14), .y(output_13_893));
wire output_15_893, output_15_14, output_14_893;
mixer gate_output_14_893(.a(output_15_893), .b(output_15_14), .y(output_14_893));
wire output_16_893, output_16_14, output_15_893;
mixer gate_output_15_893(.a(output_16_893), .b(output_16_14), .y(output_15_893));
wire output_1_894, output_1_15, output_0_894;
mixer gate_output_0_894(.a(output_1_894), .b(output_1_15), .y(output_0_894));
wire output_2_894, output_2_15, output_1_894;
mixer gate_output_1_894(.a(output_2_894), .b(output_2_15), .y(output_1_894));
wire output_3_894, output_3_15, output_2_894;
mixer gate_output_2_894(.a(output_3_894), .b(output_3_15), .y(output_2_894));
wire output_4_894, output_4_15, output_3_894;
mixer gate_output_3_894(.a(output_4_894), .b(output_4_15), .y(output_3_894));
wire output_5_894, output_5_15, output_4_894;
mixer gate_output_4_894(.a(output_5_894), .b(output_5_15), .y(output_4_894));
wire output_6_894, output_6_15, output_5_894;
mixer gate_output_5_894(.a(output_6_894), .b(output_6_15), .y(output_5_894));
wire output_7_894, output_7_15, output_6_894;
mixer gate_output_6_894(.a(output_7_894), .b(output_7_15), .y(output_6_894));
wire output_8_894, output_8_15, output_7_894;
mixer gate_output_7_894(.a(output_8_894), .b(output_8_15), .y(output_7_894));
wire output_9_894, output_9_15, output_8_894;
mixer gate_output_8_894(.a(output_9_894), .b(output_9_15), .y(output_8_894));
wire output_10_894, output_10_15, output_9_894;
mixer gate_output_9_894(.a(output_10_894), .b(output_10_15), .y(output_9_894));
wire output_11_894, output_11_15, output_10_894;
mixer gate_output_10_894(.a(output_11_894), .b(output_11_15), .y(output_10_894));
wire output_12_894, output_12_15, output_11_894;
mixer gate_output_11_894(.a(output_12_894), .b(output_12_15), .y(output_11_894));
wire output_13_894, output_13_15, output_12_894;
mixer gate_output_12_894(.a(output_13_894), .b(output_13_15), .y(output_12_894));
wire output_14_894, output_14_15, output_13_894;
mixer gate_output_13_894(.a(output_14_894), .b(output_14_15), .y(output_13_894));
wire output_15_894, output_15_15, output_14_894;
mixer gate_output_14_894(.a(output_15_894), .b(output_15_15), .y(output_14_894));
wire output_16_894, output_16_15, output_15_894;
mixer gate_output_15_894(.a(output_16_894), .b(output_16_15), .y(output_15_894));
wire output_1_895, output_1_0, output_0_895;
mixer gate_output_0_895(.a(output_1_895), .b(output_1_0), .y(output_0_895));
wire output_2_895, output_2_0, output_1_895;
mixer gate_output_1_895(.a(output_2_895), .b(output_2_0), .y(output_1_895));
wire output_3_895, output_3_0, output_2_895;
mixer gate_output_2_895(.a(output_3_895), .b(output_3_0), .y(output_2_895));
wire output_4_895, output_4_0, output_3_895;
mixer gate_output_3_895(.a(output_4_895), .b(output_4_0), .y(output_3_895));
wire output_5_895, output_5_0, output_4_895;
mixer gate_output_4_895(.a(output_5_895), .b(output_5_0), .y(output_4_895));
wire output_6_895, output_6_0, output_5_895;
mixer gate_output_5_895(.a(output_6_895), .b(output_6_0), .y(output_5_895));
wire output_7_895, output_7_0, output_6_895;
mixer gate_output_6_895(.a(output_7_895), .b(output_7_0), .y(output_6_895));
wire output_8_895, output_8_0, output_7_895;
mixer gate_output_7_895(.a(output_8_895), .b(output_8_0), .y(output_7_895));
wire output_9_895, output_9_0, output_8_895;
mixer gate_output_8_895(.a(output_9_895), .b(output_9_0), .y(output_8_895));
wire output_10_895, output_10_0, output_9_895;
mixer gate_output_9_895(.a(output_10_895), .b(output_10_0), .y(output_9_895));
wire output_11_895, output_11_0, output_10_895;
mixer gate_output_10_895(.a(output_11_895), .b(output_11_0), .y(output_10_895));
wire output_12_895, output_12_0, output_11_895;
mixer gate_output_11_895(.a(output_12_895), .b(output_12_0), .y(output_11_895));
wire output_13_895, output_13_0, output_12_895;
mixer gate_output_12_895(.a(output_13_895), .b(output_13_0), .y(output_12_895));
wire output_14_895, output_14_0, output_13_895;
mixer gate_output_13_895(.a(output_14_895), .b(output_14_0), .y(output_13_895));
wire output_15_895, output_15_0, output_14_895;
mixer gate_output_14_895(.a(output_15_895), .b(output_15_0), .y(output_14_895));
wire output_16_895, output_16_0, output_15_895;
mixer gate_output_15_895(.a(output_16_895), .b(output_16_0), .y(output_15_895));
wire output_1_896, output_1_1, output_0_896;
mixer gate_output_0_896(.a(output_1_896), .b(output_1_1), .y(output_0_896));
wire output_2_896, output_2_1, output_1_896;
mixer gate_output_1_896(.a(output_2_896), .b(output_2_1), .y(output_1_896));
wire output_3_896, output_3_1, output_2_896;
mixer gate_output_2_896(.a(output_3_896), .b(output_3_1), .y(output_2_896));
wire output_4_896, output_4_1, output_3_896;
mixer gate_output_3_896(.a(output_4_896), .b(output_4_1), .y(output_3_896));
wire output_5_896, output_5_1, output_4_896;
mixer gate_output_4_896(.a(output_5_896), .b(output_5_1), .y(output_4_896));
wire output_6_896, output_6_1, output_5_896;
mixer gate_output_5_896(.a(output_6_896), .b(output_6_1), .y(output_5_896));
wire output_7_896, output_7_1, output_6_896;
mixer gate_output_6_896(.a(output_7_896), .b(output_7_1), .y(output_6_896));
wire output_8_896, output_8_1, output_7_896;
mixer gate_output_7_896(.a(output_8_896), .b(output_8_1), .y(output_7_896));
wire output_9_896, output_9_1, output_8_896;
mixer gate_output_8_896(.a(output_9_896), .b(output_9_1), .y(output_8_896));
wire output_10_896, output_10_1, output_9_896;
mixer gate_output_9_896(.a(output_10_896), .b(output_10_1), .y(output_9_896));
wire output_11_896, output_11_1, output_10_896;
mixer gate_output_10_896(.a(output_11_896), .b(output_11_1), .y(output_10_896));
wire output_12_896, output_12_1, output_11_896;
mixer gate_output_11_896(.a(output_12_896), .b(output_12_1), .y(output_11_896));
wire output_13_896, output_13_1, output_12_896;
mixer gate_output_12_896(.a(output_13_896), .b(output_13_1), .y(output_12_896));
wire output_14_896, output_14_1, output_13_896;
mixer gate_output_13_896(.a(output_14_896), .b(output_14_1), .y(output_13_896));
wire output_15_896, output_15_1, output_14_896;
mixer gate_output_14_896(.a(output_15_896), .b(output_15_1), .y(output_14_896));
wire output_16_896, output_16_1, output_15_896;
mixer gate_output_15_896(.a(output_16_896), .b(output_16_1), .y(output_15_896));
wire output_1_897, output_1_2, output_0_897;
mixer gate_output_0_897(.a(output_1_897), .b(output_1_2), .y(output_0_897));
wire output_2_897, output_2_2, output_1_897;
mixer gate_output_1_897(.a(output_2_897), .b(output_2_2), .y(output_1_897));
wire output_3_897, output_3_2, output_2_897;
mixer gate_output_2_897(.a(output_3_897), .b(output_3_2), .y(output_2_897));
wire output_4_897, output_4_2, output_3_897;
mixer gate_output_3_897(.a(output_4_897), .b(output_4_2), .y(output_3_897));
wire output_5_897, output_5_2, output_4_897;
mixer gate_output_4_897(.a(output_5_897), .b(output_5_2), .y(output_4_897));
wire output_6_897, output_6_2, output_5_897;
mixer gate_output_5_897(.a(output_6_897), .b(output_6_2), .y(output_5_897));
wire output_7_897, output_7_2, output_6_897;
mixer gate_output_6_897(.a(output_7_897), .b(output_7_2), .y(output_6_897));
wire output_8_897, output_8_2, output_7_897;
mixer gate_output_7_897(.a(output_8_897), .b(output_8_2), .y(output_7_897));
wire output_9_897, output_9_2, output_8_897;
mixer gate_output_8_897(.a(output_9_897), .b(output_9_2), .y(output_8_897));
wire output_10_897, output_10_2, output_9_897;
mixer gate_output_9_897(.a(output_10_897), .b(output_10_2), .y(output_9_897));
wire output_11_897, output_11_2, output_10_897;
mixer gate_output_10_897(.a(output_11_897), .b(output_11_2), .y(output_10_897));
wire output_12_897, output_12_2, output_11_897;
mixer gate_output_11_897(.a(output_12_897), .b(output_12_2), .y(output_11_897));
wire output_13_897, output_13_2, output_12_897;
mixer gate_output_12_897(.a(output_13_897), .b(output_13_2), .y(output_12_897));
wire output_14_897, output_14_2, output_13_897;
mixer gate_output_13_897(.a(output_14_897), .b(output_14_2), .y(output_13_897));
wire output_15_897, output_15_2, output_14_897;
mixer gate_output_14_897(.a(output_15_897), .b(output_15_2), .y(output_14_897));
wire output_16_897, output_16_2, output_15_897;
mixer gate_output_15_897(.a(output_16_897), .b(output_16_2), .y(output_15_897));
wire output_1_898, output_1_3, output_0_898;
mixer gate_output_0_898(.a(output_1_898), .b(output_1_3), .y(output_0_898));
wire output_2_898, output_2_3, output_1_898;
mixer gate_output_1_898(.a(output_2_898), .b(output_2_3), .y(output_1_898));
wire output_3_898, output_3_3, output_2_898;
mixer gate_output_2_898(.a(output_3_898), .b(output_3_3), .y(output_2_898));
wire output_4_898, output_4_3, output_3_898;
mixer gate_output_3_898(.a(output_4_898), .b(output_4_3), .y(output_3_898));
wire output_5_898, output_5_3, output_4_898;
mixer gate_output_4_898(.a(output_5_898), .b(output_5_3), .y(output_4_898));
wire output_6_898, output_6_3, output_5_898;
mixer gate_output_5_898(.a(output_6_898), .b(output_6_3), .y(output_5_898));
wire output_7_898, output_7_3, output_6_898;
mixer gate_output_6_898(.a(output_7_898), .b(output_7_3), .y(output_6_898));
wire output_8_898, output_8_3, output_7_898;
mixer gate_output_7_898(.a(output_8_898), .b(output_8_3), .y(output_7_898));
wire output_9_898, output_9_3, output_8_898;
mixer gate_output_8_898(.a(output_9_898), .b(output_9_3), .y(output_8_898));
wire output_10_898, output_10_3, output_9_898;
mixer gate_output_9_898(.a(output_10_898), .b(output_10_3), .y(output_9_898));
wire output_11_898, output_11_3, output_10_898;
mixer gate_output_10_898(.a(output_11_898), .b(output_11_3), .y(output_10_898));
wire output_12_898, output_12_3, output_11_898;
mixer gate_output_11_898(.a(output_12_898), .b(output_12_3), .y(output_11_898));
wire output_13_898, output_13_3, output_12_898;
mixer gate_output_12_898(.a(output_13_898), .b(output_13_3), .y(output_12_898));
wire output_14_898, output_14_3, output_13_898;
mixer gate_output_13_898(.a(output_14_898), .b(output_14_3), .y(output_13_898));
wire output_15_898, output_15_3, output_14_898;
mixer gate_output_14_898(.a(output_15_898), .b(output_15_3), .y(output_14_898));
wire output_16_898, output_16_3, output_15_898;
mixer gate_output_15_898(.a(output_16_898), .b(output_16_3), .y(output_15_898));
wire output_1_899, output_1_4, output_0_899;
mixer gate_output_0_899(.a(output_1_899), .b(output_1_4), .y(output_0_899));
wire output_2_899, output_2_4, output_1_899;
mixer gate_output_1_899(.a(output_2_899), .b(output_2_4), .y(output_1_899));
wire output_3_899, output_3_4, output_2_899;
mixer gate_output_2_899(.a(output_3_899), .b(output_3_4), .y(output_2_899));
wire output_4_899, output_4_4, output_3_899;
mixer gate_output_3_899(.a(output_4_899), .b(output_4_4), .y(output_3_899));
wire output_5_899, output_5_4, output_4_899;
mixer gate_output_4_899(.a(output_5_899), .b(output_5_4), .y(output_4_899));
wire output_6_899, output_6_4, output_5_899;
mixer gate_output_5_899(.a(output_6_899), .b(output_6_4), .y(output_5_899));
wire output_7_899, output_7_4, output_6_899;
mixer gate_output_6_899(.a(output_7_899), .b(output_7_4), .y(output_6_899));
wire output_8_899, output_8_4, output_7_899;
mixer gate_output_7_899(.a(output_8_899), .b(output_8_4), .y(output_7_899));
wire output_9_899, output_9_4, output_8_899;
mixer gate_output_8_899(.a(output_9_899), .b(output_9_4), .y(output_8_899));
wire output_10_899, output_10_4, output_9_899;
mixer gate_output_9_899(.a(output_10_899), .b(output_10_4), .y(output_9_899));
wire output_11_899, output_11_4, output_10_899;
mixer gate_output_10_899(.a(output_11_899), .b(output_11_4), .y(output_10_899));
wire output_12_899, output_12_4, output_11_899;
mixer gate_output_11_899(.a(output_12_899), .b(output_12_4), .y(output_11_899));
wire output_13_899, output_13_4, output_12_899;
mixer gate_output_12_899(.a(output_13_899), .b(output_13_4), .y(output_12_899));
wire output_14_899, output_14_4, output_13_899;
mixer gate_output_13_899(.a(output_14_899), .b(output_14_4), .y(output_13_899));
wire output_15_899, output_15_4, output_14_899;
mixer gate_output_14_899(.a(output_15_899), .b(output_15_4), .y(output_14_899));
wire output_16_899, output_16_4, output_15_899;
mixer gate_output_15_899(.a(output_16_899), .b(output_16_4), .y(output_15_899));
wire output_1_900, output_1_5, output_0_900;
mixer gate_output_0_900(.a(output_1_900), .b(output_1_5), .y(output_0_900));
wire output_2_900, output_2_5, output_1_900;
mixer gate_output_1_900(.a(output_2_900), .b(output_2_5), .y(output_1_900));
wire output_3_900, output_3_5, output_2_900;
mixer gate_output_2_900(.a(output_3_900), .b(output_3_5), .y(output_2_900));
wire output_4_900, output_4_5, output_3_900;
mixer gate_output_3_900(.a(output_4_900), .b(output_4_5), .y(output_3_900));
wire output_5_900, output_5_5, output_4_900;
mixer gate_output_4_900(.a(output_5_900), .b(output_5_5), .y(output_4_900));
wire output_6_900, output_6_5, output_5_900;
mixer gate_output_5_900(.a(output_6_900), .b(output_6_5), .y(output_5_900));
wire output_7_900, output_7_5, output_6_900;
mixer gate_output_6_900(.a(output_7_900), .b(output_7_5), .y(output_6_900));
wire output_8_900, output_8_5, output_7_900;
mixer gate_output_7_900(.a(output_8_900), .b(output_8_5), .y(output_7_900));
wire output_9_900, output_9_5, output_8_900;
mixer gate_output_8_900(.a(output_9_900), .b(output_9_5), .y(output_8_900));
wire output_10_900, output_10_5, output_9_900;
mixer gate_output_9_900(.a(output_10_900), .b(output_10_5), .y(output_9_900));
wire output_11_900, output_11_5, output_10_900;
mixer gate_output_10_900(.a(output_11_900), .b(output_11_5), .y(output_10_900));
wire output_12_900, output_12_5, output_11_900;
mixer gate_output_11_900(.a(output_12_900), .b(output_12_5), .y(output_11_900));
wire output_13_900, output_13_5, output_12_900;
mixer gate_output_12_900(.a(output_13_900), .b(output_13_5), .y(output_12_900));
wire output_14_900, output_14_5, output_13_900;
mixer gate_output_13_900(.a(output_14_900), .b(output_14_5), .y(output_13_900));
wire output_15_900, output_15_5, output_14_900;
mixer gate_output_14_900(.a(output_15_900), .b(output_15_5), .y(output_14_900));
wire output_16_900, output_16_5, output_15_900;
mixer gate_output_15_900(.a(output_16_900), .b(output_16_5), .y(output_15_900));
wire output_1_901, output_1_6, output_0_901;
mixer gate_output_0_901(.a(output_1_901), .b(output_1_6), .y(output_0_901));
wire output_2_901, output_2_6, output_1_901;
mixer gate_output_1_901(.a(output_2_901), .b(output_2_6), .y(output_1_901));
wire output_3_901, output_3_6, output_2_901;
mixer gate_output_2_901(.a(output_3_901), .b(output_3_6), .y(output_2_901));
wire output_4_901, output_4_6, output_3_901;
mixer gate_output_3_901(.a(output_4_901), .b(output_4_6), .y(output_3_901));
wire output_5_901, output_5_6, output_4_901;
mixer gate_output_4_901(.a(output_5_901), .b(output_5_6), .y(output_4_901));
wire output_6_901, output_6_6, output_5_901;
mixer gate_output_5_901(.a(output_6_901), .b(output_6_6), .y(output_5_901));
wire output_7_901, output_7_6, output_6_901;
mixer gate_output_6_901(.a(output_7_901), .b(output_7_6), .y(output_6_901));
wire output_8_901, output_8_6, output_7_901;
mixer gate_output_7_901(.a(output_8_901), .b(output_8_6), .y(output_7_901));
wire output_9_901, output_9_6, output_8_901;
mixer gate_output_8_901(.a(output_9_901), .b(output_9_6), .y(output_8_901));
wire output_10_901, output_10_6, output_9_901;
mixer gate_output_9_901(.a(output_10_901), .b(output_10_6), .y(output_9_901));
wire output_11_901, output_11_6, output_10_901;
mixer gate_output_10_901(.a(output_11_901), .b(output_11_6), .y(output_10_901));
wire output_12_901, output_12_6, output_11_901;
mixer gate_output_11_901(.a(output_12_901), .b(output_12_6), .y(output_11_901));
wire output_13_901, output_13_6, output_12_901;
mixer gate_output_12_901(.a(output_13_901), .b(output_13_6), .y(output_12_901));
wire output_14_901, output_14_6, output_13_901;
mixer gate_output_13_901(.a(output_14_901), .b(output_14_6), .y(output_13_901));
wire output_15_901, output_15_6, output_14_901;
mixer gate_output_14_901(.a(output_15_901), .b(output_15_6), .y(output_14_901));
wire output_16_901, output_16_6, output_15_901;
mixer gate_output_15_901(.a(output_16_901), .b(output_16_6), .y(output_15_901));
wire output_1_902, output_1_7, output_0_902;
mixer gate_output_0_902(.a(output_1_902), .b(output_1_7), .y(output_0_902));
wire output_2_902, output_2_7, output_1_902;
mixer gate_output_1_902(.a(output_2_902), .b(output_2_7), .y(output_1_902));
wire output_3_902, output_3_7, output_2_902;
mixer gate_output_2_902(.a(output_3_902), .b(output_3_7), .y(output_2_902));
wire output_4_902, output_4_7, output_3_902;
mixer gate_output_3_902(.a(output_4_902), .b(output_4_7), .y(output_3_902));
wire output_5_902, output_5_7, output_4_902;
mixer gate_output_4_902(.a(output_5_902), .b(output_5_7), .y(output_4_902));
wire output_6_902, output_6_7, output_5_902;
mixer gate_output_5_902(.a(output_6_902), .b(output_6_7), .y(output_5_902));
wire output_7_902, output_7_7, output_6_902;
mixer gate_output_6_902(.a(output_7_902), .b(output_7_7), .y(output_6_902));
wire output_8_902, output_8_7, output_7_902;
mixer gate_output_7_902(.a(output_8_902), .b(output_8_7), .y(output_7_902));
wire output_9_902, output_9_7, output_8_902;
mixer gate_output_8_902(.a(output_9_902), .b(output_9_7), .y(output_8_902));
wire output_10_902, output_10_7, output_9_902;
mixer gate_output_9_902(.a(output_10_902), .b(output_10_7), .y(output_9_902));
wire output_11_902, output_11_7, output_10_902;
mixer gate_output_10_902(.a(output_11_902), .b(output_11_7), .y(output_10_902));
wire output_12_902, output_12_7, output_11_902;
mixer gate_output_11_902(.a(output_12_902), .b(output_12_7), .y(output_11_902));
wire output_13_902, output_13_7, output_12_902;
mixer gate_output_12_902(.a(output_13_902), .b(output_13_7), .y(output_12_902));
wire output_14_902, output_14_7, output_13_902;
mixer gate_output_13_902(.a(output_14_902), .b(output_14_7), .y(output_13_902));
wire output_15_902, output_15_7, output_14_902;
mixer gate_output_14_902(.a(output_15_902), .b(output_15_7), .y(output_14_902));
wire output_16_902, output_16_7, output_15_902;
mixer gate_output_15_902(.a(output_16_902), .b(output_16_7), .y(output_15_902));
wire output_1_903, output_1_8, output_0_903;
mixer gate_output_0_903(.a(output_1_903), .b(output_1_8), .y(output_0_903));
wire output_2_903, output_2_8, output_1_903;
mixer gate_output_1_903(.a(output_2_903), .b(output_2_8), .y(output_1_903));
wire output_3_903, output_3_8, output_2_903;
mixer gate_output_2_903(.a(output_3_903), .b(output_3_8), .y(output_2_903));
wire output_4_903, output_4_8, output_3_903;
mixer gate_output_3_903(.a(output_4_903), .b(output_4_8), .y(output_3_903));
wire output_5_903, output_5_8, output_4_903;
mixer gate_output_4_903(.a(output_5_903), .b(output_5_8), .y(output_4_903));
wire output_6_903, output_6_8, output_5_903;
mixer gate_output_5_903(.a(output_6_903), .b(output_6_8), .y(output_5_903));
wire output_7_903, output_7_8, output_6_903;
mixer gate_output_6_903(.a(output_7_903), .b(output_7_8), .y(output_6_903));
wire output_8_903, output_8_8, output_7_903;
mixer gate_output_7_903(.a(output_8_903), .b(output_8_8), .y(output_7_903));
wire output_9_903, output_9_8, output_8_903;
mixer gate_output_8_903(.a(output_9_903), .b(output_9_8), .y(output_8_903));
wire output_10_903, output_10_8, output_9_903;
mixer gate_output_9_903(.a(output_10_903), .b(output_10_8), .y(output_9_903));
wire output_11_903, output_11_8, output_10_903;
mixer gate_output_10_903(.a(output_11_903), .b(output_11_8), .y(output_10_903));
wire output_12_903, output_12_8, output_11_903;
mixer gate_output_11_903(.a(output_12_903), .b(output_12_8), .y(output_11_903));
wire output_13_903, output_13_8, output_12_903;
mixer gate_output_12_903(.a(output_13_903), .b(output_13_8), .y(output_12_903));
wire output_14_903, output_14_8, output_13_903;
mixer gate_output_13_903(.a(output_14_903), .b(output_14_8), .y(output_13_903));
wire output_15_903, output_15_8, output_14_903;
mixer gate_output_14_903(.a(output_15_903), .b(output_15_8), .y(output_14_903));
wire output_16_903, output_16_8, output_15_903;
mixer gate_output_15_903(.a(output_16_903), .b(output_16_8), .y(output_15_903));
wire output_1_904, output_1_9, output_0_904;
mixer gate_output_0_904(.a(output_1_904), .b(output_1_9), .y(output_0_904));
wire output_2_904, output_2_9, output_1_904;
mixer gate_output_1_904(.a(output_2_904), .b(output_2_9), .y(output_1_904));
wire output_3_904, output_3_9, output_2_904;
mixer gate_output_2_904(.a(output_3_904), .b(output_3_9), .y(output_2_904));
wire output_4_904, output_4_9, output_3_904;
mixer gate_output_3_904(.a(output_4_904), .b(output_4_9), .y(output_3_904));
wire output_5_904, output_5_9, output_4_904;
mixer gate_output_4_904(.a(output_5_904), .b(output_5_9), .y(output_4_904));
wire output_6_904, output_6_9, output_5_904;
mixer gate_output_5_904(.a(output_6_904), .b(output_6_9), .y(output_5_904));
wire output_7_904, output_7_9, output_6_904;
mixer gate_output_6_904(.a(output_7_904), .b(output_7_9), .y(output_6_904));
wire output_8_904, output_8_9, output_7_904;
mixer gate_output_7_904(.a(output_8_904), .b(output_8_9), .y(output_7_904));
wire output_9_904, output_9_9, output_8_904;
mixer gate_output_8_904(.a(output_9_904), .b(output_9_9), .y(output_8_904));
wire output_10_904, output_10_9, output_9_904;
mixer gate_output_9_904(.a(output_10_904), .b(output_10_9), .y(output_9_904));
wire output_11_904, output_11_9, output_10_904;
mixer gate_output_10_904(.a(output_11_904), .b(output_11_9), .y(output_10_904));
wire output_12_904, output_12_9, output_11_904;
mixer gate_output_11_904(.a(output_12_904), .b(output_12_9), .y(output_11_904));
wire output_13_904, output_13_9, output_12_904;
mixer gate_output_12_904(.a(output_13_904), .b(output_13_9), .y(output_12_904));
wire output_14_904, output_14_9, output_13_904;
mixer gate_output_13_904(.a(output_14_904), .b(output_14_9), .y(output_13_904));
wire output_15_904, output_15_9, output_14_904;
mixer gate_output_14_904(.a(output_15_904), .b(output_15_9), .y(output_14_904));
wire output_16_904, output_16_9, output_15_904;
mixer gate_output_15_904(.a(output_16_904), .b(output_16_9), .y(output_15_904));
wire output_1_905, output_1_10, output_0_905;
mixer gate_output_0_905(.a(output_1_905), .b(output_1_10), .y(output_0_905));
wire output_2_905, output_2_10, output_1_905;
mixer gate_output_1_905(.a(output_2_905), .b(output_2_10), .y(output_1_905));
wire output_3_905, output_3_10, output_2_905;
mixer gate_output_2_905(.a(output_3_905), .b(output_3_10), .y(output_2_905));
wire output_4_905, output_4_10, output_3_905;
mixer gate_output_3_905(.a(output_4_905), .b(output_4_10), .y(output_3_905));
wire output_5_905, output_5_10, output_4_905;
mixer gate_output_4_905(.a(output_5_905), .b(output_5_10), .y(output_4_905));
wire output_6_905, output_6_10, output_5_905;
mixer gate_output_5_905(.a(output_6_905), .b(output_6_10), .y(output_5_905));
wire output_7_905, output_7_10, output_6_905;
mixer gate_output_6_905(.a(output_7_905), .b(output_7_10), .y(output_6_905));
wire output_8_905, output_8_10, output_7_905;
mixer gate_output_7_905(.a(output_8_905), .b(output_8_10), .y(output_7_905));
wire output_9_905, output_9_10, output_8_905;
mixer gate_output_8_905(.a(output_9_905), .b(output_9_10), .y(output_8_905));
wire output_10_905, output_10_10, output_9_905;
mixer gate_output_9_905(.a(output_10_905), .b(output_10_10), .y(output_9_905));
wire output_11_905, output_11_10, output_10_905;
mixer gate_output_10_905(.a(output_11_905), .b(output_11_10), .y(output_10_905));
wire output_12_905, output_12_10, output_11_905;
mixer gate_output_11_905(.a(output_12_905), .b(output_12_10), .y(output_11_905));
wire output_13_905, output_13_10, output_12_905;
mixer gate_output_12_905(.a(output_13_905), .b(output_13_10), .y(output_12_905));
wire output_14_905, output_14_10, output_13_905;
mixer gate_output_13_905(.a(output_14_905), .b(output_14_10), .y(output_13_905));
wire output_15_905, output_15_10, output_14_905;
mixer gate_output_14_905(.a(output_15_905), .b(output_15_10), .y(output_14_905));
wire output_16_905, output_16_10, output_15_905;
mixer gate_output_15_905(.a(output_16_905), .b(output_16_10), .y(output_15_905));
wire output_1_906, output_1_11, output_0_906;
mixer gate_output_0_906(.a(output_1_906), .b(output_1_11), .y(output_0_906));
wire output_2_906, output_2_11, output_1_906;
mixer gate_output_1_906(.a(output_2_906), .b(output_2_11), .y(output_1_906));
wire output_3_906, output_3_11, output_2_906;
mixer gate_output_2_906(.a(output_3_906), .b(output_3_11), .y(output_2_906));
wire output_4_906, output_4_11, output_3_906;
mixer gate_output_3_906(.a(output_4_906), .b(output_4_11), .y(output_3_906));
wire output_5_906, output_5_11, output_4_906;
mixer gate_output_4_906(.a(output_5_906), .b(output_5_11), .y(output_4_906));
wire output_6_906, output_6_11, output_5_906;
mixer gate_output_5_906(.a(output_6_906), .b(output_6_11), .y(output_5_906));
wire output_7_906, output_7_11, output_6_906;
mixer gate_output_6_906(.a(output_7_906), .b(output_7_11), .y(output_6_906));
wire output_8_906, output_8_11, output_7_906;
mixer gate_output_7_906(.a(output_8_906), .b(output_8_11), .y(output_7_906));
wire output_9_906, output_9_11, output_8_906;
mixer gate_output_8_906(.a(output_9_906), .b(output_9_11), .y(output_8_906));
wire output_10_906, output_10_11, output_9_906;
mixer gate_output_9_906(.a(output_10_906), .b(output_10_11), .y(output_9_906));
wire output_11_906, output_11_11, output_10_906;
mixer gate_output_10_906(.a(output_11_906), .b(output_11_11), .y(output_10_906));
wire output_12_906, output_12_11, output_11_906;
mixer gate_output_11_906(.a(output_12_906), .b(output_12_11), .y(output_11_906));
wire output_13_906, output_13_11, output_12_906;
mixer gate_output_12_906(.a(output_13_906), .b(output_13_11), .y(output_12_906));
wire output_14_906, output_14_11, output_13_906;
mixer gate_output_13_906(.a(output_14_906), .b(output_14_11), .y(output_13_906));
wire output_15_906, output_15_11, output_14_906;
mixer gate_output_14_906(.a(output_15_906), .b(output_15_11), .y(output_14_906));
wire output_16_906, output_16_11, output_15_906;
mixer gate_output_15_906(.a(output_16_906), .b(output_16_11), .y(output_15_906));
wire output_1_907, output_1_12, output_0_907;
mixer gate_output_0_907(.a(output_1_907), .b(output_1_12), .y(output_0_907));
wire output_2_907, output_2_12, output_1_907;
mixer gate_output_1_907(.a(output_2_907), .b(output_2_12), .y(output_1_907));
wire output_3_907, output_3_12, output_2_907;
mixer gate_output_2_907(.a(output_3_907), .b(output_3_12), .y(output_2_907));
wire output_4_907, output_4_12, output_3_907;
mixer gate_output_3_907(.a(output_4_907), .b(output_4_12), .y(output_3_907));
wire output_5_907, output_5_12, output_4_907;
mixer gate_output_4_907(.a(output_5_907), .b(output_5_12), .y(output_4_907));
wire output_6_907, output_6_12, output_5_907;
mixer gate_output_5_907(.a(output_6_907), .b(output_6_12), .y(output_5_907));
wire output_7_907, output_7_12, output_6_907;
mixer gate_output_6_907(.a(output_7_907), .b(output_7_12), .y(output_6_907));
wire output_8_907, output_8_12, output_7_907;
mixer gate_output_7_907(.a(output_8_907), .b(output_8_12), .y(output_7_907));
wire output_9_907, output_9_12, output_8_907;
mixer gate_output_8_907(.a(output_9_907), .b(output_9_12), .y(output_8_907));
wire output_10_907, output_10_12, output_9_907;
mixer gate_output_9_907(.a(output_10_907), .b(output_10_12), .y(output_9_907));
wire output_11_907, output_11_12, output_10_907;
mixer gate_output_10_907(.a(output_11_907), .b(output_11_12), .y(output_10_907));
wire output_12_907, output_12_12, output_11_907;
mixer gate_output_11_907(.a(output_12_907), .b(output_12_12), .y(output_11_907));
wire output_13_907, output_13_12, output_12_907;
mixer gate_output_12_907(.a(output_13_907), .b(output_13_12), .y(output_12_907));
wire output_14_907, output_14_12, output_13_907;
mixer gate_output_13_907(.a(output_14_907), .b(output_14_12), .y(output_13_907));
wire output_15_907, output_15_12, output_14_907;
mixer gate_output_14_907(.a(output_15_907), .b(output_15_12), .y(output_14_907));
wire output_16_907, output_16_12, output_15_907;
mixer gate_output_15_907(.a(output_16_907), .b(output_16_12), .y(output_15_907));
wire output_1_908, output_1_13, output_0_908;
mixer gate_output_0_908(.a(output_1_908), .b(output_1_13), .y(output_0_908));
wire output_2_908, output_2_13, output_1_908;
mixer gate_output_1_908(.a(output_2_908), .b(output_2_13), .y(output_1_908));
wire output_3_908, output_3_13, output_2_908;
mixer gate_output_2_908(.a(output_3_908), .b(output_3_13), .y(output_2_908));
wire output_4_908, output_4_13, output_3_908;
mixer gate_output_3_908(.a(output_4_908), .b(output_4_13), .y(output_3_908));
wire output_5_908, output_5_13, output_4_908;
mixer gate_output_4_908(.a(output_5_908), .b(output_5_13), .y(output_4_908));
wire output_6_908, output_6_13, output_5_908;
mixer gate_output_5_908(.a(output_6_908), .b(output_6_13), .y(output_5_908));
wire output_7_908, output_7_13, output_6_908;
mixer gate_output_6_908(.a(output_7_908), .b(output_7_13), .y(output_6_908));
wire output_8_908, output_8_13, output_7_908;
mixer gate_output_7_908(.a(output_8_908), .b(output_8_13), .y(output_7_908));
wire output_9_908, output_9_13, output_8_908;
mixer gate_output_8_908(.a(output_9_908), .b(output_9_13), .y(output_8_908));
wire output_10_908, output_10_13, output_9_908;
mixer gate_output_9_908(.a(output_10_908), .b(output_10_13), .y(output_9_908));
wire output_11_908, output_11_13, output_10_908;
mixer gate_output_10_908(.a(output_11_908), .b(output_11_13), .y(output_10_908));
wire output_12_908, output_12_13, output_11_908;
mixer gate_output_11_908(.a(output_12_908), .b(output_12_13), .y(output_11_908));
wire output_13_908, output_13_13, output_12_908;
mixer gate_output_12_908(.a(output_13_908), .b(output_13_13), .y(output_12_908));
wire output_14_908, output_14_13, output_13_908;
mixer gate_output_13_908(.a(output_14_908), .b(output_14_13), .y(output_13_908));
wire output_15_908, output_15_13, output_14_908;
mixer gate_output_14_908(.a(output_15_908), .b(output_15_13), .y(output_14_908));
wire output_16_908, output_16_13, output_15_908;
mixer gate_output_15_908(.a(output_16_908), .b(output_16_13), .y(output_15_908));
wire output_1_909, output_1_14, output_0_909;
mixer gate_output_0_909(.a(output_1_909), .b(output_1_14), .y(output_0_909));
wire output_2_909, output_2_14, output_1_909;
mixer gate_output_1_909(.a(output_2_909), .b(output_2_14), .y(output_1_909));
wire output_3_909, output_3_14, output_2_909;
mixer gate_output_2_909(.a(output_3_909), .b(output_3_14), .y(output_2_909));
wire output_4_909, output_4_14, output_3_909;
mixer gate_output_3_909(.a(output_4_909), .b(output_4_14), .y(output_3_909));
wire output_5_909, output_5_14, output_4_909;
mixer gate_output_4_909(.a(output_5_909), .b(output_5_14), .y(output_4_909));
wire output_6_909, output_6_14, output_5_909;
mixer gate_output_5_909(.a(output_6_909), .b(output_6_14), .y(output_5_909));
wire output_7_909, output_7_14, output_6_909;
mixer gate_output_6_909(.a(output_7_909), .b(output_7_14), .y(output_6_909));
wire output_8_909, output_8_14, output_7_909;
mixer gate_output_7_909(.a(output_8_909), .b(output_8_14), .y(output_7_909));
wire output_9_909, output_9_14, output_8_909;
mixer gate_output_8_909(.a(output_9_909), .b(output_9_14), .y(output_8_909));
wire output_10_909, output_10_14, output_9_909;
mixer gate_output_9_909(.a(output_10_909), .b(output_10_14), .y(output_9_909));
wire output_11_909, output_11_14, output_10_909;
mixer gate_output_10_909(.a(output_11_909), .b(output_11_14), .y(output_10_909));
wire output_12_909, output_12_14, output_11_909;
mixer gate_output_11_909(.a(output_12_909), .b(output_12_14), .y(output_11_909));
wire output_13_909, output_13_14, output_12_909;
mixer gate_output_12_909(.a(output_13_909), .b(output_13_14), .y(output_12_909));
wire output_14_909, output_14_14, output_13_909;
mixer gate_output_13_909(.a(output_14_909), .b(output_14_14), .y(output_13_909));
wire output_15_909, output_15_14, output_14_909;
mixer gate_output_14_909(.a(output_15_909), .b(output_15_14), .y(output_14_909));
wire output_16_909, output_16_14, output_15_909;
mixer gate_output_15_909(.a(output_16_909), .b(output_16_14), .y(output_15_909));
wire output_1_910, output_1_15, output_0_910;
mixer gate_output_0_910(.a(output_1_910), .b(output_1_15), .y(output_0_910));
wire output_2_910, output_2_15, output_1_910;
mixer gate_output_1_910(.a(output_2_910), .b(output_2_15), .y(output_1_910));
wire output_3_910, output_3_15, output_2_910;
mixer gate_output_2_910(.a(output_3_910), .b(output_3_15), .y(output_2_910));
wire output_4_910, output_4_15, output_3_910;
mixer gate_output_3_910(.a(output_4_910), .b(output_4_15), .y(output_3_910));
wire output_5_910, output_5_15, output_4_910;
mixer gate_output_4_910(.a(output_5_910), .b(output_5_15), .y(output_4_910));
wire output_6_910, output_6_15, output_5_910;
mixer gate_output_5_910(.a(output_6_910), .b(output_6_15), .y(output_5_910));
wire output_7_910, output_7_15, output_6_910;
mixer gate_output_6_910(.a(output_7_910), .b(output_7_15), .y(output_6_910));
wire output_8_910, output_8_15, output_7_910;
mixer gate_output_7_910(.a(output_8_910), .b(output_8_15), .y(output_7_910));
wire output_9_910, output_9_15, output_8_910;
mixer gate_output_8_910(.a(output_9_910), .b(output_9_15), .y(output_8_910));
wire output_10_910, output_10_15, output_9_910;
mixer gate_output_9_910(.a(output_10_910), .b(output_10_15), .y(output_9_910));
wire output_11_910, output_11_15, output_10_910;
mixer gate_output_10_910(.a(output_11_910), .b(output_11_15), .y(output_10_910));
wire output_12_910, output_12_15, output_11_910;
mixer gate_output_11_910(.a(output_12_910), .b(output_12_15), .y(output_11_910));
wire output_13_910, output_13_15, output_12_910;
mixer gate_output_12_910(.a(output_13_910), .b(output_13_15), .y(output_12_910));
wire output_14_910, output_14_15, output_13_910;
mixer gate_output_13_910(.a(output_14_910), .b(output_14_15), .y(output_13_910));
wire output_15_910, output_15_15, output_14_910;
mixer gate_output_14_910(.a(output_15_910), .b(output_15_15), .y(output_14_910));
wire output_16_910, output_16_15, output_15_910;
mixer gate_output_15_910(.a(output_16_910), .b(output_16_15), .y(output_15_910));
wire output_1_911, output_1_0, output_0_911;
mixer gate_output_0_911(.a(output_1_911), .b(output_1_0), .y(output_0_911));
wire output_2_911, output_2_0, output_1_911;
mixer gate_output_1_911(.a(output_2_911), .b(output_2_0), .y(output_1_911));
wire output_3_911, output_3_0, output_2_911;
mixer gate_output_2_911(.a(output_3_911), .b(output_3_0), .y(output_2_911));
wire output_4_911, output_4_0, output_3_911;
mixer gate_output_3_911(.a(output_4_911), .b(output_4_0), .y(output_3_911));
wire output_5_911, output_5_0, output_4_911;
mixer gate_output_4_911(.a(output_5_911), .b(output_5_0), .y(output_4_911));
wire output_6_911, output_6_0, output_5_911;
mixer gate_output_5_911(.a(output_6_911), .b(output_6_0), .y(output_5_911));
wire output_7_911, output_7_0, output_6_911;
mixer gate_output_6_911(.a(output_7_911), .b(output_7_0), .y(output_6_911));
wire output_8_911, output_8_0, output_7_911;
mixer gate_output_7_911(.a(output_8_911), .b(output_8_0), .y(output_7_911));
wire output_9_911, output_9_0, output_8_911;
mixer gate_output_8_911(.a(output_9_911), .b(output_9_0), .y(output_8_911));
wire output_10_911, output_10_0, output_9_911;
mixer gate_output_9_911(.a(output_10_911), .b(output_10_0), .y(output_9_911));
wire output_11_911, output_11_0, output_10_911;
mixer gate_output_10_911(.a(output_11_911), .b(output_11_0), .y(output_10_911));
wire output_12_911, output_12_0, output_11_911;
mixer gate_output_11_911(.a(output_12_911), .b(output_12_0), .y(output_11_911));
wire output_13_911, output_13_0, output_12_911;
mixer gate_output_12_911(.a(output_13_911), .b(output_13_0), .y(output_12_911));
wire output_14_911, output_14_0, output_13_911;
mixer gate_output_13_911(.a(output_14_911), .b(output_14_0), .y(output_13_911));
wire output_15_911, output_15_0, output_14_911;
mixer gate_output_14_911(.a(output_15_911), .b(output_15_0), .y(output_14_911));
wire output_16_911, output_16_0, output_15_911;
mixer gate_output_15_911(.a(output_16_911), .b(output_16_0), .y(output_15_911));
wire output_1_912, output_1_1, output_0_912;
mixer gate_output_0_912(.a(output_1_912), .b(output_1_1), .y(output_0_912));
wire output_2_912, output_2_1, output_1_912;
mixer gate_output_1_912(.a(output_2_912), .b(output_2_1), .y(output_1_912));
wire output_3_912, output_3_1, output_2_912;
mixer gate_output_2_912(.a(output_3_912), .b(output_3_1), .y(output_2_912));
wire output_4_912, output_4_1, output_3_912;
mixer gate_output_3_912(.a(output_4_912), .b(output_4_1), .y(output_3_912));
wire output_5_912, output_5_1, output_4_912;
mixer gate_output_4_912(.a(output_5_912), .b(output_5_1), .y(output_4_912));
wire output_6_912, output_6_1, output_5_912;
mixer gate_output_5_912(.a(output_6_912), .b(output_6_1), .y(output_5_912));
wire output_7_912, output_7_1, output_6_912;
mixer gate_output_6_912(.a(output_7_912), .b(output_7_1), .y(output_6_912));
wire output_8_912, output_8_1, output_7_912;
mixer gate_output_7_912(.a(output_8_912), .b(output_8_1), .y(output_7_912));
wire output_9_912, output_9_1, output_8_912;
mixer gate_output_8_912(.a(output_9_912), .b(output_9_1), .y(output_8_912));
wire output_10_912, output_10_1, output_9_912;
mixer gate_output_9_912(.a(output_10_912), .b(output_10_1), .y(output_9_912));
wire output_11_912, output_11_1, output_10_912;
mixer gate_output_10_912(.a(output_11_912), .b(output_11_1), .y(output_10_912));
wire output_12_912, output_12_1, output_11_912;
mixer gate_output_11_912(.a(output_12_912), .b(output_12_1), .y(output_11_912));
wire output_13_912, output_13_1, output_12_912;
mixer gate_output_12_912(.a(output_13_912), .b(output_13_1), .y(output_12_912));
wire output_14_912, output_14_1, output_13_912;
mixer gate_output_13_912(.a(output_14_912), .b(output_14_1), .y(output_13_912));
wire output_15_912, output_15_1, output_14_912;
mixer gate_output_14_912(.a(output_15_912), .b(output_15_1), .y(output_14_912));
wire output_16_912, output_16_1, output_15_912;
mixer gate_output_15_912(.a(output_16_912), .b(output_16_1), .y(output_15_912));
wire output_1_913, output_1_2, output_0_913;
mixer gate_output_0_913(.a(output_1_913), .b(output_1_2), .y(output_0_913));
wire output_2_913, output_2_2, output_1_913;
mixer gate_output_1_913(.a(output_2_913), .b(output_2_2), .y(output_1_913));
wire output_3_913, output_3_2, output_2_913;
mixer gate_output_2_913(.a(output_3_913), .b(output_3_2), .y(output_2_913));
wire output_4_913, output_4_2, output_3_913;
mixer gate_output_3_913(.a(output_4_913), .b(output_4_2), .y(output_3_913));
wire output_5_913, output_5_2, output_4_913;
mixer gate_output_4_913(.a(output_5_913), .b(output_5_2), .y(output_4_913));
wire output_6_913, output_6_2, output_5_913;
mixer gate_output_5_913(.a(output_6_913), .b(output_6_2), .y(output_5_913));
wire output_7_913, output_7_2, output_6_913;
mixer gate_output_6_913(.a(output_7_913), .b(output_7_2), .y(output_6_913));
wire output_8_913, output_8_2, output_7_913;
mixer gate_output_7_913(.a(output_8_913), .b(output_8_2), .y(output_7_913));
wire output_9_913, output_9_2, output_8_913;
mixer gate_output_8_913(.a(output_9_913), .b(output_9_2), .y(output_8_913));
wire output_10_913, output_10_2, output_9_913;
mixer gate_output_9_913(.a(output_10_913), .b(output_10_2), .y(output_9_913));
wire output_11_913, output_11_2, output_10_913;
mixer gate_output_10_913(.a(output_11_913), .b(output_11_2), .y(output_10_913));
wire output_12_913, output_12_2, output_11_913;
mixer gate_output_11_913(.a(output_12_913), .b(output_12_2), .y(output_11_913));
wire output_13_913, output_13_2, output_12_913;
mixer gate_output_12_913(.a(output_13_913), .b(output_13_2), .y(output_12_913));
wire output_14_913, output_14_2, output_13_913;
mixer gate_output_13_913(.a(output_14_913), .b(output_14_2), .y(output_13_913));
wire output_15_913, output_15_2, output_14_913;
mixer gate_output_14_913(.a(output_15_913), .b(output_15_2), .y(output_14_913));
wire output_16_913, output_16_2, output_15_913;
mixer gate_output_15_913(.a(output_16_913), .b(output_16_2), .y(output_15_913));
wire output_1_914, output_1_3, output_0_914;
mixer gate_output_0_914(.a(output_1_914), .b(output_1_3), .y(output_0_914));
wire output_2_914, output_2_3, output_1_914;
mixer gate_output_1_914(.a(output_2_914), .b(output_2_3), .y(output_1_914));
wire output_3_914, output_3_3, output_2_914;
mixer gate_output_2_914(.a(output_3_914), .b(output_3_3), .y(output_2_914));
wire output_4_914, output_4_3, output_3_914;
mixer gate_output_3_914(.a(output_4_914), .b(output_4_3), .y(output_3_914));
wire output_5_914, output_5_3, output_4_914;
mixer gate_output_4_914(.a(output_5_914), .b(output_5_3), .y(output_4_914));
wire output_6_914, output_6_3, output_5_914;
mixer gate_output_5_914(.a(output_6_914), .b(output_6_3), .y(output_5_914));
wire output_7_914, output_7_3, output_6_914;
mixer gate_output_6_914(.a(output_7_914), .b(output_7_3), .y(output_6_914));
wire output_8_914, output_8_3, output_7_914;
mixer gate_output_7_914(.a(output_8_914), .b(output_8_3), .y(output_7_914));
wire output_9_914, output_9_3, output_8_914;
mixer gate_output_8_914(.a(output_9_914), .b(output_9_3), .y(output_8_914));
wire output_10_914, output_10_3, output_9_914;
mixer gate_output_9_914(.a(output_10_914), .b(output_10_3), .y(output_9_914));
wire output_11_914, output_11_3, output_10_914;
mixer gate_output_10_914(.a(output_11_914), .b(output_11_3), .y(output_10_914));
wire output_12_914, output_12_3, output_11_914;
mixer gate_output_11_914(.a(output_12_914), .b(output_12_3), .y(output_11_914));
wire output_13_914, output_13_3, output_12_914;
mixer gate_output_12_914(.a(output_13_914), .b(output_13_3), .y(output_12_914));
wire output_14_914, output_14_3, output_13_914;
mixer gate_output_13_914(.a(output_14_914), .b(output_14_3), .y(output_13_914));
wire output_15_914, output_15_3, output_14_914;
mixer gate_output_14_914(.a(output_15_914), .b(output_15_3), .y(output_14_914));
wire output_16_914, output_16_3, output_15_914;
mixer gate_output_15_914(.a(output_16_914), .b(output_16_3), .y(output_15_914));
wire output_1_915, output_1_4, output_0_915;
mixer gate_output_0_915(.a(output_1_915), .b(output_1_4), .y(output_0_915));
wire output_2_915, output_2_4, output_1_915;
mixer gate_output_1_915(.a(output_2_915), .b(output_2_4), .y(output_1_915));
wire output_3_915, output_3_4, output_2_915;
mixer gate_output_2_915(.a(output_3_915), .b(output_3_4), .y(output_2_915));
wire output_4_915, output_4_4, output_3_915;
mixer gate_output_3_915(.a(output_4_915), .b(output_4_4), .y(output_3_915));
wire output_5_915, output_5_4, output_4_915;
mixer gate_output_4_915(.a(output_5_915), .b(output_5_4), .y(output_4_915));
wire output_6_915, output_6_4, output_5_915;
mixer gate_output_5_915(.a(output_6_915), .b(output_6_4), .y(output_5_915));
wire output_7_915, output_7_4, output_6_915;
mixer gate_output_6_915(.a(output_7_915), .b(output_7_4), .y(output_6_915));
wire output_8_915, output_8_4, output_7_915;
mixer gate_output_7_915(.a(output_8_915), .b(output_8_4), .y(output_7_915));
wire output_9_915, output_9_4, output_8_915;
mixer gate_output_8_915(.a(output_9_915), .b(output_9_4), .y(output_8_915));
wire output_10_915, output_10_4, output_9_915;
mixer gate_output_9_915(.a(output_10_915), .b(output_10_4), .y(output_9_915));
wire output_11_915, output_11_4, output_10_915;
mixer gate_output_10_915(.a(output_11_915), .b(output_11_4), .y(output_10_915));
wire output_12_915, output_12_4, output_11_915;
mixer gate_output_11_915(.a(output_12_915), .b(output_12_4), .y(output_11_915));
wire output_13_915, output_13_4, output_12_915;
mixer gate_output_12_915(.a(output_13_915), .b(output_13_4), .y(output_12_915));
wire output_14_915, output_14_4, output_13_915;
mixer gate_output_13_915(.a(output_14_915), .b(output_14_4), .y(output_13_915));
wire output_15_915, output_15_4, output_14_915;
mixer gate_output_14_915(.a(output_15_915), .b(output_15_4), .y(output_14_915));
wire output_16_915, output_16_4, output_15_915;
mixer gate_output_15_915(.a(output_16_915), .b(output_16_4), .y(output_15_915));
wire output_1_916, output_1_5, output_0_916;
mixer gate_output_0_916(.a(output_1_916), .b(output_1_5), .y(output_0_916));
wire output_2_916, output_2_5, output_1_916;
mixer gate_output_1_916(.a(output_2_916), .b(output_2_5), .y(output_1_916));
wire output_3_916, output_3_5, output_2_916;
mixer gate_output_2_916(.a(output_3_916), .b(output_3_5), .y(output_2_916));
wire output_4_916, output_4_5, output_3_916;
mixer gate_output_3_916(.a(output_4_916), .b(output_4_5), .y(output_3_916));
wire output_5_916, output_5_5, output_4_916;
mixer gate_output_4_916(.a(output_5_916), .b(output_5_5), .y(output_4_916));
wire output_6_916, output_6_5, output_5_916;
mixer gate_output_5_916(.a(output_6_916), .b(output_6_5), .y(output_5_916));
wire output_7_916, output_7_5, output_6_916;
mixer gate_output_6_916(.a(output_7_916), .b(output_7_5), .y(output_6_916));
wire output_8_916, output_8_5, output_7_916;
mixer gate_output_7_916(.a(output_8_916), .b(output_8_5), .y(output_7_916));
wire output_9_916, output_9_5, output_8_916;
mixer gate_output_8_916(.a(output_9_916), .b(output_9_5), .y(output_8_916));
wire output_10_916, output_10_5, output_9_916;
mixer gate_output_9_916(.a(output_10_916), .b(output_10_5), .y(output_9_916));
wire output_11_916, output_11_5, output_10_916;
mixer gate_output_10_916(.a(output_11_916), .b(output_11_5), .y(output_10_916));
wire output_12_916, output_12_5, output_11_916;
mixer gate_output_11_916(.a(output_12_916), .b(output_12_5), .y(output_11_916));
wire output_13_916, output_13_5, output_12_916;
mixer gate_output_12_916(.a(output_13_916), .b(output_13_5), .y(output_12_916));
wire output_14_916, output_14_5, output_13_916;
mixer gate_output_13_916(.a(output_14_916), .b(output_14_5), .y(output_13_916));
wire output_15_916, output_15_5, output_14_916;
mixer gate_output_14_916(.a(output_15_916), .b(output_15_5), .y(output_14_916));
wire output_16_916, output_16_5, output_15_916;
mixer gate_output_15_916(.a(output_16_916), .b(output_16_5), .y(output_15_916));
wire output_1_917, output_1_6, output_0_917;
mixer gate_output_0_917(.a(output_1_917), .b(output_1_6), .y(output_0_917));
wire output_2_917, output_2_6, output_1_917;
mixer gate_output_1_917(.a(output_2_917), .b(output_2_6), .y(output_1_917));
wire output_3_917, output_3_6, output_2_917;
mixer gate_output_2_917(.a(output_3_917), .b(output_3_6), .y(output_2_917));
wire output_4_917, output_4_6, output_3_917;
mixer gate_output_3_917(.a(output_4_917), .b(output_4_6), .y(output_3_917));
wire output_5_917, output_5_6, output_4_917;
mixer gate_output_4_917(.a(output_5_917), .b(output_5_6), .y(output_4_917));
wire output_6_917, output_6_6, output_5_917;
mixer gate_output_5_917(.a(output_6_917), .b(output_6_6), .y(output_5_917));
wire output_7_917, output_7_6, output_6_917;
mixer gate_output_6_917(.a(output_7_917), .b(output_7_6), .y(output_6_917));
wire output_8_917, output_8_6, output_7_917;
mixer gate_output_7_917(.a(output_8_917), .b(output_8_6), .y(output_7_917));
wire output_9_917, output_9_6, output_8_917;
mixer gate_output_8_917(.a(output_9_917), .b(output_9_6), .y(output_8_917));
wire output_10_917, output_10_6, output_9_917;
mixer gate_output_9_917(.a(output_10_917), .b(output_10_6), .y(output_9_917));
wire output_11_917, output_11_6, output_10_917;
mixer gate_output_10_917(.a(output_11_917), .b(output_11_6), .y(output_10_917));
wire output_12_917, output_12_6, output_11_917;
mixer gate_output_11_917(.a(output_12_917), .b(output_12_6), .y(output_11_917));
wire output_13_917, output_13_6, output_12_917;
mixer gate_output_12_917(.a(output_13_917), .b(output_13_6), .y(output_12_917));
wire output_14_917, output_14_6, output_13_917;
mixer gate_output_13_917(.a(output_14_917), .b(output_14_6), .y(output_13_917));
wire output_15_917, output_15_6, output_14_917;
mixer gate_output_14_917(.a(output_15_917), .b(output_15_6), .y(output_14_917));
wire output_16_917, output_16_6, output_15_917;
mixer gate_output_15_917(.a(output_16_917), .b(output_16_6), .y(output_15_917));
wire output_1_918, output_1_7, output_0_918;
mixer gate_output_0_918(.a(output_1_918), .b(output_1_7), .y(output_0_918));
wire output_2_918, output_2_7, output_1_918;
mixer gate_output_1_918(.a(output_2_918), .b(output_2_7), .y(output_1_918));
wire output_3_918, output_3_7, output_2_918;
mixer gate_output_2_918(.a(output_3_918), .b(output_3_7), .y(output_2_918));
wire output_4_918, output_4_7, output_3_918;
mixer gate_output_3_918(.a(output_4_918), .b(output_4_7), .y(output_3_918));
wire output_5_918, output_5_7, output_4_918;
mixer gate_output_4_918(.a(output_5_918), .b(output_5_7), .y(output_4_918));
wire output_6_918, output_6_7, output_5_918;
mixer gate_output_5_918(.a(output_6_918), .b(output_6_7), .y(output_5_918));
wire output_7_918, output_7_7, output_6_918;
mixer gate_output_6_918(.a(output_7_918), .b(output_7_7), .y(output_6_918));
wire output_8_918, output_8_7, output_7_918;
mixer gate_output_7_918(.a(output_8_918), .b(output_8_7), .y(output_7_918));
wire output_9_918, output_9_7, output_8_918;
mixer gate_output_8_918(.a(output_9_918), .b(output_9_7), .y(output_8_918));
wire output_10_918, output_10_7, output_9_918;
mixer gate_output_9_918(.a(output_10_918), .b(output_10_7), .y(output_9_918));
wire output_11_918, output_11_7, output_10_918;
mixer gate_output_10_918(.a(output_11_918), .b(output_11_7), .y(output_10_918));
wire output_12_918, output_12_7, output_11_918;
mixer gate_output_11_918(.a(output_12_918), .b(output_12_7), .y(output_11_918));
wire output_13_918, output_13_7, output_12_918;
mixer gate_output_12_918(.a(output_13_918), .b(output_13_7), .y(output_12_918));
wire output_14_918, output_14_7, output_13_918;
mixer gate_output_13_918(.a(output_14_918), .b(output_14_7), .y(output_13_918));
wire output_15_918, output_15_7, output_14_918;
mixer gate_output_14_918(.a(output_15_918), .b(output_15_7), .y(output_14_918));
wire output_16_918, output_16_7, output_15_918;
mixer gate_output_15_918(.a(output_16_918), .b(output_16_7), .y(output_15_918));
wire output_1_919, output_1_8, output_0_919;
mixer gate_output_0_919(.a(output_1_919), .b(output_1_8), .y(output_0_919));
wire output_2_919, output_2_8, output_1_919;
mixer gate_output_1_919(.a(output_2_919), .b(output_2_8), .y(output_1_919));
wire output_3_919, output_3_8, output_2_919;
mixer gate_output_2_919(.a(output_3_919), .b(output_3_8), .y(output_2_919));
wire output_4_919, output_4_8, output_3_919;
mixer gate_output_3_919(.a(output_4_919), .b(output_4_8), .y(output_3_919));
wire output_5_919, output_5_8, output_4_919;
mixer gate_output_4_919(.a(output_5_919), .b(output_5_8), .y(output_4_919));
wire output_6_919, output_6_8, output_5_919;
mixer gate_output_5_919(.a(output_6_919), .b(output_6_8), .y(output_5_919));
wire output_7_919, output_7_8, output_6_919;
mixer gate_output_6_919(.a(output_7_919), .b(output_7_8), .y(output_6_919));
wire output_8_919, output_8_8, output_7_919;
mixer gate_output_7_919(.a(output_8_919), .b(output_8_8), .y(output_7_919));
wire output_9_919, output_9_8, output_8_919;
mixer gate_output_8_919(.a(output_9_919), .b(output_9_8), .y(output_8_919));
wire output_10_919, output_10_8, output_9_919;
mixer gate_output_9_919(.a(output_10_919), .b(output_10_8), .y(output_9_919));
wire output_11_919, output_11_8, output_10_919;
mixer gate_output_10_919(.a(output_11_919), .b(output_11_8), .y(output_10_919));
wire output_12_919, output_12_8, output_11_919;
mixer gate_output_11_919(.a(output_12_919), .b(output_12_8), .y(output_11_919));
wire output_13_919, output_13_8, output_12_919;
mixer gate_output_12_919(.a(output_13_919), .b(output_13_8), .y(output_12_919));
wire output_14_919, output_14_8, output_13_919;
mixer gate_output_13_919(.a(output_14_919), .b(output_14_8), .y(output_13_919));
wire output_15_919, output_15_8, output_14_919;
mixer gate_output_14_919(.a(output_15_919), .b(output_15_8), .y(output_14_919));
wire output_16_919, output_16_8, output_15_919;
mixer gate_output_15_919(.a(output_16_919), .b(output_16_8), .y(output_15_919));
wire output_1_920, output_1_9, output_0_920;
mixer gate_output_0_920(.a(output_1_920), .b(output_1_9), .y(output_0_920));
wire output_2_920, output_2_9, output_1_920;
mixer gate_output_1_920(.a(output_2_920), .b(output_2_9), .y(output_1_920));
wire output_3_920, output_3_9, output_2_920;
mixer gate_output_2_920(.a(output_3_920), .b(output_3_9), .y(output_2_920));
wire output_4_920, output_4_9, output_3_920;
mixer gate_output_3_920(.a(output_4_920), .b(output_4_9), .y(output_3_920));
wire output_5_920, output_5_9, output_4_920;
mixer gate_output_4_920(.a(output_5_920), .b(output_5_9), .y(output_4_920));
wire output_6_920, output_6_9, output_5_920;
mixer gate_output_5_920(.a(output_6_920), .b(output_6_9), .y(output_5_920));
wire output_7_920, output_7_9, output_6_920;
mixer gate_output_6_920(.a(output_7_920), .b(output_7_9), .y(output_6_920));
wire output_8_920, output_8_9, output_7_920;
mixer gate_output_7_920(.a(output_8_920), .b(output_8_9), .y(output_7_920));
wire output_9_920, output_9_9, output_8_920;
mixer gate_output_8_920(.a(output_9_920), .b(output_9_9), .y(output_8_920));
wire output_10_920, output_10_9, output_9_920;
mixer gate_output_9_920(.a(output_10_920), .b(output_10_9), .y(output_9_920));
wire output_11_920, output_11_9, output_10_920;
mixer gate_output_10_920(.a(output_11_920), .b(output_11_9), .y(output_10_920));
wire output_12_920, output_12_9, output_11_920;
mixer gate_output_11_920(.a(output_12_920), .b(output_12_9), .y(output_11_920));
wire output_13_920, output_13_9, output_12_920;
mixer gate_output_12_920(.a(output_13_920), .b(output_13_9), .y(output_12_920));
wire output_14_920, output_14_9, output_13_920;
mixer gate_output_13_920(.a(output_14_920), .b(output_14_9), .y(output_13_920));
wire output_15_920, output_15_9, output_14_920;
mixer gate_output_14_920(.a(output_15_920), .b(output_15_9), .y(output_14_920));
wire output_16_920, output_16_9, output_15_920;
mixer gate_output_15_920(.a(output_16_920), .b(output_16_9), .y(output_15_920));
wire output_1_921, output_1_10, output_0_921;
mixer gate_output_0_921(.a(output_1_921), .b(output_1_10), .y(output_0_921));
wire output_2_921, output_2_10, output_1_921;
mixer gate_output_1_921(.a(output_2_921), .b(output_2_10), .y(output_1_921));
wire output_3_921, output_3_10, output_2_921;
mixer gate_output_2_921(.a(output_3_921), .b(output_3_10), .y(output_2_921));
wire output_4_921, output_4_10, output_3_921;
mixer gate_output_3_921(.a(output_4_921), .b(output_4_10), .y(output_3_921));
wire output_5_921, output_5_10, output_4_921;
mixer gate_output_4_921(.a(output_5_921), .b(output_5_10), .y(output_4_921));
wire output_6_921, output_6_10, output_5_921;
mixer gate_output_5_921(.a(output_6_921), .b(output_6_10), .y(output_5_921));
wire output_7_921, output_7_10, output_6_921;
mixer gate_output_6_921(.a(output_7_921), .b(output_7_10), .y(output_6_921));
wire output_8_921, output_8_10, output_7_921;
mixer gate_output_7_921(.a(output_8_921), .b(output_8_10), .y(output_7_921));
wire output_9_921, output_9_10, output_8_921;
mixer gate_output_8_921(.a(output_9_921), .b(output_9_10), .y(output_8_921));
wire output_10_921, output_10_10, output_9_921;
mixer gate_output_9_921(.a(output_10_921), .b(output_10_10), .y(output_9_921));
wire output_11_921, output_11_10, output_10_921;
mixer gate_output_10_921(.a(output_11_921), .b(output_11_10), .y(output_10_921));
wire output_12_921, output_12_10, output_11_921;
mixer gate_output_11_921(.a(output_12_921), .b(output_12_10), .y(output_11_921));
wire output_13_921, output_13_10, output_12_921;
mixer gate_output_12_921(.a(output_13_921), .b(output_13_10), .y(output_12_921));
wire output_14_921, output_14_10, output_13_921;
mixer gate_output_13_921(.a(output_14_921), .b(output_14_10), .y(output_13_921));
wire output_15_921, output_15_10, output_14_921;
mixer gate_output_14_921(.a(output_15_921), .b(output_15_10), .y(output_14_921));
wire output_16_921, output_16_10, output_15_921;
mixer gate_output_15_921(.a(output_16_921), .b(output_16_10), .y(output_15_921));
wire output_1_922, output_1_11, output_0_922;
mixer gate_output_0_922(.a(output_1_922), .b(output_1_11), .y(output_0_922));
wire output_2_922, output_2_11, output_1_922;
mixer gate_output_1_922(.a(output_2_922), .b(output_2_11), .y(output_1_922));
wire output_3_922, output_3_11, output_2_922;
mixer gate_output_2_922(.a(output_3_922), .b(output_3_11), .y(output_2_922));
wire output_4_922, output_4_11, output_3_922;
mixer gate_output_3_922(.a(output_4_922), .b(output_4_11), .y(output_3_922));
wire output_5_922, output_5_11, output_4_922;
mixer gate_output_4_922(.a(output_5_922), .b(output_5_11), .y(output_4_922));
wire output_6_922, output_6_11, output_5_922;
mixer gate_output_5_922(.a(output_6_922), .b(output_6_11), .y(output_5_922));
wire output_7_922, output_7_11, output_6_922;
mixer gate_output_6_922(.a(output_7_922), .b(output_7_11), .y(output_6_922));
wire output_8_922, output_8_11, output_7_922;
mixer gate_output_7_922(.a(output_8_922), .b(output_8_11), .y(output_7_922));
wire output_9_922, output_9_11, output_8_922;
mixer gate_output_8_922(.a(output_9_922), .b(output_9_11), .y(output_8_922));
wire output_10_922, output_10_11, output_9_922;
mixer gate_output_9_922(.a(output_10_922), .b(output_10_11), .y(output_9_922));
wire output_11_922, output_11_11, output_10_922;
mixer gate_output_10_922(.a(output_11_922), .b(output_11_11), .y(output_10_922));
wire output_12_922, output_12_11, output_11_922;
mixer gate_output_11_922(.a(output_12_922), .b(output_12_11), .y(output_11_922));
wire output_13_922, output_13_11, output_12_922;
mixer gate_output_12_922(.a(output_13_922), .b(output_13_11), .y(output_12_922));
wire output_14_922, output_14_11, output_13_922;
mixer gate_output_13_922(.a(output_14_922), .b(output_14_11), .y(output_13_922));
wire output_15_922, output_15_11, output_14_922;
mixer gate_output_14_922(.a(output_15_922), .b(output_15_11), .y(output_14_922));
wire output_16_922, output_16_11, output_15_922;
mixer gate_output_15_922(.a(output_16_922), .b(output_16_11), .y(output_15_922));
wire output_1_923, output_1_12, output_0_923;
mixer gate_output_0_923(.a(output_1_923), .b(output_1_12), .y(output_0_923));
wire output_2_923, output_2_12, output_1_923;
mixer gate_output_1_923(.a(output_2_923), .b(output_2_12), .y(output_1_923));
wire output_3_923, output_3_12, output_2_923;
mixer gate_output_2_923(.a(output_3_923), .b(output_3_12), .y(output_2_923));
wire output_4_923, output_4_12, output_3_923;
mixer gate_output_3_923(.a(output_4_923), .b(output_4_12), .y(output_3_923));
wire output_5_923, output_5_12, output_4_923;
mixer gate_output_4_923(.a(output_5_923), .b(output_5_12), .y(output_4_923));
wire output_6_923, output_6_12, output_5_923;
mixer gate_output_5_923(.a(output_6_923), .b(output_6_12), .y(output_5_923));
wire output_7_923, output_7_12, output_6_923;
mixer gate_output_6_923(.a(output_7_923), .b(output_7_12), .y(output_6_923));
wire output_8_923, output_8_12, output_7_923;
mixer gate_output_7_923(.a(output_8_923), .b(output_8_12), .y(output_7_923));
wire output_9_923, output_9_12, output_8_923;
mixer gate_output_8_923(.a(output_9_923), .b(output_9_12), .y(output_8_923));
wire output_10_923, output_10_12, output_9_923;
mixer gate_output_9_923(.a(output_10_923), .b(output_10_12), .y(output_9_923));
wire output_11_923, output_11_12, output_10_923;
mixer gate_output_10_923(.a(output_11_923), .b(output_11_12), .y(output_10_923));
wire output_12_923, output_12_12, output_11_923;
mixer gate_output_11_923(.a(output_12_923), .b(output_12_12), .y(output_11_923));
wire output_13_923, output_13_12, output_12_923;
mixer gate_output_12_923(.a(output_13_923), .b(output_13_12), .y(output_12_923));
wire output_14_923, output_14_12, output_13_923;
mixer gate_output_13_923(.a(output_14_923), .b(output_14_12), .y(output_13_923));
wire output_15_923, output_15_12, output_14_923;
mixer gate_output_14_923(.a(output_15_923), .b(output_15_12), .y(output_14_923));
wire output_16_923, output_16_12, output_15_923;
mixer gate_output_15_923(.a(output_16_923), .b(output_16_12), .y(output_15_923));
wire output_1_924, output_1_13, output_0_924;
mixer gate_output_0_924(.a(output_1_924), .b(output_1_13), .y(output_0_924));
wire output_2_924, output_2_13, output_1_924;
mixer gate_output_1_924(.a(output_2_924), .b(output_2_13), .y(output_1_924));
wire output_3_924, output_3_13, output_2_924;
mixer gate_output_2_924(.a(output_3_924), .b(output_3_13), .y(output_2_924));
wire output_4_924, output_4_13, output_3_924;
mixer gate_output_3_924(.a(output_4_924), .b(output_4_13), .y(output_3_924));
wire output_5_924, output_5_13, output_4_924;
mixer gate_output_4_924(.a(output_5_924), .b(output_5_13), .y(output_4_924));
wire output_6_924, output_6_13, output_5_924;
mixer gate_output_5_924(.a(output_6_924), .b(output_6_13), .y(output_5_924));
wire output_7_924, output_7_13, output_6_924;
mixer gate_output_6_924(.a(output_7_924), .b(output_7_13), .y(output_6_924));
wire output_8_924, output_8_13, output_7_924;
mixer gate_output_7_924(.a(output_8_924), .b(output_8_13), .y(output_7_924));
wire output_9_924, output_9_13, output_8_924;
mixer gate_output_8_924(.a(output_9_924), .b(output_9_13), .y(output_8_924));
wire output_10_924, output_10_13, output_9_924;
mixer gate_output_9_924(.a(output_10_924), .b(output_10_13), .y(output_9_924));
wire output_11_924, output_11_13, output_10_924;
mixer gate_output_10_924(.a(output_11_924), .b(output_11_13), .y(output_10_924));
wire output_12_924, output_12_13, output_11_924;
mixer gate_output_11_924(.a(output_12_924), .b(output_12_13), .y(output_11_924));
wire output_13_924, output_13_13, output_12_924;
mixer gate_output_12_924(.a(output_13_924), .b(output_13_13), .y(output_12_924));
wire output_14_924, output_14_13, output_13_924;
mixer gate_output_13_924(.a(output_14_924), .b(output_14_13), .y(output_13_924));
wire output_15_924, output_15_13, output_14_924;
mixer gate_output_14_924(.a(output_15_924), .b(output_15_13), .y(output_14_924));
wire output_16_924, output_16_13, output_15_924;
mixer gate_output_15_924(.a(output_16_924), .b(output_16_13), .y(output_15_924));
wire output_1_925, output_1_14, output_0_925;
mixer gate_output_0_925(.a(output_1_925), .b(output_1_14), .y(output_0_925));
wire output_2_925, output_2_14, output_1_925;
mixer gate_output_1_925(.a(output_2_925), .b(output_2_14), .y(output_1_925));
wire output_3_925, output_3_14, output_2_925;
mixer gate_output_2_925(.a(output_3_925), .b(output_3_14), .y(output_2_925));
wire output_4_925, output_4_14, output_3_925;
mixer gate_output_3_925(.a(output_4_925), .b(output_4_14), .y(output_3_925));
wire output_5_925, output_5_14, output_4_925;
mixer gate_output_4_925(.a(output_5_925), .b(output_5_14), .y(output_4_925));
wire output_6_925, output_6_14, output_5_925;
mixer gate_output_5_925(.a(output_6_925), .b(output_6_14), .y(output_5_925));
wire output_7_925, output_7_14, output_6_925;
mixer gate_output_6_925(.a(output_7_925), .b(output_7_14), .y(output_6_925));
wire output_8_925, output_8_14, output_7_925;
mixer gate_output_7_925(.a(output_8_925), .b(output_8_14), .y(output_7_925));
wire output_9_925, output_9_14, output_8_925;
mixer gate_output_8_925(.a(output_9_925), .b(output_9_14), .y(output_8_925));
wire output_10_925, output_10_14, output_9_925;
mixer gate_output_9_925(.a(output_10_925), .b(output_10_14), .y(output_9_925));
wire output_11_925, output_11_14, output_10_925;
mixer gate_output_10_925(.a(output_11_925), .b(output_11_14), .y(output_10_925));
wire output_12_925, output_12_14, output_11_925;
mixer gate_output_11_925(.a(output_12_925), .b(output_12_14), .y(output_11_925));
wire output_13_925, output_13_14, output_12_925;
mixer gate_output_12_925(.a(output_13_925), .b(output_13_14), .y(output_12_925));
wire output_14_925, output_14_14, output_13_925;
mixer gate_output_13_925(.a(output_14_925), .b(output_14_14), .y(output_13_925));
wire output_15_925, output_15_14, output_14_925;
mixer gate_output_14_925(.a(output_15_925), .b(output_15_14), .y(output_14_925));
wire output_16_925, output_16_14, output_15_925;
mixer gate_output_15_925(.a(output_16_925), .b(output_16_14), .y(output_15_925));
wire output_1_926, output_1_15, output_0_926;
mixer gate_output_0_926(.a(output_1_926), .b(output_1_15), .y(output_0_926));
wire output_2_926, output_2_15, output_1_926;
mixer gate_output_1_926(.a(output_2_926), .b(output_2_15), .y(output_1_926));
wire output_3_926, output_3_15, output_2_926;
mixer gate_output_2_926(.a(output_3_926), .b(output_3_15), .y(output_2_926));
wire output_4_926, output_4_15, output_3_926;
mixer gate_output_3_926(.a(output_4_926), .b(output_4_15), .y(output_3_926));
wire output_5_926, output_5_15, output_4_926;
mixer gate_output_4_926(.a(output_5_926), .b(output_5_15), .y(output_4_926));
wire output_6_926, output_6_15, output_5_926;
mixer gate_output_5_926(.a(output_6_926), .b(output_6_15), .y(output_5_926));
wire output_7_926, output_7_15, output_6_926;
mixer gate_output_6_926(.a(output_7_926), .b(output_7_15), .y(output_6_926));
wire output_8_926, output_8_15, output_7_926;
mixer gate_output_7_926(.a(output_8_926), .b(output_8_15), .y(output_7_926));
wire output_9_926, output_9_15, output_8_926;
mixer gate_output_8_926(.a(output_9_926), .b(output_9_15), .y(output_8_926));
wire output_10_926, output_10_15, output_9_926;
mixer gate_output_9_926(.a(output_10_926), .b(output_10_15), .y(output_9_926));
wire output_11_926, output_11_15, output_10_926;
mixer gate_output_10_926(.a(output_11_926), .b(output_11_15), .y(output_10_926));
wire output_12_926, output_12_15, output_11_926;
mixer gate_output_11_926(.a(output_12_926), .b(output_12_15), .y(output_11_926));
wire output_13_926, output_13_15, output_12_926;
mixer gate_output_12_926(.a(output_13_926), .b(output_13_15), .y(output_12_926));
wire output_14_926, output_14_15, output_13_926;
mixer gate_output_13_926(.a(output_14_926), .b(output_14_15), .y(output_13_926));
wire output_15_926, output_15_15, output_14_926;
mixer gate_output_14_926(.a(output_15_926), .b(output_15_15), .y(output_14_926));
wire output_16_926, output_16_15, output_15_926;
mixer gate_output_15_926(.a(output_16_926), .b(output_16_15), .y(output_15_926));
wire output_1_927, output_1_0, output_0_927;
mixer gate_output_0_927(.a(output_1_927), .b(output_1_0), .y(output_0_927));
wire output_2_927, output_2_0, output_1_927;
mixer gate_output_1_927(.a(output_2_927), .b(output_2_0), .y(output_1_927));
wire output_3_927, output_3_0, output_2_927;
mixer gate_output_2_927(.a(output_3_927), .b(output_3_0), .y(output_2_927));
wire output_4_927, output_4_0, output_3_927;
mixer gate_output_3_927(.a(output_4_927), .b(output_4_0), .y(output_3_927));
wire output_5_927, output_5_0, output_4_927;
mixer gate_output_4_927(.a(output_5_927), .b(output_5_0), .y(output_4_927));
wire output_6_927, output_6_0, output_5_927;
mixer gate_output_5_927(.a(output_6_927), .b(output_6_0), .y(output_5_927));
wire output_7_927, output_7_0, output_6_927;
mixer gate_output_6_927(.a(output_7_927), .b(output_7_0), .y(output_6_927));
wire output_8_927, output_8_0, output_7_927;
mixer gate_output_7_927(.a(output_8_927), .b(output_8_0), .y(output_7_927));
wire output_9_927, output_9_0, output_8_927;
mixer gate_output_8_927(.a(output_9_927), .b(output_9_0), .y(output_8_927));
wire output_10_927, output_10_0, output_9_927;
mixer gate_output_9_927(.a(output_10_927), .b(output_10_0), .y(output_9_927));
wire output_11_927, output_11_0, output_10_927;
mixer gate_output_10_927(.a(output_11_927), .b(output_11_0), .y(output_10_927));
wire output_12_927, output_12_0, output_11_927;
mixer gate_output_11_927(.a(output_12_927), .b(output_12_0), .y(output_11_927));
wire output_13_927, output_13_0, output_12_927;
mixer gate_output_12_927(.a(output_13_927), .b(output_13_0), .y(output_12_927));
wire output_14_927, output_14_0, output_13_927;
mixer gate_output_13_927(.a(output_14_927), .b(output_14_0), .y(output_13_927));
wire output_15_927, output_15_0, output_14_927;
mixer gate_output_14_927(.a(output_15_927), .b(output_15_0), .y(output_14_927));
wire output_16_927, output_16_0, output_15_927;
mixer gate_output_15_927(.a(output_16_927), .b(output_16_0), .y(output_15_927));
wire output_1_928, output_1_1, output_0_928;
mixer gate_output_0_928(.a(output_1_928), .b(output_1_1), .y(output_0_928));
wire output_2_928, output_2_1, output_1_928;
mixer gate_output_1_928(.a(output_2_928), .b(output_2_1), .y(output_1_928));
wire output_3_928, output_3_1, output_2_928;
mixer gate_output_2_928(.a(output_3_928), .b(output_3_1), .y(output_2_928));
wire output_4_928, output_4_1, output_3_928;
mixer gate_output_3_928(.a(output_4_928), .b(output_4_1), .y(output_3_928));
wire output_5_928, output_5_1, output_4_928;
mixer gate_output_4_928(.a(output_5_928), .b(output_5_1), .y(output_4_928));
wire output_6_928, output_6_1, output_5_928;
mixer gate_output_5_928(.a(output_6_928), .b(output_6_1), .y(output_5_928));
wire output_7_928, output_7_1, output_6_928;
mixer gate_output_6_928(.a(output_7_928), .b(output_7_1), .y(output_6_928));
wire output_8_928, output_8_1, output_7_928;
mixer gate_output_7_928(.a(output_8_928), .b(output_8_1), .y(output_7_928));
wire output_9_928, output_9_1, output_8_928;
mixer gate_output_8_928(.a(output_9_928), .b(output_9_1), .y(output_8_928));
wire output_10_928, output_10_1, output_9_928;
mixer gate_output_9_928(.a(output_10_928), .b(output_10_1), .y(output_9_928));
wire output_11_928, output_11_1, output_10_928;
mixer gate_output_10_928(.a(output_11_928), .b(output_11_1), .y(output_10_928));
wire output_12_928, output_12_1, output_11_928;
mixer gate_output_11_928(.a(output_12_928), .b(output_12_1), .y(output_11_928));
wire output_13_928, output_13_1, output_12_928;
mixer gate_output_12_928(.a(output_13_928), .b(output_13_1), .y(output_12_928));
wire output_14_928, output_14_1, output_13_928;
mixer gate_output_13_928(.a(output_14_928), .b(output_14_1), .y(output_13_928));
wire output_15_928, output_15_1, output_14_928;
mixer gate_output_14_928(.a(output_15_928), .b(output_15_1), .y(output_14_928));
wire output_16_928, output_16_1, output_15_928;
mixer gate_output_15_928(.a(output_16_928), .b(output_16_1), .y(output_15_928));
wire output_1_929, output_1_2, output_0_929;
mixer gate_output_0_929(.a(output_1_929), .b(output_1_2), .y(output_0_929));
wire output_2_929, output_2_2, output_1_929;
mixer gate_output_1_929(.a(output_2_929), .b(output_2_2), .y(output_1_929));
wire output_3_929, output_3_2, output_2_929;
mixer gate_output_2_929(.a(output_3_929), .b(output_3_2), .y(output_2_929));
wire output_4_929, output_4_2, output_3_929;
mixer gate_output_3_929(.a(output_4_929), .b(output_4_2), .y(output_3_929));
wire output_5_929, output_5_2, output_4_929;
mixer gate_output_4_929(.a(output_5_929), .b(output_5_2), .y(output_4_929));
wire output_6_929, output_6_2, output_5_929;
mixer gate_output_5_929(.a(output_6_929), .b(output_6_2), .y(output_5_929));
wire output_7_929, output_7_2, output_6_929;
mixer gate_output_6_929(.a(output_7_929), .b(output_7_2), .y(output_6_929));
wire output_8_929, output_8_2, output_7_929;
mixer gate_output_7_929(.a(output_8_929), .b(output_8_2), .y(output_7_929));
wire output_9_929, output_9_2, output_8_929;
mixer gate_output_8_929(.a(output_9_929), .b(output_9_2), .y(output_8_929));
wire output_10_929, output_10_2, output_9_929;
mixer gate_output_9_929(.a(output_10_929), .b(output_10_2), .y(output_9_929));
wire output_11_929, output_11_2, output_10_929;
mixer gate_output_10_929(.a(output_11_929), .b(output_11_2), .y(output_10_929));
wire output_12_929, output_12_2, output_11_929;
mixer gate_output_11_929(.a(output_12_929), .b(output_12_2), .y(output_11_929));
wire output_13_929, output_13_2, output_12_929;
mixer gate_output_12_929(.a(output_13_929), .b(output_13_2), .y(output_12_929));
wire output_14_929, output_14_2, output_13_929;
mixer gate_output_13_929(.a(output_14_929), .b(output_14_2), .y(output_13_929));
wire output_15_929, output_15_2, output_14_929;
mixer gate_output_14_929(.a(output_15_929), .b(output_15_2), .y(output_14_929));
wire output_16_929, output_16_2, output_15_929;
mixer gate_output_15_929(.a(output_16_929), .b(output_16_2), .y(output_15_929));
wire output_1_930, output_1_3, output_0_930;
mixer gate_output_0_930(.a(output_1_930), .b(output_1_3), .y(output_0_930));
wire output_2_930, output_2_3, output_1_930;
mixer gate_output_1_930(.a(output_2_930), .b(output_2_3), .y(output_1_930));
wire output_3_930, output_3_3, output_2_930;
mixer gate_output_2_930(.a(output_3_930), .b(output_3_3), .y(output_2_930));
wire output_4_930, output_4_3, output_3_930;
mixer gate_output_3_930(.a(output_4_930), .b(output_4_3), .y(output_3_930));
wire output_5_930, output_5_3, output_4_930;
mixer gate_output_4_930(.a(output_5_930), .b(output_5_3), .y(output_4_930));
wire output_6_930, output_6_3, output_5_930;
mixer gate_output_5_930(.a(output_6_930), .b(output_6_3), .y(output_5_930));
wire output_7_930, output_7_3, output_6_930;
mixer gate_output_6_930(.a(output_7_930), .b(output_7_3), .y(output_6_930));
wire output_8_930, output_8_3, output_7_930;
mixer gate_output_7_930(.a(output_8_930), .b(output_8_3), .y(output_7_930));
wire output_9_930, output_9_3, output_8_930;
mixer gate_output_8_930(.a(output_9_930), .b(output_9_3), .y(output_8_930));
wire output_10_930, output_10_3, output_9_930;
mixer gate_output_9_930(.a(output_10_930), .b(output_10_3), .y(output_9_930));
wire output_11_930, output_11_3, output_10_930;
mixer gate_output_10_930(.a(output_11_930), .b(output_11_3), .y(output_10_930));
wire output_12_930, output_12_3, output_11_930;
mixer gate_output_11_930(.a(output_12_930), .b(output_12_3), .y(output_11_930));
wire output_13_930, output_13_3, output_12_930;
mixer gate_output_12_930(.a(output_13_930), .b(output_13_3), .y(output_12_930));
wire output_14_930, output_14_3, output_13_930;
mixer gate_output_13_930(.a(output_14_930), .b(output_14_3), .y(output_13_930));
wire output_15_930, output_15_3, output_14_930;
mixer gate_output_14_930(.a(output_15_930), .b(output_15_3), .y(output_14_930));
wire output_16_930, output_16_3, output_15_930;
mixer gate_output_15_930(.a(output_16_930), .b(output_16_3), .y(output_15_930));
wire output_1_931, output_1_4, output_0_931;
mixer gate_output_0_931(.a(output_1_931), .b(output_1_4), .y(output_0_931));
wire output_2_931, output_2_4, output_1_931;
mixer gate_output_1_931(.a(output_2_931), .b(output_2_4), .y(output_1_931));
wire output_3_931, output_3_4, output_2_931;
mixer gate_output_2_931(.a(output_3_931), .b(output_3_4), .y(output_2_931));
wire output_4_931, output_4_4, output_3_931;
mixer gate_output_3_931(.a(output_4_931), .b(output_4_4), .y(output_3_931));
wire output_5_931, output_5_4, output_4_931;
mixer gate_output_4_931(.a(output_5_931), .b(output_5_4), .y(output_4_931));
wire output_6_931, output_6_4, output_5_931;
mixer gate_output_5_931(.a(output_6_931), .b(output_6_4), .y(output_5_931));
wire output_7_931, output_7_4, output_6_931;
mixer gate_output_6_931(.a(output_7_931), .b(output_7_4), .y(output_6_931));
wire output_8_931, output_8_4, output_7_931;
mixer gate_output_7_931(.a(output_8_931), .b(output_8_4), .y(output_7_931));
wire output_9_931, output_9_4, output_8_931;
mixer gate_output_8_931(.a(output_9_931), .b(output_9_4), .y(output_8_931));
wire output_10_931, output_10_4, output_9_931;
mixer gate_output_9_931(.a(output_10_931), .b(output_10_4), .y(output_9_931));
wire output_11_931, output_11_4, output_10_931;
mixer gate_output_10_931(.a(output_11_931), .b(output_11_4), .y(output_10_931));
wire output_12_931, output_12_4, output_11_931;
mixer gate_output_11_931(.a(output_12_931), .b(output_12_4), .y(output_11_931));
wire output_13_931, output_13_4, output_12_931;
mixer gate_output_12_931(.a(output_13_931), .b(output_13_4), .y(output_12_931));
wire output_14_931, output_14_4, output_13_931;
mixer gate_output_13_931(.a(output_14_931), .b(output_14_4), .y(output_13_931));
wire output_15_931, output_15_4, output_14_931;
mixer gate_output_14_931(.a(output_15_931), .b(output_15_4), .y(output_14_931));
wire output_16_931, output_16_4, output_15_931;
mixer gate_output_15_931(.a(output_16_931), .b(output_16_4), .y(output_15_931));
wire output_1_932, output_1_5, output_0_932;
mixer gate_output_0_932(.a(output_1_932), .b(output_1_5), .y(output_0_932));
wire output_2_932, output_2_5, output_1_932;
mixer gate_output_1_932(.a(output_2_932), .b(output_2_5), .y(output_1_932));
wire output_3_932, output_3_5, output_2_932;
mixer gate_output_2_932(.a(output_3_932), .b(output_3_5), .y(output_2_932));
wire output_4_932, output_4_5, output_3_932;
mixer gate_output_3_932(.a(output_4_932), .b(output_4_5), .y(output_3_932));
wire output_5_932, output_5_5, output_4_932;
mixer gate_output_4_932(.a(output_5_932), .b(output_5_5), .y(output_4_932));
wire output_6_932, output_6_5, output_5_932;
mixer gate_output_5_932(.a(output_6_932), .b(output_6_5), .y(output_5_932));
wire output_7_932, output_7_5, output_6_932;
mixer gate_output_6_932(.a(output_7_932), .b(output_7_5), .y(output_6_932));
wire output_8_932, output_8_5, output_7_932;
mixer gate_output_7_932(.a(output_8_932), .b(output_8_5), .y(output_7_932));
wire output_9_932, output_9_5, output_8_932;
mixer gate_output_8_932(.a(output_9_932), .b(output_9_5), .y(output_8_932));
wire output_10_932, output_10_5, output_9_932;
mixer gate_output_9_932(.a(output_10_932), .b(output_10_5), .y(output_9_932));
wire output_11_932, output_11_5, output_10_932;
mixer gate_output_10_932(.a(output_11_932), .b(output_11_5), .y(output_10_932));
wire output_12_932, output_12_5, output_11_932;
mixer gate_output_11_932(.a(output_12_932), .b(output_12_5), .y(output_11_932));
wire output_13_932, output_13_5, output_12_932;
mixer gate_output_12_932(.a(output_13_932), .b(output_13_5), .y(output_12_932));
wire output_14_932, output_14_5, output_13_932;
mixer gate_output_13_932(.a(output_14_932), .b(output_14_5), .y(output_13_932));
wire output_15_932, output_15_5, output_14_932;
mixer gate_output_14_932(.a(output_15_932), .b(output_15_5), .y(output_14_932));
wire output_16_932, output_16_5, output_15_932;
mixer gate_output_15_932(.a(output_16_932), .b(output_16_5), .y(output_15_932));
wire output_1_933, output_1_6, output_0_933;
mixer gate_output_0_933(.a(output_1_933), .b(output_1_6), .y(output_0_933));
wire output_2_933, output_2_6, output_1_933;
mixer gate_output_1_933(.a(output_2_933), .b(output_2_6), .y(output_1_933));
wire output_3_933, output_3_6, output_2_933;
mixer gate_output_2_933(.a(output_3_933), .b(output_3_6), .y(output_2_933));
wire output_4_933, output_4_6, output_3_933;
mixer gate_output_3_933(.a(output_4_933), .b(output_4_6), .y(output_3_933));
wire output_5_933, output_5_6, output_4_933;
mixer gate_output_4_933(.a(output_5_933), .b(output_5_6), .y(output_4_933));
wire output_6_933, output_6_6, output_5_933;
mixer gate_output_5_933(.a(output_6_933), .b(output_6_6), .y(output_5_933));
wire output_7_933, output_7_6, output_6_933;
mixer gate_output_6_933(.a(output_7_933), .b(output_7_6), .y(output_6_933));
wire output_8_933, output_8_6, output_7_933;
mixer gate_output_7_933(.a(output_8_933), .b(output_8_6), .y(output_7_933));
wire output_9_933, output_9_6, output_8_933;
mixer gate_output_8_933(.a(output_9_933), .b(output_9_6), .y(output_8_933));
wire output_10_933, output_10_6, output_9_933;
mixer gate_output_9_933(.a(output_10_933), .b(output_10_6), .y(output_9_933));
wire output_11_933, output_11_6, output_10_933;
mixer gate_output_10_933(.a(output_11_933), .b(output_11_6), .y(output_10_933));
wire output_12_933, output_12_6, output_11_933;
mixer gate_output_11_933(.a(output_12_933), .b(output_12_6), .y(output_11_933));
wire output_13_933, output_13_6, output_12_933;
mixer gate_output_12_933(.a(output_13_933), .b(output_13_6), .y(output_12_933));
wire output_14_933, output_14_6, output_13_933;
mixer gate_output_13_933(.a(output_14_933), .b(output_14_6), .y(output_13_933));
wire output_15_933, output_15_6, output_14_933;
mixer gate_output_14_933(.a(output_15_933), .b(output_15_6), .y(output_14_933));
wire output_16_933, output_16_6, output_15_933;
mixer gate_output_15_933(.a(output_16_933), .b(output_16_6), .y(output_15_933));
wire output_1_934, output_1_7, output_0_934;
mixer gate_output_0_934(.a(output_1_934), .b(output_1_7), .y(output_0_934));
wire output_2_934, output_2_7, output_1_934;
mixer gate_output_1_934(.a(output_2_934), .b(output_2_7), .y(output_1_934));
wire output_3_934, output_3_7, output_2_934;
mixer gate_output_2_934(.a(output_3_934), .b(output_3_7), .y(output_2_934));
wire output_4_934, output_4_7, output_3_934;
mixer gate_output_3_934(.a(output_4_934), .b(output_4_7), .y(output_3_934));
wire output_5_934, output_5_7, output_4_934;
mixer gate_output_4_934(.a(output_5_934), .b(output_5_7), .y(output_4_934));
wire output_6_934, output_6_7, output_5_934;
mixer gate_output_5_934(.a(output_6_934), .b(output_6_7), .y(output_5_934));
wire output_7_934, output_7_7, output_6_934;
mixer gate_output_6_934(.a(output_7_934), .b(output_7_7), .y(output_6_934));
wire output_8_934, output_8_7, output_7_934;
mixer gate_output_7_934(.a(output_8_934), .b(output_8_7), .y(output_7_934));
wire output_9_934, output_9_7, output_8_934;
mixer gate_output_8_934(.a(output_9_934), .b(output_9_7), .y(output_8_934));
wire output_10_934, output_10_7, output_9_934;
mixer gate_output_9_934(.a(output_10_934), .b(output_10_7), .y(output_9_934));
wire output_11_934, output_11_7, output_10_934;
mixer gate_output_10_934(.a(output_11_934), .b(output_11_7), .y(output_10_934));
wire output_12_934, output_12_7, output_11_934;
mixer gate_output_11_934(.a(output_12_934), .b(output_12_7), .y(output_11_934));
wire output_13_934, output_13_7, output_12_934;
mixer gate_output_12_934(.a(output_13_934), .b(output_13_7), .y(output_12_934));
wire output_14_934, output_14_7, output_13_934;
mixer gate_output_13_934(.a(output_14_934), .b(output_14_7), .y(output_13_934));
wire output_15_934, output_15_7, output_14_934;
mixer gate_output_14_934(.a(output_15_934), .b(output_15_7), .y(output_14_934));
wire output_16_934, output_16_7, output_15_934;
mixer gate_output_15_934(.a(output_16_934), .b(output_16_7), .y(output_15_934));
wire output_1_935, output_1_8, output_0_935;
mixer gate_output_0_935(.a(output_1_935), .b(output_1_8), .y(output_0_935));
wire output_2_935, output_2_8, output_1_935;
mixer gate_output_1_935(.a(output_2_935), .b(output_2_8), .y(output_1_935));
wire output_3_935, output_3_8, output_2_935;
mixer gate_output_2_935(.a(output_3_935), .b(output_3_8), .y(output_2_935));
wire output_4_935, output_4_8, output_3_935;
mixer gate_output_3_935(.a(output_4_935), .b(output_4_8), .y(output_3_935));
wire output_5_935, output_5_8, output_4_935;
mixer gate_output_4_935(.a(output_5_935), .b(output_5_8), .y(output_4_935));
wire output_6_935, output_6_8, output_5_935;
mixer gate_output_5_935(.a(output_6_935), .b(output_6_8), .y(output_5_935));
wire output_7_935, output_7_8, output_6_935;
mixer gate_output_6_935(.a(output_7_935), .b(output_7_8), .y(output_6_935));
wire output_8_935, output_8_8, output_7_935;
mixer gate_output_7_935(.a(output_8_935), .b(output_8_8), .y(output_7_935));
wire output_9_935, output_9_8, output_8_935;
mixer gate_output_8_935(.a(output_9_935), .b(output_9_8), .y(output_8_935));
wire output_10_935, output_10_8, output_9_935;
mixer gate_output_9_935(.a(output_10_935), .b(output_10_8), .y(output_9_935));
wire output_11_935, output_11_8, output_10_935;
mixer gate_output_10_935(.a(output_11_935), .b(output_11_8), .y(output_10_935));
wire output_12_935, output_12_8, output_11_935;
mixer gate_output_11_935(.a(output_12_935), .b(output_12_8), .y(output_11_935));
wire output_13_935, output_13_8, output_12_935;
mixer gate_output_12_935(.a(output_13_935), .b(output_13_8), .y(output_12_935));
wire output_14_935, output_14_8, output_13_935;
mixer gate_output_13_935(.a(output_14_935), .b(output_14_8), .y(output_13_935));
wire output_15_935, output_15_8, output_14_935;
mixer gate_output_14_935(.a(output_15_935), .b(output_15_8), .y(output_14_935));
wire output_16_935, output_16_8, output_15_935;
mixer gate_output_15_935(.a(output_16_935), .b(output_16_8), .y(output_15_935));
wire output_1_936, output_1_9, output_0_936;
mixer gate_output_0_936(.a(output_1_936), .b(output_1_9), .y(output_0_936));
wire output_2_936, output_2_9, output_1_936;
mixer gate_output_1_936(.a(output_2_936), .b(output_2_9), .y(output_1_936));
wire output_3_936, output_3_9, output_2_936;
mixer gate_output_2_936(.a(output_3_936), .b(output_3_9), .y(output_2_936));
wire output_4_936, output_4_9, output_3_936;
mixer gate_output_3_936(.a(output_4_936), .b(output_4_9), .y(output_3_936));
wire output_5_936, output_5_9, output_4_936;
mixer gate_output_4_936(.a(output_5_936), .b(output_5_9), .y(output_4_936));
wire output_6_936, output_6_9, output_5_936;
mixer gate_output_5_936(.a(output_6_936), .b(output_6_9), .y(output_5_936));
wire output_7_936, output_7_9, output_6_936;
mixer gate_output_6_936(.a(output_7_936), .b(output_7_9), .y(output_6_936));
wire output_8_936, output_8_9, output_7_936;
mixer gate_output_7_936(.a(output_8_936), .b(output_8_9), .y(output_7_936));
wire output_9_936, output_9_9, output_8_936;
mixer gate_output_8_936(.a(output_9_936), .b(output_9_9), .y(output_8_936));
wire output_10_936, output_10_9, output_9_936;
mixer gate_output_9_936(.a(output_10_936), .b(output_10_9), .y(output_9_936));
wire output_11_936, output_11_9, output_10_936;
mixer gate_output_10_936(.a(output_11_936), .b(output_11_9), .y(output_10_936));
wire output_12_936, output_12_9, output_11_936;
mixer gate_output_11_936(.a(output_12_936), .b(output_12_9), .y(output_11_936));
wire output_13_936, output_13_9, output_12_936;
mixer gate_output_12_936(.a(output_13_936), .b(output_13_9), .y(output_12_936));
wire output_14_936, output_14_9, output_13_936;
mixer gate_output_13_936(.a(output_14_936), .b(output_14_9), .y(output_13_936));
wire output_15_936, output_15_9, output_14_936;
mixer gate_output_14_936(.a(output_15_936), .b(output_15_9), .y(output_14_936));
wire output_16_936, output_16_9, output_15_936;
mixer gate_output_15_936(.a(output_16_936), .b(output_16_9), .y(output_15_936));
wire output_1_937, output_1_10, output_0_937;
mixer gate_output_0_937(.a(output_1_937), .b(output_1_10), .y(output_0_937));
wire output_2_937, output_2_10, output_1_937;
mixer gate_output_1_937(.a(output_2_937), .b(output_2_10), .y(output_1_937));
wire output_3_937, output_3_10, output_2_937;
mixer gate_output_2_937(.a(output_3_937), .b(output_3_10), .y(output_2_937));
wire output_4_937, output_4_10, output_3_937;
mixer gate_output_3_937(.a(output_4_937), .b(output_4_10), .y(output_3_937));
wire output_5_937, output_5_10, output_4_937;
mixer gate_output_4_937(.a(output_5_937), .b(output_5_10), .y(output_4_937));
wire output_6_937, output_6_10, output_5_937;
mixer gate_output_5_937(.a(output_6_937), .b(output_6_10), .y(output_5_937));
wire output_7_937, output_7_10, output_6_937;
mixer gate_output_6_937(.a(output_7_937), .b(output_7_10), .y(output_6_937));
wire output_8_937, output_8_10, output_7_937;
mixer gate_output_7_937(.a(output_8_937), .b(output_8_10), .y(output_7_937));
wire output_9_937, output_9_10, output_8_937;
mixer gate_output_8_937(.a(output_9_937), .b(output_9_10), .y(output_8_937));
wire output_10_937, output_10_10, output_9_937;
mixer gate_output_9_937(.a(output_10_937), .b(output_10_10), .y(output_9_937));
wire output_11_937, output_11_10, output_10_937;
mixer gate_output_10_937(.a(output_11_937), .b(output_11_10), .y(output_10_937));
wire output_12_937, output_12_10, output_11_937;
mixer gate_output_11_937(.a(output_12_937), .b(output_12_10), .y(output_11_937));
wire output_13_937, output_13_10, output_12_937;
mixer gate_output_12_937(.a(output_13_937), .b(output_13_10), .y(output_12_937));
wire output_14_937, output_14_10, output_13_937;
mixer gate_output_13_937(.a(output_14_937), .b(output_14_10), .y(output_13_937));
wire output_15_937, output_15_10, output_14_937;
mixer gate_output_14_937(.a(output_15_937), .b(output_15_10), .y(output_14_937));
wire output_16_937, output_16_10, output_15_937;
mixer gate_output_15_937(.a(output_16_937), .b(output_16_10), .y(output_15_937));
wire output_1_938, output_1_11, output_0_938;
mixer gate_output_0_938(.a(output_1_938), .b(output_1_11), .y(output_0_938));
wire output_2_938, output_2_11, output_1_938;
mixer gate_output_1_938(.a(output_2_938), .b(output_2_11), .y(output_1_938));
wire output_3_938, output_3_11, output_2_938;
mixer gate_output_2_938(.a(output_3_938), .b(output_3_11), .y(output_2_938));
wire output_4_938, output_4_11, output_3_938;
mixer gate_output_3_938(.a(output_4_938), .b(output_4_11), .y(output_3_938));
wire output_5_938, output_5_11, output_4_938;
mixer gate_output_4_938(.a(output_5_938), .b(output_5_11), .y(output_4_938));
wire output_6_938, output_6_11, output_5_938;
mixer gate_output_5_938(.a(output_6_938), .b(output_6_11), .y(output_5_938));
wire output_7_938, output_7_11, output_6_938;
mixer gate_output_6_938(.a(output_7_938), .b(output_7_11), .y(output_6_938));
wire output_8_938, output_8_11, output_7_938;
mixer gate_output_7_938(.a(output_8_938), .b(output_8_11), .y(output_7_938));
wire output_9_938, output_9_11, output_8_938;
mixer gate_output_8_938(.a(output_9_938), .b(output_9_11), .y(output_8_938));
wire output_10_938, output_10_11, output_9_938;
mixer gate_output_9_938(.a(output_10_938), .b(output_10_11), .y(output_9_938));
wire output_11_938, output_11_11, output_10_938;
mixer gate_output_10_938(.a(output_11_938), .b(output_11_11), .y(output_10_938));
wire output_12_938, output_12_11, output_11_938;
mixer gate_output_11_938(.a(output_12_938), .b(output_12_11), .y(output_11_938));
wire output_13_938, output_13_11, output_12_938;
mixer gate_output_12_938(.a(output_13_938), .b(output_13_11), .y(output_12_938));
wire output_14_938, output_14_11, output_13_938;
mixer gate_output_13_938(.a(output_14_938), .b(output_14_11), .y(output_13_938));
wire output_15_938, output_15_11, output_14_938;
mixer gate_output_14_938(.a(output_15_938), .b(output_15_11), .y(output_14_938));
wire output_16_938, output_16_11, output_15_938;
mixer gate_output_15_938(.a(output_16_938), .b(output_16_11), .y(output_15_938));
wire output_1_939, output_1_12, output_0_939;
mixer gate_output_0_939(.a(output_1_939), .b(output_1_12), .y(output_0_939));
wire output_2_939, output_2_12, output_1_939;
mixer gate_output_1_939(.a(output_2_939), .b(output_2_12), .y(output_1_939));
wire output_3_939, output_3_12, output_2_939;
mixer gate_output_2_939(.a(output_3_939), .b(output_3_12), .y(output_2_939));
wire output_4_939, output_4_12, output_3_939;
mixer gate_output_3_939(.a(output_4_939), .b(output_4_12), .y(output_3_939));
wire output_5_939, output_5_12, output_4_939;
mixer gate_output_4_939(.a(output_5_939), .b(output_5_12), .y(output_4_939));
wire output_6_939, output_6_12, output_5_939;
mixer gate_output_5_939(.a(output_6_939), .b(output_6_12), .y(output_5_939));
wire output_7_939, output_7_12, output_6_939;
mixer gate_output_6_939(.a(output_7_939), .b(output_7_12), .y(output_6_939));
wire output_8_939, output_8_12, output_7_939;
mixer gate_output_7_939(.a(output_8_939), .b(output_8_12), .y(output_7_939));
wire output_9_939, output_9_12, output_8_939;
mixer gate_output_8_939(.a(output_9_939), .b(output_9_12), .y(output_8_939));
wire output_10_939, output_10_12, output_9_939;
mixer gate_output_9_939(.a(output_10_939), .b(output_10_12), .y(output_9_939));
wire output_11_939, output_11_12, output_10_939;
mixer gate_output_10_939(.a(output_11_939), .b(output_11_12), .y(output_10_939));
wire output_12_939, output_12_12, output_11_939;
mixer gate_output_11_939(.a(output_12_939), .b(output_12_12), .y(output_11_939));
wire output_13_939, output_13_12, output_12_939;
mixer gate_output_12_939(.a(output_13_939), .b(output_13_12), .y(output_12_939));
wire output_14_939, output_14_12, output_13_939;
mixer gate_output_13_939(.a(output_14_939), .b(output_14_12), .y(output_13_939));
wire output_15_939, output_15_12, output_14_939;
mixer gate_output_14_939(.a(output_15_939), .b(output_15_12), .y(output_14_939));
wire output_16_939, output_16_12, output_15_939;
mixer gate_output_15_939(.a(output_16_939), .b(output_16_12), .y(output_15_939));
wire output_1_940, output_1_13, output_0_940;
mixer gate_output_0_940(.a(output_1_940), .b(output_1_13), .y(output_0_940));
wire output_2_940, output_2_13, output_1_940;
mixer gate_output_1_940(.a(output_2_940), .b(output_2_13), .y(output_1_940));
wire output_3_940, output_3_13, output_2_940;
mixer gate_output_2_940(.a(output_3_940), .b(output_3_13), .y(output_2_940));
wire output_4_940, output_4_13, output_3_940;
mixer gate_output_3_940(.a(output_4_940), .b(output_4_13), .y(output_3_940));
wire output_5_940, output_5_13, output_4_940;
mixer gate_output_4_940(.a(output_5_940), .b(output_5_13), .y(output_4_940));
wire output_6_940, output_6_13, output_5_940;
mixer gate_output_5_940(.a(output_6_940), .b(output_6_13), .y(output_5_940));
wire output_7_940, output_7_13, output_6_940;
mixer gate_output_6_940(.a(output_7_940), .b(output_7_13), .y(output_6_940));
wire output_8_940, output_8_13, output_7_940;
mixer gate_output_7_940(.a(output_8_940), .b(output_8_13), .y(output_7_940));
wire output_9_940, output_9_13, output_8_940;
mixer gate_output_8_940(.a(output_9_940), .b(output_9_13), .y(output_8_940));
wire output_10_940, output_10_13, output_9_940;
mixer gate_output_9_940(.a(output_10_940), .b(output_10_13), .y(output_9_940));
wire output_11_940, output_11_13, output_10_940;
mixer gate_output_10_940(.a(output_11_940), .b(output_11_13), .y(output_10_940));
wire output_12_940, output_12_13, output_11_940;
mixer gate_output_11_940(.a(output_12_940), .b(output_12_13), .y(output_11_940));
wire output_13_940, output_13_13, output_12_940;
mixer gate_output_12_940(.a(output_13_940), .b(output_13_13), .y(output_12_940));
wire output_14_940, output_14_13, output_13_940;
mixer gate_output_13_940(.a(output_14_940), .b(output_14_13), .y(output_13_940));
wire output_15_940, output_15_13, output_14_940;
mixer gate_output_14_940(.a(output_15_940), .b(output_15_13), .y(output_14_940));
wire output_16_940, output_16_13, output_15_940;
mixer gate_output_15_940(.a(output_16_940), .b(output_16_13), .y(output_15_940));
wire output_1_941, output_1_14, output_0_941;
mixer gate_output_0_941(.a(output_1_941), .b(output_1_14), .y(output_0_941));
wire output_2_941, output_2_14, output_1_941;
mixer gate_output_1_941(.a(output_2_941), .b(output_2_14), .y(output_1_941));
wire output_3_941, output_3_14, output_2_941;
mixer gate_output_2_941(.a(output_3_941), .b(output_3_14), .y(output_2_941));
wire output_4_941, output_4_14, output_3_941;
mixer gate_output_3_941(.a(output_4_941), .b(output_4_14), .y(output_3_941));
wire output_5_941, output_5_14, output_4_941;
mixer gate_output_4_941(.a(output_5_941), .b(output_5_14), .y(output_4_941));
wire output_6_941, output_6_14, output_5_941;
mixer gate_output_5_941(.a(output_6_941), .b(output_6_14), .y(output_5_941));
wire output_7_941, output_7_14, output_6_941;
mixer gate_output_6_941(.a(output_7_941), .b(output_7_14), .y(output_6_941));
wire output_8_941, output_8_14, output_7_941;
mixer gate_output_7_941(.a(output_8_941), .b(output_8_14), .y(output_7_941));
wire output_9_941, output_9_14, output_8_941;
mixer gate_output_8_941(.a(output_9_941), .b(output_9_14), .y(output_8_941));
wire output_10_941, output_10_14, output_9_941;
mixer gate_output_9_941(.a(output_10_941), .b(output_10_14), .y(output_9_941));
wire output_11_941, output_11_14, output_10_941;
mixer gate_output_10_941(.a(output_11_941), .b(output_11_14), .y(output_10_941));
wire output_12_941, output_12_14, output_11_941;
mixer gate_output_11_941(.a(output_12_941), .b(output_12_14), .y(output_11_941));
wire output_13_941, output_13_14, output_12_941;
mixer gate_output_12_941(.a(output_13_941), .b(output_13_14), .y(output_12_941));
wire output_14_941, output_14_14, output_13_941;
mixer gate_output_13_941(.a(output_14_941), .b(output_14_14), .y(output_13_941));
wire output_15_941, output_15_14, output_14_941;
mixer gate_output_14_941(.a(output_15_941), .b(output_15_14), .y(output_14_941));
wire output_16_941, output_16_14, output_15_941;
mixer gate_output_15_941(.a(output_16_941), .b(output_16_14), .y(output_15_941));
wire output_1_942, output_1_15, output_0_942;
mixer gate_output_0_942(.a(output_1_942), .b(output_1_15), .y(output_0_942));
wire output_2_942, output_2_15, output_1_942;
mixer gate_output_1_942(.a(output_2_942), .b(output_2_15), .y(output_1_942));
wire output_3_942, output_3_15, output_2_942;
mixer gate_output_2_942(.a(output_3_942), .b(output_3_15), .y(output_2_942));
wire output_4_942, output_4_15, output_3_942;
mixer gate_output_3_942(.a(output_4_942), .b(output_4_15), .y(output_3_942));
wire output_5_942, output_5_15, output_4_942;
mixer gate_output_4_942(.a(output_5_942), .b(output_5_15), .y(output_4_942));
wire output_6_942, output_6_15, output_5_942;
mixer gate_output_5_942(.a(output_6_942), .b(output_6_15), .y(output_5_942));
wire output_7_942, output_7_15, output_6_942;
mixer gate_output_6_942(.a(output_7_942), .b(output_7_15), .y(output_6_942));
wire output_8_942, output_8_15, output_7_942;
mixer gate_output_7_942(.a(output_8_942), .b(output_8_15), .y(output_7_942));
wire output_9_942, output_9_15, output_8_942;
mixer gate_output_8_942(.a(output_9_942), .b(output_9_15), .y(output_8_942));
wire output_10_942, output_10_15, output_9_942;
mixer gate_output_9_942(.a(output_10_942), .b(output_10_15), .y(output_9_942));
wire output_11_942, output_11_15, output_10_942;
mixer gate_output_10_942(.a(output_11_942), .b(output_11_15), .y(output_10_942));
wire output_12_942, output_12_15, output_11_942;
mixer gate_output_11_942(.a(output_12_942), .b(output_12_15), .y(output_11_942));
wire output_13_942, output_13_15, output_12_942;
mixer gate_output_12_942(.a(output_13_942), .b(output_13_15), .y(output_12_942));
wire output_14_942, output_14_15, output_13_942;
mixer gate_output_13_942(.a(output_14_942), .b(output_14_15), .y(output_13_942));
wire output_15_942, output_15_15, output_14_942;
mixer gate_output_14_942(.a(output_15_942), .b(output_15_15), .y(output_14_942));
wire output_16_942, output_16_15, output_15_942;
mixer gate_output_15_942(.a(output_16_942), .b(output_16_15), .y(output_15_942));
wire output_1_943, output_1_0, output_0_943;
mixer gate_output_0_943(.a(output_1_943), .b(output_1_0), .y(output_0_943));
wire output_2_943, output_2_0, output_1_943;
mixer gate_output_1_943(.a(output_2_943), .b(output_2_0), .y(output_1_943));
wire output_3_943, output_3_0, output_2_943;
mixer gate_output_2_943(.a(output_3_943), .b(output_3_0), .y(output_2_943));
wire output_4_943, output_4_0, output_3_943;
mixer gate_output_3_943(.a(output_4_943), .b(output_4_0), .y(output_3_943));
wire output_5_943, output_5_0, output_4_943;
mixer gate_output_4_943(.a(output_5_943), .b(output_5_0), .y(output_4_943));
wire output_6_943, output_6_0, output_5_943;
mixer gate_output_5_943(.a(output_6_943), .b(output_6_0), .y(output_5_943));
wire output_7_943, output_7_0, output_6_943;
mixer gate_output_6_943(.a(output_7_943), .b(output_7_0), .y(output_6_943));
wire output_8_943, output_8_0, output_7_943;
mixer gate_output_7_943(.a(output_8_943), .b(output_8_0), .y(output_7_943));
wire output_9_943, output_9_0, output_8_943;
mixer gate_output_8_943(.a(output_9_943), .b(output_9_0), .y(output_8_943));
wire output_10_943, output_10_0, output_9_943;
mixer gate_output_9_943(.a(output_10_943), .b(output_10_0), .y(output_9_943));
wire output_11_943, output_11_0, output_10_943;
mixer gate_output_10_943(.a(output_11_943), .b(output_11_0), .y(output_10_943));
wire output_12_943, output_12_0, output_11_943;
mixer gate_output_11_943(.a(output_12_943), .b(output_12_0), .y(output_11_943));
wire output_13_943, output_13_0, output_12_943;
mixer gate_output_12_943(.a(output_13_943), .b(output_13_0), .y(output_12_943));
wire output_14_943, output_14_0, output_13_943;
mixer gate_output_13_943(.a(output_14_943), .b(output_14_0), .y(output_13_943));
wire output_15_943, output_15_0, output_14_943;
mixer gate_output_14_943(.a(output_15_943), .b(output_15_0), .y(output_14_943));
wire output_16_943, output_16_0, output_15_943;
mixer gate_output_15_943(.a(output_16_943), .b(output_16_0), .y(output_15_943));
wire output_1_944, output_1_1, output_0_944;
mixer gate_output_0_944(.a(output_1_944), .b(output_1_1), .y(output_0_944));
wire output_2_944, output_2_1, output_1_944;
mixer gate_output_1_944(.a(output_2_944), .b(output_2_1), .y(output_1_944));
wire output_3_944, output_3_1, output_2_944;
mixer gate_output_2_944(.a(output_3_944), .b(output_3_1), .y(output_2_944));
wire output_4_944, output_4_1, output_3_944;
mixer gate_output_3_944(.a(output_4_944), .b(output_4_1), .y(output_3_944));
wire output_5_944, output_5_1, output_4_944;
mixer gate_output_4_944(.a(output_5_944), .b(output_5_1), .y(output_4_944));
wire output_6_944, output_6_1, output_5_944;
mixer gate_output_5_944(.a(output_6_944), .b(output_6_1), .y(output_5_944));
wire output_7_944, output_7_1, output_6_944;
mixer gate_output_6_944(.a(output_7_944), .b(output_7_1), .y(output_6_944));
wire output_8_944, output_8_1, output_7_944;
mixer gate_output_7_944(.a(output_8_944), .b(output_8_1), .y(output_7_944));
wire output_9_944, output_9_1, output_8_944;
mixer gate_output_8_944(.a(output_9_944), .b(output_9_1), .y(output_8_944));
wire output_10_944, output_10_1, output_9_944;
mixer gate_output_9_944(.a(output_10_944), .b(output_10_1), .y(output_9_944));
wire output_11_944, output_11_1, output_10_944;
mixer gate_output_10_944(.a(output_11_944), .b(output_11_1), .y(output_10_944));
wire output_12_944, output_12_1, output_11_944;
mixer gate_output_11_944(.a(output_12_944), .b(output_12_1), .y(output_11_944));
wire output_13_944, output_13_1, output_12_944;
mixer gate_output_12_944(.a(output_13_944), .b(output_13_1), .y(output_12_944));
wire output_14_944, output_14_1, output_13_944;
mixer gate_output_13_944(.a(output_14_944), .b(output_14_1), .y(output_13_944));
wire output_15_944, output_15_1, output_14_944;
mixer gate_output_14_944(.a(output_15_944), .b(output_15_1), .y(output_14_944));
wire output_16_944, output_16_1, output_15_944;
mixer gate_output_15_944(.a(output_16_944), .b(output_16_1), .y(output_15_944));
wire output_1_945, output_1_2, output_0_945;
mixer gate_output_0_945(.a(output_1_945), .b(output_1_2), .y(output_0_945));
wire output_2_945, output_2_2, output_1_945;
mixer gate_output_1_945(.a(output_2_945), .b(output_2_2), .y(output_1_945));
wire output_3_945, output_3_2, output_2_945;
mixer gate_output_2_945(.a(output_3_945), .b(output_3_2), .y(output_2_945));
wire output_4_945, output_4_2, output_3_945;
mixer gate_output_3_945(.a(output_4_945), .b(output_4_2), .y(output_3_945));
wire output_5_945, output_5_2, output_4_945;
mixer gate_output_4_945(.a(output_5_945), .b(output_5_2), .y(output_4_945));
wire output_6_945, output_6_2, output_5_945;
mixer gate_output_5_945(.a(output_6_945), .b(output_6_2), .y(output_5_945));
wire output_7_945, output_7_2, output_6_945;
mixer gate_output_6_945(.a(output_7_945), .b(output_7_2), .y(output_6_945));
wire output_8_945, output_8_2, output_7_945;
mixer gate_output_7_945(.a(output_8_945), .b(output_8_2), .y(output_7_945));
wire output_9_945, output_9_2, output_8_945;
mixer gate_output_8_945(.a(output_9_945), .b(output_9_2), .y(output_8_945));
wire output_10_945, output_10_2, output_9_945;
mixer gate_output_9_945(.a(output_10_945), .b(output_10_2), .y(output_9_945));
wire output_11_945, output_11_2, output_10_945;
mixer gate_output_10_945(.a(output_11_945), .b(output_11_2), .y(output_10_945));
wire output_12_945, output_12_2, output_11_945;
mixer gate_output_11_945(.a(output_12_945), .b(output_12_2), .y(output_11_945));
wire output_13_945, output_13_2, output_12_945;
mixer gate_output_12_945(.a(output_13_945), .b(output_13_2), .y(output_12_945));
wire output_14_945, output_14_2, output_13_945;
mixer gate_output_13_945(.a(output_14_945), .b(output_14_2), .y(output_13_945));
wire output_15_945, output_15_2, output_14_945;
mixer gate_output_14_945(.a(output_15_945), .b(output_15_2), .y(output_14_945));
wire output_16_945, output_16_2, output_15_945;
mixer gate_output_15_945(.a(output_16_945), .b(output_16_2), .y(output_15_945));
wire output_1_946, output_1_3, output_0_946;
mixer gate_output_0_946(.a(output_1_946), .b(output_1_3), .y(output_0_946));
wire output_2_946, output_2_3, output_1_946;
mixer gate_output_1_946(.a(output_2_946), .b(output_2_3), .y(output_1_946));
wire output_3_946, output_3_3, output_2_946;
mixer gate_output_2_946(.a(output_3_946), .b(output_3_3), .y(output_2_946));
wire output_4_946, output_4_3, output_3_946;
mixer gate_output_3_946(.a(output_4_946), .b(output_4_3), .y(output_3_946));
wire output_5_946, output_5_3, output_4_946;
mixer gate_output_4_946(.a(output_5_946), .b(output_5_3), .y(output_4_946));
wire output_6_946, output_6_3, output_5_946;
mixer gate_output_5_946(.a(output_6_946), .b(output_6_3), .y(output_5_946));
wire output_7_946, output_7_3, output_6_946;
mixer gate_output_6_946(.a(output_7_946), .b(output_7_3), .y(output_6_946));
wire output_8_946, output_8_3, output_7_946;
mixer gate_output_7_946(.a(output_8_946), .b(output_8_3), .y(output_7_946));
wire output_9_946, output_9_3, output_8_946;
mixer gate_output_8_946(.a(output_9_946), .b(output_9_3), .y(output_8_946));
wire output_10_946, output_10_3, output_9_946;
mixer gate_output_9_946(.a(output_10_946), .b(output_10_3), .y(output_9_946));
wire output_11_946, output_11_3, output_10_946;
mixer gate_output_10_946(.a(output_11_946), .b(output_11_3), .y(output_10_946));
wire output_12_946, output_12_3, output_11_946;
mixer gate_output_11_946(.a(output_12_946), .b(output_12_3), .y(output_11_946));
wire output_13_946, output_13_3, output_12_946;
mixer gate_output_12_946(.a(output_13_946), .b(output_13_3), .y(output_12_946));
wire output_14_946, output_14_3, output_13_946;
mixer gate_output_13_946(.a(output_14_946), .b(output_14_3), .y(output_13_946));
wire output_15_946, output_15_3, output_14_946;
mixer gate_output_14_946(.a(output_15_946), .b(output_15_3), .y(output_14_946));
wire output_16_946, output_16_3, output_15_946;
mixer gate_output_15_946(.a(output_16_946), .b(output_16_3), .y(output_15_946));
wire output_1_947, output_1_4, output_0_947;
mixer gate_output_0_947(.a(output_1_947), .b(output_1_4), .y(output_0_947));
wire output_2_947, output_2_4, output_1_947;
mixer gate_output_1_947(.a(output_2_947), .b(output_2_4), .y(output_1_947));
wire output_3_947, output_3_4, output_2_947;
mixer gate_output_2_947(.a(output_3_947), .b(output_3_4), .y(output_2_947));
wire output_4_947, output_4_4, output_3_947;
mixer gate_output_3_947(.a(output_4_947), .b(output_4_4), .y(output_3_947));
wire output_5_947, output_5_4, output_4_947;
mixer gate_output_4_947(.a(output_5_947), .b(output_5_4), .y(output_4_947));
wire output_6_947, output_6_4, output_5_947;
mixer gate_output_5_947(.a(output_6_947), .b(output_6_4), .y(output_5_947));
wire output_7_947, output_7_4, output_6_947;
mixer gate_output_6_947(.a(output_7_947), .b(output_7_4), .y(output_6_947));
wire output_8_947, output_8_4, output_7_947;
mixer gate_output_7_947(.a(output_8_947), .b(output_8_4), .y(output_7_947));
wire output_9_947, output_9_4, output_8_947;
mixer gate_output_8_947(.a(output_9_947), .b(output_9_4), .y(output_8_947));
wire output_10_947, output_10_4, output_9_947;
mixer gate_output_9_947(.a(output_10_947), .b(output_10_4), .y(output_9_947));
wire output_11_947, output_11_4, output_10_947;
mixer gate_output_10_947(.a(output_11_947), .b(output_11_4), .y(output_10_947));
wire output_12_947, output_12_4, output_11_947;
mixer gate_output_11_947(.a(output_12_947), .b(output_12_4), .y(output_11_947));
wire output_13_947, output_13_4, output_12_947;
mixer gate_output_12_947(.a(output_13_947), .b(output_13_4), .y(output_12_947));
wire output_14_947, output_14_4, output_13_947;
mixer gate_output_13_947(.a(output_14_947), .b(output_14_4), .y(output_13_947));
wire output_15_947, output_15_4, output_14_947;
mixer gate_output_14_947(.a(output_15_947), .b(output_15_4), .y(output_14_947));
wire output_16_947, output_16_4, output_15_947;
mixer gate_output_15_947(.a(output_16_947), .b(output_16_4), .y(output_15_947));
wire output_1_948, output_1_5, output_0_948;
mixer gate_output_0_948(.a(output_1_948), .b(output_1_5), .y(output_0_948));
wire output_2_948, output_2_5, output_1_948;
mixer gate_output_1_948(.a(output_2_948), .b(output_2_5), .y(output_1_948));
wire output_3_948, output_3_5, output_2_948;
mixer gate_output_2_948(.a(output_3_948), .b(output_3_5), .y(output_2_948));
wire output_4_948, output_4_5, output_3_948;
mixer gate_output_3_948(.a(output_4_948), .b(output_4_5), .y(output_3_948));
wire output_5_948, output_5_5, output_4_948;
mixer gate_output_4_948(.a(output_5_948), .b(output_5_5), .y(output_4_948));
wire output_6_948, output_6_5, output_5_948;
mixer gate_output_5_948(.a(output_6_948), .b(output_6_5), .y(output_5_948));
wire output_7_948, output_7_5, output_6_948;
mixer gate_output_6_948(.a(output_7_948), .b(output_7_5), .y(output_6_948));
wire output_8_948, output_8_5, output_7_948;
mixer gate_output_7_948(.a(output_8_948), .b(output_8_5), .y(output_7_948));
wire output_9_948, output_9_5, output_8_948;
mixer gate_output_8_948(.a(output_9_948), .b(output_9_5), .y(output_8_948));
wire output_10_948, output_10_5, output_9_948;
mixer gate_output_9_948(.a(output_10_948), .b(output_10_5), .y(output_9_948));
wire output_11_948, output_11_5, output_10_948;
mixer gate_output_10_948(.a(output_11_948), .b(output_11_5), .y(output_10_948));
wire output_12_948, output_12_5, output_11_948;
mixer gate_output_11_948(.a(output_12_948), .b(output_12_5), .y(output_11_948));
wire output_13_948, output_13_5, output_12_948;
mixer gate_output_12_948(.a(output_13_948), .b(output_13_5), .y(output_12_948));
wire output_14_948, output_14_5, output_13_948;
mixer gate_output_13_948(.a(output_14_948), .b(output_14_5), .y(output_13_948));
wire output_15_948, output_15_5, output_14_948;
mixer gate_output_14_948(.a(output_15_948), .b(output_15_5), .y(output_14_948));
wire output_16_948, output_16_5, output_15_948;
mixer gate_output_15_948(.a(output_16_948), .b(output_16_5), .y(output_15_948));
wire output_1_949, output_1_6, output_0_949;
mixer gate_output_0_949(.a(output_1_949), .b(output_1_6), .y(output_0_949));
wire output_2_949, output_2_6, output_1_949;
mixer gate_output_1_949(.a(output_2_949), .b(output_2_6), .y(output_1_949));
wire output_3_949, output_3_6, output_2_949;
mixer gate_output_2_949(.a(output_3_949), .b(output_3_6), .y(output_2_949));
wire output_4_949, output_4_6, output_3_949;
mixer gate_output_3_949(.a(output_4_949), .b(output_4_6), .y(output_3_949));
wire output_5_949, output_5_6, output_4_949;
mixer gate_output_4_949(.a(output_5_949), .b(output_5_6), .y(output_4_949));
wire output_6_949, output_6_6, output_5_949;
mixer gate_output_5_949(.a(output_6_949), .b(output_6_6), .y(output_5_949));
wire output_7_949, output_7_6, output_6_949;
mixer gate_output_6_949(.a(output_7_949), .b(output_7_6), .y(output_6_949));
wire output_8_949, output_8_6, output_7_949;
mixer gate_output_7_949(.a(output_8_949), .b(output_8_6), .y(output_7_949));
wire output_9_949, output_9_6, output_8_949;
mixer gate_output_8_949(.a(output_9_949), .b(output_9_6), .y(output_8_949));
wire output_10_949, output_10_6, output_9_949;
mixer gate_output_9_949(.a(output_10_949), .b(output_10_6), .y(output_9_949));
wire output_11_949, output_11_6, output_10_949;
mixer gate_output_10_949(.a(output_11_949), .b(output_11_6), .y(output_10_949));
wire output_12_949, output_12_6, output_11_949;
mixer gate_output_11_949(.a(output_12_949), .b(output_12_6), .y(output_11_949));
wire output_13_949, output_13_6, output_12_949;
mixer gate_output_12_949(.a(output_13_949), .b(output_13_6), .y(output_12_949));
wire output_14_949, output_14_6, output_13_949;
mixer gate_output_13_949(.a(output_14_949), .b(output_14_6), .y(output_13_949));
wire output_15_949, output_15_6, output_14_949;
mixer gate_output_14_949(.a(output_15_949), .b(output_15_6), .y(output_14_949));
wire output_16_949, output_16_6, output_15_949;
mixer gate_output_15_949(.a(output_16_949), .b(output_16_6), .y(output_15_949));
wire output_1_950, output_1_7, output_0_950;
mixer gate_output_0_950(.a(output_1_950), .b(output_1_7), .y(output_0_950));
wire output_2_950, output_2_7, output_1_950;
mixer gate_output_1_950(.a(output_2_950), .b(output_2_7), .y(output_1_950));
wire output_3_950, output_3_7, output_2_950;
mixer gate_output_2_950(.a(output_3_950), .b(output_3_7), .y(output_2_950));
wire output_4_950, output_4_7, output_3_950;
mixer gate_output_3_950(.a(output_4_950), .b(output_4_7), .y(output_3_950));
wire output_5_950, output_5_7, output_4_950;
mixer gate_output_4_950(.a(output_5_950), .b(output_5_7), .y(output_4_950));
wire output_6_950, output_6_7, output_5_950;
mixer gate_output_5_950(.a(output_6_950), .b(output_6_7), .y(output_5_950));
wire output_7_950, output_7_7, output_6_950;
mixer gate_output_6_950(.a(output_7_950), .b(output_7_7), .y(output_6_950));
wire output_8_950, output_8_7, output_7_950;
mixer gate_output_7_950(.a(output_8_950), .b(output_8_7), .y(output_7_950));
wire output_9_950, output_9_7, output_8_950;
mixer gate_output_8_950(.a(output_9_950), .b(output_9_7), .y(output_8_950));
wire output_10_950, output_10_7, output_9_950;
mixer gate_output_9_950(.a(output_10_950), .b(output_10_7), .y(output_9_950));
wire output_11_950, output_11_7, output_10_950;
mixer gate_output_10_950(.a(output_11_950), .b(output_11_7), .y(output_10_950));
wire output_12_950, output_12_7, output_11_950;
mixer gate_output_11_950(.a(output_12_950), .b(output_12_7), .y(output_11_950));
wire output_13_950, output_13_7, output_12_950;
mixer gate_output_12_950(.a(output_13_950), .b(output_13_7), .y(output_12_950));
wire output_14_950, output_14_7, output_13_950;
mixer gate_output_13_950(.a(output_14_950), .b(output_14_7), .y(output_13_950));
wire output_15_950, output_15_7, output_14_950;
mixer gate_output_14_950(.a(output_15_950), .b(output_15_7), .y(output_14_950));
wire output_16_950, output_16_7, output_15_950;
mixer gate_output_15_950(.a(output_16_950), .b(output_16_7), .y(output_15_950));
wire output_1_951, output_1_8, output_0_951;
mixer gate_output_0_951(.a(output_1_951), .b(output_1_8), .y(output_0_951));
wire output_2_951, output_2_8, output_1_951;
mixer gate_output_1_951(.a(output_2_951), .b(output_2_8), .y(output_1_951));
wire output_3_951, output_3_8, output_2_951;
mixer gate_output_2_951(.a(output_3_951), .b(output_3_8), .y(output_2_951));
wire output_4_951, output_4_8, output_3_951;
mixer gate_output_3_951(.a(output_4_951), .b(output_4_8), .y(output_3_951));
wire output_5_951, output_5_8, output_4_951;
mixer gate_output_4_951(.a(output_5_951), .b(output_5_8), .y(output_4_951));
wire output_6_951, output_6_8, output_5_951;
mixer gate_output_5_951(.a(output_6_951), .b(output_6_8), .y(output_5_951));
wire output_7_951, output_7_8, output_6_951;
mixer gate_output_6_951(.a(output_7_951), .b(output_7_8), .y(output_6_951));
wire output_8_951, output_8_8, output_7_951;
mixer gate_output_7_951(.a(output_8_951), .b(output_8_8), .y(output_7_951));
wire output_9_951, output_9_8, output_8_951;
mixer gate_output_8_951(.a(output_9_951), .b(output_9_8), .y(output_8_951));
wire output_10_951, output_10_8, output_9_951;
mixer gate_output_9_951(.a(output_10_951), .b(output_10_8), .y(output_9_951));
wire output_11_951, output_11_8, output_10_951;
mixer gate_output_10_951(.a(output_11_951), .b(output_11_8), .y(output_10_951));
wire output_12_951, output_12_8, output_11_951;
mixer gate_output_11_951(.a(output_12_951), .b(output_12_8), .y(output_11_951));
wire output_13_951, output_13_8, output_12_951;
mixer gate_output_12_951(.a(output_13_951), .b(output_13_8), .y(output_12_951));
wire output_14_951, output_14_8, output_13_951;
mixer gate_output_13_951(.a(output_14_951), .b(output_14_8), .y(output_13_951));
wire output_15_951, output_15_8, output_14_951;
mixer gate_output_14_951(.a(output_15_951), .b(output_15_8), .y(output_14_951));
wire output_16_951, output_16_8, output_15_951;
mixer gate_output_15_951(.a(output_16_951), .b(output_16_8), .y(output_15_951));
wire output_1_952, output_1_9, output_0_952;
mixer gate_output_0_952(.a(output_1_952), .b(output_1_9), .y(output_0_952));
wire output_2_952, output_2_9, output_1_952;
mixer gate_output_1_952(.a(output_2_952), .b(output_2_9), .y(output_1_952));
wire output_3_952, output_3_9, output_2_952;
mixer gate_output_2_952(.a(output_3_952), .b(output_3_9), .y(output_2_952));
wire output_4_952, output_4_9, output_3_952;
mixer gate_output_3_952(.a(output_4_952), .b(output_4_9), .y(output_3_952));
wire output_5_952, output_5_9, output_4_952;
mixer gate_output_4_952(.a(output_5_952), .b(output_5_9), .y(output_4_952));
wire output_6_952, output_6_9, output_5_952;
mixer gate_output_5_952(.a(output_6_952), .b(output_6_9), .y(output_5_952));
wire output_7_952, output_7_9, output_6_952;
mixer gate_output_6_952(.a(output_7_952), .b(output_7_9), .y(output_6_952));
wire output_8_952, output_8_9, output_7_952;
mixer gate_output_7_952(.a(output_8_952), .b(output_8_9), .y(output_7_952));
wire output_9_952, output_9_9, output_8_952;
mixer gate_output_8_952(.a(output_9_952), .b(output_9_9), .y(output_8_952));
wire output_10_952, output_10_9, output_9_952;
mixer gate_output_9_952(.a(output_10_952), .b(output_10_9), .y(output_9_952));
wire output_11_952, output_11_9, output_10_952;
mixer gate_output_10_952(.a(output_11_952), .b(output_11_9), .y(output_10_952));
wire output_12_952, output_12_9, output_11_952;
mixer gate_output_11_952(.a(output_12_952), .b(output_12_9), .y(output_11_952));
wire output_13_952, output_13_9, output_12_952;
mixer gate_output_12_952(.a(output_13_952), .b(output_13_9), .y(output_12_952));
wire output_14_952, output_14_9, output_13_952;
mixer gate_output_13_952(.a(output_14_952), .b(output_14_9), .y(output_13_952));
wire output_15_952, output_15_9, output_14_952;
mixer gate_output_14_952(.a(output_15_952), .b(output_15_9), .y(output_14_952));
wire output_16_952, output_16_9, output_15_952;
mixer gate_output_15_952(.a(output_16_952), .b(output_16_9), .y(output_15_952));
wire output_1_953, output_1_10, output_0_953;
mixer gate_output_0_953(.a(output_1_953), .b(output_1_10), .y(output_0_953));
wire output_2_953, output_2_10, output_1_953;
mixer gate_output_1_953(.a(output_2_953), .b(output_2_10), .y(output_1_953));
wire output_3_953, output_3_10, output_2_953;
mixer gate_output_2_953(.a(output_3_953), .b(output_3_10), .y(output_2_953));
wire output_4_953, output_4_10, output_3_953;
mixer gate_output_3_953(.a(output_4_953), .b(output_4_10), .y(output_3_953));
wire output_5_953, output_5_10, output_4_953;
mixer gate_output_4_953(.a(output_5_953), .b(output_5_10), .y(output_4_953));
wire output_6_953, output_6_10, output_5_953;
mixer gate_output_5_953(.a(output_6_953), .b(output_6_10), .y(output_5_953));
wire output_7_953, output_7_10, output_6_953;
mixer gate_output_6_953(.a(output_7_953), .b(output_7_10), .y(output_6_953));
wire output_8_953, output_8_10, output_7_953;
mixer gate_output_7_953(.a(output_8_953), .b(output_8_10), .y(output_7_953));
wire output_9_953, output_9_10, output_8_953;
mixer gate_output_8_953(.a(output_9_953), .b(output_9_10), .y(output_8_953));
wire output_10_953, output_10_10, output_9_953;
mixer gate_output_9_953(.a(output_10_953), .b(output_10_10), .y(output_9_953));
wire output_11_953, output_11_10, output_10_953;
mixer gate_output_10_953(.a(output_11_953), .b(output_11_10), .y(output_10_953));
wire output_12_953, output_12_10, output_11_953;
mixer gate_output_11_953(.a(output_12_953), .b(output_12_10), .y(output_11_953));
wire output_13_953, output_13_10, output_12_953;
mixer gate_output_12_953(.a(output_13_953), .b(output_13_10), .y(output_12_953));
wire output_14_953, output_14_10, output_13_953;
mixer gate_output_13_953(.a(output_14_953), .b(output_14_10), .y(output_13_953));
wire output_15_953, output_15_10, output_14_953;
mixer gate_output_14_953(.a(output_15_953), .b(output_15_10), .y(output_14_953));
wire output_16_953, output_16_10, output_15_953;
mixer gate_output_15_953(.a(output_16_953), .b(output_16_10), .y(output_15_953));
wire output_1_954, output_1_11, output_0_954;
mixer gate_output_0_954(.a(output_1_954), .b(output_1_11), .y(output_0_954));
wire output_2_954, output_2_11, output_1_954;
mixer gate_output_1_954(.a(output_2_954), .b(output_2_11), .y(output_1_954));
wire output_3_954, output_3_11, output_2_954;
mixer gate_output_2_954(.a(output_3_954), .b(output_3_11), .y(output_2_954));
wire output_4_954, output_4_11, output_3_954;
mixer gate_output_3_954(.a(output_4_954), .b(output_4_11), .y(output_3_954));
wire output_5_954, output_5_11, output_4_954;
mixer gate_output_4_954(.a(output_5_954), .b(output_5_11), .y(output_4_954));
wire output_6_954, output_6_11, output_5_954;
mixer gate_output_5_954(.a(output_6_954), .b(output_6_11), .y(output_5_954));
wire output_7_954, output_7_11, output_6_954;
mixer gate_output_6_954(.a(output_7_954), .b(output_7_11), .y(output_6_954));
wire output_8_954, output_8_11, output_7_954;
mixer gate_output_7_954(.a(output_8_954), .b(output_8_11), .y(output_7_954));
wire output_9_954, output_9_11, output_8_954;
mixer gate_output_8_954(.a(output_9_954), .b(output_9_11), .y(output_8_954));
wire output_10_954, output_10_11, output_9_954;
mixer gate_output_9_954(.a(output_10_954), .b(output_10_11), .y(output_9_954));
wire output_11_954, output_11_11, output_10_954;
mixer gate_output_10_954(.a(output_11_954), .b(output_11_11), .y(output_10_954));
wire output_12_954, output_12_11, output_11_954;
mixer gate_output_11_954(.a(output_12_954), .b(output_12_11), .y(output_11_954));
wire output_13_954, output_13_11, output_12_954;
mixer gate_output_12_954(.a(output_13_954), .b(output_13_11), .y(output_12_954));
wire output_14_954, output_14_11, output_13_954;
mixer gate_output_13_954(.a(output_14_954), .b(output_14_11), .y(output_13_954));
wire output_15_954, output_15_11, output_14_954;
mixer gate_output_14_954(.a(output_15_954), .b(output_15_11), .y(output_14_954));
wire output_16_954, output_16_11, output_15_954;
mixer gate_output_15_954(.a(output_16_954), .b(output_16_11), .y(output_15_954));
wire output_1_955, output_1_12, output_0_955;
mixer gate_output_0_955(.a(output_1_955), .b(output_1_12), .y(output_0_955));
wire output_2_955, output_2_12, output_1_955;
mixer gate_output_1_955(.a(output_2_955), .b(output_2_12), .y(output_1_955));
wire output_3_955, output_3_12, output_2_955;
mixer gate_output_2_955(.a(output_3_955), .b(output_3_12), .y(output_2_955));
wire output_4_955, output_4_12, output_3_955;
mixer gate_output_3_955(.a(output_4_955), .b(output_4_12), .y(output_3_955));
wire output_5_955, output_5_12, output_4_955;
mixer gate_output_4_955(.a(output_5_955), .b(output_5_12), .y(output_4_955));
wire output_6_955, output_6_12, output_5_955;
mixer gate_output_5_955(.a(output_6_955), .b(output_6_12), .y(output_5_955));
wire output_7_955, output_7_12, output_6_955;
mixer gate_output_6_955(.a(output_7_955), .b(output_7_12), .y(output_6_955));
wire output_8_955, output_8_12, output_7_955;
mixer gate_output_7_955(.a(output_8_955), .b(output_8_12), .y(output_7_955));
wire output_9_955, output_9_12, output_8_955;
mixer gate_output_8_955(.a(output_9_955), .b(output_9_12), .y(output_8_955));
wire output_10_955, output_10_12, output_9_955;
mixer gate_output_9_955(.a(output_10_955), .b(output_10_12), .y(output_9_955));
wire output_11_955, output_11_12, output_10_955;
mixer gate_output_10_955(.a(output_11_955), .b(output_11_12), .y(output_10_955));
wire output_12_955, output_12_12, output_11_955;
mixer gate_output_11_955(.a(output_12_955), .b(output_12_12), .y(output_11_955));
wire output_13_955, output_13_12, output_12_955;
mixer gate_output_12_955(.a(output_13_955), .b(output_13_12), .y(output_12_955));
wire output_14_955, output_14_12, output_13_955;
mixer gate_output_13_955(.a(output_14_955), .b(output_14_12), .y(output_13_955));
wire output_15_955, output_15_12, output_14_955;
mixer gate_output_14_955(.a(output_15_955), .b(output_15_12), .y(output_14_955));
wire output_16_955, output_16_12, output_15_955;
mixer gate_output_15_955(.a(output_16_955), .b(output_16_12), .y(output_15_955));
wire output_1_956, output_1_13, output_0_956;
mixer gate_output_0_956(.a(output_1_956), .b(output_1_13), .y(output_0_956));
wire output_2_956, output_2_13, output_1_956;
mixer gate_output_1_956(.a(output_2_956), .b(output_2_13), .y(output_1_956));
wire output_3_956, output_3_13, output_2_956;
mixer gate_output_2_956(.a(output_3_956), .b(output_3_13), .y(output_2_956));
wire output_4_956, output_4_13, output_3_956;
mixer gate_output_3_956(.a(output_4_956), .b(output_4_13), .y(output_3_956));
wire output_5_956, output_5_13, output_4_956;
mixer gate_output_4_956(.a(output_5_956), .b(output_5_13), .y(output_4_956));
wire output_6_956, output_6_13, output_5_956;
mixer gate_output_5_956(.a(output_6_956), .b(output_6_13), .y(output_5_956));
wire output_7_956, output_7_13, output_6_956;
mixer gate_output_6_956(.a(output_7_956), .b(output_7_13), .y(output_6_956));
wire output_8_956, output_8_13, output_7_956;
mixer gate_output_7_956(.a(output_8_956), .b(output_8_13), .y(output_7_956));
wire output_9_956, output_9_13, output_8_956;
mixer gate_output_8_956(.a(output_9_956), .b(output_9_13), .y(output_8_956));
wire output_10_956, output_10_13, output_9_956;
mixer gate_output_9_956(.a(output_10_956), .b(output_10_13), .y(output_9_956));
wire output_11_956, output_11_13, output_10_956;
mixer gate_output_10_956(.a(output_11_956), .b(output_11_13), .y(output_10_956));
wire output_12_956, output_12_13, output_11_956;
mixer gate_output_11_956(.a(output_12_956), .b(output_12_13), .y(output_11_956));
wire output_13_956, output_13_13, output_12_956;
mixer gate_output_12_956(.a(output_13_956), .b(output_13_13), .y(output_12_956));
wire output_14_956, output_14_13, output_13_956;
mixer gate_output_13_956(.a(output_14_956), .b(output_14_13), .y(output_13_956));
wire output_15_956, output_15_13, output_14_956;
mixer gate_output_14_956(.a(output_15_956), .b(output_15_13), .y(output_14_956));
wire output_16_956, output_16_13, output_15_956;
mixer gate_output_15_956(.a(output_16_956), .b(output_16_13), .y(output_15_956));
wire output_1_957, output_1_14, output_0_957;
mixer gate_output_0_957(.a(output_1_957), .b(output_1_14), .y(output_0_957));
wire output_2_957, output_2_14, output_1_957;
mixer gate_output_1_957(.a(output_2_957), .b(output_2_14), .y(output_1_957));
wire output_3_957, output_3_14, output_2_957;
mixer gate_output_2_957(.a(output_3_957), .b(output_3_14), .y(output_2_957));
wire output_4_957, output_4_14, output_3_957;
mixer gate_output_3_957(.a(output_4_957), .b(output_4_14), .y(output_3_957));
wire output_5_957, output_5_14, output_4_957;
mixer gate_output_4_957(.a(output_5_957), .b(output_5_14), .y(output_4_957));
wire output_6_957, output_6_14, output_5_957;
mixer gate_output_5_957(.a(output_6_957), .b(output_6_14), .y(output_5_957));
wire output_7_957, output_7_14, output_6_957;
mixer gate_output_6_957(.a(output_7_957), .b(output_7_14), .y(output_6_957));
wire output_8_957, output_8_14, output_7_957;
mixer gate_output_7_957(.a(output_8_957), .b(output_8_14), .y(output_7_957));
wire output_9_957, output_9_14, output_8_957;
mixer gate_output_8_957(.a(output_9_957), .b(output_9_14), .y(output_8_957));
wire output_10_957, output_10_14, output_9_957;
mixer gate_output_9_957(.a(output_10_957), .b(output_10_14), .y(output_9_957));
wire output_11_957, output_11_14, output_10_957;
mixer gate_output_10_957(.a(output_11_957), .b(output_11_14), .y(output_10_957));
wire output_12_957, output_12_14, output_11_957;
mixer gate_output_11_957(.a(output_12_957), .b(output_12_14), .y(output_11_957));
wire output_13_957, output_13_14, output_12_957;
mixer gate_output_12_957(.a(output_13_957), .b(output_13_14), .y(output_12_957));
wire output_14_957, output_14_14, output_13_957;
mixer gate_output_13_957(.a(output_14_957), .b(output_14_14), .y(output_13_957));
wire output_15_957, output_15_14, output_14_957;
mixer gate_output_14_957(.a(output_15_957), .b(output_15_14), .y(output_14_957));
wire output_16_957, output_16_14, output_15_957;
mixer gate_output_15_957(.a(output_16_957), .b(output_16_14), .y(output_15_957));
wire output_1_958, output_1_15, output_0_958;
mixer gate_output_0_958(.a(output_1_958), .b(output_1_15), .y(output_0_958));
wire output_2_958, output_2_15, output_1_958;
mixer gate_output_1_958(.a(output_2_958), .b(output_2_15), .y(output_1_958));
wire output_3_958, output_3_15, output_2_958;
mixer gate_output_2_958(.a(output_3_958), .b(output_3_15), .y(output_2_958));
wire output_4_958, output_4_15, output_3_958;
mixer gate_output_3_958(.a(output_4_958), .b(output_4_15), .y(output_3_958));
wire output_5_958, output_5_15, output_4_958;
mixer gate_output_4_958(.a(output_5_958), .b(output_5_15), .y(output_4_958));
wire output_6_958, output_6_15, output_5_958;
mixer gate_output_5_958(.a(output_6_958), .b(output_6_15), .y(output_5_958));
wire output_7_958, output_7_15, output_6_958;
mixer gate_output_6_958(.a(output_7_958), .b(output_7_15), .y(output_6_958));
wire output_8_958, output_8_15, output_7_958;
mixer gate_output_7_958(.a(output_8_958), .b(output_8_15), .y(output_7_958));
wire output_9_958, output_9_15, output_8_958;
mixer gate_output_8_958(.a(output_9_958), .b(output_9_15), .y(output_8_958));
wire output_10_958, output_10_15, output_9_958;
mixer gate_output_9_958(.a(output_10_958), .b(output_10_15), .y(output_9_958));
wire output_11_958, output_11_15, output_10_958;
mixer gate_output_10_958(.a(output_11_958), .b(output_11_15), .y(output_10_958));
wire output_12_958, output_12_15, output_11_958;
mixer gate_output_11_958(.a(output_12_958), .b(output_12_15), .y(output_11_958));
wire output_13_958, output_13_15, output_12_958;
mixer gate_output_12_958(.a(output_13_958), .b(output_13_15), .y(output_12_958));
wire output_14_958, output_14_15, output_13_958;
mixer gate_output_13_958(.a(output_14_958), .b(output_14_15), .y(output_13_958));
wire output_15_958, output_15_15, output_14_958;
mixer gate_output_14_958(.a(output_15_958), .b(output_15_15), .y(output_14_958));
wire output_16_958, output_16_15, output_15_958;
mixer gate_output_15_958(.a(output_16_958), .b(output_16_15), .y(output_15_958));
wire output_1_959, output_1_0, output_0_959;
mixer gate_output_0_959(.a(output_1_959), .b(output_1_0), .y(output_0_959));
wire output_2_959, output_2_0, output_1_959;
mixer gate_output_1_959(.a(output_2_959), .b(output_2_0), .y(output_1_959));
wire output_3_959, output_3_0, output_2_959;
mixer gate_output_2_959(.a(output_3_959), .b(output_3_0), .y(output_2_959));
wire output_4_959, output_4_0, output_3_959;
mixer gate_output_3_959(.a(output_4_959), .b(output_4_0), .y(output_3_959));
wire output_5_959, output_5_0, output_4_959;
mixer gate_output_4_959(.a(output_5_959), .b(output_5_0), .y(output_4_959));
wire output_6_959, output_6_0, output_5_959;
mixer gate_output_5_959(.a(output_6_959), .b(output_6_0), .y(output_5_959));
wire output_7_959, output_7_0, output_6_959;
mixer gate_output_6_959(.a(output_7_959), .b(output_7_0), .y(output_6_959));
wire output_8_959, output_8_0, output_7_959;
mixer gate_output_7_959(.a(output_8_959), .b(output_8_0), .y(output_7_959));
wire output_9_959, output_9_0, output_8_959;
mixer gate_output_8_959(.a(output_9_959), .b(output_9_0), .y(output_8_959));
wire output_10_959, output_10_0, output_9_959;
mixer gate_output_9_959(.a(output_10_959), .b(output_10_0), .y(output_9_959));
wire output_11_959, output_11_0, output_10_959;
mixer gate_output_10_959(.a(output_11_959), .b(output_11_0), .y(output_10_959));
wire output_12_959, output_12_0, output_11_959;
mixer gate_output_11_959(.a(output_12_959), .b(output_12_0), .y(output_11_959));
wire output_13_959, output_13_0, output_12_959;
mixer gate_output_12_959(.a(output_13_959), .b(output_13_0), .y(output_12_959));
wire output_14_959, output_14_0, output_13_959;
mixer gate_output_13_959(.a(output_14_959), .b(output_14_0), .y(output_13_959));
wire output_15_959, output_15_0, output_14_959;
mixer gate_output_14_959(.a(output_15_959), .b(output_15_0), .y(output_14_959));
wire output_16_959, output_16_0, output_15_959;
mixer gate_output_15_959(.a(output_16_959), .b(output_16_0), .y(output_15_959));
wire output_1_960, output_1_1, output_0_960;
mixer gate_output_0_960(.a(output_1_960), .b(output_1_1), .y(output_0_960));
wire output_2_960, output_2_1, output_1_960;
mixer gate_output_1_960(.a(output_2_960), .b(output_2_1), .y(output_1_960));
wire output_3_960, output_3_1, output_2_960;
mixer gate_output_2_960(.a(output_3_960), .b(output_3_1), .y(output_2_960));
wire output_4_960, output_4_1, output_3_960;
mixer gate_output_3_960(.a(output_4_960), .b(output_4_1), .y(output_3_960));
wire output_5_960, output_5_1, output_4_960;
mixer gate_output_4_960(.a(output_5_960), .b(output_5_1), .y(output_4_960));
wire output_6_960, output_6_1, output_5_960;
mixer gate_output_5_960(.a(output_6_960), .b(output_6_1), .y(output_5_960));
wire output_7_960, output_7_1, output_6_960;
mixer gate_output_6_960(.a(output_7_960), .b(output_7_1), .y(output_6_960));
wire output_8_960, output_8_1, output_7_960;
mixer gate_output_7_960(.a(output_8_960), .b(output_8_1), .y(output_7_960));
wire output_9_960, output_9_1, output_8_960;
mixer gate_output_8_960(.a(output_9_960), .b(output_9_1), .y(output_8_960));
wire output_10_960, output_10_1, output_9_960;
mixer gate_output_9_960(.a(output_10_960), .b(output_10_1), .y(output_9_960));
wire output_11_960, output_11_1, output_10_960;
mixer gate_output_10_960(.a(output_11_960), .b(output_11_1), .y(output_10_960));
wire output_12_960, output_12_1, output_11_960;
mixer gate_output_11_960(.a(output_12_960), .b(output_12_1), .y(output_11_960));
wire output_13_960, output_13_1, output_12_960;
mixer gate_output_12_960(.a(output_13_960), .b(output_13_1), .y(output_12_960));
wire output_14_960, output_14_1, output_13_960;
mixer gate_output_13_960(.a(output_14_960), .b(output_14_1), .y(output_13_960));
wire output_15_960, output_15_1, output_14_960;
mixer gate_output_14_960(.a(output_15_960), .b(output_15_1), .y(output_14_960));
wire output_16_960, output_16_1, output_15_960;
mixer gate_output_15_960(.a(output_16_960), .b(output_16_1), .y(output_15_960));
wire output_1_961, output_1_2, output_0_961;
mixer gate_output_0_961(.a(output_1_961), .b(output_1_2), .y(output_0_961));
wire output_2_961, output_2_2, output_1_961;
mixer gate_output_1_961(.a(output_2_961), .b(output_2_2), .y(output_1_961));
wire output_3_961, output_3_2, output_2_961;
mixer gate_output_2_961(.a(output_3_961), .b(output_3_2), .y(output_2_961));
wire output_4_961, output_4_2, output_3_961;
mixer gate_output_3_961(.a(output_4_961), .b(output_4_2), .y(output_3_961));
wire output_5_961, output_5_2, output_4_961;
mixer gate_output_4_961(.a(output_5_961), .b(output_5_2), .y(output_4_961));
wire output_6_961, output_6_2, output_5_961;
mixer gate_output_5_961(.a(output_6_961), .b(output_6_2), .y(output_5_961));
wire output_7_961, output_7_2, output_6_961;
mixer gate_output_6_961(.a(output_7_961), .b(output_7_2), .y(output_6_961));
wire output_8_961, output_8_2, output_7_961;
mixer gate_output_7_961(.a(output_8_961), .b(output_8_2), .y(output_7_961));
wire output_9_961, output_9_2, output_8_961;
mixer gate_output_8_961(.a(output_9_961), .b(output_9_2), .y(output_8_961));
wire output_10_961, output_10_2, output_9_961;
mixer gate_output_9_961(.a(output_10_961), .b(output_10_2), .y(output_9_961));
wire output_11_961, output_11_2, output_10_961;
mixer gate_output_10_961(.a(output_11_961), .b(output_11_2), .y(output_10_961));
wire output_12_961, output_12_2, output_11_961;
mixer gate_output_11_961(.a(output_12_961), .b(output_12_2), .y(output_11_961));
wire output_13_961, output_13_2, output_12_961;
mixer gate_output_12_961(.a(output_13_961), .b(output_13_2), .y(output_12_961));
wire output_14_961, output_14_2, output_13_961;
mixer gate_output_13_961(.a(output_14_961), .b(output_14_2), .y(output_13_961));
wire output_15_961, output_15_2, output_14_961;
mixer gate_output_14_961(.a(output_15_961), .b(output_15_2), .y(output_14_961));
wire output_16_961, output_16_2, output_15_961;
mixer gate_output_15_961(.a(output_16_961), .b(output_16_2), .y(output_15_961));
wire output_1_962, output_1_3, output_0_962;
mixer gate_output_0_962(.a(output_1_962), .b(output_1_3), .y(output_0_962));
wire output_2_962, output_2_3, output_1_962;
mixer gate_output_1_962(.a(output_2_962), .b(output_2_3), .y(output_1_962));
wire output_3_962, output_3_3, output_2_962;
mixer gate_output_2_962(.a(output_3_962), .b(output_3_3), .y(output_2_962));
wire output_4_962, output_4_3, output_3_962;
mixer gate_output_3_962(.a(output_4_962), .b(output_4_3), .y(output_3_962));
wire output_5_962, output_5_3, output_4_962;
mixer gate_output_4_962(.a(output_5_962), .b(output_5_3), .y(output_4_962));
wire output_6_962, output_6_3, output_5_962;
mixer gate_output_5_962(.a(output_6_962), .b(output_6_3), .y(output_5_962));
wire output_7_962, output_7_3, output_6_962;
mixer gate_output_6_962(.a(output_7_962), .b(output_7_3), .y(output_6_962));
wire output_8_962, output_8_3, output_7_962;
mixer gate_output_7_962(.a(output_8_962), .b(output_8_3), .y(output_7_962));
wire output_9_962, output_9_3, output_8_962;
mixer gate_output_8_962(.a(output_9_962), .b(output_9_3), .y(output_8_962));
wire output_10_962, output_10_3, output_9_962;
mixer gate_output_9_962(.a(output_10_962), .b(output_10_3), .y(output_9_962));
wire output_11_962, output_11_3, output_10_962;
mixer gate_output_10_962(.a(output_11_962), .b(output_11_3), .y(output_10_962));
wire output_12_962, output_12_3, output_11_962;
mixer gate_output_11_962(.a(output_12_962), .b(output_12_3), .y(output_11_962));
wire output_13_962, output_13_3, output_12_962;
mixer gate_output_12_962(.a(output_13_962), .b(output_13_3), .y(output_12_962));
wire output_14_962, output_14_3, output_13_962;
mixer gate_output_13_962(.a(output_14_962), .b(output_14_3), .y(output_13_962));
wire output_15_962, output_15_3, output_14_962;
mixer gate_output_14_962(.a(output_15_962), .b(output_15_3), .y(output_14_962));
wire output_16_962, output_16_3, output_15_962;
mixer gate_output_15_962(.a(output_16_962), .b(output_16_3), .y(output_15_962));
wire output_1_963, output_1_4, output_0_963;
mixer gate_output_0_963(.a(output_1_963), .b(output_1_4), .y(output_0_963));
wire output_2_963, output_2_4, output_1_963;
mixer gate_output_1_963(.a(output_2_963), .b(output_2_4), .y(output_1_963));
wire output_3_963, output_3_4, output_2_963;
mixer gate_output_2_963(.a(output_3_963), .b(output_3_4), .y(output_2_963));
wire output_4_963, output_4_4, output_3_963;
mixer gate_output_3_963(.a(output_4_963), .b(output_4_4), .y(output_3_963));
wire output_5_963, output_5_4, output_4_963;
mixer gate_output_4_963(.a(output_5_963), .b(output_5_4), .y(output_4_963));
wire output_6_963, output_6_4, output_5_963;
mixer gate_output_5_963(.a(output_6_963), .b(output_6_4), .y(output_5_963));
wire output_7_963, output_7_4, output_6_963;
mixer gate_output_6_963(.a(output_7_963), .b(output_7_4), .y(output_6_963));
wire output_8_963, output_8_4, output_7_963;
mixer gate_output_7_963(.a(output_8_963), .b(output_8_4), .y(output_7_963));
wire output_9_963, output_9_4, output_8_963;
mixer gate_output_8_963(.a(output_9_963), .b(output_9_4), .y(output_8_963));
wire output_10_963, output_10_4, output_9_963;
mixer gate_output_9_963(.a(output_10_963), .b(output_10_4), .y(output_9_963));
wire output_11_963, output_11_4, output_10_963;
mixer gate_output_10_963(.a(output_11_963), .b(output_11_4), .y(output_10_963));
wire output_12_963, output_12_4, output_11_963;
mixer gate_output_11_963(.a(output_12_963), .b(output_12_4), .y(output_11_963));
wire output_13_963, output_13_4, output_12_963;
mixer gate_output_12_963(.a(output_13_963), .b(output_13_4), .y(output_12_963));
wire output_14_963, output_14_4, output_13_963;
mixer gate_output_13_963(.a(output_14_963), .b(output_14_4), .y(output_13_963));
wire output_15_963, output_15_4, output_14_963;
mixer gate_output_14_963(.a(output_15_963), .b(output_15_4), .y(output_14_963));
wire output_16_963, output_16_4, output_15_963;
mixer gate_output_15_963(.a(output_16_963), .b(output_16_4), .y(output_15_963));
wire output_1_964, output_1_5, output_0_964;
mixer gate_output_0_964(.a(output_1_964), .b(output_1_5), .y(output_0_964));
wire output_2_964, output_2_5, output_1_964;
mixer gate_output_1_964(.a(output_2_964), .b(output_2_5), .y(output_1_964));
wire output_3_964, output_3_5, output_2_964;
mixer gate_output_2_964(.a(output_3_964), .b(output_3_5), .y(output_2_964));
wire output_4_964, output_4_5, output_3_964;
mixer gate_output_3_964(.a(output_4_964), .b(output_4_5), .y(output_3_964));
wire output_5_964, output_5_5, output_4_964;
mixer gate_output_4_964(.a(output_5_964), .b(output_5_5), .y(output_4_964));
wire output_6_964, output_6_5, output_5_964;
mixer gate_output_5_964(.a(output_6_964), .b(output_6_5), .y(output_5_964));
wire output_7_964, output_7_5, output_6_964;
mixer gate_output_6_964(.a(output_7_964), .b(output_7_5), .y(output_6_964));
wire output_8_964, output_8_5, output_7_964;
mixer gate_output_7_964(.a(output_8_964), .b(output_8_5), .y(output_7_964));
wire output_9_964, output_9_5, output_8_964;
mixer gate_output_8_964(.a(output_9_964), .b(output_9_5), .y(output_8_964));
wire output_10_964, output_10_5, output_9_964;
mixer gate_output_9_964(.a(output_10_964), .b(output_10_5), .y(output_9_964));
wire output_11_964, output_11_5, output_10_964;
mixer gate_output_10_964(.a(output_11_964), .b(output_11_5), .y(output_10_964));
wire output_12_964, output_12_5, output_11_964;
mixer gate_output_11_964(.a(output_12_964), .b(output_12_5), .y(output_11_964));
wire output_13_964, output_13_5, output_12_964;
mixer gate_output_12_964(.a(output_13_964), .b(output_13_5), .y(output_12_964));
wire output_14_964, output_14_5, output_13_964;
mixer gate_output_13_964(.a(output_14_964), .b(output_14_5), .y(output_13_964));
wire output_15_964, output_15_5, output_14_964;
mixer gate_output_14_964(.a(output_15_964), .b(output_15_5), .y(output_14_964));
wire output_16_964, output_16_5, output_15_964;
mixer gate_output_15_964(.a(output_16_964), .b(output_16_5), .y(output_15_964));
wire output_1_965, output_1_6, output_0_965;
mixer gate_output_0_965(.a(output_1_965), .b(output_1_6), .y(output_0_965));
wire output_2_965, output_2_6, output_1_965;
mixer gate_output_1_965(.a(output_2_965), .b(output_2_6), .y(output_1_965));
wire output_3_965, output_3_6, output_2_965;
mixer gate_output_2_965(.a(output_3_965), .b(output_3_6), .y(output_2_965));
wire output_4_965, output_4_6, output_3_965;
mixer gate_output_3_965(.a(output_4_965), .b(output_4_6), .y(output_3_965));
wire output_5_965, output_5_6, output_4_965;
mixer gate_output_4_965(.a(output_5_965), .b(output_5_6), .y(output_4_965));
wire output_6_965, output_6_6, output_5_965;
mixer gate_output_5_965(.a(output_6_965), .b(output_6_6), .y(output_5_965));
wire output_7_965, output_7_6, output_6_965;
mixer gate_output_6_965(.a(output_7_965), .b(output_7_6), .y(output_6_965));
wire output_8_965, output_8_6, output_7_965;
mixer gate_output_7_965(.a(output_8_965), .b(output_8_6), .y(output_7_965));
wire output_9_965, output_9_6, output_8_965;
mixer gate_output_8_965(.a(output_9_965), .b(output_9_6), .y(output_8_965));
wire output_10_965, output_10_6, output_9_965;
mixer gate_output_9_965(.a(output_10_965), .b(output_10_6), .y(output_9_965));
wire output_11_965, output_11_6, output_10_965;
mixer gate_output_10_965(.a(output_11_965), .b(output_11_6), .y(output_10_965));
wire output_12_965, output_12_6, output_11_965;
mixer gate_output_11_965(.a(output_12_965), .b(output_12_6), .y(output_11_965));
wire output_13_965, output_13_6, output_12_965;
mixer gate_output_12_965(.a(output_13_965), .b(output_13_6), .y(output_12_965));
wire output_14_965, output_14_6, output_13_965;
mixer gate_output_13_965(.a(output_14_965), .b(output_14_6), .y(output_13_965));
wire output_15_965, output_15_6, output_14_965;
mixer gate_output_14_965(.a(output_15_965), .b(output_15_6), .y(output_14_965));
wire output_16_965, output_16_6, output_15_965;
mixer gate_output_15_965(.a(output_16_965), .b(output_16_6), .y(output_15_965));
wire output_1_966, output_1_7, output_0_966;
mixer gate_output_0_966(.a(output_1_966), .b(output_1_7), .y(output_0_966));
wire output_2_966, output_2_7, output_1_966;
mixer gate_output_1_966(.a(output_2_966), .b(output_2_7), .y(output_1_966));
wire output_3_966, output_3_7, output_2_966;
mixer gate_output_2_966(.a(output_3_966), .b(output_3_7), .y(output_2_966));
wire output_4_966, output_4_7, output_3_966;
mixer gate_output_3_966(.a(output_4_966), .b(output_4_7), .y(output_3_966));
wire output_5_966, output_5_7, output_4_966;
mixer gate_output_4_966(.a(output_5_966), .b(output_5_7), .y(output_4_966));
wire output_6_966, output_6_7, output_5_966;
mixer gate_output_5_966(.a(output_6_966), .b(output_6_7), .y(output_5_966));
wire output_7_966, output_7_7, output_6_966;
mixer gate_output_6_966(.a(output_7_966), .b(output_7_7), .y(output_6_966));
wire output_8_966, output_8_7, output_7_966;
mixer gate_output_7_966(.a(output_8_966), .b(output_8_7), .y(output_7_966));
wire output_9_966, output_9_7, output_8_966;
mixer gate_output_8_966(.a(output_9_966), .b(output_9_7), .y(output_8_966));
wire output_10_966, output_10_7, output_9_966;
mixer gate_output_9_966(.a(output_10_966), .b(output_10_7), .y(output_9_966));
wire output_11_966, output_11_7, output_10_966;
mixer gate_output_10_966(.a(output_11_966), .b(output_11_7), .y(output_10_966));
wire output_12_966, output_12_7, output_11_966;
mixer gate_output_11_966(.a(output_12_966), .b(output_12_7), .y(output_11_966));
wire output_13_966, output_13_7, output_12_966;
mixer gate_output_12_966(.a(output_13_966), .b(output_13_7), .y(output_12_966));
wire output_14_966, output_14_7, output_13_966;
mixer gate_output_13_966(.a(output_14_966), .b(output_14_7), .y(output_13_966));
wire output_15_966, output_15_7, output_14_966;
mixer gate_output_14_966(.a(output_15_966), .b(output_15_7), .y(output_14_966));
wire output_16_966, output_16_7, output_15_966;
mixer gate_output_15_966(.a(output_16_966), .b(output_16_7), .y(output_15_966));
wire output_1_967, output_1_8, output_0_967;
mixer gate_output_0_967(.a(output_1_967), .b(output_1_8), .y(output_0_967));
wire output_2_967, output_2_8, output_1_967;
mixer gate_output_1_967(.a(output_2_967), .b(output_2_8), .y(output_1_967));
wire output_3_967, output_3_8, output_2_967;
mixer gate_output_2_967(.a(output_3_967), .b(output_3_8), .y(output_2_967));
wire output_4_967, output_4_8, output_3_967;
mixer gate_output_3_967(.a(output_4_967), .b(output_4_8), .y(output_3_967));
wire output_5_967, output_5_8, output_4_967;
mixer gate_output_4_967(.a(output_5_967), .b(output_5_8), .y(output_4_967));
wire output_6_967, output_6_8, output_5_967;
mixer gate_output_5_967(.a(output_6_967), .b(output_6_8), .y(output_5_967));
wire output_7_967, output_7_8, output_6_967;
mixer gate_output_6_967(.a(output_7_967), .b(output_7_8), .y(output_6_967));
wire output_8_967, output_8_8, output_7_967;
mixer gate_output_7_967(.a(output_8_967), .b(output_8_8), .y(output_7_967));
wire output_9_967, output_9_8, output_8_967;
mixer gate_output_8_967(.a(output_9_967), .b(output_9_8), .y(output_8_967));
wire output_10_967, output_10_8, output_9_967;
mixer gate_output_9_967(.a(output_10_967), .b(output_10_8), .y(output_9_967));
wire output_11_967, output_11_8, output_10_967;
mixer gate_output_10_967(.a(output_11_967), .b(output_11_8), .y(output_10_967));
wire output_12_967, output_12_8, output_11_967;
mixer gate_output_11_967(.a(output_12_967), .b(output_12_8), .y(output_11_967));
wire output_13_967, output_13_8, output_12_967;
mixer gate_output_12_967(.a(output_13_967), .b(output_13_8), .y(output_12_967));
wire output_14_967, output_14_8, output_13_967;
mixer gate_output_13_967(.a(output_14_967), .b(output_14_8), .y(output_13_967));
wire output_15_967, output_15_8, output_14_967;
mixer gate_output_14_967(.a(output_15_967), .b(output_15_8), .y(output_14_967));
wire output_16_967, output_16_8, output_15_967;
mixer gate_output_15_967(.a(output_16_967), .b(output_16_8), .y(output_15_967));
wire output_1_968, output_1_9, output_0_968;
mixer gate_output_0_968(.a(output_1_968), .b(output_1_9), .y(output_0_968));
wire output_2_968, output_2_9, output_1_968;
mixer gate_output_1_968(.a(output_2_968), .b(output_2_9), .y(output_1_968));
wire output_3_968, output_3_9, output_2_968;
mixer gate_output_2_968(.a(output_3_968), .b(output_3_9), .y(output_2_968));
wire output_4_968, output_4_9, output_3_968;
mixer gate_output_3_968(.a(output_4_968), .b(output_4_9), .y(output_3_968));
wire output_5_968, output_5_9, output_4_968;
mixer gate_output_4_968(.a(output_5_968), .b(output_5_9), .y(output_4_968));
wire output_6_968, output_6_9, output_5_968;
mixer gate_output_5_968(.a(output_6_968), .b(output_6_9), .y(output_5_968));
wire output_7_968, output_7_9, output_6_968;
mixer gate_output_6_968(.a(output_7_968), .b(output_7_9), .y(output_6_968));
wire output_8_968, output_8_9, output_7_968;
mixer gate_output_7_968(.a(output_8_968), .b(output_8_9), .y(output_7_968));
wire output_9_968, output_9_9, output_8_968;
mixer gate_output_8_968(.a(output_9_968), .b(output_9_9), .y(output_8_968));
wire output_10_968, output_10_9, output_9_968;
mixer gate_output_9_968(.a(output_10_968), .b(output_10_9), .y(output_9_968));
wire output_11_968, output_11_9, output_10_968;
mixer gate_output_10_968(.a(output_11_968), .b(output_11_9), .y(output_10_968));
wire output_12_968, output_12_9, output_11_968;
mixer gate_output_11_968(.a(output_12_968), .b(output_12_9), .y(output_11_968));
wire output_13_968, output_13_9, output_12_968;
mixer gate_output_12_968(.a(output_13_968), .b(output_13_9), .y(output_12_968));
wire output_14_968, output_14_9, output_13_968;
mixer gate_output_13_968(.a(output_14_968), .b(output_14_9), .y(output_13_968));
wire output_15_968, output_15_9, output_14_968;
mixer gate_output_14_968(.a(output_15_968), .b(output_15_9), .y(output_14_968));
wire output_16_968, output_16_9, output_15_968;
mixer gate_output_15_968(.a(output_16_968), .b(output_16_9), .y(output_15_968));
wire output_1_969, output_1_10, output_0_969;
mixer gate_output_0_969(.a(output_1_969), .b(output_1_10), .y(output_0_969));
wire output_2_969, output_2_10, output_1_969;
mixer gate_output_1_969(.a(output_2_969), .b(output_2_10), .y(output_1_969));
wire output_3_969, output_3_10, output_2_969;
mixer gate_output_2_969(.a(output_3_969), .b(output_3_10), .y(output_2_969));
wire output_4_969, output_4_10, output_3_969;
mixer gate_output_3_969(.a(output_4_969), .b(output_4_10), .y(output_3_969));
wire output_5_969, output_5_10, output_4_969;
mixer gate_output_4_969(.a(output_5_969), .b(output_5_10), .y(output_4_969));
wire output_6_969, output_6_10, output_5_969;
mixer gate_output_5_969(.a(output_6_969), .b(output_6_10), .y(output_5_969));
wire output_7_969, output_7_10, output_6_969;
mixer gate_output_6_969(.a(output_7_969), .b(output_7_10), .y(output_6_969));
wire output_8_969, output_8_10, output_7_969;
mixer gate_output_7_969(.a(output_8_969), .b(output_8_10), .y(output_7_969));
wire output_9_969, output_9_10, output_8_969;
mixer gate_output_8_969(.a(output_9_969), .b(output_9_10), .y(output_8_969));
wire output_10_969, output_10_10, output_9_969;
mixer gate_output_9_969(.a(output_10_969), .b(output_10_10), .y(output_9_969));
wire output_11_969, output_11_10, output_10_969;
mixer gate_output_10_969(.a(output_11_969), .b(output_11_10), .y(output_10_969));
wire output_12_969, output_12_10, output_11_969;
mixer gate_output_11_969(.a(output_12_969), .b(output_12_10), .y(output_11_969));
wire output_13_969, output_13_10, output_12_969;
mixer gate_output_12_969(.a(output_13_969), .b(output_13_10), .y(output_12_969));
wire output_14_969, output_14_10, output_13_969;
mixer gate_output_13_969(.a(output_14_969), .b(output_14_10), .y(output_13_969));
wire output_15_969, output_15_10, output_14_969;
mixer gate_output_14_969(.a(output_15_969), .b(output_15_10), .y(output_14_969));
wire output_16_969, output_16_10, output_15_969;
mixer gate_output_15_969(.a(output_16_969), .b(output_16_10), .y(output_15_969));
wire output_1_970, output_1_11, output_0_970;
mixer gate_output_0_970(.a(output_1_970), .b(output_1_11), .y(output_0_970));
wire output_2_970, output_2_11, output_1_970;
mixer gate_output_1_970(.a(output_2_970), .b(output_2_11), .y(output_1_970));
wire output_3_970, output_3_11, output_2_970;
mixer gate_output_2_970(.a(output_3_970), .b(output_3_11), .y(output_2_970));
wire output_4_970, output_4_11, output_3_970;
mixer gate_output_3_970(.a(output_4_970), .b(output_4_11), .y(output_3_970));
wire output_5_970, output_5_11, output_4_970;
mixer gate_output_4_970(.a(output_5_970), .b(output_5_11), .y(output_4_970));
wire output_6_970, output_6_11, output_5_970;
mixer gate_output_5_970(.a(output_6_970), .b(output_6_11), .y(output_5_970));
wire output_7_970, output_7_11, output_6_970;
mixer gate_output_6_970(.a(output_7_970), .b(output_7_11), .y(output_6_970));
wire output_8_970, output_8_11, output_7_970;
mixer gate_output_7_970(.a(output_8_970), .b(output_8_11), .y(output_7_970));
wire output_9_970, output_9_11, output_8_970;
mixer gate_output_8_970(.a(output_9_970), .b(output_9_11), .y(output_8_970));
wire output_10_970, output_10_11, output_9_970;
mixer gate_output_9_970(.a(output_10_970), .b(output_10_11), .y(output_9_970));
wire output_11_970, output_11_11, output_10_970;
mixer gate_output_10_970(.a(output_11_970), .b(output_11_11), .y(output_10_970));
wire output_12_970, output_12_11, output_11_970;
mixer gate_output_11_970(.a(output_12_970), .b(output_12_11), .y(output_11_970));
wire output_13_970, output_13_11, output_12_970;
mixer gate_output_12_970(.a(output_13_970), .b(output_13_11), .y(output_12_970));
wire output_14_970, output_14_11, output_13_970;
mixer gate_output_13_970(.a(output_14_970), .b(output_14_11), .y(output_13_970));
wire output_15_970, output_15_11, output_14_970;
mixer gate_output_14_970(.a(output_15_970), .b(output_15_11), .y(output_14_970));
wire output_16_970, output_16_11, output_15_970;
mixer gate_output_15_970(.a(output_16_970), .b(output_16_11), .y(output_15_970));
wire output_1_971, output_1_12, output_0_971;
mixer gate_output_0_971(.a(output_1_971), .b(output_1_12), .y(output_0_971));
wire output_2_971, output_2_12, output_1_971;
mixer gate_output_1_971(.a(output_2_971), .b(output_2_12), .y(output_1_971));
wire output_3_971, output_3_12, output_2_971;
mixer gate_output_2_971(.a(output_3_971), .b(output_3_12), .y(output_2_971));
wire output_4_971, output_4_12, output_3_971;
mixer gate_output_3_971(.a(output_4_971), .b(output_4_12), .y(output_3_971));
wire output_5_971, output_5_12, output_4_971;
mixer gate_output_4_971(.a(output_5_971), .b(output_5_12), .y(output_4_971));
wire output_6_971, output_6_12, output_5_971;
mixer gate_output_5_971(.a(output_6_971), .b(output_6_12), .y(output_5_971));
wire output_7_971, output_7_12, output_6_971;
mixer gate_output_6_971(.a(output_7_971), .b(output_7_12), .y(output_6_971));
wire output_8_971, output_8_12, output_7_971;
mixer gate_output_7_971(.a(output_8_971), .b(output_8_12), .y(output_7_971));
wire output_9_971, output_9_12, output_8_971;
mixer gate_output_8_971(.a(output_9_971), .b(output_9_12), .y(output_8_971));
wire output_10_971, output_10_12, output_9_971;
mixer gate_output_9_971(.a(output_10_971), .b(output_10_12), .y(output_9_971));
wire output_11_971, output_11_12, output_10_971;
mixer gate_output_10_971(.a(output_11_971), .b(output_11_12), .y(output_10_971));
wire output_12_971, output_12_12, output_11_971;
mixer gate_output_11_971(.a(output_12_971), .b(output_12_12), .y(output_11_971));
wire output_13_971, output_13_12, output_12_971;
mixer gate_output_12_971(.a(output_13_971), .b(output_13_12), .y(output_12_971));
wire output_14_971, output_14_12, output_13_971;
mixer gate_output_13_971(.a(output_14_971), .b(output_14_12), .y(output_13_971));
wire output_15_971, output_15_12, output_14_971;
mixer gate_output_14_971(.a(output_15_971), .b(output_15_12), .y(output_14_971));
wire output_16_971, output_16_12, output_15_971;
mixer gate_output_15_971(.a(output_16_971), .b(output_16_12), .y(output_15_971));
wire output_1_972, output_1_13, output_0_972;
mixer gate_output_0_972(.a(output_1_972), .b(output_1_13), .y(output_0_972));
wire output_2_972, output_2_13, output_1_972;
mixer gate_output_1_972(.a(output_2_972), .b(output_2_13), .y(output_1_972));
wire output_3_972, output_3_13, output_2_972;
mixer gate_output_2_972(.a(output_3_972), .b(output_3_13), .y(output_2_972));
wire output_4_972, output_4_13, output_3_972;
mixer gate_output_3_972(.a(output_4_972), .b(output_4_13), .y(output_3_972));
wire output_5_972, output_5_13, output_4_972;
mixer gate_output_4_972(.a(output_5_972), .b(output_5_13), .y(output_4_972));
wire output_6_972, output_6_13, output_5_972;
mixer gate_output_5_972(.a(output_6_972), .b(output_6_13), .y(output_5_972));
wire output_7_972, output_7_13, output_6_972;
mixer gate_output_6_972(.a(output_7_972), .b(output_7_13), .y(output_6_972));
wire output_8_972, output_8_13, output_7_972;
mixer gate_output_7_972(.a(output_8_972), .b(output_8_13), .y(output_7_972));
wire output_9_972, output_9_13, output_8_972;
mixer gate_output_8_972(.a(output_9_972), .b(output_9_13), .y(output_8_972));
wire output_10_972, output_10_13, output_9_972;
mixer gate_output_9_972(.a(output_10_972), .b(output_10_13), .y(output_9_972));
wire output_11_972, output_11_13, output_10_972;
mixer gate_output_10_972(.a(output_11_972), .b(output_11_13), .y(output_10_972));
wire output_12_972, output_12_13, output_11_972;
mixer gate_output_11_972(.a(output_12_972), .b(output_12_13), .y(output_11_972));
wire output_13_972, output_13_13, output_12_972;
mixer gate_output_12_972(.a(output_13_972), .b(output_13_13), .y(output_12_972));
wire output_14_972, output_14_13, output_13_972;
mixer gate_output_13_972(.a(output_14_972), .b(output_14_13), .y(output_13_972));
wire output_15_972, output_15_13, output_14_972;
mixer gate_output_14_972(.a(output_15_972), .b(output_15_13), .y(output_14_972));
wire output_16_972, output_16_13, output_15_972;
mixer gate_output_15_972(.a(output_16_972), .b(output_16_13), .y(output_15_972));
wire output_1_973, output_1_14, output_0_973;
mixer gate_output_0_973(.a(output_1_973), .b(output_1_14), .y(output_0_973));
wire output_2_973, output_2_14, output_1_973;
mixer gate_output_1_973(.a(output_2_973), .b(output_2_14), .y(output_1_973));
wire output_3_973, output_3_14, output_2_973;
mixer gate_output_2_973(.a(output_3_973), .b(output_3_14), .y(output_2_973));
wire output_4_973, output_4_14, output_3_973;
mixer gate_output_3_973(.a(output_4_973), .b(output_4_14), .y(output_3_973));
wire output_5_973, output_5_14, output_4_973;
mixer gate_output_4_973(.a(output_5_973), .b(output_5_14), .y(output_4_973));
wire output_6_973, output_6_14, output_5_973;
mixer gate_output_5_973(.a(output_6_973), .b(output_6_14), .y(output_5_973));
wire output_7_973, output_7_14, output_6_973;
mixer gate_output_6_973(.a(output_7_973), .b(output_7_14), .y(output_6_973));
wire output_8_973, output_8_14, output_7_973;
mixer gate_output_7_973(.a(output_8_973), .b(output_8_14), .y(output_7_973));
wire output_9_973, output_9_14, output_8_973;
mixer gate_output_8_973(.a(output_9_973), .b(output_9_14), .y(output_8_973));
wire output_10_973, output_10_14, output_9_973;
mixer gate_output_9_973(.a(output_10_973), .b(output_10_14), .y(output_9_973));
wire output_11_973, output_11_14, output_10_973;
mixer gate_output_10_973(.a(output_11_973), .b(output_11_14), .y(output_10_973));
wire output_12_973, output_12_14, output_11_973;
mixer gate_output_11_973(.a(output_12_973), .b(output_12_14), .y(output_11_973));
wire output_13_973, output_13_14, output_12_973;
mixer gate_output_12_973(.a(output_13_973), .b(output_13_14), .y(output_12_973));
wire output_14_973, output_14_14, output_13_973;
mixer gate_output_13_973(.a(output_14_973), .b(output_14_14), .y(output_13_973));
wire output_15_973, output_15_14, output_14_973;
mixer gate_output_14_973(.a(output_15_973), .b(output_15_14), .y(output_14_973));
wire output_16_973, output_16_14, output_15_973;
mixer gate_output_15_973(.a(output_16_973), .b(output_16_14), .y(output_15_973));
wire output_1_974, output_1_15, output_0_974;
mixer gate_output_0_974(.a(output_1_974), .b(output_1_15), .y(output_0_974));
wire output_2_974, output_2_15, output_1_974;
mixer gate_output_1_974(.a(output_2_974), .b(output_2_15), .y(output_1_974));
wire output_3_974, output_3_15, output_2_974;
mixer gate_output_2_974(.a(output_3_974), .b(output_3_15), .y(output_2_974));
wire output_4_974, output_4_15, output_3_974;
mixer gate_output_3_974(.a(output_4_974), .b(output_4_15), .y(output_3_974));
wire output_5_974, output_5_15, output_4_974;
mixer gate_output_4_974(.a(output_5_974), .b(output_5_15), .y(output_4_974));
wire output_6_974, output_6_15, output_5_974;
mixer gate_output_5_974(.a(output_6_974), .b(output_6_15), .y(output_5_974));
wire output_7_974, output_7_15, output_6_974;
mixer gate_output_6_974(.a(output_7_974), .b(output_7_15), .y(output_6_974));
wire output_8_974, output_8_15, output_7_974;
mixer gate_output_7_974(.a(output_8_974), .b(output_8_15), .y(output_7_974));
wire output_9_974, output_9_15, output_8_974;
mixer gate_output_8_974(.a(output_9_974), .b(output_9_15), .y(output_8_974));
wire output_10_974, output_10_15, output_9_974;
mixer gate_output_9_974(.a(output_10_974), .b(output_10_15), .y(output_9_974));
wire output_11_974, output_11_15, output_10_974;
mixer gate_output_10_974(.a(output_11_974), .b(output_11_15), .y(output_10_974));
wire output_12_974, output_12_15, output_11_974;
mixer gate_output_11_974(.a(output_12_974), .b(output_12_15), .y(output_11_974));
wire output_13_974, output_13_15, output_12_974;
mixer gate_output_12_974(.a(output_13_974), .b(output_13_15), .y(output_12_974));
wire output_14_974, output_14_15, output_13_974;
mixer gate_output_13_974(.a(output_14_974), .b(output_14_15), .y(output_13_974));
wire output_15_974, output_15_15, output_14_974;
mixer gate_output_14_974(.a(output_15_974), .b(output_15_15), .y(output_14_974));
wire output_16_974, output_16_15, output_15_974;
mixer gate_output_15_974(.a(output_16_974), .b(output_16_15), .y(output_15_974));
wire output_1_975, output_1_0, output_0_975;
mixer gate_output_0_975(.a(output_1_975), .b(output_1_0), .y(output_0_975));
wire output_2_975, output_2_0, output_1_975;
mixer gate_output_1_975(.a(output_2_975), .b(output_2_0), .y(output_1_975));
wire output_3_975, output_3_0, output_2_975;
mixer gate_output_2_975(.a(output_3_975), .b(output_3_0), .y(output_2_975));
wire output_4_975, output_4_0, output_3_975;
mixer gate_output_3_975(.a(output_4_975), .b(output_4_0), .y(output_3_975));
wire output_5_975, output_5_0, output_4_975;
mixer gate_output_4_975(.a(output_5_975), .b(output_5_0), .y(output_4_975));
wire output_6_975, output_6_0, output_5_975;
mixer gate_output_5_975(.a(output_6_975), .b(output_6_0), .y(output_5_975));
wire output_7_975, output_7_0, output_6_975;
mixer gate_output_6_975(.a(output_7_975), .b(output_7_0), .y(output_6_975));
wire output_8_975, output_8_0, output_7_975;
mixer gate_output_7_975(.a(output_8_975), .b(output_8_0), .y(output_7_975));
wire output_9_975, output_9_0, output_8_975;
mixer gate_output_8_975(.a(output_9_975), .b(output_9_0), .y(output_8_975));
wire output_10_975, output_10_0, output_9_975;
mixer gate_output_9_975(.a(output_10_975), .b(output_10_0), .y(output_9_975));
wire output_11_975, output_11_0, output_10_975;
mixer gate_output_10_975(.a(output_11_975), .b(output_11_0), .y(output_10_975));
wire output_12_975, output_12_0, output_11_975;
mixer gate_output_11_975(.a(output_12_975), .b(output_12_0), .y(output_11_975));
wire output_13_975, output_13_0, output_12_975;
mixer gate_output_12_975(.a(output_13_975), .b(output_13_0), .y(output_12_975));
wire output_14_975, output_14_0, output_13_975;
mixer gate_output_13_975(.a(output_14_975), .b(output_14_0), .y(output_13_975));
wire output_15_975, output_15_0, output_14_975;
mixer gate_output_14_975(.a(output_15_975), .b(output_15_0), .y(output_14_975));
wire output_16_975, output_16_0, output_15_975;
mixer gate_output_15_975(.a(output_16_975), .b(output_16_0), .y(output_15_975));
wire output_1_976, output_1_1, output_0_976;
mixer gate_output_0_976(.a(output_1_976), .b(output_1_1), .y(output_0_976));
wire output_2_976, output_2_1, output_1_976;
mixer gate_output_1_976(.a(output_2_976), .b(output_2_1), .y(output_1_976));
wire output_3_976, output_3_1, output_2_976;
mixer gate_output_2_976(.a(output_3_976), .b(output_3_1), .y(output_2_976));
wire output_4_976, output_4_1, output_3_976;
mixer gate_output_3_976(.a(output_4_976), .b(output_4_1), .y(output_3_976));
wire output_5_976, output_5_1, output_4_976;
mixer gate_output_4_976(.a(output_5_976), .b(output_5_1), .y(output_4_976));
wire output_6_976, output_6_1, output_5_976;
mixer gate_output_5_976(.a(output_6_976), .b(output_6_1), .y(output_5_976));
wire output_7_976, output_7_1, output_6_976;
mixer gate_output_6_976(.a(output_7_976), .b(output_7_1), .y(output_6_976));
wire output_8_976, output_8_1, output_7_976;
mixer gate_output_7_976(.a(output_8_976), .b(output_8_1), .y(output_7_976));
wire output_9_976, output_9_1, output_8_976;
mixer gate_output_8_976(.a(output_9_976), .b(output_9_1), .y(output_8_976));
wire output_10_976, output_10_1, output_9_976;
mixer gate_output_9_976(.a(output_10_976), .b(output_10_1), .y(output_9_976));
wire output_11_976, output_11_1, output_10_976;
mixer gate_output_10_976(.a(output_11_976), .b(output_11_1), .y(output_10_976));
wire output_12_976, output_12_1, output_11_976;
mixer gate_output_11_976(.a(output_12_976), .b(output_12_1), .y(output_11_976));
wire output_13_976, output_13_1, output_12_976;
mixer gate_output_12_976(.a(output_13_976), .b(output_13_1), .y(output_12_976));
wire output_14_976, output_14_1, output_13_976;
mixer gate_output_13_976(.a(output_14_976), .b(output_14_1), .y(output_13_976));
wire output_15_976, output_15_1, output_14_976;
mixer gate_output_14_976(.a(output_15_976), .b(output_15_1), .y(output_14_976));
wire output_16_976, output_16_1, output_15_976;
mixer gate_output_15_976(.a(output_16_976), .b(output_16_1), .y(output_15_976));
wire output_1_977, output_1_2, output_0_977;
mixer gate_output_0_977(.a(output_1_977), .b(output_1_2), .y(output_0_977));
wire output_2_977, output_2_2, output_1_977;
mixer gate_output_1_977(.a(output_2_977), .b(output_2_2), .y(output_1_977));
wire output_3_977, output_3_2, output_2_977;
mixer gate_output_2_977(.a(output_3_977), .b(output_3_2), .y(output_2_977));
wire output_4_977, output_4_2, output_3_977;
mixer gate_output_3_977(.a(output_4_977), .b(output_4_2), .y(output_3_977));
wire output_5_977, output_5_2, output_4_977;
mixer gate_output_4_977(.a(output_5_977), .b(output_5_2), .y(output_4_977));
wire output_6_977, output_6_2, output_5_977;
mixer gate_output_5_977(.a(output_6_977), .b(output_6_2), .y(output_5_977));
wire output_7_977, output_7_2, output_6_977;
mixer gate_output_6_977(.a(output_7_977), .b(output_7_2), .y(output_6_977));
wire output_8_977, output_8_2, output_7_977;
mixer gate_output_7_977(.a(output_8_977), .b(output_8_2), .y(output_7_977));
wire output_9_977, output_9_2, output_8_977;
mixer gate_output_8_977(.a(output_9_977), .b(output_9_2), .y(output_8_977));
wire output_10_977, output_10_2, output_9_977;
mixer gate_output_9_977(.a(output_10_977), .b(output_10_2), .y(output_9_977));
wire output_11_977, output_11_2, output_10_977;
mixer gate_output_10_977(.a(output_11_977), .b(output_11_2), .y(output_10_977));
wire output_12_977, output_12_2, output_11_977;
mixer gate_output_11_977(.a(output_12_977), .b(output_12_2), .y(output_11_977));
wire output_13_977, output_13_2, output_12_977;
mixer gate_output_12_977(.a(output_13_977), .b(output_13_2), .y(output_12_977));
wire output_14_977, output_14_2, output_13_977;
mixer gate_output_13_977(.a(output_14_977), .b(output_14_2), .y(output_13_977));
wire output_15_977, output_15_2, output_14_977;
mixer gate_output_14_977(.a(output_15_977), .b(output_15_2), .y(output_14_977));
wire output_16_977, output_16_2, output_15_977;
mixer gate_output_15_977(.a(output_16_977), .b(output_16_2), .y(output_15_977));
wire output_1_978, output_1_3, output_0_978;
mixer gate_output_0_978(.a(output_1_978), .b(output_1_3), .y(output_0_978));
wire output_2_978, output_2_3, output_1_978;
mixer gate_output_1_978(.a(output_2_978), .b(output_2_3), .y(output_1_978));
wire output_3_978, output_3_3, output_2_978;
mixer gate_output_2_978(.a(output_3_978), .b(output_3_3), .y(output_2_978));
wire output_4_978, output_4_3, output_3_978;
mixer gate_output_3_978(.a(output_4_978), .b(output_4_3), .y(output_3_978));
wire output_5_978, output_5_3, output_4_978;
mixer gate_output_4_978(.a(output_5_978), .b(output_5_3), .y(output_4_978));
wire output_6_978, output_6_3, output_5_978;
mixer gate_output_5_978(.a(output_6_978), .b(output_6_3), .y(output_5_978));
wire output_7_978, output_7_3, output_6_978;
mixer gate_output_6_978(.a(output_7_978), .b(output_7_3), .y(output_6_978));
wire output_8_978, output_8_3, output_7_978;
mixer gate_output_7_978(.a(output_8_978), .b(output_8_3), .y(output_7_978));
wire output_9_978, output_9_3, output_8_978;
mixer gate_output_8_978(.a(output_9_978), .b(output_9_3), .y(output_8_978));
wire output_10_978, output_10_3, output_9_978;
mixer gate_output_9_978(.a(output_10_978), .b(output_10_3), .y(output_9_978));
wire output_11_978, output_11_3, output_10_978;
mixer gate_output_10_978(.a(output_11_978), .b(output_11_3), .y(output_10_978));
wire output_12_978, output_12_3, output_11_978;
mixer gate_output_11_978(.a(output_12_978), .b(output_12_3), .y(output_11_978));
wire output_13_978, output_13_3, output_12_978;
mixer gate_output_12_978(.a(output_13_978), .b(output_13_3), .y(output_12_978));
wire output_14_978, output_14_3, output_13_978;
mixer gate_output_13_978(.a(output_14_978), .b(output_14_3), .y(output_13_978));
wire output_15_978, output_15_3, output_14_978;
mixer gate_output_14_978(.a(output_15_978), .b(output_15_3), .y(output_14_978));
wire output_16_978, output_16_3, output_15_978;
mixer gate_output_15_978(.a(output_16_978), .b(output_16_3), .y(output_15_978));
wire output_1_979, output_1_4, output_0_979;
mixer gate_output_0_979(.a(output_1_979), .b(output_1_4), .y(output_0_979));
wire output_2_979, output_2_4, output_1_979;
mixer gate_output_1_979(.a(output_2_979), .b(output_2_4), .y(output_1_979));
wire output_3_979, output_3_4, output_2_979;
mixer gate_output_2_979(.a(output_3_979), .b(output_3_4), .y(output_2_979));
wire output_4_979, output_4_4, output_3_979;
mixer gate_output_3_979(.a(output_4_979), .b(output_4_4), .y(output_3_979));
wire output_5_979, output_5_4, output_4_979;
mixer gate_output_4_979(.a(output_5_979), .b(output_5_4), .y(output_4_979));
wire output_6_979, output_6_4, output_5_979;
mixer gate_output_5_979(.a(output_6_979), .b(output_6_4), .y(output_5_979));
wire output_7_979, output_7_4, output_6_979;
mixer gate_output_6_979(.a(output_7_979), .b(output_7_4), .y(output_6_979));
wire output_8_979, output_8_4, output_7_979;
mixer gate_output_7_979(.a(output_8_979), .b(output_8_4), .y(output_7_979));
wire output_9_979, output_9_4, output_8_979;
mixer gate_output_8_979(.a(output_9_979), .b(output_9_4), .y(output_8_979));
wire output_10_979, output_10_4, output_9_979;
mixer gate_output_9_979(.a(output_10_979), .b(output_10_4), .y(output_9_979));
wire output_11_979, output_11_4, output_10_979;
mixer gate_output_10_979(.a(output_11_979), .b(output_11_4), .y(output_10_979));
wire output_12_979, output_12_4, output_11_979;
mixer gate_output_11_979(.a(output_12_979), .b(output_12_4), .y(output_11_979));
wire output_13_979, output_13_4, output_12_979;
mixer gate_output_12_979(.a(output_13_979), .b(output_13_4), .y(output_12_979));
wire output_14_979, output_14_4, output_13_979;
mixer gate_output_13_979(.a(output_14_979), .b(output_14_4), .y(output_13_979));
wire output_15_979, output_15_4, output_14_979;
mixer gate_output_14_979(.a(output_15_979), .b(output_15_4), .y(output_14_979));
wire output_16_979, output_16_4, output_15_979;
mixer gate_output_15_979(.a(output_16_979), .b(output_16_4), .y(output_15_979));
wire output_1_980, output_1_5, output_0_980;
mixer gate_output_0_980(.a(output_1_980), .b(output_1_5), .y(output_0_980));
wire output_2_980, output_2_5, output_1_980;
mixer gate_output_1_980(.a(output_2_980), .b(output_2_5), .y(output_1_980));
wire output_3_980, output_3_5, output_2_980;
mixer gate_output_2_980(.a(output_3_980), .b(output_3_5), .y(output_2_980));
wire output_4_980, output_4_5, output_3_980;
mixer gate_output_3_980(.a(output_4_980), .b(output_4_5), .y(output_3_980));
wire output_5_980, output_5_5, output_4_980;
mixer gate_output_4_980(.a(output_5_980), .b(output_5_5), .y(output_4_980));
wire output_6_980, output_6_5, output_5_980;
mixer gate_output_5_980(.a(output_6_980), .b(output_6_5), .y(output_5_980));
wire output_7_980, output_7_5, output_6_980;
mixer gate_output_6_980(.a(output_7_980), .b(output_7_5), .y(output_6_980));
wire output_8_980, output_8_5, output_7_980;
mixer gate_output_7_980(.a(output_8_980), .b(output_8_5), .y(output_7_980));
wire output_9_980, output_9_5, output_8_980;
mixer gate_output_8_980(.a(output_9_980), .b(output_9_5), .y(output_8_980));
wire output_10_980, output_10_5, output_9_980;
mixer gate_output_9_980(.a(output_10_980), .b(output_10_5), .y(output_9_980));
wire output_11_980, output_11_5, output_10_980;
mixer gate_output_10_980(.a(output_11_980), .b(output_11_5), .y(output_10_980));
wire output_12_980, output_12_5, output_11_980;
mixer gate_output_11_980(.a(output_12_980), .b(output_12_5), .y(output_11_980));
wire output_13_980, output_13_5, output_12_980;
mixer gate_output_12_980(.a(output_13_980), .b(output_13_5), .y(output_12_980));
wire output_14_980, output_14_5, output_13_980;
mixer gate_output_13_980(.a(output_14_980), .b(output_14_5), .y(output_13_980));
wire output_15_980, output_15_5, output_14_980;
mixer gate_output_14_980(.a(output_15_980), .b(output_15_5), .y(output_14_980));
wire output_16_980, output_16_5, output_15_980;
mixer gate_output_15_980(.a(output_16_980), .b(output_16_5), .y(output_15_980));
wire output_1_981, output_1_6, output_0_981;
mixer gate_output_0_981(.a(output_1_981), .b(output_1_6), .y(output_0_981));
wire output_2_981, output_2_6, output_1_981;
mixer gate_output_1_981(.a(output_2_981), .b(output_2_6), .y(output_1_981));
wire output_3_981, output_3_6, output_2_981;
mixer gate_output_2_981(.a(output_3_981), .b(output_3_6), .y(output_2_981));
wire output_4_981, output_4_6, output_3_981;
mixer gate_output_3_981(.a(output_4_981), .b(output_4_6), .y(output_3_981));
wire output_5_981, output_5_6, output_4_981;
mixer gate_output_4_981(.a(output_5_981), .b(output_5_6), .y(output_4_981));
wire output_6_981, output_6_6, output_5_981;
mixer gate_output_5_981(.a(output_6_981), .b(output_6_6), .y(output_5_981));
wire output_7_981, output_7_6, output_6_981;
mixer gate_output_6_981(.a(output_7_981), .b(output_7_6), .y(output_6_981));
wire output_8_981, output_8_6, output_7_981;
mixer gate_output_7_981(.a(output_8_981), .b(output_8_6), .y(output_7_981));
wire output_9_981, output_9_6, output_8_981;
mixer gate_output_8_981(.a(output_9_981), .b(output_9_6), .y(output_8_981));
wire output_10_981, output_10_6, output_9_981;
mixer gate_output_9_981(.a(output_10_981), .b(output_10_6), .y(output_9_981));
wire output_11_981, output_11_6, output_10_981;
mixer gate_output_10_981(.a(output_11_981), .b(output_11_6), .y(output_10_981));
wire output_12_981, output_12_6, output_11_981;
mixer gate_output_11_981(.a(output_12_981), .b(output_12_6), .y(output_11_981));
wire output_13_981, output_13_6, output_12_981;
mixer gate_output_12_981(.a(output_13_981), .b(output_13_6), .y(output_12_981));
wire output_14_981, output_14_6, output_13_981;
mixer gate_output_13_981(.a(output_14_981), .b(output_14_6), .y(output_13_981));
wire output_15_981, output_15_6, output_14_981;
mixer gate_output_14_981(.a(output_15_981), .b(output_15_6), .y(output_14_981));
wire output_16_981, output_16_6, output_15_981;
mixer gate_output_15_981(.a(output_16_981), .b(output_16_6), .y(output_15_981));
wire output_1_982, output_1_7, output_0_982;
mixer gate_output_0_982(.a(output_1_982), .b(output_1_7), .y(output_0_982));
wire output_2_982, output_2_7, output_1_982;
mixer gate_output_1_982(.a(output_2_982), .b(output_2_7), .y(output_1_982));
wire output_3_982, output_3_7, output_2_982;
mixer gate_output_2_982(.a(output_3_982), .b(output_3_7), .y(output_2_982));
wire output_4_982, output_4_7, output_3_982;
mixer gate_output_3_982(.a(output_4_982), .b(output_4_7), .y(output_3_982));
wire output_5_982, output_5_7, output_4_982;
mixer gate_output_4_982(.a(output_5_982), .b(output_5_7), .y(output_4_982));
wire output_6_982, output_6_7, output_5_982;
mixer gate_output_5_982(.a(output_6_982), .b(output_6_7), .y(output_5_982));
wire output_7_982, output_7_7, output_6_982;
mixer gate_output_6_982(.a(output_7_982), .b(output_7_7), .y(output_6_982));
wire output_8_982, output_8_7, output_7_982;
mixer gate_output_7_982(.a(output_8_982), .b(output_8_7), .y(output_7_982));
wire output_9_982, output_9_7, output_8_982;
mixer gate_output_8_982(.a(output_9_982), .b(output_9_7), .y(output_8_982));
wire output_10_982, output_10_7, output_9_982;
mixer gate_output_9_982(.a(output_10_982), .b(output_10_7), .y(output_9_982));
wire output_11_982, output_11_7, output_10_982;
mixer gate_output_10_982(.a(output_11_982), .b(output_11_7), .y(output_10_982));
wire output_12_982, output_12_7, output_11_982;
mixer gate_output_11_982(.a(output_12_982), .b(output_12_7), .y(output_11_982));
wire output_13_982, output_13_7, output_12_982;
mixer gate_output_12_982(.a(output_13_982), .b(output_13_7), .y(output_12_982));
wire output_14_982, output_14_7, output_13_982;
mixer gate_output_13_982(.a(output_14_982), .b(output_14_7), .y(output_13_982));
wire output_15_982, output_15_7, output_14_982;
mixer gate_output_14_982(.a(output_15_982), .b(output_15_7), .y(output_14_982));
wire output_16_982, output_16_7, output_15_982;
mixer gate_output_15_982(.a(output_16_982), .b(output_16_7), .y(output_15_982));
wire output_1_983, output_1_8, output_0_983;
mixer gate_output_0_983(.a(output_1_983), .b(output_1_8), .y(output_0_983));
wire output_2_983, output_2_8, output_1_983;
mixer gate_output_1_983(.a(output_2_983), .b(output_2_8), .y(output_1_983));
wire output_3_983, output_3_8, output_2_983;
mixer gate_output_2_983(.a(output_3_983), .b(output_3_8), .y(output_2_983));
wire output_4_983, output_4_8, output_3_983;
mixer gate_output_3_983(.a(output_4_983), .b(output_4_8), .y(output_3_983));
wire output_5_983, output_5_8, output_4_983;
mixer gate_output_4_983(.a(output_5_983), .b(output_5_8), .y(output_4_983));
wire output_6_983, output_6_8, output_5_983;
mixer gate_output_5_983(.a(output_6_983), .b(output_6_8), .y(output_5_983));
wire output_7_983, output_7_8, output_6_983;
mixer gate_output_6_983(.a(output_7_983), .b(output_7_8), .y(output_6_983));
wire output_8_983, output_8_8, output_7_983;
mixer gate_output_7_983(.a(output_8_983), .b(output_8_8), .y(output_7_983));
wire output_9_983, output_9_8, output_8_983;
mixer gate_output_8_983(.a(output_9_983), .b(output_9_8), .y(output_8_983));
wire output_10_983, output_10_8, output_9_983;
mixer gate_output_9_983(.a(output_10_983), .b(output_10_8), .y(output_9_983));
wire output_11_983, output_11_8, output_10_983;
mixer gate_output_10_983(.a(output_11_983), .b(output_11_8), .y(output_10_983));
wire output_12_983, output_12_8, output_11_983;
mixer gate_output_11_983(.a(output_12_983), .b(output_12_8), .y(output_11_983));
wire output_13_983, output_13_8, output_12_983;
mixer gate_output_12_983(.a(output_13_983), .b(output_13_8), .y(output_12_983));
wire output_14_983, output_14_8, output_13_983;
mixer gate_output_13_983(.a(output_14_983), .b(output_14_8), .y(output_13_983));
wire output_15_983, output_15_8, output_14_983;
mixer gate_output_14_983(.a(output_15_983), .b(output_15_8), .y(output_14_983));
wire output_16_983, output_16_8, output_15_983;
mixer gate_output_15_983(.a(output_16_983), .b(output_16_8), .y(output_15_983));
wire output_1_984, output_1_9, output_0_984;
mixer gate_output_0_984(.a(output_1_984), .b(output_1_9), .y(output_0_984));
wire output_2_984, output_2_9, output_1_984;
mixer gate_output_1_984(.a(output_2_984), .b(output_2_9), .y(output_1_984));
wire output_3_984, output_3_9, output_2_984;
mixer gate_output_2_984(.a(output_3_984), .b(output_3_9), .y(output_2_984));
wire output_4_984, output_4_9, output_3_984;
mixer gate_output_3_984(.a(output_4_984), .b(output_4_9), .y(output_3_984));
wire output_5_984, output_5_9, output_4_984;
mixer gate_output_4_984(.a(output_5_984), .b(output_5_9), .y(output_4_984));
wire output_6_984, output_6_9, output_5_984;
mixer gate_output_5_984(.a(output_6_984), .b(output_6_9), .y(output_5_984));
wire output_7_984, output_7_9, output_6_984;
mixer gate_output_6_984(.a(output_7_984), .b(output_7_9), .y(output_6_984));
wire output_8_984, output_8_9, output_7_984;
mixer gate_output_7_984(.a(output_8_984), .b(output_8_9), .y(output_7_984));
wire output_9_984, output_9_9, output_8_984;
mixer gate_output_8_984(.a(output_9_984), .b(output_9_9), .y(output_8_984));
wire output_10_984, output_10_9, output_9_984;
mixer gate_output_9_984(.a(output_10_984), .b(output_10_9), .y(output_9_984));
wire output_11_984, output_11_9, output_10_984;
mixer gate_output_10_984(.a(output_11_984), .b(output_11_9), .y(output_10_984));
wire output_12_984, output_12_9, output_11_984;
mixer gate_output_11_984(.a(output_12_984), .b(output_12_9), .y(output_11_984));
wire output_13_984, output_13_9, output_12_984;
mixer gate_output_12_984(.a(output_13_984), .b(output_13_9), .y(output_12_984));
wire output_14_984, output_14_9, output_13_984;
mixer gate_output_13_984(.a(output_14_984), .b(output_14_9), .y(output_13_984));
wire output_15_984, output_15_9, output_14_984;
mixer gate_output_14_984(.a(output_15_984), .b(output_15_9), .y(output_14_984));
wire output_16_984, output_16_9, output_15_984;
mixer gate_output_15_984(.a(output_16_984), .b(output_16_9), .y(output_15_984));
wire output_1_985, output_1_10, output_0_985;
mixer gate_output_0_985(.a(output_1_985), .b(output_1_10), .y(output_0_985));
wire output_2_985, output_2_10, output_1_985;
mixer gate_output_1_985(.a(output_2_985), .b(output_2_10), .y(output_1_985));
wire output_3_985, output_3_10, output_2_985;
mixer gate_output_2_985(.a(output_3_985), .b(output_3_10), .y(output_2_985));
wire output_4_985, output_4_10, output_3_985;
mixer gate_output_3_985(.a(output_4_985), .b(output_4_10), .y(output_3_985));
wire output_5_985, output_5_10, output_4_985;
mixer gate_output_4_985(.a(output_5_985), .b(output_5_10), .y(output_4_985));
wire output_6_985, output_6_10, output_5_985;
mixer gate_output_5_985(.a(output_6_985), .b(output_6_10), .y(output_5_985));
wire output_7_985, output_7_10, output_6_985;
mixer gate_output_6_985(.a(output_7_985), .b(output_7_10), .y(output_6_985));
wire output_8_985, output_8_10, output_7_985;
mixer gate_output_7_985(.a(output_8_985), .b(output_8_10), .y(output_7_985));
wire output_9_985, output_9_10, output_8_985;
mixer gate_output_8_985(.a(output_9_985), .b(output_9_10), .y(output_8_985));
wire output_10_985, output_10_10, output_9_985;
mixer gate_output_9_985(.a(output_10_985), .b(output_10_10), .y(output_9_985));
wire output_11_985, output_11_10, output_10_985;
mixer gate_output_10_985(.a(output_11_985), .b(output_11_10), .y(output_10_985));
wire output_12_985, output_12_10, output_11_985;
mixer gate_output_11_985(.a(output_12_985), .b(output_12_10), .y(output_11_985));
wire output_13_985, output_13_10, output_12_985;
mixer gate_output_12_985(.a(output_13_985), .b(output_13_10), .y(output_12_985));
wire output_14_985, output_14_10, output_13_985;
mixer gate_output_13_985(.a(output_14_985), .b(output_14_10), .y(output_13_985));
wire output_15_985, output_15_10, output_14_985;
mixer gate_output_14_985(.a(output_15_985), .b(output_15_10), .y(output_14_985));
wire output_16_985, output_16_10, output_15_985;
mixer gate_output_15_985(.a(output_16_985), .b(output_16_10), .y(output_15_985));
wire output_1_986, output_1_11, output_0_986;
mixer gate_output_0_986(.a(output_1_986), .b(output_1_11), .y(output_0_986));
wire output_2_986, output_2_11, output_1_986;
mixer gate_output_1_986(.a(output_2_986), .b(output_2_11), .y(output_1_986));
wire output_3_986, output_3_11, output_2_986;
mixer gate_output_2_986(.a(output_3_986), .b(output_3_11), .y(output_2_986));
wire output_4_986, output_4_11, output_3_986;
mixer gate_output_3_986(.a(output_4_986), .b(output_4_11), .y(output_3_986));
wire output_5_986, output_5_11, output_4_986;
mixer gate_output_4_986(.a(output_5_986), .b(output_5_11), .y(output_4_986));
wire output_6_986, output_6_11, output_5_986;
mixer gate_output_5_986(.a(output_6_986), .b(output_6_11), .y(output_5_986));
wire output_7_986, output_7_11, output_6_986;
mixer gate_output_6_986(.a(output_7_986), .b(output_7_11), .y(output_6_986));
wire output_8_986, output_8_11, output_7_986;
mixer gate_output_7_986(.a(output_8_986), .b(output_8_11), .y(output_7_986));
wire output_9_986, output_9_11, output_8_986;
mixer gate_output_8_986(.a(output_9_986), .b(output_9_11), .y(output_8_986));
wire output_10_986, output_10_11, output_9_986;
mixer gate_output_9_986(.a(output_10_986), .b(output_10_11), .y(output_9_986));
wire output_11_986, output_11_11, output_10_986;
mixer gate_output_10_986(.a(output_11_986), .b(output_11_11), .y(output_10_986));
wire output_12_986, output_12_11, output_11_986;
mixer gate_output_11_986(.a(output_12_986), .b(output_12_11), .y(output_11_986));
wire output_13_986, output_13_11, output_12_986;
mixer gate_output_12_986(.a(output_13_986), .b(output_13_11), .y(output_12_986));
wire output_14_986, output_14_11, output_13_986;
mixer gate_output_13_986(.a(output_14_986), .b(output_14_11), .y(output_13_986));
wire output_15_986, output_15_11, output_14_986;
mixer gate_output_14_986(.a(output_15_986), .b(output_15_11), .y(output_14_986));
wire output_16_986, output_16_11, output_15_986;
mixer gate_output_15_986(.a(output_16_986), .b(output_16_11), .y(output_15_986));
wire output_1_987, output_1_12, output_0_987;
mixer gate_output_0_987(.a(output_1_987), .b(output_1_12), .y(output_0_987));
wire output_2_987, output_2_12, output_1_987;
mixer gate_output_1_987(.a(output_2_987), .b(output_2_12), .y(output_1_987));
wire output_3_987, output_3_12, output_2_987;
mixer gate_output_2_987(.a(output_3_987), .b(output_3_12), .y(output_2_987));
wire output_4_987, output_4_12, output_3_987;
mixer gate_output_3_987(.a(output_4_987), .b(output_4_12), .y(output_3_987));
wire output_5_987, output_5_12, output_4_987;
mixer gate_output_4_987(.a(output_5_987), .b(output_5_12), .y(output_4_987));
wire output_6_987, output_6_12, output_5_987;
mixer gate_output_5_987(.a(output_6_987), .b(output_6_12), .y(output_5_987));
wire output_7_987, output_7_12, output_6_987;
mixer gate_output_6_987(.a(output_7_987), .b(output_7_12), .y(output_6_987));
wire output_8_987, output_8_12, output_7_987;
mixer gate_output_7_987(.a(output_8_987), .b(output_8_12), .y(output_7_987));
wire output_9_987, output_9_12, output_8_987;
mixer gate_output_8_987(.a(output_9_987), .b(output_9_12), .y(output_8_987));
wire output_10_987, output_10_12, output_9_987;
mixer gate_output_9_987(.a(output_10_987), .b(output_10_12), .y(output_9_987));
wire output_11_987, output_11_12, output_10_987;
mixer gate_output_10_987(.a(output_11_987), .b(output_11_12), .y(output_10_987));
wire output_12_987, output_12_12, output_11_987;
mixer gate_output_11_987(.a(output_12_987), .b(output_12_12), .y(output_11_987));
wire output_13_987, output_13_12, output_12_987;
mixer gate_output_12_987(.a(output_13_987), .b(output_13_12), .y(output_12_987));
wire output_14_987, output_14_12, output_13_987;
mixer gate_output_13_987(.a(output_14_987), .b(output_14_12), .y(output_13_987));
wire output_15_987, output_15_12, output_14_987;
mixer gate_output_14_987(.a(output_15_987), .b(output_15_12), .y(output_14_987));
wire output_16_987, output_16_12, output_15_987;
mixer gate_output_15_987(.a(output_16_987), .b(output_16_12), .y(output_15_987));
wire output_1_988, output_1_13, output_0_988;
mixer gate_output_0_988(.a(output_1_988), .b(output_1_13), .y(output_0_988));
wire output_2_988, output_2_13, output_1_988;
mixer gate_output_1_988(.a(output_2_988), .b(output_2_13), .y(output_1_988));
wire output_3_988, output_3_13, output_2_988;
mixer gate_output_2_988(.a(output_3_988), .b(output_3_13), .y(output_2_988));
wire output_4_988, output_4_13, output_3_988;
mixer gate_output_3_988(.a(output_4_988), .b(output_4_13), .y(output_3_988));
wire output_5_988, output_5_13, output_4_988;
mixer gate_output_4_988(.a(output_5_988), .b(output_5_13), .y(output_4_988));
wire output_6_988, output_6_13, output_5_988;
mixer gate_output_5_988(.a(output_6_988), .b(output_6_13), .y(output_5_988));
wire output_7_988, output_7_13, output_6_988;
mixer gate_output_6_988(.a(output_7_988), .b(output_7_13), .y(output_6_988));
wire output_8_988, output_8_13, output_7_988;
mixer gate_output_7_988(.a(output_8_988), .b(output_8_13), .y(output_7_988));
wire output_9_988, output_9_13, output_8_988;
mixer gate_output_8_988(.a(output_9_988), .b(output_9_13), .y(output_8_988));
wire output_10_988, output_10_13, output_9_988;
mixer gate_output_9_988(.a(output_10_988), .b(output_10_13), .y(output_9_988));
wire output_11_988, output_11_13, output_10_988;
mixer gate_output_10_988(.a(output_11_988), .b(output_11_13), .y(output_10_988));
wire output_12_988, output_12_13, output_11_988;
mixer gate_output_11_988(.a(output_12_988), .b(output_12_13), .y(output_11_988));
wire output_13_988, output_13_13, output_12_988;
mixer gate_output_12_988(.a(output_13_988), .b(output_13_13), .y(output_12_988));
wire output_14_988, output_14_13, output_13_988;
mixer gate_output_13_988(.a(output_14_988), .b(output_14_13), .y(output_13_988));
wire output_15_988, output_15_13, output_14_988;
mixer gate_output_14_988(.a(output_15_988), .b(output_15_13), .y(output_14_988));
wire output_16_988, output_16_13, output_15_988;
mixer gate_output_15_988(.a(output_16_988), .b(output_16_13), .y(output_15_988));
wire output_1_989, output_1_14, output_0_989;
mixer gate_output_0_989(.a(output_1_989), .b(output_1_14), .y(output_0_989));
wire output_2_989, output_2_14, output_1_989;
mixer gate_output_1_989(.a(output_2_989), .b(output_2_14), .y(output_1_989));
wire output_3_989, output_3_14, output_2_989;
mixer gate_output_2_989(.a(output_3_989), .b(output_3_14), .y(output_2_989));
wire output_4_989, output_4_14, output_3_989;
mixer gate_output_3_989(.a(output_4_989), .b(output_4_14), .y(output_3_989));
wire output_5_989, output_5_14, output_4_989;
mixer gate_output_4_989(.a(output_5_989), .b(output_5_14), .y(output_4_989));
wire output_6_989, output_6_14, output_5_989;
mixer gate_output_5_989(.a(output_6_989), .b(output_6_14), .y(output_5_989));
wire output_7_989, output_7_14, output_6_989;
mixer gate_output_6_989(.a(output_7_989), .b(output_7_14), .y(output_6_989));
wire output_8_989, output_8_14, output_7_989;
mixer gate_output_7_989(.a(output_8_989), .b(output_8_14), .y(output_7_989));
wire output_9_989, output_9_14, output_8_989;
mixer gate_output_8_989(.a(output_9_989), .b(output_9_14), .y(output_8_989));
wire output_10_989, output_10_14, output_9_989;
mixer gate_output_9_989(.a(output_10_989), .b(output_10_14), .y(output_9_989));
wire output_11_989, output_11_14, output_10_989;
mixer gate_output_10_989(.a(output_11_989), .b(output_11_14), .y(output_10_989));
wire output_12_989, output_12_14, output_11_989;
mixer gate_output_11_989(.a(output_12_989), .b(output_12_14), .y(output_11_989));
wire output_13_989, output_13_14, output_12_989;
mixer gate_output_12_989(.a(output_13_989), .b(output_13_14), .y(output_12_989));
wire output_14_989, output_14_14, output_13_989;
mixer gate_output_13_989(.a(output_14_989), .b(output_14_14), .y(output_13_989));
wire output_15_989, output_15_14, output_14_989;
mixer gate_output_14_989(.a(output_15_989), .b(output_15_14), .y(output_14_989));
wire output_16_989, output_16_14, output_15_989;
mixer gate_output_15_989(.a(output_16_989), .b(output_16_14), .y(output_15_989));
wire output_1_990, output_1_15, output_0_990;
mixer gate_output_0_990(.a(output_1_990), .b(output_1_15), .y(output_0_990));
wire output_2_990, output_2_15, output_1_990;
mixer gate_output_1_990(.a(output_2_990), .b(output_2_15), .y(output_1_990));
wire output_3_990, output_3_15, output_2_990;
mixer gate_output_2_990(.a(output_3_990), .b(output_3_15), .y(output_2_990));
wire output_4_990, output_4_15, output_3_990;
mixer gate_output_3_990(.a(output_4_990), .b(output_4_15), .y(output_3_990));
wire output_5_990, output_5_15, output_4_990;
mixer gate_output_4_990(.a(output_5_990), .b(output_5_15), .y(output_4_990));
wire output_6_990, output_6_15, output_5_990;
mixer gate_output_5_990(.a(output_6_990), .b(output_6_15), .y(output_5_990));
wire output_7_990, output_7_15, output_6_990;
mixer gate_output_6_990(.a(output_7_990), .b(output_7_15), .y(output_6_990));
wire output_8_990, output_8_15, output_7_990;
mixer gate_output_7_990(.a(output_8_990), .b(output_8_15), .y(output_7_990));
wire output_9_990, output_9_15, output_8_990;
mixer gate_output_8_990(.a(output_9_990), .b(output_9_15), .y(output_8_990));
wire output_10_990, output_10_15, output_9_990;
mixer gate_output_9_990(.a(output_10_990), .b(output_10_15), .y(output_9_990));
wire output_11_990, output_11_15, output_10_990;
mixer gate_output_10_990(.a(output_11_990), .b(output_11_15), .y(output_10_990));
wire output_12_990, output_12_15, output_11_990;
mixer gate_output_11_990(.a(output_12_990), .b(output_12_15), .y(output_11_990));
wire output_13_990, output_13_15, output_12_990;
mixer gate_output_12_990(.a(output_13_990), .b(output_13_15), .y(output_12_990));
wire output_14_990, output_14_15, output_13_990;
mixer gate_output_13_990(.a(output_14_990), .b(output_14_15), .y(output_13_990));
wire output_15_990, output_15_15, output_14_990;
mixer gate_output_14_990(.a(output_15_990), .b(output_15_15), .y(output_14_990));
wire output_16_990, output_16_15, output_15_990;
mixer gate_output_15_990(.a(output_16_990), .b(output_16_15), .y(output_15_990));
wire output_1_991, output_1_0, output_0_991;
mixer gate_output_0_991(.a(output_1_991), .b(output_1_0), .y(output_0_991));
wire output_2_991, output_2_0, output_1_991;
mixer gate_output_1_991(.a(output_2_991), .b(output_2_0), .y(output_1_991));
wire output_3_991, output_3_0, output_2_991;
mixer gate_output_2_991(.a(output_3_991), .b(output_3_0), .y(output_2_991));
wire output_4_991, output_4_0, output_3_991;
mixer gate_output_3_991(.a(output_4_991), .b(output_4_0), .y(output_3_991));
wire output_5_991, output_5_0, output_4_991;
mixer gate_output_4_991(.a(output_5_991), .b(output_5_0), .y(output_4_991));
wire output_6_991, output_6_0, output_5_991;
mixer gate_output_5_991(.a(output_6_991), .b(output_6_0), .y(output_5_991));
wire output_7_991, output_7_0, output_6_991;
mixer gate_output_6_991(.a(output_7_991), .b(output_7_0), .y(output_6_991));
wire output_8_991, output_8_0, output_7_991;
mixer gate_output_7_991(.a(output_8_991), .b(output_8_0), .y(output_7_991));
wire output_9_991, output_9_0, output_8_991;
mixer gate_output_8_991(.a(output_9_991), .b(output_9_0), .y(output_8_991));
wire output_10_991, output_10_0, output_9_991;
mixer gate_output_9_991(.a(output_10_991), .b(output_10_0), .y(output_9_991));
wire output_11_991, output_11_0, output_10_991;
mixer gate_output_10_991(.a(output_11_991), .b(output_11_0), .y(output_10_991));
wire output_12_991, output_12_0, output_11_991;
mixer gate_output_11_991(.a(output_12_991), .b(output_12_0), .y(output_11_991));
wire output_13_991, output_13_0, output_12_991;
mixer gate_output_12_991(.a(output_13_991), .b(output_13_0), .y(output_12_991));
wire output_14_991, output_14_0, output_13_991;
mixer gate_output_13_991(.a(output_14_991), .b(output_14_0), .y(output_13_991));
wire output_15_991, output_15_0, output_14_991;
mixer gate_output_14_991(.a(output_15_991), .b(output_15_0), .y(output_14_991));
wire output_16_991, output_16_0, output_15_991;
mixer gate_output_15_991(.a(output_16_991), .b(output_16_0), .y(output_15_991));
wire output_1_992, output_1_1, output_0_992;
mixer gate_output_0_992(.a(output_1_992), .b(output_1_1), .y(output_0_992));
wire output_2_992, output_2_1, output_1_992;
mixer gate_output_1_992(.a(output_2_992), .b(output_2_1), .y(output_1_992));
wire output_3_992, output_3_1, output_2_992;
mixer gate_output_2_992(.a(output_3_992), .b(output_3_1), .y(output_2_992));
wire output_4_992, output_4_1, output_3_992;
mixer gate_output_3_992(.a(output_4_992), .b(output_4_1), .y(output_3_992));
wire output_5_992, output_5_1, output_4_992;
mixer gate_output_4_992(.a(output_5_992), .b(output_5_1), .y(output_4_992));
wire output_6_992, output_6_1, output_5_992;
mixer gate_output_5_992(.a(output_6_992), .b(output_6_1), .y(output_5_992));
wire output_7_992, output_7_1, output_6_992;
mixer gate_output_6_992(.a(output_7_992), .b(output_7_1), .y(output_6_992));
wire output_8_992, output_8_1, output_7_992;
mixer gate_output_7_992(.a(output_8_992), .b(output_8_1), .y(output_7_992));
wire output_9_992, output_9_1, output_8_992;
mixer gate_output_8_992(.a(output_9_992), .b(output_9_1), .y(output_8_992));
wire output_10_992, output_10_1, output_9_992;
mixer gate_output_9_992(.a(output_10_992), .b(output_10_1), .y(output_9_992));
wire output_11_992, output_11_1, output_10_992;
mixer gate_output_10_992(.a(output_11_992), .b(output_11_1), .y(output_10_992));
wire output_12_992, output_12_1, output_11_992;
mixer gate_output_11_992(.a(output_12_992), .b(output_12_1), .y(output_11_992));
wire output_13_992, output_13_1, output_12_992;
mixer gate_output_12_992(.a(output_13_992), .b(output_13_1), .y(output_12_992));
wire output_14_992, output_14_1, output_13_992;
mixer gate_output_13_992(.a(output_14_992), .b(output_14_1), .y(output_13_992));
wire output_15_992, output_15_1, output_14_992;
mixer gate_output_14_992(.a(output_15_992), .b(output_15_1), .y(output_14_992));
wire output_16_992, output_16_1, output_15_992;
mixer gate_output_15_992(.a(output_16_992), .b(output_16_1), .y(output_15_992));
wire output_1_993, output_1_2, output_0_993;
mixer gate_output_0_993(.a(output_1_993), .b(output_1_2), .y(output_0_993));
wire output_2_993, output_2_2, output_1_993;
mixer gate_output_1_993(.a(output_2_993), .b(output_2_2), .y(output_1_993));
wire output_3_993, output_3_2, output_2_993;
mixer gate_output_2_993(.a(output_3_993), .b(output_3_2), .y(output_2_993));
wire output_4_993, output_4_2, output_3_993;
mixer gate_output_3_993(.a(output_4_993), .b(output_4_2), .y(output_3_993));
wire output_5_993, output_5_2, output_4_993;
mixer gate_output_4_993(.a(output_5_993), .b(output_5_2), .y(output_4_993));
wire output_6_993, output_6_2, output_5_993;
mixer gate_output_5_993(.a(output_6_993), .b(output_6_2), .y(output_5_993));
wire output_7_993, output_7_2, output_6_993;
mixer gate_output_6_993(.a(output_7_993), .b(output_7_2), .y(output_6_993));
wire output_8_993, output_8_2, output_7_993;
mixer gate_output_7_993(.a(output_8_993), .b(output_8_2), .y(output_7_993));
wire output_9_993, output_9_2, output_8_993;
mixer gate_output_8_993(.a(output_9_993), .b(output_9_2), .y(output_8_993));
wire output_10_993, output_10_2, output_9_993;
mixer gate_output_9_993(.a(output_10_993), .b(output_10_2), .y(output_9_993));
wire output_11_993, output_11_2, output_10_993;
mixer gate_output_10_993(.a(output_11_993), .b(output_11_2), .y(output_10_993));
wire output_12_993, output_12_2, output_11_993;
mixer gate_output_11_993(.a(output_12_993), .b(output_12_2), .y(output_11_993));
wire output_13_993, output_13_2, output_12_993;
mixer gate_output_12_993(.a(output_13_993), .b(output_13_2), .y(output_12_993));
wire output_14_993, output_14_2, output_13_993;
mixer gate_output_13_993(.a(output_14_993), .b(output_14_2), .y(output_13_993));
wire output_15_993, output_15_2, output_14_993;
mixer gate_output_14_993(.a(output_15_993), .b(output_15_2), .y(output_14_993));
wire output_16_993, output_16_2, output_15_993;
mixer gate_output_15_993(.a(output_16_993), .b(output_16_2), .y(output_15_993));
wire output_1_994, output_1_3, output_0_994;
mixer gate_output_0_994(.a(output_1_994), .b(output_1_3), .y(output_0_994));
wire output_2_994, output_2_3, output_1_994;
mixer gate_output_1_994(.a(output_2_994), .b(output_2_3), .y(output_1_994));
wire output_3_994, output_3_3, output_2_994;
mixer gate_output_2_994(.a(output_3_994), .b(output_3_3), .y(output_2_994));
wire output_4_994, output_4_3, output_3_994;
mixer gate_output_3_994(.a(output_4_994), .b(output_4_3), .y(output_3_994));
wire output_5_994, output_5_3, output_4_994;
mixer gate_output_4_994(.a(output_5_994), .b(output_5_3), .y(output_4_994));
wire output_6_994, output_6_3, output_5_994;
mixer gate_output_5_994(.a(output_6_994), .b(output_6_3), .y(output_5_994));
wire output_7_994, output_7_3, output_6_994;
mixer gate_output_6_994(.a(output_7_994), .b(output_7_3), .y(output_6_994));
wire output_8_994, output_8_3, output_7_994;
mixer gate_output_7_994(.a(output_8_994), .b(output_8_3), .y(output_7_994));
wire output_9_994, output_9_3, output_8_994;
mixer gate_output_8_994(.a(output_9_994), .b(output_9_3), .y(output_8_994));
wire output_10_994, output_10_3, output_9_994;
mixer gate_output_9_994(.a(output_10_994), .b(output_10_3), .y(output_9_994));
wire output_11_994, output_11_3, output_10_994;
mixer gate_output_10_994(.a(output_11_994), .b(output_11_3), .y(output_10_994));
wire output_12_994, output_12_3, output_11_994;
mixer gate_output_11_994(.a(output_12_994), .b(output_12_3), .y(output_11_994));
wire output_13_994, output_13_3, output_12_994;
mixer gate_output_12_994(.a(output_13_994), .b(output_13_3), .y(output_12_994));
wire output_14_994, output_14_3, output_13_994;
mixer gate_output_13_994(.a(output_14_994), .b(output_14_3), .y(output_13_994));
wire output_15_994, output_15_3, output_14_994;
mixer gate_output_14_994(.a(output_15_994), .b(output_15_3), .y(output_14_994));
wire output_16_994, output_16_3, output_15_994;
mixer gate_output_15_994(.a(output_16_994), .b(output_16_3), .y(output_15_994));
wire output_1_995, output_1_4, output_0_995;
mixer gate_output_0_995(.a(output_1_995), .b(output_1_4), .y(output_0_995));
wire output_2_995, output_2_4, output_1_995;
mixer gate_output_1_995(.a(output_2_995), .b(output_2_4), .y(output_1_995));
wire output_3_995, output_3_4, output_2_995;
mixer gate_output_2_995(.a(output_3_995), .b(output_3_4), .y(output_2_995));
wire output_4_995, output_4_4, output_3_995;
mixer gate_output_3_995(.a(output_4_995), .b(output_4_4), .y(output_3_995));
wire output_5_995, output_5_4, output_4_995;
mixer gate_output_4_995(.a(output_5_995), .b(output_5_4), .y(output_4_995));
wire output_6_995, output_6_4, output_5_995;
mixer gate_output_5_995(.a(output_6_995), .b(output_6_4), .y(output_5_995));
wire output_7_995, output_7_4, output_6_995;
mixer gate_output_6_995(.a(output_7_995), .b(output_7_4), .y(output_6_995));
wire output_8_995, output_8_4, output_7_995;
mixer gate_output_7_995(.a(output_8_995), .b(output_8_4), .y(output_7_995));
wire output_9_995, output_9_4, output_8_995;
mixer gate_output_8_995(.a(output_9_995), .b(output_9_4), .y(output_8_995));
wire output_10_995, output_10_4, output_9_995;
mixer gate_output_9_995(.a(output_10_995), .b(output_10_4), .y(output_9_995));
wire output_11_995, output_11_4, output_10_995;
mixer gate_output_10_995(.a(output_11_995), .b(output_11_4), .y(output_10_995));
wire output_12_995, output_12_4, output_11_995;
mixer gate_output_11_995(.a(output_12_995), .b(output_12_4), .y(output_11_995));
wire output_13_995, output_13_4, output_12_995;
mixer gate_output_12_995(.a(output_13_995), .b(output_13_4), .y(output_12_995));
wire output_14_995, output_14_4, output_13_995;
mixer gate_output_13_995(.a(output_14_995), .b(output_14_4), .y(output_13_995));
wire output_15_995, output_15_4, output_14_995;
mixer gate_output_14_995(.a(output_15_995), .b(output_15_4), .y(output_14_995));
wire output_16_995, output_16_4, output_15_995;
mixer gate_output_15_995(.a(output_16_995), .b(output_16_4), .y(output_15_995));
wire output_1_996, output_1_5, output_0_996;
mixer gate_output_0_996(.a(output_1_996), .b(output_1_5), .y(output_0_996));
wire output_2_996, output_2_5, output_1_996;
mixer gate_output_1_996(.a(output_2_996), .b(output_2_5), .y(output_1_996));
wire output_3_996, output_3_5, output_2_996;
mixer gate_output_2_996(.a(output_3_996), .b(output_3_5), .y(output_2_996));
wire output_4_996, output_4_5, output_3_996;
mixer gate_output_3_996(.a(output_4_996), .b(output_4_5), .y(output_3_996));
wire output_5_996, output_5_5, output_4_996;
mixer gate_output_4_996(.a(output_5_996), .b(output_5_5), .y(output_4_996));
wire output_6_996, output_6_5, output_5_996;
mixer gate_output_5_996(.a(output_6_996), .b(output_6_5), .y(output_5_996));
wire output_7_996, output_7_5, output_6_996;
mixer gate_output_6_996(.a(output_7_996), .b(output_7_5), .y(output_6_996));
wire output_8_996, output_8_5, output_7_996;
mixer gate_output_7_996(.a(output_8_996), .b(output_8_5), .y(output_7_996));
wire output_9_996, output_9_5, output_8_996;
mixer gate_output_8_996(.a(output_9_996), .b(output_9_5), .y(output_8_996));
wire output_10_996, output_10_5, output_9_996;
mixer gate_output_9_996(.a(output_10_996), .b(output_10_5), .y(output_9_996));
wire output_11_996, output_11_5, output_10_996;
mixer gate_output_10_996(.a(output_11_996), .b(output_11_5), .y(output_10_996));
wire output_12_996, output_12_5, output_11_996;
mixer gate_output_11_996(.a(output_12_996), .b(output_12_5), .y(output_11_996));
wire output_13_996, output_13_5, output_12_996;
mixer gate_output_12_996(.a(output_13_996), .b(output_13_5), .y(output_12_996));
wire output_14_996, output_14_5, output_13_996;
mixer gate_output_13_996(.a(output_14_996), .b(output_14_5), .y(output_13_996));
wire output_15_996, output_15_5, output_14_996;
mixer gate_output_14_996(.a(output_15_996), .b(output_15_5), .y(output_14_996));
wire output_16_996, output_16_5, output_15_996;
mixer gate_output_15_996(.a(output_16_996), .b(output_16_5), .y(output_15_996));
wire output_1_997, output_1_6, output_0_997;
mixer gate_output_0_997(.a(output_1_997), .b(output_1_6), .y(output_0_997));
wire output_2_997, output_2_6, output_1_997;
mixer gate_output_1_997(.a(output_2_997), .b(output_2_6), .y(output_1_997));
wire output_3_997, output_3_6, output_2_997;
mixer gate_output_2_997(.a(output_3_997), .b(output_3_6), .y(output_2_997));
wire output_4_997, output_4_6, output_3_997;
mixer gate_output_3_997(.a(output_4_997), .b(output_4_6), .y(output_3_997));
wire output_5_997, output_5_6, output_4_997;
mixer gate_output_4_997(.a(output_5_997), .b(output_5_6), .y(output_4_997));
wire output_6_997, output_6_6, output_5_997;
mixer gate_output_5_997(.a(output_6_997), .b(output_6_6), .y(output_5_997));
wire output_7_997, output_7_6, output_6_997;
mixer gate_output_6_997(.a(output_7_997), .b(output_7_6), .y(output_6_997));
wire output_8_997, output_8_6, output_7_997;
mixer gate_output_7_997(.a(output_8_997), .b(output_8_6), .y(output_7_997));
wire output_9_997, output_9_6, output_8_997;
mixer gate_output_8_997(.a(output_9_997), .b(output_9_6), .y(output_8_997));
wire output_10_997, output_10_6, output_9_997;
mixer gate_output_9_997(.a(output_10_997), .b(output_10_6), .y(output_9_997));
wire output_11_997, output_11_6, output_10_997;
mixer gate_output_10_997(.a(output_11_997), .b(output_11_6), .y(output_10_997));
wire output_12_997, output_12_6, output_11_997;
mixer gate_output_11_997(.a(output_12_997), .b(output_12_6), .y(output_11_997));
wire output_13_997, output_13_6, output_12_997;
mixer gate_output_12_997(.a(output_13_997), .b(output_13_6), .y(output_12_997));
wire output_14_997, output_14_6, output_13_997;
mixer gate_output_13_997(.a(output_14_997), .b(output_14_6), .y(output_13_997));
wire output_15_997, output_15_6, output_14_997;
mixer gate_output_14_997(.a(output_15_997), .b(output_15_6), .y(output_14_997));
wire output_16_997, output_16_6, output_15_997;
mixer gate_output_15_997(.a(output_16_997), .b(output_16_6), .y(output_15_997));
wire output_1_998, output_1_7, output_0_998;
mixer gate_output_0_998(.a(output_1_998), .b(output_1_7), .y(output_0_998));
wire output_2_998, output_2_7, output_1_998;
mixer gate_output_1_998(.a(output_2_998), .b(output_2_7), .y(output_1_998));
wire output_3_998, output_3_7, output_2_998;
mixer gate_output_2_998(.a(output_3_998), .b(output_3_7), .y(output_2_998));
wire output_4_998, output_4_7, output_3_998;
mixer gate_output_3_998(.a(output_4_998), .b(output_4_7), .y(output_3_998));
wire output_5_998, output_5_7, output_4_998;
mixer gate_output_4_998(.a(output_5_998), .b(output_5_7), .y(output_4_998));
wire output_6_998, output_6_7, output_5_998;
mixer gate_output_5_998(.a(output_6_998), .b(output_6_7), .y(output_5_998));
wire output_7_998, output_7_7, output_6_998;
mixer gate_output_6_998(.a(output_7_998), .b(output_7_7), .y(output_6_998));
wire output_8_998, output_8_7, output_7_998;
mixer gate_output_7_998(.a(output_8_998), .b(output_8_7), .y(output_7_998));
wire output_9_998, output_9_7, output_8_998;
mixer gate_output_8_998(.a(output_9_998), .b(output_9_7), .y(output_8_998));
wire output_10_998, output_10_7, output_9_998;
mixer gate_output_9_998(.a(output_10_998), .b(output_10_7), .y(output_9_998));
wire output_11_998, output_11_7, output_10_998;
mixer gate_output_10_998(.a(output_11_998), .b(output_11_7), .y(output_10_998));
wire output_12_998, output_12_7, output_11_998;
mixer gate_output_11_998(.a(output_12_998), .b(output_12_7), .y(output_11_998));
wire output_13_998, output_13_7, output_12_998;
mixer gate_output_12_998(.a(output_13_998), .b(output_13_7), .y(output_12_998));
wire output_14_998, output_14_7, output_13_998;
mixer gate_output_13_998(.a(output_14_998), .b(output_14_7), .y(output_13_998));
wire output_15_998, output_15_7, output_14_998;
mixer gate_output_14_998(.a(output_15_998), .b(output_15_7), .y(output_14_998));
wire output_16_998, output_16_7, output_15_998;
mixer gate_output_15_998(.a(output_16_998), .b(output_16_7), .y(output_15_998));
wire output_1_999, output_1_8, output_0_999;
mixer gate_output_0_999(.a(output_1_999), .b(output_1_8), .y(output_0_999));
wire output_2_999, output_2_8, output_1_999;
mixer gate_output_1_999(.a(output_2_999), .b(output_2_8), .y(output_1_999));
wire output_3_999, output_3_8, output_2_999;
mixer gate_output_2_999(.a(output_3_999), .b(output_3_8), .y(output_2_999));
wire output_4_999, output_4_8, output_3_999;
mixer gate_output_3_999(.a(output_4_999), .b(output_4_8), .y(output_3_999));
wire output_5_999, output_5_8, output_4_999;
mixer gate_output_4_999(.a(output_5_999), .b(output_5_8), .y(output_4_999));
wire output_6_999, output_6_8, output_5_999;
mixer gate_output_5_999(.a(output_6_999), .b(output_6_8), .y(output_5_999));
wire output_7_999, output_7_8, output_6_999;
mixer gate_output_6_999(.a(output_7_999), .b(output_7_8), .y(output_6_999));
wire output_8_999, output_8_8, output_7_999;
mixer gate_output_7_999(.a(output_8_999), .b(output_8_8), .y(output_7_999));
wire output_9_999, output_9_8, output_8_999;
mixer gate_output_8_999(.a(output_9_999), .b(output_9_8), .y(output_8_999));
wire output_10_999, output_10_8, output_9_999;
mixer gate_output_9_999(.a(output_10_999), .b(output_10_8), .y(output_9_999));
wire output_11_999, output_11_8, output_10_999;
mixer gate_output_10_999(.a(output_11_999), .b(output_11_8), .y(output_10_999));
wire output_12_999, output_12_8, output_11_999;
mixer gate_output_11_999(.a(output_12_999), .b(output_12_8), .y(output_11_999));
wire output_13_999, output_13_8, output_12_999;
mixer gate_output_12_999(.a(output_13_999), .b(output_13_8), .y(output_12_999));
wire output_14_999, output_14_8, output_13_999;
mixer gate_output_13_999(.a(output_14_999), .b(output_14_8), .y(output_13_999));
wire output_15_999, output_15_8, output_14_999;
mixer gate_output_14_999(.a(output_15_999), .b(output_15_8), .y(output_14_999));
wire output_16_999, output_16_8, output_15_999;
mixer gate_output_15_999(.a(output_16_999), .b(output_16_8), .y(output_15_999));
wire output_1_1000, output_1_9, output_0_1000;
mixer gate_output_0_1000(.a(output_1_1000), .b(output_1_9), .y(output_0_1000));
wire output_2_1000, output_2_9, output_1_1000;
mixer gate_output_1_1000(.a(output_2_1000), .b(output_2_9), .y(output_1_1000));
wire output_3_1000, output_3_9, output_2_1000;
mixer gate_output_2_1000(.a(output_3_1000), .b(output_3_9), .y(output_2_1000));
wire output_4_1000, output_4_9, output_3_1000;
mixer gate_output_3_1000(.a(output_4_1000), .b(output_4_9), .y(output_3_1000));
wire output_5_1000, output_5_9, output_4_1000;
mixer gate_output_4_1000(.a(output_5_1000), .b(output_5_9), .y(output_4_1000));
wire output_6_1000, output_6_9, output_5_1000;
mixer gate_output_5_1000(.a(output_6_1000), .b(output_6_9), .y(output_5_1000));
wire output_7_1000, output_7_9, output_6_1000;
mixer gate_output_6_1000(.a(output_7_1000), .b(output_7_9), .y(output_6_1000));
wire output_8_1000, output_8_9, output_7_1000;
mixer gate_output_7_1000(.a(output_8_1000), .b(output_8_9), .y(output_7_1000));
wire output_9_1000, output_9_9, output_8_1000;
mixer gate_output_8_1000(.a(output_9_1000), .b(output_9_9), .y(output_8_1000));
wire output_10_1000, output_10_9, output_9_1000;
mixer gate_output_9_1000(.a(output_10_1000), .b(output_10_9), .y(output_9_1000));
wire output_11_1000, output_11_9, output_10_1000;
mixer gate_output_10_1000(.a(output_11_1000), .b(output_11_9), .y(output_10_1000));
wire output_12_1000, output_12_9, output_11_1000;
mixer gate_output_11_1000(.a(output_12_1000), .b(output_12_9), .y(output_11_1000));
wire output_13_1000, output_13_9, output_12_1000;
mixer gate_output_12_1000(.a(output_13_1000), .b(output_13_9), .y(output_12_1000));
wire output_14_1000, output_14_9, output_13_1000;
mixer gate_output_13_1000(.a(output_14_1000), .b(output_14_9), .y(output_13_1000));
wire output_15_1000, output_15_9, output_14_1000;
mixer gate_output_14_1000(.a(output_15_1000), .b(output_15_9), .y(output_14_1000));
wire output_16_1000, output_16_9, output_15_1000;
mixer gate_output_15_1000(.a(output_16_1000), .b(output_16_9), .y(output_15_1000));
wire output_1_1001, output_1_10, output_0_1001;
mixer gate_output_0_1001(.a(output_1_1001), .b(output_1_10), .y(output_0_1001));
wire output_2_1001, output_2_10, output_1_1001;
mixer gate_output_1_1001(.a(output_2_1001), .b(output_2_10), .y(output_1_1001));
wire output_3_1001, output_3_10, output_2_1001;
mixer gate_output_2_1001(.a(output_3_1001), .b(output_3_10), .y(output_2_1001));
wire output_4_1001, output_4_10, output_3_1001;
mixer gate_output_3_1001(.a(output_4_1001), .b(output_4_10), .y(output_3_1001));
wire output_5_1001, output_5_10, output_4_1001;
mixer gate_output_4_1001(.a(output_5_1001), .b(output_5_10), .y(output_4_1001));
wire output_6_1001, output_6_10, output_5_1001;
mixer gate_output_5_1001(.a(output_6_1001), .b(output_6_10), .y(output_5_1001));
wire output_7_1001, output_7_10, output_6_1001;
mixer gate_output_6_1001(.a(output_7_1001), .b(output_7_10), .y(output_6_1001));
wire output_8_1001, output_8_10, output_7_1001;
mixer gate_output_7_1001(.a(output_8_1001), .b(output_8_10), .y(output_7_1001));
wire output_9_1001, output_9_10, output_8_1001;
mixer gate_output_8_1001(.a(output_9_1001), .b(output_9_10), .y(output_8_1001));
wire output_10_1001, output_10_10, output_9_1001;
mixer gate_output_9_1001(.a(output_10_1001), .b(output_10_10), .y(output_9_1001));
wire output_11_1001, output_11_10, output_10_1001;
mixer gate_output_10_1001(.a(output_11_1001), .b(output_11_10), .y(output_10_1001));
wire output_12_1001, output_12_10, output_11_1001;
mixer gate_output_11_1001(.a(output_12_1001), .b(output_12_10), .y(output_11_1001));
wire output_13_1001, output_13_10, output_12_1001;
mixer gate_output_12_1001(.a(output_13_1001), .b(output_13_10), .y(output_12_1001));
wire output_14_1001, output_14_10, output_13_1001;
mixer gate_output_13_1001(.a(output_14_1001), .b(output_14_10), .y(output_13_1001));
wire output_15_1001, output_15_10, output_14_1001;
mixer gate_output_14_1001(.a(output_15_1001), .b(output_15_10), .y(output_14_1001));
wire output_16_1001, output_16_10, output_15_1001;
mixer gate_output_15_1001(.a(output_16_1001), .b(output_16_10), .y(output_15_1001));
wire output_1_1002, output_1_11, output_0_1002;
mixer gate_output_0_1002(.a(output_1_1002), .b(output_1_11), .y(output_0_1002));
wire output_2_1002, output_2_11, output_1_1002;
mixer gate_output_1_1002(.a(output_2_1002), .b(output_2_11), .y(output_1_1002));
wire output_3_1002, output_3_11, output_2_1002;
mixer gate_output_2_1002(.a(output_3_1002), .b(output_3_11), .y(output_2_1002));
wire output_4_1002, output_4_11, output_3_1002;
mixer gate_output_3_1002(.a(output_4_1002), .b(output_4_11), .y(output_3_1002));
wire output_5_1002, output_5_11, output_4_1002;
mixer gate_output_4_1002(.a(output_5_1002), .b(output_5_11), .y(output_4_1002));
wire output_6_1002, output_6_11, output_5_1002;
mixer gate_output_5_1002(.a(output_6_1002), .b(output_6_11), .y(output_5_1002));
wire output_7_1002, output_7_11, output_6_1002;
mixer gate_output_6_1002(.a(output_7_1002), .b(output_7_11), .y(output_6_1002));
wire output_8_1002, output_8_11, output_7_1002;
mixer gate_output_7_1002(.a(output_8_1002), .b(output_8_11), .y(output_7_1002));
wire output_9_1002, output_9_11, output_8_1002;
mixer gate_output_8_1002(.a(output_9_1002), .b(output_9_11), .y(output_8_1002));
wire output_10_1002, output_10_11, output_9_1002;
mixer gate_output_9_1002(.a(output_10_1002), .b(output_10_11), .y(output_9_1002));
wire output_11_1002, output_11_11, output_10_1002;
mixer gate_output_10_1002(.a(output_11_1002), .b(output_11_11), .y(output_10_1002));
wire output_12_1002, output_12_11, output_11_1002;
mixer gate_output_11_1002(.a(output_12_1002), .b(output_12_11), .y(output_11_1002));
wire output_13_1002, output_13_11, output_12_1002;
mixer gate_output_12_1002(.a(output_13_1002), .b(output_13_11), .y(output_12_1002));
wire output_14_1002, output_14_11, output_13_1002;
mixer gate_output_13_1002(.a(output_14_1002), .b(output_14_11), .y(output_13_1002));
wire output_15_1002, output_15_11, output_14_1002;
mixer gate_output_14_1002(.a(output_15_1002), .b(output_15_11), .y(output_14_1002));
wire output_16_1002, output_16_11, output_15_1002;
mixer gate_output_15_1002(.a(output_16_1002), .b(output_16_11), .y(output_15_1002));
wire output_1_1003, output_1_12, output_0_1003;
mixer gate_output_0_1003(.a(output_1_1003), .b(output_1_12), .y(output_0_1003));
wire output_2_1003, output_2_12, output_1_1003;
mixer gate_output_1_1003(.a(output_2_1003), .b(output_2_12), .y(output_1_1003));
wire output_3_1003, output_3_12, output_2_1003;
mixer gate_output_2_1003(.a(output_3_1003), .b(output_3_12), .y(output_2_1003));
wire output_4_1003, output_4_12, output_3_1003;
mixer gate_output_3_1003(.a(output_4_1003), .b(output_4_12), .y(output_3_1003));
wire output_5_1003, output_5_12, output_4_1003;
mixer gate_output_4_1003(.a(output_5_1003), .b(output_5_12), .y(output_4_1003));
wire output_6_1003, output_6_12, output_5_1003;
mixer gate_output_5_1003(.a(output_6_1003), .b(output_6_12), .y(output_5_1003));
wire output_7_1003, output_7_12, output_6_1003;
mixer gate_output_6_1003(.a(output_7_1003), .b(output_7_12), .y(output_6_1003));
wire output_8_1003, output_8_12, output_7_1003;
mixer gate_output_7_1003(.a(output_8_1003), .b(output_8_12), .y(output_7_1003));
wire output_9_1003, output_9_12, output_8_1003;
mixer gate_output_8_1003(.a(output_9_1003), .b(output_9_12), .y(output_8_1003));
wire output_10_1003, output_10_12, output_9_1003;
mixer gate_output_9_1003(.a(output_10_1003), .b(output_10_12), .y(output_9_1003));
wire output_11_1003, output_11_12, output_10_1003;
mixer gate_output_10_1003(.a(output_11_1003), .b(output_11_12), .y(output_10_1003));
wire output_12_1003, output_12_12, output_11_1003;
mixer gate_output_11_1003(.a(output_12_1003), .b(output_12_12), .y(output_11_1003));
wire output_13_1003, output_13_12, output_12_1003;
mixer gate_output_12_1003(.a(output_13_1003), .b(output_13_12), .y(output_12_1003));
wire output_14_1003, output_14_12, output_13_1003;
mixer gate_output_13_1003(.a(output_14_1003), .b(output_14_12), .y(output_13_1003));
wire output_15_1003, output_15_12, output_14_1003;
mixer gate_output_14_1003(.a(output_15_1003), .b(output_15_12), .y(output_14_1003));
wire output_16_1003, output_16_12, output_15_1003;
mixer gate_output_15_1003(.a(output_16_1003), .b(output_16_12), .y(output_15_1003));
wire output_1_1004, output_1_13, output_0_1004;
mixer gate_output_0_1004(.a(output_1_1004), .b(output_1_13), .y(output_0_1004));
wire output_2_1004, output_2_13, output_1_1004;
mixer gate_output_1_1004(.a(output_2_1004), .b(output_2_13), .y(output_1_1004));
wire output_3_1004, output_3_13, output_2_1004;
mixer gate_output_2_1004(.a(output_3_1004), .b(output_3_13), .y(output_2_1004));
wire output_4_1004, output_4_13, output_3_1004;
mixer gate_output_3_1004(.a(output_4_1004), .b(output_4_13), .y(output_3_1004));
wire output_5_1004, output_5_13, output_4_1004;
mixer gate_output_4_1004(.a(output_5_1004), .b(output_5_13), .y(output_4_1004));
wire output_6_1004, output_6_13, output_5_1004;
mixer gate_output_5_1004(.a(output_6_1004), .b(output_6_13), .y(output_5_1004));
wire output_7_1004, output_7_13, output_6_1004;
mixer gate_output_6_1004(.a(output_7_1004), .b(output_7_13), .y(output_6_1004));
wire output_8_1004, output_8_13, output_7_1004;
mixer gate_output_7_1004(.a(output_8_1004), .b(output_8_13), .y(output_7_1004));
wire output_9_1004, output_9_13, output_8_1004;
mixer gate_output_8_1004(.a(output_9_1004), .b(output_9_13), .y(output_8_1004));
wire output_10_1004, output_10_13, output_9_1004;
mixer gate_output_9_1004(.a(output_10_1004), .b(output_10_13), .y(output_9_1004));
wire output_11_1004, output_11_13, output_10_1004;
mixer gate_output_10_1004(.a(output_11_1004), .b(output_11_13), .y(output_10_1004));
wire output_12_1004, output_12_13, output_11_1004;
mixer gate_output_11_1004(.a(output_12_1004), .b(output_12_13), .y(output_11_1004));
wire output_13_1004, output_13_13, output_12_1004;
mixer gate_output_12_1004(.a(output_13_1004), .b(output_13_13), .y(output_12_1004));
wire output_14_1004, output_14_13, output_13_1004;
mixer gate_output_13_1004(.a(output_14_1004), .b(output_14_13), .y(output_13_1004));
wire output_15_1004, output_15_13, output_14_1004;
mixer gate_output_14_1004(.a(output_15_1004), .b(output_15_13), .y(output_14_1004));
wire output_16_1004, output_16_13, output_15_1004;
mixer gate_output_15_1004(.a(output_16_1004), .b(output_16_13), .y(output_15_1004));
wire output_1_1005, output_1_14, output_0_1005;
mixer gate_output_0_1005(.a(output_1_1005), .b(output_1_14), .y(output_0_1005));
wire output_2_1005, output_2_14, output_1_1005;
mixer gate_output_1_1005(.a(output_2_1005), .b(output_2_14), .y(output_1_1005));
wire output_3_1005, output_3_14, output_2_1005;
mixer gate_output_2_1005(.a(output_3_1005), .b(output_3_14), .y(output_2_1005));
wire output_4_1005, output_4_14, output_3_1005;
mixer gate_output_3_1005(.a(output_4_1005), .b(output_4_14), .y(output_3_1005));
wire output_5_1005, output_5_14, output_4_1005;
mixer gate_output_4_1005(.a(output_5_1005), .b(output_5_14), .y(output_4_1005));
wire output_6_1005, output_6_14, output_5_1005;
mixer gate_output_5_1005(.a(output_6_1005), .b(output_6_14), .y(output_5_1005));
wire output_7_1005, output_7_14, output_6_1005;
mixer gate_output_6_1005(.a(output_7_1005), .b(output_7_14), .y(output_6_1005));
wire output_8_1005, output_8_14, output_7_1005;
mixer gate_output_7_1005(.a(output_8_1005), .b(output_8_14), .y(output_7_1005));
wire output_9_1005, output_9_14, output_8_1005;
mixer gate_output_8_1005(.a(output_9_1005), .b(output_9_14), .y(output_8_1005));
wire output_10_1005, output_10_14, output_9_1005;
mixer gate_output_9_1005(.a(output_10_1005), .b(output_10_14), .y(output_9_1005));
wire output_11_1005, output_11_14, output_10_1005;
mixer gate_output_10_1005(.a(output_11_1005), .b(output_11_14), .y(output_10_1005));
wire output_12_1005, output_12_14, output_11_1005;
mixer gate_output_11_1005(.a(output_12_1005), .b(output_12_14), .y(output_11_1005));
wire output_13_1005, output_13_14, output_12_1005;
mixer gate_output_12_1005(.a(output_13_1005), .b(output_13_14), .y(output_12_1005));
wire output_14_1005, output_14_14, output_13_1005;
mixer gate_output_13_1005(.a(output_14_1005), .b(output_14_14), .y(output_13_1005));
wire output_15_1005, output_15_14, output_14_1005;
mixer gate_output_14_1005(.a(output_15_1005), .b(output_15_14), .y(output_14_1005));
wire output_16_1005, output_16_14, output_15_1005;
mixer gate_output_15_1005(.a(output_16_1005), .b(output_16_14), .y(output_15_1005));
wire output_1_1006, output_1_15, output_0_1006;
mixer gate_output_0_1006(.a(output_1_1006), .b(output_1_15), .y(output_0_1006));
wire output_2_1006, output_2_15, output_1_1006;
mixer gate_output_1_1006(.a(output_2_1006), .b(output_2_15), .y(output_1_1006));
wire output_3_1006, output_3_15, output_2_1006;
mixer gate_output_2_1006(.a(output_3_1006), .b(output_3_15), .y(output_2_1006));
wire output_4_1006, output_4_15, output_3_1006;
mixer gate_output_3_1006(.a(output_4_1006), .b(output_4_15), .y(output_3_1006));
wire output_5_1006, output_5_15, output_4_1006;
mixer gate_output_4_1006(.a(output_5_1006), .b(output_5_15), .y(output_4_1006));
wire output_6_1006, output_6_15, output_5_1006;
mixer gate_output_5_1006(.a(output_6_1006), .b(output_6_15), .y(output_5_1006));
wire output_7_1006, output_7_15, output_6_1006;
mixer gate_output_6_1006(.a(output_7_1006), .b(output_7_15), .y(output_6_1006));
wire output_8_1006, output_8_15, output_7_1006;
mixer gate_output_7_1006(.a(output_8_1006), .b(output_8_15), .y(output_7_1006));
wire output_9_1006, output_9_15, output_8_1006;
mixer gate_output_8_1006(.a(output_9_1006), .b(output_9_15), .y(output_8_1006));
wire output_10_1006, output_10_15, output_9_1006;
mixer gate_output_9_1006(.a(output_10_1006), .b(output_10_15), .y(output_9_1006));
wire output_11_1006, output_11_15, output_10_1006;
mixer gate_output_10_1006(.a(output_11_1006), .b(output_11_15), .y(output_10_1006));
wire output_12_1006, output_12_15, output_11_1006;
mixer gate_output_11_1006(.a(output_12_1006), .b(output_12_15), .y(output_11_1006));
wire output_13_1006, output_13_15, output_12_1006;
mixer gate_output_12_1006(.a(output_13_1006), .b(output_13_15), .y(output_12_1006));
wire output_14_1006, output_14_15, output_13_1006;
mixer gate_output_13_1006(.a(output_14_1006), .b(output_14_15), .y(output_13_1006));
wire output_15_1006, output_15_15, output_14_1006;
mixer gate_output_14_1006(.a(output_15_1006), .b(output_15_15), .y(output_14_1006));
wire output_16_1006, output_16_15, output_15_1006;
mixer gate_output_15_1006(.a(output_16_1006), .b(output_16_15), .y(output_15_1006));
wire output_1_1007, output_1_0, output_0_1007;
mixer gate_output_0_1007(.a(output_1_1007), .b(output_1_0), .y(output_0_1007));
wire output_2_1007, output_2_0, output_1_1007;
mixer gate_output_1_1007(.a(output_2_1007), .b(output_2_0), .y(output_1_1007));
wire output_3_1007, output_3_0, output_2_1007;
mixer gate_output_2_1007(.a(output_3_1007), .b(output_3_0), .y(output_2_1007));
wire output_4_1007, output_4_0, output_3_1007;
mixer gate_output_3_1007(.a(output_4_1007), .b(output_4_0), .y(output_3_1007));
wire output_5_1007, output_5_0, output_4_1007;
mixer gate_output_4_1007(.a(output_5_1007), .b(output_5_0), .y(output_4_1007));
wire output_6_1007, output_6_0, output_5_1007;
mixer gate_output_5_1007(.a(output_6_1007), .b(output_6_0), .y(output_5_1007));
wire output_7_1007, output_7_0, output_6_1007;
mixer gate_output_6_1007(.a(output_7_1007), .b(output_7_0), .y(output_6_1007));
wire output_8_1007, output_8_0, output_7_1007;
mixer gate_output_7_1007(.a(output_8_1007), .b(output_8_0), .y(output_7_1007));
wire output_9_1007, output_9_0, output_8_1007;
mixer gate_output_8_1007(.a(output_9_1007), .b(output_9_0), .y(output_8_1007));
wire output_10_1007, output_10_0, output_9_1007;
mixer gate_output_9_1007(.a(output_10_1007), .b(output_10_0), .y(output_9_1007));
wire output_11_1007, output_11_0, output_10_1007;
mixer gate_output_10_1007(.a(output_11_1007), .b(output_11_0), .y(output_10_1007));
wire output_12_1007, output_12_0, output_11_1007;
mixer gate_output_11_1007(.a(output_12_1007), .b(output_12_0), .y(output_11_1007));
wire output_13_1007, output_13_0, output_12_1007;
mixer gate_output_12_1007(.a(output_13_1007), .b(output_13_0), .y(output_12_1007));
wire output_14_1007, output_14_0, output_13_1007;
mixer gate_output_13_1007(.a(output_14_1007), .b(output_14_0), .y(output_13_1007));
wire output_15_1007, output_15_0, output_14_1007;
mixer gate_output_14_1007(.a(output_15_1007), .b(output_15_0), .y(output_14_1007));
wire output_16_1007, output_16_0, output_15_1007;
mixer gate_output_15_1007(.a(output_16_1007), .b(output_16_0), .y(output_15_1007));
wire output_1_1008, output_1_1, output_0_1008;
mixer gate_output_0_1008(.a(output_1_1008), .b(output_1_1), .y(output_0_1008));
wire output_2_1008, output_2_1, output_1_1008;
mixer gate_output_1_1008(.a(output_2_1008), .b(output_2_1), .y(output_1_1008));
wire output_3_1008, output_3_1, output_2_1008;
mixer gate_output_2_1008(.a(output_3_1008), .b(output_3_1), .y(output_2_1008));
wire output_4_1008, output_4_1, output_3_1008;
mixer gate_output_3_1008(.a(output_4_1008), .b(output_4_1), .y(output_3_1008));
wire output_5_1008, output_5_1, output_4_1008;
mixer gate_output_4_1008(.a(output_5_1008), .b(output_5_1), .y(output_4_1008));
wire output_6_1008, output_6_1, output_5_1008;
mixer gate_output_5_1008(.a(output_6_1008), .b(output_6_1), .y(output_5_1008));
wire output_7_1008, output_7_1, output_6_1008;
mixer gate_output_6_1008(.a(output_7_1008), .b(output_7_1), .y(output_6_1008));
wire output_8_1008, output_8_1, output_7_1008;
mixer gate_output_7_1008(.a(output_8_1008), .b(output_8_1), .y(output_7_1008));
wire output_9_1008, output_9_1, output_8_1008;
mixer gate_output_8_1008(.a(output_9_1008), .b(output_9_1), .y(output_8_1008));
wire output_10_1008, output_10_1, output_9_1008;
mixer gate_output_9_1008(.a(output_10_1008), .b(output_10_1), .y(output_9_1008));
wire output_11_1008, output_11_1, output_10_1008;
mixer gate_output_10_1008(.a(output_11_1008), .b(output_11_1), .y(output_10_1008));
wire output_12_1008, output_12_1, output_11_1008;
mixer gate_output_11_1008(.a(output_12_1008), .b(output_12_1), .y(output_11_1008));
wire output_13_1008, output_13_1, output_12_1008;
mixer gate_output_12_1008(.a(output_13_1008), .b(output_13_1), .y(output_12_1008));
wire output_14_1008, output_14_1, output_13_1008;
mixer gate_output_13_1008(.a(output_14_1008), .b(output_14_1), .y(output_13_1008));
wire output_15_1008, output_15_1, output_14_1008;
mixer gate_output_14_1008(.a(output_15_1008), .b(output_15_1), .y(output_14_1008));
wire output_16_1008, output_16_1, output_15_1008;
mixer gate_output_15_1008(.a(output_16_1008), .b(output_16_1), .y(output_15_1008));
wire output_1_1009, output_1_2, output_0_1009;
mixer gate_output_0_1009(.a(output_1_1009), .b(output_1_2), .y(output_0_1009));
wire output_2_1009, output_2_2, output_1_1009;
mixer gate_output_1_1009(.a(output_2_1009), .b(output_2_2), .y(output_1_1009));
wire output_3_1009, output_3_2, output_2_1009;
mixer gate_output_2_1009(.a(output_3_1009), .b(output_3_2), .y(output_2_1009));
wire output_4_1009, output_4_2, output_3_1009;
mixer gate_output_3_1009(.a(output_4_1009), .b(output_4_2), .y(output_3_1009));
wire output_5_1009, output_5_2, output_4_1009;
mixer gate_output_4_1009(.a(output_5_1009), .b(output_5_2), .y(output_4_1009));
wire output_6_1009, output_6_2, output_5_1009;
mixer gate_output_5_1009(.a(output_6_1009), .b(output_6_2), .y(output_5_1009));
wire output_7_1009, output_7_2, output_6_1009;
mixer gate_output_6_1009(.a(output_7_1009), .b(output_7_2), .y(output_6_1009));
wire output_8_1009, output_8_2, output_7_1009;
mixer gate_output_7_1009(.a(output_8_1009), .b(output_8_2), .y(output_7_1009));
wire output_9_1009, output_9_2, output_8_1009;
mixer gate_output_8_1009(.a(output_9_1009), .b(output_9_2), .y(output_8_1009));
wire output_10_1009, output_10_2, output_9_1009;
mixer gate_output_9_1009(.a(output_10_1009), .b(output_10_2), .y(output_9_1009));
wire output_11_1009, output_11_2, output_10_1009;
mixer gate_output_10_1009(.a(output_11_1009), .b(output_11_2), .y(output_10_1009));
wire output_12_1009, output_12_2, output_11_1009;
mixer gate_output_11_1009(.a(output_12_1009), .b(output_12_2), .y(output_11_1009));
wire output_13_1009, output_13_2, output_12_1009;
mixer gate_output_12_1009(.a(output_13_1009), .b(output_13_2), .y(output_12_1009));
wire output_14_1009, output_14_2, output_13_1009;
mixer gate_output_13_1009(.a(output_14_1009), .b(output_14_2), .y(output_13_1009));
wire output_15_1009, output_15_2, output_14_1009;
mixer gate_output_14_1009(.a(output_15_1009), .b(output_15_2), .y(output_14_1009));
wire output_16_1009, output_16_2, output_15_1009;
mixer gate_output_15_1009(.a(output_16_1009), .b(output_16_2), .y(output_15_1009));
wire output_1_1010, output_1_3, output_0_1010;
mixer gate_output_0_1010(.a(output_1_1010), .b(output_1_3), .y(output_0_1010));
wire output_2_1010, output_2_3, output_1_1010;
mixer gate_output_1_1010(.a(output_2_1010), .b(output_2_3), .y(output_1_1010));
wire output_3_1010, output_3_3, output_2_1010;
mixer gate_output_2_1010(.a(output_3_1010), .b(output_3_3), .y(output_2_1010));
wire output_4_1010, output_4_3, output_3_1010;
mixer gate_output_3_1010(.a(output_4_1010), .b(output_4_3), .y(output_3_1010));
wire output_5_1010, output_5_3, output_4_1010;
mixer gate_output_4_1010(.a(output_5_1010), .b(output_5_3), .y(output_4_1010));
wire output_6_1010, output_6_3, output_5_1010;
mixer gate_output_5_1010(.a(output_6_1010), .b(output_6_3), .y(output_5_1010));
wire output_7_1010, output_7_3, output_6_1010;
mixer gate_output_6_1010(.a(output_7_1010), .b(output_7_3), .y(output_6_1010));
wire output_8_1010, output_8_3, output_7_1010;
mixer gate_output_7_1010(.a(output_8_1010), .b(output_8_3), .y(output_7_1010));
wire output_9_1010, output_9_3, output_8_1010;
mixer gate_output_8_1010(.a(output_9_1010), .b(output_9_3), .y(output_8_1010));
wire output_10_1010, output_10_3, output_9_1010;
mixer gate_output_9_1010(.a(output_10_1010), .b(output_10_3), .y(output_9_1010));
wire output_11_1010, output_11_3, output_10_1010;
mixer gate_output_10_1010(.a(output_11_1010), .b(output_11_3), .y(output_10_1010));
wire output_12_1010, output_12_3, output_11_1010;
mixer gate_output_11_1010(.a(output_12_1010), .b(output_12_3), .y(output_11_1010));
wire output_13_1010, output_13_3, output_12_1010;
mixer gate_output_12_1010(.a(output_13_1010), .b(output_13_3), .y(output_12_1010));
wire output_14_1010, output_14_3, output_13_1010;
mixer gate_output_13_1010(.a(output_14_1010), .b(output_14_3), .y(output_13_1010));
wire output_15_1010, output_15_3, output_14_1010;
mixer gate_output_14_1010(.a(output_15_1010), .b(output_15_3), .y(output_14_1010));
wire output_16_1010, output_16_3, output_15_1010;
mixer gate_output_15_1010(.a(output_16_1010), .b(output_16_3), .y(output_15_1010));
wire output_1_1011, output_1_4, output_0_1011;
mixer gate_output_0_1011(.a(output_1_1011), .b(output_1_4), .y(output_0_1011));
wire output_2_1011, output_2_4, output_1_1011;
mixer gate_output_1_1011(.a(output_2_1011), .b(output_2_4), .y(output_1_1011));
wire output_3_1011, output_3_4, output_2_1011;
mixer gate_output_2_1011(.a(output_3_1011), .b(output_3_4), .y(output_2_1011));
wire output_4_1011, output_4_4, output_3_1011;
mixer gate_output_3_1011(.a(output_4_1011), .b(output_4_4), .y(output_3_1011));
wire output_5_1011, output_5_4, output_4_1011;
mixer gate_output_4_1011(.a(output_5_1011), .b(output_5_4), .y(output_4_1011));
wire output_6_1011, output_6_4, output_5_1011;
mixer gate_output_5_1011(.a(output_6_1011), .b(output_6_4), .y(output_5_1011));
wire output_7_1011, output_7_4, output_6_1011;
mixer gate_output_6_1011(.a(output_7_1011), .b(output_7_4), .y(output_6_1011));
wire output_8_1011, output_8_4, output_7_1011;
mixer gate_output_7_1011(.a(output_8_1011), .b(output_8_4), .y(output_7_1011));
wire output_9_1011, output_9_4, output_8_1011;
mixer gate_output_8_1011(.a(output_9_1011), .b(output_9_4), .y(output_8_1011));
wire output_10_1011, output_10_4, output_9_1011;
mixer gate_output_9_1011(.a(output_10_1011), .b(output_10_4), .y(output_9_1011));
wire output_11_1011, output_11_4, output_10_1011;
mixer gate_output_10_1011(.a(output_11_1011), .b(output_11_4), .y(output_10_1011));
wire output_12_1011, output_12_4, output_11_1011;
mixer gate_output_11_1011(.a(output_12_1011), .b(output_12_4), .y(output_11_1011));
wire output_13_1011, output_13_4, output_12_1011;
mixer gate_output_12_1011(.a(output_13_1011), .b(output_13_4), .y(output_12_1011));
wire output_14_1011, output_14_4, output_13_1011;
mixer gate_output_13_1011(.a(output_14_1011), .b(output_14_4), .y(output_13_1011));
wire output_15_1011, output_15_4, output_14_1011;
mixer gate_output_14_1011(.a(output_15_1011), .b(output_15_4), .y(output_14_1011));
wire output_16_1011, output_16_4, output_15_1011;
mixer gate_output_15_1011(.a(output_16_1011), .b(output_16_4), .y(output_15_1011));
wire output_1_1012, output_1_5, output_0_1012;
mixer gate_output_0_1012(.a(output_1_1012), .b(output_1_5), .y(output_0_1012));
wire output_2_1012, output_2_5, output_1_1012;
mixer gate_output_1_1012(.a(output_2_1012), .b(output_2_5), .y(output_1_1012));
wire output_3_1012, output_3_5, output_2_1012;
mixer gate_output_2_1012(.a(output_3_1012), .b(output_3_5), .y(output_2_1012));
wire output_4_1012, output_4_5, output_3_1012;
mixer gate_output_3_1012(.a(output_4_1012), .b(output_4_5), .y(output_3_1012));
wire output_5_1012, output_5_5, output_4_1012;
mixer gate_output_4_1012(.a(output_5_1012), .b(output_5_5), .y(output_4_1012));
wire output_6_1012, output_6_5, output_5_1012;
mixer gate_output_5_1012(.a(output_6_1012), .b(output_6_5), .y(output_5_1012));
wire output_7_1012, output_7_5, output_6_1012;
mixer gate_output_6_1012(.a(output_7_1012), .b(output_7_5), .y(output_6_1012));
wire output_8_1012, output_8_5, output_7_1012;
mixer gate_output_7_1012(.a(output_8_1012), .b(output_8_5), .y(output_7_1012));
wire output_9_1012, output_9_5, output_8_1012;
mixer gate_output_8_1012(.a(output_9_1012), .b(output_9_5), .y(output_8_1012));
wire output_10_1012, output_10_5, output_9_1012;
mixer gate_output_9_1012(.a(output_10_1012), .b(output_10_5), .y(output_9_1012));
wire output_11_1012, output_11_5, output_10_1012;
mixer gate_output_10_1012(.a(output_11_1012), .b(output_11_5), .y(output_10_1012));
wire output_12_1012, output_12_5, output_11_1012;
mixer gate_output_11_1012(.a(output_12_1012), .b(output_12_5), .y(output_11_1012));
wire output_13_1012, output_13_5, output_12_1012;
mixer gate_output_12_1012(.a(output_13_1012), .b(output_13_5), .y(output_12_1012));
wire output_14_1012, output_14_5, output_13_1012;
mixer gate_output_13_1012(.a(output_14_1012), .b(output_14_5), .y(output_13_1012));
wire output_15_1012, output_15_5, output_14_1012;
mixer gate_output_14_1012(.a(output_15_1012), .b(output_15_5), .y(output_14_1012));
wire output_16_1012, output_16_5, output_15_1012;
mixer gate_output_15_1012(.a(output_16_1012), .b(output_16_5), .y(output_15_1012));
wire output_1_1013, output_1_6, output_0_1013;
mixer gate_output_0_1013(.a(output_1_1013), .b(output_1_6), .y(output_0_1013));
wire output_2_1013, output_2_6, output_1_1013;
mixer gate_output_1_1013(.a(output_2_1013), .b(output_2_6), .y(output_1_1013));
wire output_3_1013, output_3_6, output_2_1013;
mixer gate_output_2_1013(.a(output_3_1013), .b(output_3_6), .y(output_2_1013));
wire output_4_1013, output_4_6, output_3_1013;
mixer gate_output_3_1013(.a(output_4_1013), .b(output_4_6), .y(output_3_1013));
wire output_5_1013, output_5_6, output_4_1013;
mixer gate_output_4_1013(.a(output_5_1013), .b(output_5_6), .y(output_4_1013));
wire output_6_1013, output_6_6, output_5_1013;
mixer gate_output_5_1013(.a(output_6_1013), .b(output_6_6), .y(output_5_1013));
wire output_7_1013, output_7_6, output_6_1013;
mixer gate_output_6_1013(.a(output_7_1013), .b(output_7_6), .y(output_6_1013));
wire output_8_1013, output_8_6, output_7_1013;
mixer gate_output_7_1013(.a(output_8_1013), .b(output_8_6), .y(output_7_1013));
wire output_9_1013, output_9_6, output_8_1013;
mixer gate_output_8_1013(.a(output_9_1013), .b(output_9_6), .y(output_8_1013));
wire output_10_1013, output_10_6, output_9_1013;
mixer gate_output_9_1013(.a(output_10_1013), .b(output_10_6), .y(output_9_1013));
wire output_11_1013, output_11_6, output_10_1013;
mixer gate_output_10_1013(.a(output_11_1013), .b(output_11_6), .y(output_10_1013));
wire output_12_1013, output_12_6, output_11_1013;
mixer gate_output_11_1013(.a(output_12_1013), .b(output_12_6), .y(output_11_1013));
wire output_13_1013, output_13_6, output_12_1013;
mixer gate_output_12_1013(.a(output_13_1013), .b(output_13_6), .y(output_12_1013));
wire output_14_1013, output_14_6, output_13_1013;
mixer gate_output_13_1013(.a(output_14_1013), .b(output_14_6), .y(output_13_1013));
wire output_15_1013, output_15_6, output_14_1013;
mixer gate_output_14_1013(.a(output_15_1013), .b(output_15_6), .y(output_14_1013));
wire output_16_1013, output_16_6, output_15_1013;
mixer gate_output_15_1013(.a(output_16_1013), .b(output_16_6), .y(output_15_1013));
wire output_1_1014, output_1_7, output_0_1014;
mixer gate_output_0_1014(.a(output_1_1014), .b(output_1_7), .y(output_0_1014));
wire output_2_1014, output_2_7, output_1_1014;
mixer gate_output_1_1014(.a(output_2_1014), .b(output_2_7), .y(output_1_1014));
wire output_3_1014, output_3_7, output_2_1014;
mixer gate_output_2_1014(.a(output_3_1014), .b(output_3_7), .y(output_2_1014));
wire output_4_1014, output_4_7, output_3_1014;
mixer gate_output_3_1014(.a(output_4_1014), .b(output_4_7), .y(output_3_1014));
wire output_5_1014, output_5_7, output_4_1014;
mixer gate_output_4_1014(.a(output_5_1014), .b(output_5_7), .y(output_4_1014));
wire output_6_1014, output_6_7, output_5_1014;
mixer gate_output_5_1014(.a(output_6_1014), .b(output_6_7), .y(output_5_1014));
wire output_7_1014, output_7_7, output_6_1014;
mixer gate_output_6_1014(.a(output_7_1014), .b(output_7_7), .y(output_6_1014));
wire output_8_1014, output_8_7, output_7_1014;
mixer gate_output_7_1014(.a(output_8_1014), .b(output_8_7), .y(output_7_1014));
wire output_9_1014, output_9_7, output_8_1014;
mixer gate_output_8_1014(.a(output_9_1014), .b(output_9_7), .y(output_8_1014));
wire output_10_1014, output_10_7, output_9_1014;
mixer gate_output_9_1014(.a(output_10_1014), .b(output_10_7), .y(output_9_1014));
wire output_11_1014, output_11_7, output_10_1014;
mixer gate_output_10_1014(.a(output_11_1014), .b(output_11_7), .y(output_10_1014));
wire output_12_1014, output_12_7, output_11_1014;
mixer gate_output_11_1014(.a(output_12_1014), .b(output_12_7), .y(output_11_1014));
wire output_13_1014, output_13_7, output_12_1014;
mixer gate_output_12_1014(.a(output_13_1014), .b(output_13_7), .y(output_12_1014));
wire output_14_1014, output_14_7, output_13_1014;
mixer gate_output_13_1014(.a(output_14_1014), .b(output_14_7), .y(output_13_1014));
wire output_15_1014, output_15_7, output_14_1014;
mixer gate_output_14_1014(.a(output_15_1014), .b(output_15_7), .y(output_14_1014));
wire output_16_1014, output_16_7, output_15_1014;
mixer gate_output_15_1014(.a(output_16_1014), .b(output_16_7), .y(output_15_1014));
wire output_1_1015, output_1_8, output_0_1015;
mixer gate_output_0_1015(.a(output_1_1015), .b(output_1_8), .y(output_0_1015));
wire output_2_1015, output_2_8, output_1_1015;
mixer gate_output_1_1015(.a(output_2_1015), .b(output_2_8), .y(output_1_1015));
wire output_3_1015, output_3_8, output_2_1015;
mixer gate_output_2_1015(.a(output_3_1015), .b(output_3_8), .y(output_2_1015));
wire output_4_1015, output_4_8, output_3_1015;
mixer gate_output_3_1015(.a(output_4_1015), .b(output_4_8), .y(output_3_1015));
wire output_5_1015, output_5_8, output_4_1015;
mixer gate_output_4_1015(.a(output_5_1015), .b(output_5_8), .y(output_4_1015));
wire output_6_1015, output_6_8, output_5_1015;
mixer gate_output_5_1015(.a(output_6_1015), .b(output_6_8), .y(output_5_1015));
wire output_7_1015, output_7_8, output_6_1015;
mixer gate_output_6_1015(.a(output_7_1015), .b(output_7_8), .y(output_6_1015));
wire output_8_1015, output_8_8, output_7_1015;
mixer gate_output_7_1015(.a(output_8_1015), .b(output_8_8), .y(output_7_1015));
wire output_9_1015, output_9_8, output_8_1015;
mixer gate_output_8_1015(.a(output_9_1015), .b(output_9_8), .y(output_8_1015));
wire output_10_1015, output_10_8, output_9_1015;
mixer gate_output_9_1015(.a(output_10_1015), .b(output_10_8), .y(output_9_1015));
wire output_11_1015, output_11_8, output_10_1015;
mixer gate_output_10_1015(.a(output_11_1015), .b(output_11_8), .y(output_10_1015));
wire output_12_1015, output_12_8, output_11_1015;
mixer gate_output_11_1015(.a(output_12_1015), .b(output_12_8), .y(output_11_1015));
wire output_13_1015, output_13_8, output_12_1015;
mixer gate_output_12_1015(.a(output_13_1015), .b(output_13_8), .y(output_12_1015));
wire output_14_1015, output_14_8, output_13_1015;
mixer gate_output_13_1015(.a(output_14_1015), .b(output_14_8), .y(output_13_1015));
wire output_15_1015, output_15_8, output_14_1015;
mixer gate_output_14_1015(.a(output_15_1015), .b(output_15_8), .y(output_14_1015));
wire output_16_1015, output_16_8, output_15_1015;
mixer gate_output_15_1015(.a(output_16_1015), .b(output_16_8), .y(output_15_1015));
wire output_1_1016, output_1_9, output_0_1016;
mixer gate_output_0_1016(.a(output_1_1016), .b(output_1_9), .y(output_0_1016));
wire output_2_1016, output_2_9, output_1_1016;
mixer gate_output_1_1016(.a(output_2_1016), .b(output_2_9), .y(output_1_1016));
wire output_3_1016, output_3_9, output_2_1016;
mixer gate_output_2_1016(.a(output_3_1016), .b(output_3_9), .y(output_2_1016));
wire output_4_1016, output_4_9, output_3_1016;
mixer gate_output_3_1016(.a(output_4_1016), .b(output_4_9), .y(output_3_1016));
wire output_5_1016, output_5_9, output_4_1016;
mixer gate_output_4_1016(.a(output_5_1016), .b(output_5_9), .y(output_4_1016));
wire output_6_1016, output_6_9, output_5_1016;
mixer gate_output_5_1016(.a(output_6_1016), .b(output_6_9), .y(output_5_1016));
wire output_7_1016, output_7_9, output_6_1016;
mixer gate_output_6_1016(.a(output_7_1016), .b(output_7_9), .y(output_6_1016));
wire output_8_1016, output_8_9, output_7_1016;
mixer gate_output_7_1016(.a(output_8_1016), .b(output_8_9), .y(output_7_1016));
wire output_9_1016, output_9_9, output_8_1016;
mixer gate_output_8_1016(.a(output_9_1016), .b(output_9_9), .y(output_8_1016));
wire output_10_1016, output_10_9, output_9_1016;
mixer gate_output_9_1016(.a(output_10_1016), .b(output_10_9), .y(output_9_1016));
wire output_11_1016, output_11_9, output_10_1016;
mixer gate_output_10_1016(.a(output_11_1016), .b(output_11_9), .y(output_10_1016));
wire output_12_1016, output_12_9, output_11_1016;
mixer gate_output_11_1016(.a(output_12_1016), .b(output_12_9), .y(output_11_1016));
wire output_13_1016, output_13_9, output_12_1016;
mixer gate_output_12_1016(.a(output_13_1016), .b(output_13_9), .y(output_12_1016));
wire output_14_1016, output_14_9, output_13_1016;
mixer gate_output_13_1016(.a(output_14_1016), .b(output_14_9), .y(output_13_1016));
wire output_15_1016, output_15_9, output_14_1016;
mixer gate_output_14_1016(.a(output_15_1016), .b(output_15_9), .y(output_14_1016));
wire output_16_1016, output_16_9, output_15_1016;
mixer gate_output_15_1016(.a(output_16_1016), .b(output_16_9), .y(output_15_1016));
wire output_1_1017, output_1_10, output_0_1017;
mixer gate_output_0_1017(.a(output_1_1017), .b(output_1_10), .y(output_0_1017));
wire output_2_1017, output_2_10, output_1_1017;
mixer gate_output_1_1017(.a(output_2_1017), .b(output_2_10), .y(output_1_1017));
wire output_3_1017, output_3_10, output_2_1017;
mixer gate_output_2_1017(.a(output_3_1017), .b(output_3_10), .y(output_2_1017));
wire output_4_1017, output_4_10, output_3_1017;
mixer gate_output_3_1017(.a(output_4_1017), .b(output_4_10), .y(output_3_1017));
wire output_5_1017, output_5_10, output_4_1017;
mixer gate_output_4_1017(.a(output_5_1017), .b(output_5_10), .y(output_4_1017));
wire output_6_1017, output_6_10, output_5_1017;
mixer gate_output_5_1017(.a(output_6_1017), .b(output_6_10), .y(output_5_1017));
wire output_7_1017, output_7_10, output_6_1017;
mixer gate_output_6_1017(.a(output_7_1017), .b(output_7_10), .y(output_6_1017));
wire output_8_1017, output_8_10, output_7_1017;
mixer gate_output_7_1017(.a(output_8_1017), .b(output_8_10), .y(output_7_1017));
wire output_9_1017, output_9_10, output_8_1017;
mixer gate_output_8_1017(.a(output_9_1017), .b(output_9_10), .y(output_8_1017));
wire output_10_1017, output_10_10, output_9_1017;
mixer gate_output_9_1017(.a(output_10_1017), .b(output_10_10), .y(output_9_1017));
wire output_11_1017, output_11_10, output_10_1017;
mixer gate_output_10_1017(.a(output_11_1017), .b(output_11_10), .y(output_10_1017));
wire output_12_1017, output_12_10, output_11_1017;
mixer gate_output_11_1017(.a(output_12_1017), .b(output_12_10), .y(output_11_1017));
wire output_13_1017, output_13_10, output_12_1017;
mixer gate_output_12_1017(.a(output_13_1017), .b(output_13_10), .y(output_12_1017));
wire output_14_1017, output_14_10, output_13_1017;
mixer gate_output_13_1017(.a(output_14_1017), .b(output_14_10), .y(output_13_1017));
wire output_15_1017, output_15_10, output_14_1017;
mixer gate_output_14_1017(.a(output_15_1017), .b(output_15_10), .y(output_14_1017));
wire output_16_1017, output_16_10, output_15_1017;
mixer gate_output_15_1017(.a(output_16_1017), .b(output_16_10), .y(output_15_1017));
wire output_1_1018, output_1_11, output_0_1018;
mixer gate_output_0_1018(.a(output_1_1018), .b(output_1_11), .y(output_0_1018));
wire output_2_1018, output_2_11, output_1_1018;
mixer gate_output_1_1018(.a(output_2_1018), .b(output_2_11), .y(output_1_1018));
wire output_3_1018, output_3_11, output_2_1018;
mixer gate_output_2_1018(.a(output_3_1018), .b(output_3_11), .y(output_2_1018));
wire output_4_1018, output_4_11, output_3_1018;
mixer gate_output_3_1018(.a(output_4_1018), .b(output_4_11), .y(output_3_1018));
wire output_5_1018, output_5_11, output_4_1018;
mixer gate_output_4_1018(.a(output_5_1018), .b(output_5_11), .y(output_4_1018));
wire output_6_1018, output_6_11, output_5_1018;
mixer gate_output_5_1018(.a(output_6_1018), .b(output_6_11), .y(output_5_1018));
wire output_7_1018, output_7_11, output_6_1018;
mixer gate_output_6_1018(.a(output_7_1018), .b(output_7_11), .y(output_6_1018));
wire output_8_1018, output_8_11, output_7_1018;
mixer gate_output_7_1018(.a(output_8_1018), .b(output_8_11), .y(output_7_1018));
wire output_9_1018, output_9_11, output_8_1018;
mixer gate_output_8_1018(.a(output_9_1018), .b(output_9_11), .y(output_8_1018));
wire output_10_1018, output_10_11, output_9_1018;
mixer gate_output_9_1018(.a(output_10_1018), .b(output_10_11), .y(output_9_1018));
wire output_11_1018, output_11_11, output_10_1018;
mixer gate_output_10_1018(.a(output_11_1018), .b(output_11_11), .y(output_10_1018));
wire output_12_1018, output_12_11, output_11_1018;
mixer gate_output_11_1018(.a(output_12_1018), .b(output_12_11), .y(output_11_1018));
wire output_13_1018, output_13_11, output_12_1018;
mixer gate_output_12_1018(.a(output_13_1018), .b(output_13_11), .y(output_12_1018));
wire output_14_1018, output_14_11, output_13_1018;
mixer gate_output_13_1018(.a(output_14_1018), .b(output_14_11), .y(output_13_1018));
wire output_15_1018, output_15_11, output_14_1018;
mixer gate_output_14_1018(.a(output_15_1018), .b(output_15_11), .y(output_14_1018));
wire output_16_1018, output_16_11, output_15_1018;
mixer gate_output_15_1018(.a(output_16_1018), .b(output_16_11), .y(output_15_1018));
wire output_1_1019, output_1_12, output_0_1019;
mixer gate_output_0_1019(.a(output_1_1019), .b(output_1_12), .y(output_0_1019));
wire output_2_1019, output_2_12, output_1_1019;
mixer gate_output_1_1019(.a(output_2_1019), .b(output_2_12), .y(output_1_1019));
wire output_3_1019, output_3_12, output_2_1019;
mixer gate_output_2_1019(.a(output_3_1019), .b(output_3_12), .y(output_2_1019));
wire output_4_1019, output_4_12, output_3_1019;
mixer gate_output_3_1019(.a(output_4_1019), .b(output_4_12), .y(output_3_1019));
wire output_5_1019, output_5_12, output_4_1019;
mixer gate_output_4_1019(.a(output_5_1019), .b(output_5_12), .y(output_4_1019));
wire output_6_1019, output_6_12, output_5_1019;
mixer gate_output_5_1019(.a(output_6_1019), .b(output_6_12), .y(output_5_1019));
wire output_7_1019, output_7_12, output_6_1019;
mixer gate_output_6_1019(.a(output_7_1019), .b(output_7_12), .y(output_6_1019));
wire output_8_1019, output_8_12, output_7_1019;
mixer gate_output_7_1019(.a(output_8_1019), .b(output_8_12), .y(output_7_1019));
wire output_9_1019, output_9_12, output_8_1019;
mixer gate_output_8_1019(.a(output_9_1019), .b(output_9_12), .y(output_8_1019));
wire output_10_1019, output_10_12, output_9_1019;
mixer gate_output_9_1019(.a(output_10_1019), .b(output_10_12), .y(output_9_1019));
wire output_11_1019, output_11_12, output_10_1019;
mixer gate_output_10_1019(.a(output_11_1019), .b(output_11_12), .y(output_10_1019));
wire output_12_1019, output_12_12, output_11_1019;
mixer gate_output_11_1019(.a(output_12_1019), .b(output_12_12), .y(output_11_1019));
wire output_13_1019, output_13_12, output_12_1019;
mixer gate_output_12_1019(.a(output_13_1019), .b(output_13_12), .y(output_12_1019));
wire output_14_1019, output_14_12, output_13_1019;
mixer gate_output_13_1019(.a(output_14_1019), .b(output_14_12), .y(output_13_1019));
wire output_15_1019, output_15_12, output_14_1019;
mixer gate_output_14_1019(.a(output_15_1019), .b(output_15_12), .y(output_14_1019));
wire output_16_1019, output_16_12, output_15_1019;
mixer gate_output_15_1019(.a(output_16_1019), .b(output_16_12), .y(output_15_1019));
wire output_1_1020, output_1_13, output_0_1020;
mixer gate_output_0_1020(.a(output_1_1020), .b(output_1_13), .y(output_0_1020));
wire output_2_1020, output_2_13, output_1_1020;
mixer gate_output_1_1020(.a(output_2_1020), .b(output_2_13), .y(output_1_1020));
wire output_3_1020, output_3_13, output_2_1020;
mixer gate_output_2_1020(.a(output_3_1020), .b(output_3_13), .y(output_2_1020));
wire output_4_1020, output_4_13, output_3_1020;
mixer gate_output_3_1020(.a(output_4_1020), .b(output_4_13), .y(output_3_1020));
wire output_5_1020, output_5_13, output_4_1020;
mixer gate_output_4_1020(.a(output_5_1020), .b(output_5_13), .y(output_4_1020));
wire output_6_1020, output_6_13, output_5_1020;
mixer gate_output_5_1020(.a(output_6_1020), .b(output_6_13), .y(output_5_1020));
wire output_7_1020, output_7_13, output_6_1020;
mixer gate_output_6_1020(.a(output_7_1020), .b(output_7_13), .y(output_6_1020));
wire output_8_1020, output_8_13, output_7_1020;
mixer gate_output_7_1020(.a(output_8_1020), .b(output_8_13), .y(output_7_1020));
wire output_9_1020, output_9_13, output_8_1020;
mixer gate_output_8_1020(.a(output_9_1020), .b(output_9_13), .y(output_8_1020));
wire output_10_1020, output_10_13, output_9_1020;
mixer gate_output_9_1020(.a(output_10_1020), .b(output_10_13), .y(output_9_1020));
wire output_11_1020, output_11_13, output_10_1020;
mixer gate_output_10_1020(.a(output_11_1020), .b(output_11_13), .y(output_10_1020));
wire output_12_1020, output_12_13, output_11_1020;
mixer gate_output_11_1020(.a(output_12_1020), .b(output_12_13), .y(output_11_1020));
wire output_13_1020, output_13_13, output_12_1020;
mixer gate_output_12_1020(.a(output_13_1020), .b(output_13_13), .y(output_12_1020));
wire output_14_1020, output_14_13, output_13_1020;
mixer gate_output_13_1020(.a(output_14_1020), .b(output_14_13), .y(output_13_1020));
wire output_15_1020, output_15_13, output_14_1020;
mixer gate_output_14_1020(.a(output_15_1020), .b(output_15_13), .y(output_14_1020));
wire output_16_1020, output_16_13, output_15_1020;
mixer gate_output_15_1020(.a(output_16_1020), .b(output_16_13), .y(output_15_1020));
wire output_1_1021, output_1_14, output_0_1021;
mixer gate_output_0_1021(.a(output_1_1021), .b(output_1_14), .y(output_0_1021));
wire output_2_1021, output_2_14, output_1_1021;
mixer gate_output_1_1021(.a(output_2_1021), .b(output_2_14), .y(output_1_1021));
wire output_3_1021, output_3_14, output_2_1021;
mixer gate_output_2_1021(.a(output_3_1021), .b(output_3_14), .y(output_2_1021));
wire output_4_1021, output_4_14, output_3_1021;
mixer gate_output_3_1021(.a(output_4_1021), .b(output_4_14), .y(output_3_1021));
wire output_5_1021, output_5_14, output_4_1021;
mixer gate_output_4_1021(.a(output_5_1021), .b(output_5_14), .y(output_4_1021));
wire output_6_1021, output_6_14, output_5_1021;
mixer gate_output_5_1021(.a(output_6_1021), .b(output_6_14), .y(output_5_1021));
wire output_7_1021, output_7_14, output_6_1021;
mixer gate_output_6_1021(.a(output_7_1021), .b(output_7_14), .y(output_6_1021));
wire output_8_1021, output_8_14, output_7_1021;
mixer gate_output_7_1021(.a(output_8_1021), .b(output_8_14), .y(output_7_1021));
wire output_9_1021, output_9_14, output_8_1021;
mixer gate_output_8_1021(.a(output_9_1021), .b(output_9_14), .y(output_8_1021));
wire output_10_1021, output_10_14, output_9_1021;
mixer gate_output_9_1021(.a(output_10_1021), .b(output_10_14), .y(output_9_1021));
wire output_11_1021, output_11_14, output_10_1021;
mixer gate_output_10_1021(.a(output_11_1021), .b(output_11_14), .y(output_10_1021));
wire output_12_1021, output_12_14, output_11_1021;
mixer gate_output_11_1021(.a(output_12_1021), .b(output_12_14), .y(output_11_1021));
wire output_13_1021, output_13_14, output_12_1021;
mixer gate_output_12_1021(.a(output_13_1021), .b(output_13_14), .y(output_12_1021));
wire output_14_1021, output_14_14, output_13_1021;
mixer gate_output_13_1021(.a(output_14_1021), .b(output_14_14), .y(output_13_1021));
wire output_15_1021, output_15_14, output_14_1021;
mixer gate_output_14_1021(.a(output_15_1021), .b(output_15_14), .y(output_14_1021));
wire output_16_1021, output_16_14, output_15_1021;
mixer gate_output_15_1021(.a(output_16_1021), .b(output_16_14), .y(output_15_1021));
wire output_1_1022, output_1_15, output_0_1022;
mixer gate_output_0_1022(.a(output_1_1022), .b(output_1_15), .y(output_0_1022));
wire output_2_1022, output_2_15, output_1_1022;
mixer gate_output_1_1022(.a(output_2_1022), .b(output_2_15), .y(output_1_1022));
wire output_3_1022, output_3_15, output_2_1022;
mixer gate_output_2_1022(.a(output_3_1022), .b(output_3_15), .y(output_2_1022));
wire output_4_1022, output_4_15, output_3_1022;
mixer gate_output_3_1022(.a(output_4_1022), .b(output_4_15), .y(output_3_1022));
wire output_5_1022, output_5_15, output_4_1022;
mixer gate_output_4_1022(.a(output_5_1022), .b(output_5_15), .y(output_4_1022));
wire output_6_1022, output_6_15, output_5_1022;
mixer gate_output_5_1022(.a(output_6_1022), .b(output_6_15), .y(output_5_1022));
wire output_7_1022, output_7_15, output_6_1022;
mixer gate_output_6_1022(.a(output_7_1022), .b(output_7_15), .y(output_6_1022));
wire output_8_1022, output_8_15, output_7_1022;
mixer gate_output_7_1022(.a(output_8_1022), .b(output_8_15), .y(output_7_1022));
wire output_9_1022, output_9_15, output_8_1022;
mixer gate_output_8_1022(.a(output_9_1022), .b(output_9_15), .y(output_8_1022));
wire output_10_1022, output_10_15, output_9_1022;
mixer gate_output_9_1022(.a(output_10_1022), .b(output_10_15), .y(output_9_1022));
wire output_11_1022, output_11_15, output_10_1022;
mixer gate_output_10_1022(.a(output_11_1022), .b(output_11_15), .y(output_10_1022));
wire output_12_1022, output_12_15, output_11_1022;
mixer gate_output_11_1022(.a(output_12_1022), .b(output_12_15), .y(output_11_1022));
wire output_13_1022, output_13_15, output_12_1022;
mixer gate_output_12_1022(.a(output_13_1022), .b(output_13_15), .y(output_12_1022));
wire output_14_1022, output_14_15, output_13_1022;
mixer gate_output_13_1022(.a(output_14_1022), .b(output_14_15), .y(output_13_1022));
wire output_15_1022, output_15_15, output_14_1022;
mixer gate_output_14_1022(.a(output_15_1022), .b(output_15_15), .y(output_14_1022));
wire output_16_1022, output_16_15, output_15_1022;
mixer gate_output_15_1022(.a(output_16_1022), .b(output_16_15), .y(output_15_1022));
wire output_1_1023, output_1_0, output_0_1023;
mixer gate_output_0_1023(.a(output_1_1023), .b(output_1_0), .y(output_0_1023));
wire output_2_1023, output_2_0, output_1_1023;
mixer gate_output_1_1023(.a(output_2_1023), .b(output_2_0), .y(output_1_1023));
wire output_3_1023, output_3_0, output_2_1023;
mixer gate_output_2_1023(.a(output_3_1023), .b(output_3_0), .y(output_2_1023));
wire output_4_1023, output_4_0, output_3_1023;
mixer gate_output_3_1023(.a(output_4_1023), .b(output_4_0), .y(output_3_1023));
wire output_5_1023, output_5_0, output_4_1023;
mixer gate_output_4_1023(.a(output_5_1023), .b(output_5_0), .y(output_4_1023));
wire output_6_1023, output_6_0, output_5_1023;
mixer gate_output_5_1023(.a(output_6_1023), .b(output_6_0), .y(output_5_1023));
wire output_7_1023, output_7_0, output_6_1023;
mixer gate_output_6_1023(.a(output_7_1023), .b(output_7_0), .y(output_6_1023));
wire output_8_1023, output_8_0, output_7_1023;
mixer gate_output_7_1023(.a(output_8_1023), .b(output_8_0), .y(output_7_1023));
wire output_9_1023, output_9_0, output_8_1023;
mixer gate_output_8_1023(.a(output_9_1023), .b(output_9_0), .y(output_8_1023));
wire output_10_1023, output_10_0, output_9_1023;
mixer gate_output_9_1023(.a(output_10_1023), .b(output_10_0), .y(output_9_1023));
wire output_11_1023, output_11_0, output_10_1023;
mixer gate_output_10_1023(.a(output_11_1023), .b(output_11_0), .y(output_10_1023));
wire output_12_1023, output_12_0, output_11_1023;
mixer gate_output_11_1023(.a(output_12_1023), .b(output_12_0), .y(output_11_1023));
wire output_13_1023, output_13_0, output_12_1023;
mixer gate_output_12_1023(.a(output_13_1023), .b(output_13_0), .y(output_12_1023));
wire output_14_1023, output_14_0, output_13_1023;
mixer gate_output_13_1023(.a(output_14_1023), .b(output_14_0), .y(output_13_1023));
wire output_15_1023, output_15_0, output_14_1023;
mixer gate_output_14_1023(.a(output_15_1023), .b(output_15_0), .y(output_14_1023));
wire output_16_1023, output_16_0, output_15_1023;
mixer gate_output_15_1023(.a(output_16_1023), .b(output_16_0), .y(output_15_1023));
assign output_0 = output_0_0;
wire output_0_1024;
assign output_0_1024 = input_0;
assign output_1 = output_1_0;
wire output_1_1024;
assign output_1_1024 = input_1;
assign output_2 = output_2_0;
wire output_2_1024;
assign output_2_1024 = input_2;
assign output_3 = output_3_0;
wire output_3_1024;
assign output_3_1024 = input_3;
assign output_4 = output_4_0;
wire output_4_1024;
assign output_4_1024 = input_4;
assign output_5 = output_5_0;
wire output_5_1024;
assign output_5_1024 = input_5;
assign output_6 = output_6_0;
wire output_6_1024;
assign output_6_1024 = input_6;
assign output_7 = output_7_0;
wire output_7_1024;
assign output_7_1024 = input_7;
assign output_8 = output_8_0;
wire output_8_1024;
assign output_8_1024 = input_8;
assign output_9 = output_9_0;
wire output_9_1024;
assign output_9_1024 = input_9;
assign output_10 = output_10_0;
wire output_10_1024;
assign output_10_1024 = input_10;
assign output_11 = output_11_0;
wire output_11_1024;
assign output_11_1024 = input_11;
assign output_12 = output_12_0;
wire output_12_1024;
assign output_12_1024 = input_12;
assign output_13 = output_13_0;
wire output_13_1024;
assign output_13_1024 = input_13;
assign output_14 = output_14_0;
wire output_14_1024;
assign output_14_1024 = input_14;
assign output_15 = output_15_0;
wire output_15_1024;
assign output_15_1024 = input_15;
endmodule
