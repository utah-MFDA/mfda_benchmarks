module chain_64 (
inout k0, k64
);
wire {wires};
chamber ch0 (.in(k0), .out(k1)
chamber ch1 (.in(k1), .out(k2)
chamber ch2 (.in(k2), .out(k3)
chamber ch3 (.in(k3), .out(k4)
chamber ch4 (.in(k4), .out(k5)
chamber ch5 (.in(k5), .out(k6)
chamber ch6 (.in(k6), .out(k7)
chamber ch7 (.in(k7), .out(k8)
chamber ch8 (.in(k8), .out(k9)
chamber ch9 (.in(k9), .out(k10)
chamber ch10 (.in(k10), .out(k11)
chamber ch11 (.in(k11), .out(k12)
chamber ch12 (.in(k12), .out(k13)
chamber ch13 (.in(k13), .out(k14)
chamber ch14 (.in(k14), .out(k15)
chamber ch15 (.in(k15), .out(k16)
chamber ch16 (.in(k16), .out(k17)
chamber ch17 (.in(k17), .out(k18)
chamber ch18 (.in(k18), .out(k19)
chamber ch19 (.in(k19), .out(k20)
chamber ch20 (.in(k20), .out(k21)
chamber ch21 (.in(k21), .out(k22)
chamber ch22 (.in(k22), .out(k23)
chamber ch23 (.in(k23), .out(k24)
chamber ch24 (.in(k24), .out(k25)
chamber ch25 (.in(k25), .out(k26)
chamber ch26 (.in(k26), .out(k27)
chamber ch27 (.in(k27), .out(k28)
chamber ch28 (.in(k28), .out(k29)
chamber ch29 (.in(k29), .out(k30)
chamber ch30 (.in(k30), .out(k31)
chamber ch31 (.in(k31), .out(k32)
chamber ch32 (.in(k32), .out(k33)
chamber ch33 (.in(k33), .out(k34)
chamber ch34 (.in(k34), .out(k35)
chamber ch35 (.in(k35), .out(k36)
chamber ch36 (.in(k36), .out(k37)
chamber ch37 (.in(k37), .out(k38)
chamber ch38 (.in(k38), .out(k39)
chamber ch39 (.in(k39), .out(k40)
chamber ch40 (.in(k40), .out(k41)
chamber ch41 (.in(k41), .out(k42)
chamber ch42 (.in(k42), .out(k43)
chamber ch43 (.in(k43), .out(k44)
chamber ch44 (.in(k44), .out(k45)
chamber ch45 (.in(k45), .out(k46)
chamber ch46 (.in(k46), .out(k47)
chamber ch47 (.in(k47), .out(k48)
chamber ch48 (.in(k48), .out(k49)
chamber ch49 (.in(k49), .out(k50)
chamber ch50 (.in(k50), .out(k51)
chamber ch51 (.in(k51), .out(k52)
chamber ch52 (.in(k52), .out(k53)
chamber ch53 (.in(k53), .out(k54)
chamber ch54 (.in(k54), .out(k55)
chamber ch55 (.in(k55), .out(k56)
chamber ch56 (.in(k56), .out(k57)
chamber ch57 (.in(k57), .out(k58)
chamber ch58 (.in(k58), .out(k59)
chamber ch59 (.in(k59), .out(k60)
chamber ch60 (.in(k60), .out(k61)
chamber ch61 (.in(k61), .out(k62)
chamber ch62 (.in(k62), .out(k63)
chamber ch63 (.in(k63), .out(k64)
endmodule
