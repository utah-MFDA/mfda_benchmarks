module multiplexer_10 (
inout k_0_0,k_10_0,k_10_1,k_10_2,k_10_3,k_10_4,k_10_5,k_10_6,k_10_7,k_10_8,k_10_9,k_10_10,k_10_11,k_10_12,k_10_13,k_10_14,k_10_15,k_10_16,k_10_17,k_10_18,k_10_19,k_10_20,k_10_21,k_10_22,k_10_23,k_10_24,k_10_25,k_10_26,k_10_27,k_10_28,k_10_29,k_10_30,k_10_31,k_10_32,k_10_33,k_10_34,k_10_35,k_10_36,k_10_37,k_10_38,k_10_39,k_10_40,k_10_41,k_10_42,k_10_43,k_10_44,k_10_45,k_10_46,k_10_47,k_10_48,k_10_49,k_10_50,k_10_51,k_10_52,k_10_53,k_10_54,k_10_55,k_10_56,k_10_57,k_10_58,k_10_59,k_10_60,k_10_61,k_10_62,k_10_63,k_10_64,k_10_65,k_10_66,k_10_67,k_10_68,k_10_69,k_10_70,k_10_71,k_10_72,k_10_73,k_10_74,k_10_75,k_10_76,k_10_77,k_10_78,k_10_79,k_10_80,k_10_81,k_10_82,k_10_83,k_10_84,k_10_85,k_10_86,k_10_87,k_10_88,k_10_89,k_10_90,k_10_91,k_10_92,k_10_93,k_10_94,k_10_95,k_10_96,k_10_97,k_10_98,k_10_99,k_10_100,k_10_101,k_10_102,k_10_103,k_10_104,k_10_105,k_10_106,k_10_107,k_10_108,k_10_109,k_10_110,k_10_111,k_10_112,k_10_113,k_10_114,k_10_115,k_10_116,k_10_117,k_10_118,k_10_119,k_10_120,k_10_121,k_10_122,k_10_123,k_10_124,k_10_125,k_10_126,k_10_127,k_10_128,k_10_129,k_10_130,k_10_131,k_10_132,k_10_133,k_10_134,k_10_135,k_10_136,k_10_137,k_10_138,k_10_139,k_10_140,k_10_141,k_10_142,k_10_143,k_10_144,k_10_145,k_10_146,k_10_147,k_10_148,k_10_149,k_10_150,k_10_151,k_10_152,k_10_153,k_10_154,k_10_155,k_10_156,k_10_157,k_10_158,k_10_159,k_10_160,k_10_161,k_10_162,k_10_163,k_10_164,k_10_165,k_10_166,k_10_167,k_10_168,k_10_169,k_10_170,k_10_171,k_10_172,k_10_173,k_10_174,k_10_175,k_10_176,k_10_177,k_10_178,k_10_179,k_10_180,k_10_181,k_10_182,k_10_183,k_10_184,k_10_185,k_10_186,k_10_187,k_10_188,k_10_189,k_10_190,k_10_191,k_10_192,k_10_193,k_10_194,k_10_195,k_10_196,k_10_197,k_10_198,k_10_199,k_10_200,k_10_201,k_10_202,k_10_203,k_10_204,k_10_205,k_10_206,k_10_207,k_10_208,k_10_209,k_10_210,k_10_211,k_10_212,k_10_213,k_10_214,k_10_215,k_10_216,k_10_217,k_10_218,k_10_219,k_10_220,k_10_221,k_10_222,k_10_223,k_10_224,k_10_225,k_10_226,k_10_227,k_10_228,k_10_229,k_10_230,k_10_231,k_10_232,k_10_233,k_10_234,k_10_235,k_10_236,k_10_237,k_10_238,k_10_239,k_10_240,k_10_241,k_10_242,k_10_243,k_10_244,k_10_245,k_10_246,k_10_247,k_10_248,k_10_249,k_10_250,k_10_251,k_10_252,k_10_253,k_10_254,k_10_255,k_10_256,k_10_257,k_10_258,k_10_259,k_10_260,k_10_261,k_10_262,k_10_263,k_10_264,k_10_265,k_10_266,k_10_267,k_10_268,k_10_269,k_10_270,k_10_271,k_10_272,k_10_273,k_10_274,k_10_275,k_10_276,k_10_277,k_10_278,k_10_279,k_10_280,k_10_281,k_10_282,k_10_283,k_10_284,k_10_285,k_10_286,k_10_287,k_10_288,k_10_289,k_10_290,k_10_291,k_10_292,k_10_293,k_10_294,k_10_295,k_10_296,k_10_297,k_10_298,k_10_299,k_10_300,k_10_301,k_10_302,k_10_303,k_10_304,k_10_305,k_10_306,k_10_307,k_10_308,k_10_309,k_10_310,k_10_311,k_10_312,k_10_313,k_10_314,k_10_315,k_10_316,k_10_317,k_10_318,k_10_319,k_10_320,k_10_321,k_10_322,k_10_323,k_10_324,k_10_325,k_10_326,k_10_327,k_10_328,k_10_329,k_10_330,k_10_331,k_10_332,k_10_333,k_10_334,k_10_335,k_10_336,k_10_337,k_10_338,k_10_339,k_10_340,k_10_341,k_10_342,k_10_343,k_10_344,k_10_345,k_10_346,k_10_347,k_10_348,k_10_349,k_10_350,k_10_351,k_10_352,k_10_353,k_10_354,k_10_355,k_10_356,k_10_357,k_10_358,k_10_359,k_10_360,k_10_361,k_10_362,k_10_363,k_10_364,k_10_365,k_10_366,k_10_367,k_10_368,k_10_369,k_10_370,k_10_371,k_10_372,k_10_373,k_10_374,k_10_375,k_10_376,k_10_377,k_10_378,k_10_379,k_10_380,k_10_381,k_10_382,k_10_383,k_10_384,k_10_385,k_10_386,k_10_387,k_10_388,k_10_389,k_10_390,k_10_391,k_10_392,k_10_393,k_10_394,k_10_395,k_10_396,k_10_397,k_10_398,k_10_399,k_10_400,k_10_401,k_10_402,k_10_403,k_10_404,k_10_405,k_10_406,k_10_407,k_10_408,k_10_409,k_10_410,k_10_411,k_10_412,k_10_413,k_10_414,k_10_415,k_10_416,k_10_417,k_10_418,k_10_419,k_10_420,k_10_421,k_10_422,k_10_423,k_10_424,k_10_425,k_10_426,k_10_427,k_10_428,k_10_429,k_10_430,k_10_431,k_10_432,k_10_433,k_10_434,k_10_435,k_10_436,k_10_437,k_10_438,k_10_439,k_10_440,k_10_441,k_10_442,k_10_443,k_10_444,k_10_445,k_10_446,k_10_447,k_10_448,k_10_449,k_10_450,k_10_451,k_10_452,k_10_453,k_10_454,k_10_455,k_10_456,k_10_457,k_10_458,k_10_459,k_10_460,k_10_461,k_10_462,k_10_463,k_10_464,k_10_465,k_10_466,k_10_467,k_10_468,k_10_469,k_10_470,k_10_471,k_10_472,k_10_473,k_10_474,k_10_475,k_10_476,k_10_477,k_10_478,k_10_479,k_10_480,k_10_481,k_10_482,k_10_483,k_10_484,k_10_485,k_10_486,k_10_487,k_10_488,k_10_489,k_10_490,k_10_491,k_10_492,k_10_493,k_10_494,k_10_495,k_10_496,k_10_497,k_10_498,k_10_499,k_10_500,k_10_501,k_10_502,k_10_503,k_10_504,k_10_505,k_10_506,k_10_507,k_10_508,k_10_509,k_10_510,k_10_511,k_10_512,k_10_513,k_10_514,k_10_515,k_10_516,k_10_517,k_10_518,k_10_519,k_10_520,k_10_521,k_10_522,k_10_523,k_10_524,k_10_525,k_10_526,k_10_527,k_10_528,k_10_529,k_10_530,k_10_531,k_10_532,k_10_533,k_10_534,k_10_535,k_10_536,k_10_537,k_10_538,k_10_539,k_10_540,k_10_541,k_10_542,k_10_543,k_10_544,k_10_545,k_10_546,k_10_547,k_10_548,k_10_549,k_10_550,k_10_551,k_10_552,k_10_553,k_10_554,k_10_555,k_10_556,k_10_557,k_10_558,k_10_559,k_10_560,k_10_561,k_10_562,k_10_563,k_10_564,k_10_565,k_10_566,k_10_567,k_10_568,k_10_569,k_10_570,k_10_571,k_10_572,k_10_573,k_10_574,k_10_575,k_10_576,k_10_577,k_10_578,k_10_579,k_10_580,k_10_581,k_10_582,k_10_583,k_10_584,k_10_585,k_10_586,k_10_587,k_10_588,k_10_589,k_10_590,k_10_591,k_10_592,k_10_593,k_10_594,k_10_595,k_10_596,k_10_597,k_10_598,k_10_599,k_10_600,k_10_601,k_10_602,k_10_603,k_10_604,k_10_605,k_10_606,k_10_607,k_10_608,k_10_609,k_10_610,k_10_611,k_10_612,k_10_613,k_10_614,k_10_615,k_10_616,k_10_617,k_10_618,k_10_619,k_10_620,k_10_621,k_10_622,k_10_623,k_10_624,k_10_625,k_10_626,k_10_627,k_10_628,k_10_629,k_10_630,k_10_631,k_10_632,k_10_633,k_10_634,k_10_635,k_10_636,k_10_637,k_10_638,k_10_639,k_10_640,k_10_641,k_10_642,k_10_643,k_10_644,k_10_645,k_10_646,k_10_647,k_10_648,k_10_649,k_10_650,k_10_651,k_10_652,k_10_653,k_10_654,k_10_655,k_10_656,k_10_657,k_10_658,k_10_659,k_10_660,k_10_661,k_10_662,k_10_663,k_10_664,k_10_665,k_10_666,k_10_667,k_10_668,k_10_669,k_10_670,k_10_671,k_10_672,k_10_673,k_10_674,k_10_675,k_10_676,k_10_677,k_10_678,k_10_679,k_10_680,k_10_681,k_10_682,k_10_683,k_10_684,k_10_685,k_10_686,k_10_687,k_10_688,k_10_689,k_10_690,k_10_691,k_10_692,k_10_693,k_10_694,k_10_695,k_10_696,k_10_697,k_10_698,k_10_699,k_10_700,k_10_701,k_10_702,k_10_703,k_10_704,k_10_705,k_10_706,k_10_707,k_10_708,k_10_709,k_10_710,k_10_711,k_10_712,k_10_713,k_10_714,k_10_715,k_10_716,k_10_717,k_10_718,k_10_719,k_10_720,k_10_721,k_10_722,k_10_723,k_10_724,k_10_725,k_10_726,k_10_727,k_10_728,k_10_729,k_10_730,k_10_731,k_10_732,k_10_733,k_10_734,k_10_735,k_10_736,k_10_737,k_10_738,k_10_739,k_10_740,k_10_741,k_10_742,k_10_743,k_10_744,k_10_745,k_10_746,k_10_747,k_10_748,k_10_749,k_10_750,k_10_751,k_10_752,k_10_753,k_10_754,k_10_755,k_10_756,k_10_757,k_10_758,k_10_759,k_10_760,k_10_761,k_10_762,k_10_763,k_10_764,k_10_765,k_10_766,k_10_767,k_10_768,k_10_769,k_10_770,k_10_771,k_10_772,k_10_773,k_10_774,k_10_775,k_10_776,k_10_777,k_10_778,k_10_779,k_10_780,k_10_781,k_10_782,k_10_783,k_10_784,k_10_785,k_10_786,k_10_787,k_10_788,k_10_789,k_10_790,k_10_791,k_10_792,k_10_793,k_10_794,k_10_795,k_10_796,k_10_797,k_10_798,k_10_799,k_10_800,k_10_801,k_10_802,k_10_803,k_10_804,k_10_805,k_10_806,k_10_807,k_10_808,k_10_809,k_10_810,k_10_811,k_10_812,k_10_813,k_10_814,k_10_815,k_10_816,k_10_817,k_10_818,k_10_819,k_10_820,k_10_821,k_10_822,k_10_823,k_10_824,k_10_825,k_10_826,k_10_827,k_10_828,k_10_829,k_10_830,k_10_831,k_10_832,k_10_833,k_10_834,k_10_835,k_10_836,k_10_837,k_10_838,k_10_839,k_10_840,k_10_841,k_10_842,k_10_843,k_10_844,k_10_845,k_10_846,k_10_847,k_10_848,k_10_849,k_10_850,k_10_851,k_10_852,k_10_853,k_10_854,k_10_855,k_10_856,k_10_857,k_10_858,k_10_859,k_10_860,k_10_861,k_10_862,k_10_863,k_10_864,k_10_865,k_10_866,k_10_867,k_10_868,k_10_869,k_10_870,k_10_871,k_10_872,k_10_873,k_10_874,k_10_875,k_10_876,k_10_877,k_10_878,k_10_879,k_10_880,k_10_881,k_10_882,k_10_883,k_10_884,k_10_885,k_10_886,k_10_887,k_10_888,k_10_889,k_10_890,k_10_891,k_10_892,k_10_893,k_10_894,k_10_895,k_10_896,k_10_897,k_10_898,k_10_899,k_10_900,k_10_901,k_10_902,k_10_903,k_10_904,k_10_905,k_10_906,k_10_907,k_10_908,k_10_909,k_10_910,k_10_911,k_10_912,k_10_913,k_10_914,k_10_915,k_10_916,k_10_917,k_10_918,k_10_919,k_10_920,k_10_921,k_10_922,k_10_923,k_10_924,k_10_925,k_10_926,k_10_927,k_10_928,k_10_929,k_10_930,k_10_931,k_10_932,k_10_933,k_10_934,k_10_935,k_10_936,k_10_937,k_10_938,k_10_939,k_10_940,k_10_941,k_10_942,k_10_943,k_10_944,k_10_945,k_10_946,k_10_947,k_10_948,k_10_949,k_10_950,k_10_951,k_10_952,k_10_953,k_10_954,k_10_955,k_10_956,k_10_957,k_10_958,k_10_959,k_10_960,k_10_961,k_10_962,k_10_963,k_10_964,k_10_965,k_10_966,k_10_967,k_10_968,k_10_969,k_10_970,k_10_971,k_10_972,k_10_973,k_10_974,k_10_975,k_10_976,k_10_977,k_10_978,k_10_979,k_10_980,k_10_981,k_10_982,k_10_983,k_10_984,k_10_985,k_10_986,k_10_987,k_10_988,k_10_989,k_10_990,k_10_991,k_10_992,k_10_993,k_10_994,k_10_995,k_10_996,k_10_997,k_10_998,k_10_999,k_10_1000,k_10_1001,k_10_1002,k_10_1003,k_10_1004,k_10_1005,k_10_1006,k_10_1007,k_10_1008,k_10_1009,k_10_1010,k_10_1011,k_10_1012,k_10_1013,k_10_1014,k_10_1015,k_10_1016,k_10_1017,k_10_1018,k_10_1019,k_10_1020,k_10_1021,k_10_1022,k_10_1023,
input c_0_0, c_0_1,
input c_1_0, c_1_1,
input c_2_0, c_2_1,
input c_3_0, c_3_1,
input c_4_0, c_4_1,
input c_5_0, c_5_1,
input c_6_0, c_6_1,
input c_7_0, c_7_1,
input c_8_0, c_8_1,
input c_9_0, c_9_1,
input c_10_0, c_10_1
);
wire k_1_0,k_1_1;
wire k_2_0,k_2_1,k_2_2,k_2_3;
wire k_3_0,k_3_1,k_3_2,k_3_3,k_3_4,k_3_5,k_3_6,k_3_7;
wire k_4_0,k_4_1,k_4_2,k_4_3,k_4_4,k_4_5,k_4_6,k_4_7,k_4_8,k_4_9,k_4_10,k_4_11,k_4_12,k_4_13,k_4_14,k_4_15;
wire k_5_0,k_5_1,k_5_2,k_5_3,k_5_4,k_5_5,k_5_6,k_5_7,k_5_8,k_5_9,k_5_10,k_5_11,k_5_12,k_5_13,k_5_14,k_5_15,k_5_16,k_5_17,k_5_18,k_5_19,k_5_20,k_5_21,k_5_22,k_5_23,k_5_24,k_5_25,k_5_26,k_5_27,k_5_28,k_5_29,k_5_30,k_5_31;
wire k_6_0,k_6_1,k_6_2,k_6_3,k_6_4,k_6_5,k_6_6,k_6_7,k_6_8,k_6_9,k_6_10,k_6_11,k_6_12,k_6_13,k_6_14,k_6_15,k_6_16,k_6_17,k_6_18,k_6_19,k_6_20,k_6_21,k_6_22,k_6_23,k_6_24,k_6_25,k_6_26,k_6_27,k_6_28,k_6_29,k_6_30,k_6_31,k_6_32,k_6_33,k_6_34,k_6_35,k_6_36,k_6_37,k_6_38,k_6_39,k_6_40,k_6_41,k_6_42,k_6_43,k_6_44,k_6_45,k_6_46,k_6_47,k_6_48,k_6_49,k_6_50,k_6_51,k_6_52,k_6_53,k_6_54,k_6_55,k_6_56,k_6_57,k_6_58,k_6_59,k_6_60,k_6_61,k_6_62,k_6_63;
wire k_7_0,k_7_1,k_7_2,k_7_3,k_7_4,k_7_5,k_7_6,k_7_7,k_7_8,k_7_9,k_7_10,k_7_11,k_7_12,k_7_13,k_7_14,k_7_15,k_7_16,k_7_17,k_7_18,k_7_19,k_7_20,k_7_21,k_7_22,k_7_23,k_7_24,k_7_25,k_7_26,k_7_27,k_7_28,k_7_29,k_7_30,k_7_31,k_7_32,k_7_33,k_7_34,k_7_35,k_7_36,k_7_37,k_7_38,k_7_39,k_7_40,k_7_41,k_7_42,k_7_43,k_7_44,k_7_45,k_7_46,k_7_47,k_7_48,k_7_49,k_7_50,k_7_51,k_7_52,k_7_53,k_7_54,k_7_55,k_7_56,k_7_57,k_7_58,k_7_59,k_7_60,k_7_61,k_7_62,k_7_63,k_7_64,k_7_65,k_7_66,k_7_67,k_7_68,k_7_69,k_7_70,k_7_71,k_7_72,k_7_73,k_7_74,k_7_75,k_7_76,k_7_77,k_7_78,k_7_79,k_7_80,k_7_81,k_7_82,k_7_83,k_7_84,k_7_85,k_7_86,k_7_87,k_7_88,k_7_89,k_7_90,k_7_91,k_7_92,k_7_93,k_7_94,k_7_95,k_7_96,k_7_97,k_7_98,k_7_99,k_7_100,k_7_101,k_7_102,k_7_103,k_7_104,k_7_105,k_7_106,k_7_107,k_7_108,k_7_109,k_7_110,k_7_111,k_7_112,k_7_113,k_7_114,k_7_115,k_7_116,k_7_117,k_7_118,k_7_119,k_7_120,k_7_121,k_7_122,k_7_123,k_7_124,k_7_125,k_7_126,k_7_127;
wire k_8_0,k_8_1,k_8_2,k_8_3,k_8_4,k_8_5,k_8_6,k_8_7,k_8_8,k_8_9,k_8_10,k_8_11,k_8_12,k_8_13,k_8_14,k_8_15,k_8_16,k_8_17,k_8_18,k_8_19,k_8_20,k_8_21,k_8_22,k_8_23,k_8_24,k_8_25,k_8_26,k_8_27,k_8_28,k_8_29,k_8_30,k_8_31,k_8_32,k_8_33,k_8_34,k_8_35,k_8_36,k_8_37,k_8_38,k_8_39,k_8_40,k_8_41,k_8_42,k_8_43,k_8_44,k_8_45,k_8_46,k_8_47,k_8_48,k_8_49,k_8_50,k_8_51,k_8_52,k_8_53,k_8_54,k_8_55,k_8_56,k_8_57,k_8_58,k_8_59,k_8_60,k_8_61,k_8_62,k_8_63,k_8_64,k_8_65,k_8_66,k_8_67,k_8_68,k_8_69,k_8_70,k_8_71,k_8_72,k_8_73,k_8_74,k_8_75,k_8_76,k_8_77,k_8_78,k_8_79,k_8_80,k_8_81,k_8_82,k_8_83,k_8_84,k_8_85,k_8_86,k_8_87,k_8_88,k_8_89,k_8_90,k_8_91,k_8_92,k_8_93,k_8_94,k_8_95,k_8_96,k_8_97,k_8_98,k_8_99,k_8_100,k_8_101,k_8_102,k_8_103,k_8_104,k_8_105,k_8_106,k_8_107,k_8_108,k_8_109,k_8_110,k_8_111,k_8_112,k_8_113,k_8_114,k_8_115,k_8_116,k_8_117,k_8_118,k_8_119,k_8_120,k_8_121,k_8_122,k_8_123,k_8_124,k_8_125,k_8_126,k_8_127,k_8_128,k_8_129,k_8_130,k_8_131,k_8_132,k_8_133,k_8_134,k_8_135,k_8_136,k_8_137,k_8_138,k_8_139,k_8_140,k_8_141,k_8_142,k_8_143,k_8_144,k_8_145,k_8_146,k_8_147,k_8_148,k_8_149,k_8_150,k_8_151,k_8_152,k_8_153,k_8_154,k_8_155,k_8_156,k_8_157,k_8_158,k_8_159,k_8_160,k_8_161,k_8_162,k_8_163,k_8_164,k_8_165,k_8_166,k_8_167,k_8_168,k_8_169,k_8_170,k_8_171,k_8_172,k_8_173,k_8_174,k_8_175,k_8_176,k_8_177,k_8_178,k_8_179,k_8_180,k_8_181,k_8_182,k_8_183,k_8_184,k_8_185,k_8_186,k_8_187,k_8_188,k_8_189,k_8_190,k_8_191,k_8_192,k_8_193,k_8_194,k_8_195,k_8_196,k_8_197,k_8_198,k_8_199,k_8_200,k_8_201,k_8_202,k_8_203,k_8_204,k_8_205,k_8_206,k_8_207,k_8_208,k_8_209,k_8_210,k_8_211,k_8_212,k_8_213,k_8_214,k_8_215,k_8_216,k_8_217,k_8_218,k_8_219,k_8_220,k_8_221,k_8_222,k_8_223,k_8_224,k_8_225,k_8_226,k_8_227,k_8_228,k_8_229,k_8_230,k_8_231,k_8_232,k_8_233,k_8_234,k_8_235,k_8_236,k_8_237,k_8_238,k_8_239,k_8_240,k_8_241,k_8_242,k_8_243,k_8_244,k_8_245,k_8_246,k_8_247,k_8_248,k_8_249,k_8_250,k_8_251,k_8_252,k_8_253,k_8_254,k_8_255;
wire k_9_0,k_9_1,k_9_2,k_9_3,k_9_4,k_9_5,k_9_6,k_9_7,k_9_8,k_9_9,k_9_10,k_9_11,k_9_12,k_9_13,k_9_14,k_9_15,k_9_16,k_9_17,k_9_18,k_9_19,k_9_20,k_9_21,k_9_22,k_9_23,k_9_24,k_9_25,k_9_26,k_9_27,k_9_28,k_9_29,k_9_30,k_9_31,k_9_32,k_9_33,k_9_34,k_9_35,k_9_36,k_9_37,k_9_38,k_9_39,k_9_40,k_9_41,k_9_42,k_9_43,k_9_44,k_9_45,k_9_46,k_9_47,k_9_48,k_9_49,k_9_50,k_9_51,k_9_52,k_9_53,k_9_54,k_9_55,k_9_56,k_9_57,k_9_58,k_9_59,k_9_60,k_9_61,k_9_62,k_9_63,k_9_64,k_9_65,k_9_66,k_9_67,k_9_68,k_9_69,k_9_70,k_9_71,k_9_72,k_9_73,k_9_74,k_9_75,k_9_76,k_9_77,k_9_78,k_9_79,k_9_80,k_9_81,k_9_82,k_9_83,k_9_84,k_9_85,k_9_86,k_9_87,k_9_88,k_9_89,k_9_90,k_9_91,k_9_92,k_9_93,k_9_94,k_9_95,k_9_96,k_9_97,k_9_98,k_9_99,k_9_100,k_9_101,k_9_102,k_9_103,k_9_104,k_9_105,k_9_106,k_9_107,k_9_108,k_9_109,k_9_110,k_9_111,k_9_112,k_9_113,k_9_114,k_9_115,k_9_116,k_9_117,k_9_118,k_9_119,k_9_120,k_9_121,k_9_122,k_9_123,k_9_124,k_9_125,k_9_126,k_9_127,k_9_128,k_9_129,k_9_130,k_9_131,k_9_132,k_9_133,k_9_134,k_9_135,k_9_136,k_9_137,k_9_138,k_9_139,k_9_140,k_9_141,k_9_142,k_9_143,k_9_144,k_9_145,k_9_146,k_9_147,k_9_148,k_9_149,k_9_150,k_9_151,k_9_152,k_9_153,k_9_154,k_9_155,k_9_156,k_9_157,k_9_158,k_9_159,k_9_160,k_9_161,k_9_162,k_9_163,k_9_164,k_9_165,k_9_166,k_9_167,k_9_168,k_9_169,k_9_170,k_9_171,k_9_172,k_9_173,k_9_174,k_9_175,k_9_176,k_9_177,k_9_178,k_9_179,k_9_180,k_9_181,k_9_182,k_9_183,k_9_184,k_9_185,k_9_186,k_9_187,k_9_188,k_9_189,k_9_190,k_9_191,k_9_192,k_9_193,k_9_194,k_9_195,k_9_196,k_9_197,k_9_198,k_9_199,k_9_200,k_9_201,k_9_202,k_9_203,k_9_204,k_9_205,k_9_206,k_9_207,k_9_208,k_9_209,k_9_210,k_9_211,k_9_212,k_9_213,k_9_214,k_9_215,k_9_216,k_9_217,k_9_218,k_9_219,k_9_220,k_9_221,k_9_222,k_9_223,k_9_224,k_9_225,k_9_226,k_9_227,k_9_228,k_9_229,k_9_230,k_9_231,k_9_232,k_9_233,k_9_234,k_9_235,k_9_236,k_9_237,k_9_238,k_9_239,k_9_240,k_9_241,k_9_242,k_9_243,k_9_244,k_9_245,k_9_246,k_9_247,k_9_248,k_9_249,k_9_250,k_9_251,k_9_252,k_9_253,k_9_254,k_9_255,k_9_256,k_9_257,k_9_258,k_9_259,k_9_260,k_9_261,k_9_262,k_9_263,k_9_264,k_9_265,k_9_266,k_9_267,k_9_268,k_9_269,k_9_270,k_9_271,k_9_272,k_9_273,k_9_274,k_9_275,k_9_276,k_9_277,k_9_278,k_9_279,k_9_280,k_9_281,k_9_282,k_9_283,k_9_284,k_9_285,k_9_286,k_9_287,k_9_288,k_9_289,k_9_290,k_9_291,k_9_292,k_9_293,k_9_294,k_9_295,k_9_296,k_9_297,k_9_298,k_9_299,k_9_300,k_9_301,k_9_302,k_9_303,k_9_304,k_9_305,k_9_306,k_9_307,k_9_308,k_9_309,k_9_310,k_9_311,k_9_312,k_9_313,k_9_314,k_9_315,k_9_316,k_9_317,k_9_318,k_9_319,k_9_320,k_9_321,k_9_322,k_9_323,k_9_324,k_9_325,k_9_326,k_9_327,k_9_328,k_9_329,k_9_330,k_9_331,k_9_332,k_9_333,k_9_334,k_9_335,k_9_336,k_9_337,k_9_338,k_9_339,k_9_340,k_9_341,k_9_342,k_9_343,k_9_344,k_9_345,k_9_346,k_9_347,k_9_348,k_9_349,k_9_350,k_9_351,k_9_352,k_9_353,k_9_354,k_9_355,k_9_356,k_9_357,k_9_358,k_9_359,k_9_360,k_9_361,k_9_362,k_9_363,k_9_364,k_9_365,k_9_366,k_9_367,k_9_368,k_9_369,k_9_370,k_9_371,k_9_372,k_9_373,k_9_374,k_9_375,k_9_376,k_9_377,k_9_378,k_9_379,k_9_380,k_9_381,k_9_382,k_9_383,k_9_384,k_9_385,k_9_386,k_9_387,k_9_388,k_9_389,k_9_390,k_9_391,k_9_392,k_9_393,k_9_394,k_9_395,k_9_396,k_9_397,k_9_398,k_9_399,k_9_400,k_9_401,k_9_402,k_9_403,k_9_404,k_9_405,k_9_406,k_9_407,k_9_408,k_9_409,k_9_410,k_9_411,k_9_412,k_9_413,k_9_414,k_9_415,k_9_416,k_9_417,k_9_418,k_9_419,k_9_420,k_9_421,k_9_422,k_9_423,k_9_424,k_9_425,k_9_426,k_9_427,k_9_428,k_9_429,k_9_430,k_9_431,k_9_432,k_9_433,k_9_434,k_9_435,k_9_436,k_9_437,k_9_438,k_9_439,k_9_440,k_9_441,k_9_442,k_9_443,k_9_444,k_9_445,k_9_446,k_9_447,k_9_448,k_9_449,k_9_450,k_9_451,k_9_452,k_9_453,k_9_454,k_9_455,k_9_456,k_9_457,k_9_458,k_9_459,k_9_460,k_9_461,k_9_462,k_9_463,k_9_464,k_9_465,k_9_466,k_9_467,k_9_468,k_9_469,k_9_470,k_9_471,k_9_472,k_9_473,k_9_474,k_9_475,k_9_476,k_9_477,k_9_478,k_9_479,k_9_480,k_9_481,k_9_482,k_9_483,k_9_484,k_9_485,k_9_486,k_9_487,k_9_488,k_9_489,k_9_490,k_9_491,k_9_492,k_9_493,k_9_494,k_9_495,k_9_496,k_9_497,k_9_498,k_9_499,k_9_500,k_9_501,k_9_502,k_9_503,k_9_504,k_9_505,k_9_506,k_9_507,k_9_508,k_9_509,k_9_510,k_9_511;
valve v_1_0 (.fluid_in(k_1_0), .fluid_out(k_0_0), .air_in(c_1_0));
valve v_1_1 (.fluid_in(k_1_1), .fluid_out(k_0_0), .air_in(c_1_1));
valve v_2_0 (.fluid_in(k_2_0), .fluid_out(k_1_0), .air_in(c_2_0));
valve v_2_1 (.fluid_in(k_2_1), .fluid_out(k_1_0), .air_in(c_2_1));
valve v_2_2 (.fluid_in(k_2_2), .fluid_out(k_1_1), .air_in(c_2_0));
valve v_2_3 (.fluid_in(k_2_3), .fluid_out(k_1_1), .air_in(c_2_1));
valve v_3_0 (.fluid_in(k_3_0), .fluid_out(k_2_0), .air_in(c_3_0));
valve v_3_1 (.fluid_in(k_3_1), .fluid_out(k_2_0), .air_in(c_3_1));
valve v_3_2 (.fluid_in(k_3_2), .fluid_out(k_2_1), .air_in(c_3_0));
valve v_3_3 (.fluid_in(k_3_3), .fluid_out(k_2_1), .air_in(c_3_1));
valve v_3_4 (.fluid_in(k_3_4), .fluid_out(k_2_2), .air_in(c_3_0));
valve v_3_5 (.fluid_in(k_3_5), .fluid_out(k_2_2), .air_in(c_3_1));
valve v_3_6 (.fluid_in(k_3_6), .fluid_out(k_2_3), .air_in(c_3_0));
valve v_3_7 (.fluid_in(k_3_7), .fluid_out(k_2_3), .air_in(c_3_1));
valve v_4_0 (.fluid_in(k_4_0), .fluid_out(k_3_0), .air_in(c_4_0));
valve v_4_1 (.fluid_in(k_4_1), .fluid_out(k_3_0), .air_in(c_4_1));
valve v_4_2 (.fluid_in(k_4_2), .fluid_out(k_3_1), .air_in(c_4_0));
valve v_4_3 (.fluid_in(k_4_3), .fluid_out(k_3_1), .air_in(c_4_1));
valve v_4_4 (.fluid_in(k_4_4), .fluid_out(k_3_2), .air_in(c_4_0));
valve v_4_5 (.fluid_in(k_4_5), .fluid_out(k_3_2), .air_in(c_4_1));
valve v_4_6 (.fluid_in(k_4_6), .fluid_out(k_3_3), .air_in(c_4_0));
valve v_4_7 (.fluid_in(k_4_7), .fluid_out(k_3_3), .air_in(c_4_1));
valve v_4_8 (.fluid_in(k_4_8), .fluid_out(k_3_4), .air_in(c_4_0));
valve v_4_9 (.fluid_in(k_4_9), .fluid_out(k_3_4), .air_in(c_4_1));
valve v_4_10 (.fluid_in(k_4_10), .fluid_out(k_3_5), .air_in(c_4_0));
valve v_4_11 (.fluid_in(k_4_11), .fluid_out(k_3_5), .air_in(c_4_1));
valve v_4_12 (.fluid_in(k_4_12), .fluid_out(k_3_6), .air_in(c_4_0));
valve v_4_13 (.fluid_in(k_4_13), .fluid_out(k_3_6), .air_in(c_4_1));
valve v_4_14 (.fluid_in(k_4_14), .fluid_out(k_3_7), .air_in(c_4_0));
valve v_4_15 (.fluid_in(k_4_15), .fluid_out(k_3_7), .air_in(c_4_1));
valve v_5_0 (.fluid_in(k_5_0), .fluid_out(k_4_0), .air_in(c_5_0));
valve v_5_1 (.fluid_in(k_5_1), .fluid_out(k_4_0), .air_in(c_5_1));
valve v_5_2 (.fluid_in(k_5_2), .fluid_out(k_4_1), .air_in(c_5_0));
valve v_5_3 (.fluid_in(k_5_3), .fluid_out(k_4_1), .air_in(c_5_1));
valve v_5_4 (.fluid_in(k_5_4), .fluid_out(k_4_2), .air_in(c_5_0));
valve v_5_5 (.fluid_in(k_5_5), .fluid_out(k_4_2), .air_in(c_5_1));
valve v_5_6 (.fluid_in(k_5_6), .fluid_out(k_4_3), .air_in(c_5_0));
valve v_5_7 (.fluid_in(k_5_7), .fluid_out(k_4_3), .air_in(c_5_1));
valve v_5_8 (.fluid_in(k_5_8), .fluid_out(k_4_4), .air_in(c_5_0));
valve v_5_9 (.fluid_in(k_5_9), .fluid_out(k_4_4), .air_in(c_5_1));
valve v_5_10 (.fluid_in(k_5_10), .fluid_out(k_4_5), .air_in(c_5_0));
valve v_5_11 (.fluid_in(k_5_11), .fluid_out(k_4_5), .air_in(c_5_1));
valve v_5_12 (.fluid_in(k_5_12), .fluid_out(k_4_6), .air_in(c_5_0));
valve v_5_13 (.fluid_in(k_5_13), .fluid_out(k_4_6), .air_in(c_5_1));
valve v_5_14 (.fluid_in(k_5_14), .fluid_out(k_4_7), .air_in(c_5_0));
valve v_5_15 (.fluid_in(k_5_15), .fluid_out(k_4_7), .air_in(c_5_1));
valve v_5_16 (.fluid_in(k_5_16), .fluid_out(k_4_8), .air_in(c_5_0));
valve v_5_17 (.fluid_in(k_5_17), .fluid_out(k_4_8), .air_in(c_5_1));
valve v_5_18 (.fluid_in(k_5_18), .fluid_out(k_4_9), .air_in(c_5_0));
valve v_5_19 (.fluid_in(k_5_19), .fluid_out(k_4_9), .air_in(c_5_1));
valve v_5_20 (.fluid_in(k_5_20), .fluid_out(k_4_10), .air_in(c_5_0));
valve v_5_21 (.fluid_in(k_5_21), .fluid_out(k_4_10), .air_in(c_5_1));
valve v_5_22 (.fluid_in(k_5_22), .fluid_out(k_4_11), .air_in(c_5_0));
valve v_5_23 (.fluid_in(k_5_23), .fluid_out(k_4_11), .air_in(c_5_1));
valve v_5_24 (.fluid_in(k_5_24), .fluid_out(k_4_12), .air_in(c_5_0));
valve v_5_25 (.fluid_in(k_5_25), .fluid_out(k_4_12), .air_in(c_5_1));
valve v_5_26 (.fluid_in(k_5_26), .fluid_out(k_4_13), .air_in(c_5_0));
valve v_5_27 (.fluid_in(k_5_27), .fluid_out(k_4_13), .air_in(c_5_1));
valve v_5_28 (.fluid_in(k_5_28), .fluid_out(k_4_14), .air_in(c_5_0));
valve v_5_29 (.fluid_in(k_5_29), .fluid_out(k_4_14), .air_in(c_5_1));
valve v_5_30 (.fluid_in(k_5_30), .fluid_out(k_4_15), .air_in(c_5_0));
valve v_5_31 (.fluid_in(k_5_31), .fluid_out(k_4_15), .air_in(c_5_1));
valve v_6_0 (.fluid_in(k_6_0), .fluid_out(k_5_0), .air_in(c_6_0));
valve v_6_1 (.fluid_in(k_6_1), .fluid_out(k_5_0), .air_in(c_6_1));
valve v_6_2 (.fluid_in(k_6_2), .fluid_out(k_5_1), .air_in(c_6_0));
valve v_6_3 (.fluid_in(k_6_3), .fluid_out(k_5_1), .air_in(c_6_1));
valve v_6_4 (.fluid_in(k_6_4), .fluid_out(k_5_2), .air_in(c_6_0));
valve v_6_5 (.fluid_in(k_6_5), .fluid_out(k_5_2), .air_in(c_6_1));
valve v_6_6 (.fluid_in(k_6_6), .fluid_out(k_5_3), .air_in(c_6_0));
valve v_6_7 (.fluid_in(k_6_7), .fluid_out(k_5_3), .air_in(c_6_1));
valve v_6_8 (.fluid_in(k_6_8), .fluid_out(k_5_4), .air_in(c_6_0));
valve v_6_9 (.fluid_in(k_6_9), .fluid_out(k_5_4), .air_in(c_6_1));
valve v_6_10 (.fluid_in(k_6_10), .fluid_out(k_5_5), .air_in(c_6_0));
valve v_6_11 (.fluid_in(k_6_11), .fluid_out(k_5_5), .air_in(c_6_1));
valve v_6_12 (.fluid_in(k_6_12), .fluid_out(k_5_6), .air_in(c_6_0));
valve v_6_13 (.fluid_in(k_6_13), .fluid_out(k_5_6), .air_in(c_6_1));
valve v_6_14 (.fluid_in(k_6_14), .fluid_out(k_5_7), .air_in(c_6_0));
valve v_6_15 (.fluid_in(k_6_15), .fluid_out(k_5_7), .air_in(c_6_1));
valve v_6_16 (.fluid_in(k_6_16), .fluid_out(k_5_8), .air_in(c_6_0));
valve v_6_17 (.fluid_in(k_6_17), .fluid_out(k_5_8), .air_in(c_6_1));
valve v_6_18 (.fluid_in(k_6_18), .fluid_out(k_5_9), .air_in(c_6_0));
valve v_6_19 (.fluid_in(k_6_19), .fluid_out(k_5_9), .air_in(c_6_1));
valve v_6_20 (.fluid_in(k_6_20), .fluid_out(k_5_10), .air_in(c_6_0));
valve v_6_21 (.fluid_in(k_6_21), .fluid_out(k_5_10), .air_in(c_6_1));
valve v_6_22 (.fluid_in(k_6_22), .fluid_out(k_5_11), .air_in(c_6_0));
valve v_6_23 (.fluid_in(k_6_23), .fluid_out(k_5_11), .air_in(c_6_1));
valve v_6_24 (.fluid_in(k_6_24), .fluid_out(k_5_12), .air_in(c_6_0));
valve v_6_25 (.fluid_in(k_6_25), .fluid_out(k_5_12), .air_in(c_6_1));
valve v_6_26 (.fluid_in(k_6_26), .fluid_out(k_5_13), .air_in(c_6_0));
valve v_6_27 (.fluid_in(k_6_27), .fluid_out(k_5_13), .air_in(c_6_1));
valve v_6_28 (.fluid_in(k_6_28), .fluid_out(k_5_14), .air_in(c_6_0));
valve v_6_29 (.fluid_in(k_6_29), .fluid_out(k_5_14), .air_in(c_6_1));
valve v_6_30 (.fluid_in(k_6_30), .fluid_out(k_5_15), .air_in(c_6_0));
valve v_6_31 (.fluid_in(k_6_31), .fluid_out(k_5_15), .air_in(c_6_1));
valve v_6_32 (.fluid_in(k_6_32), .fluid_out(k_5_16), .air_in(c_6_0));
valve v_6_33 (.fluid_in(k_6_33), .fluid_out(k_5_16), .air_in(c_6_1));
valve v_6_34 (.fluid_in(k_6_34), .fluid_out(k_5_17), .air_in(c_6_0));
valve v_6_35 (.fluid_in(k_6_35), .fluid_out(k_5_17), .air_in(c_6_1));
valve v_6_36 (.fluid_in(k_6_36), .fluid_out(k_5_18), .air_in(c_6_0));
valve v_6_37 (.fluid_in(k_6_37), .fluid_out(k_5_18), .air_in(c_6_1));
valve v_6_38 (.fluid_in(k_6_38), .fluid_out(k_5_19), .air_in(c_6_0));
valve v_6_39 (.fluid_in(k_6_39), .fluid_out(k_5_19), .air_in(c_6_1));
valve v_6_40 (.fluid_in(k_6_40), .fluid_out(k_5_20), .air_in(c_6_0));
valve v_6_41 (.fluid_in(k_6_41), .fluid_out(k_5_20), .air_in(c_6_1));
valve v_6_42 (.fluid_in(k_6_42), .fluid_out(k_5_21), .air_in(c_6_0));
valve v_6_43 (.fluid_in(k_6_43), .fluid_out(k_5_21), .air_in(c_6_1));
valve v_6_44 (.fluid_in(k_6_44), .fluid_out(k_5_22), .air_in(c_6_0));
valve v_6_45 (.fluid_in(k_6_45), .fluid_out(k_5_22), .air_in(c_6_1));
valve v_6_46 (.fluid_in(k_6_46), .fluid_out(k_5_23), .air_in(c_6_0));
valve v_6_47 (.fluid_in(k_6_47), .fluid_out(k_5_23), .air_in(c_6_1));
valve v_6_48 (.fluid_in(k_6_48), .fluid_out(k_5_24), .air_in(c_6_0));
valve v_6_49 (.fluid_in(k_6_49), .fluid_out(k_5_24), .air_in(c_6_1));
valve v_6_50 (.fluid_in(k_6_50), .fluid_out(k_5_25), .air_in(c_6_0));
valve v_6_51 (.fluid_in(k_6_51), .fluid_out(k_5_25), .air_in(c_6_1));
valve v_6_52 (.fluid_in(k_6_52), .fluid_out(k_5_26), .air_in(c_6_0));
valve v_6_53 (.fluid_in(k_6_53), .fluid_out(k_5_26), .air_in(c_6_1));
valve v_6_54 (.fluid_in(k_6_54), .fluid_out(k_5_27), .air_in(c_6_0));
valve v_6_55 (.fluid_in(k_6_55), .fluid_out(k_5_27), .air_in(c_6_1));
valve v_6_56 (.fluid_in(k_6_56), .fluid_out(k_5_28), .air_in(c_6_0));
valve v_6_57 (.fluid_in(k_6_57), .fluid_out(k_5_28), .air_in(c_6_1));
valve v_6_58 (.fluid_in(k_6_58), .fluid_out(k_5_29), .air_in(c_6_0));
valve v_6_59 (.fluid_in(k_6_59), .fluid_out(k_5_29), .air_in(c_6_1));
valve v_6_60 (.fluid_in(k_6_60), .fluid_out(k_5_30), .air_in(c_6_0));
valve v_6_61 (.fluid_in(k_6_61), .fluid_out(k_5_30), .air_in(c_6_1));
valve v_6_62 (.fluid_in(k_6_62), .fluid_out(k_5_31), .air_in(c_6_0));
valve v_6_63 (.fluid_in(k_6_63), .fluid_out(k_5_31), .air_in(c_6_1));
valve v_7_0 (.fluid_in(k_7_0), .fluid_out(k_6_0), .air_in(c_7_0));
valve v_7_1 (.fluid_in(k_7_1), .fluid_out(k_6_0), .air_in(c_7_1));
valve v_7_2 (.fluid_in(k_7_2), .fluid_out(k_6_1), .air_in(c_7_0));
valve v_7_3 (.fluid_in(k_7_3), .fluid_out(k_6_1), .air_in(c_7_1));
valve v_7_4 (.fluid_in(k_7_4), .fluid_out(k_6_2), .air_in(c_7_0));
valve v_7_5 (.fluid_in(k_7_5), .fluid_out(k_6_2), .air_in(c_7_1));
valve v_7_6 (.fluid_in(k_7_6), .fluid_out(k_6_3), .air_in(c_7_0));
valve v_7_7 (.fluid_in(k_7_7), .fluid_out(k_6_3), .air_in(c_7_1));
valve v_7_8 (.fluid_in(k_7_8), .fluid_out(k_6_4), .air_in(c_7_0));
valve v_7_9 (.fluid_in(k_7_9), .fluid_out(k_6_4), .air_in(c_7_1));
valve v_7_10 (.fluid_in(k_7_10), .fluid_out(k_6_5), .air_in(c_7_0));
valve v_7_11 (.fluid_in(k_7_11), .fluid_out(k_6_5), .air_in(c_7_1));
valve v_7_12 (.fluid_in(k_7_12), .fluid_out(k_6_6), .air_in(c_7_0));
valve v_7_13 (.fluid_in(k_7_13), .fluid_out(k_6_6), .air_in(c_7_1));
valve v_7_14 (.fluid_in(k_7_14), .fluid_out(k_6_7), .air_in(c_7_0));
valve v_7_15 (.fluid_in(k_7_15), .fluid_out(k_6_7), .air_in(c_7_1));
valve v_7_16 (.fluid_in(k_7_16), .fluid_out(k_6_8), .air_in(c_7_0));
valve v_7_17 (.fluid_in(k_7_17), .fluid_out(k_6_8), .air_in(c_7_1));
valve v_7_18 (.fluid_in(k_7_18), .fluid_out(k_6_9), .air_in(c_7_0));
valve v_7_19 (.fluid_in(k_7_19), .fluid_out(k_6_9), .air_in(c_7_1));
valve v_7_20 (.fluid_in(k_7_20), .fluid_out(k_6_10), .air_in(c_7_0));
valve v_7_21 (.fluid_in(k_7_21), .fluid_out(k_6_10), .air_in(c_7_1));
valve v_7_22 (.fluid_in(k_7_22), .fluid_out(k_6_11), .air_in(c_7_0));
valve v_7_23 (.fluid_in(k_7_23), .fluid_out(k_6_11), .air_in(c_7_1));
valve v_7_24 (.fluid_in(k_7_24), .fluid_out(k_6_12), .air_in(c_7_0));
valve v_7_25 (.fluid_in(k_7_25), .fluid_out(k_6_12), .air_in(c_7_1));
valve v_7_26 (.fluid_in(k_7_26), .fluid_out(k_6_13), .air_in(c_7_0));
valve v_7_27 (.fluid_in(k_7_27), .fluid_out(k_6_13), .air_in(c_7_1));
valve v_7_28 (.fluid_in(k_7_28), .fluid_out(k_6_14), .air_in(c_7_0));
valve v_7_29 (.fluid_in(k_7_29), .fluid_out(k_6_14), .air_in(c_7_1));
valve v_7_30 (.fluid_in(k_7_30), .fluid_out(k_6_15), .air_in(c_7_0));
valve v_7_31 (.fluid_in(k_7_31), .fluid_out(k_6_15), .air_in(c_7_1));
valve v_7_32 (.fluid_in(k_7_32), .fluid_out(k_6_16), .air_in(c_7_0));
valve v_7_33 (.fluid_in(k_7_33), .fluid_out(k_6_16), .air_in(c_7_1));
valve v_7_34 (.fluid_in(k_7_34), .fluid_out(k_6_17), .air_in(c_7_0));
valve v_7_35 (.fluid_in(k_7_35), .fluid_out(k_6_17), .air_in(c_7_1));
valve v_7_36 (.fluid_in(k_7_36), .fluid_out(k_6_18), .air_in(c_7_0));
valve v_7_37 (.fluid_in(k_7_37), .fluid_out(k_6_18), .air_in(c_7_1));
valve v_7_38 (.fluid_in(k_7_38), .fluid_out(k_6_19), .air_in(c_7_0));
valve v_7_39 (.fluid_in(k_7_39), .fluid_out(k_6_19), .air_in(c_7_1));
valve v_7_40 (.fluid_in(k_7_40), .fluid_out(k_6_20), .air_in(c_7_0));
valve v_7_41 (.fluid_in(k_7_41), .fluid_out(k_6_20), .air_in(c_7_1));
valve v_7_42 (.fluid_in(k_7_42), .fluid_out(k_6_21), .air_in(c_7_0));
valve v_7_43 (.fluid_in(k_7_43), .fluid_out(k_6_21), .air_in(c_7_1));
valve v_7_44 (.fluid_in(k_7_44), .fluid_out(k_6_22), .air_in(c_7_0));
valve v_7_45 (.fluid_in(k_7_45), .fluid_out(k_6_22), .air_in(c_7_1));
valve v_7_46 (.fluid_in(k_7_46), .fluid_out(k_6_23), .air_in(c_7_0));
valve v_7_47 (.fluid_in(k_7_47), .fluid_out(k_6_23), .air_in(c_7_1));
valve v_7_48 (.fluid_in(k_7_48), .fluid_out(k_6_24), .air_in(c_7_0));
valve v_7_49 (.fluid_in(k_7_49), .fluid_out(k_6_24), .air_in(c_7_1));
valve v_7_50 (.fluid_in(k_7_50), .fluid_out(k_6_25), .air_in(c_7_0));
valve v_7_51 (.fluid_in(k_7_51), .fluid_out(k_6_25), .air_in(c_7_1));
valve v_7_52 (.fluid_in(k_7_52), .fluid_out(k_6_26), .air_in(c_7_0));
valve v_7_53 (.fluid_in(k_7_53), .fluid_out(k_6_26), .air_in(c_7_1));
valve v_7_54 (.fluid_in(k_7_54), .fluid_out(k_6_27), .air_in(c_7_0));
valve v_7_55 (.fluid_in(k_7_55), .fluid_out(k_6_27), .air_in(c_7_1));
valve v_7_56 (.fluid_in(k_7_56), .fluid_out(k_6_28), .air_in(c_7_0));
valve v_7_57 (.fluid_in(k_7_57), .fluid_out(k_6_28), .air_in(c_7_1));
valve v_7_58 (.fluid_in(k_7_58), .fluid_out(k_6_29), .air_in(c_7_0));
valve v_7_59 (.fluid_in(k_7_59), .fluid_out(k_6_29), .air_in(c_7_1));
valve v_7_60 (.fluid_in(k_7_60), .fluid_out(k_6_30), .air_in(c_7_0));
valve v_7_61 (.fluid_in(k_7_61), .fluid_out(k_6_30), .air_in(c_7_1));
valve v_7_62 (.fluid_in(k_7_62), .fluid_out(k_6_31), .air_in(c_7_0));
valve v_7_63 (.fluid_in(k_7_63), .fluid_out(k_6_31), .air_in(c_7_1));
valve v_7_64 (.fluid_in(k_7_64), .fluid_out(k_6_32), .air_in(c_7_0));
valve v_7_65 (.fluid_in(k_7_65), .fluid_out(k_6_32), .air_in(c_7_1));
valve v_7_66 (.fluid_in(k_7_66), .fluid_out(k_6_33), .air_in(c_7_0));
valve v_7_67 (.fluid_in(k_7_67), .fluid_out(k_6_33), .air_in(c_7_1));
valve v_7_68 (.fluid_in(k_7_68), .fluid_out(k_6_34), .air_in(c_7_0));
valve v_7_69 (.fluid_in(k_7_69), .fluid_out(k_6_34), .air_in(c_7_1));
valve v_7_70 (.fluid_in(k_7_70), .fluid_out(k_6_35), .air_in(c_7_0));
valve v_7_71 (.fluid_in(k_7_71), .fluid_out(k_6_35), .air_in(c_7_1));
valve v_7_72 (.fluid_in(k_7_72), .fluid_out(k_6_36), .air_in(c_7_0));
valve v_7_73 (.fluid_in(k_7_73), .fluid_out(k_6_36), .air_in(c_7_1));
valve v_7_74 (.fluid_in(k_7_74), .fluid_out(k_6_37), .air_in(c_7_0));
valve v_7_75 (.fluid_in(k_7_75), .fluid_out(k_6_37), .air_in(c_7_1));
valve v_7_76 (.fluid_in(k_7_76), .fluid_out(k_6_38), .air_in(c_7_0));
valve v_7_77 (.fluid_in(k_7_77), .fluid_out(k_6_38), .air_in(c_7_1));
valve v_7_78 (.fluid_in(k_7_78), .fluid_out(k_6_39), .air_in(c_7_0));
valve v_7_79 (.fluid_in(k_7_79), .fluid_out(k_6_39), .air_in(c_7_1));
valve v_7_80 (.fluid_in(k_7_80), .fluid_out(k_6_40), .air_in(c_7_0));
valve v_7_81 (.fluid_in(k_7_81), .fluid_out(k_6_40), .air_in(c_7_1));
valve v_7_82 (.fluid_in(k_7_82), .fluid_out(k_6_41), .air_in(c_7_0));
valve v_7_83 (.fluid_in(k_7_83), .fluid_out(k_6_41), .air_in(c_7_1));
valve v_7_84 (.fluid_in(k_7_84), .fluid_out(k_6_42), .air_in(c_7_0));
valve v_7_85 (.fluid_in(k_7_85), .fluid_out(k_6_42), .air_in(c_7_1));
valve v_7_86 (.fluid_in(k_7_86), .fluid_out(k_6_43), .air_in(c_7_0));
valve v_7_87 (.fluid_in(k_7_87), .fluid_out(k_6_43), .air_in(c_7_1));
valve v_7_88 (.fluid_in(k_7_88), .fluid_out(k_6_44), .air_in(c_7_0));
valve v_7_89 (.fluid_in(k_7_89), .fluid_out(k_6_44), .air_in(c_7_1));
valve v_7_90 (.fluid_in(k_7_90), .fluid_out(k_6_45), .air_in(c_7_0));
valve v_7_91 (.fluid_in(k_7_91), .fluid_out(k_6_45), .air_in(c_7_1));
valve v_7_92 (.fluid_in(k_7_92), .fluid_out(k_6_46), .air_in(c_7_0));
valve v_7_93 (.fluid_in(k_7_93), .fluid_out(k_6_46), .air_in(c_7_1));
valve v_7_94 (.fluid_in(k_7_94), .fluid_out(k_6_47), .air_in(c_7_0));
valve v_7_95 (.fluid_in(k_7_95), .fluid_out(k_6_47), .air_in(c_7_1));
valve v_7_96 (.fluid_in(k_7_96), .fluid_out(k_6_48), .air_in(c_7_0));
valve v_7_97 (.fluid_in(k_7_97), .fluid_out(k_6_48), .air_in(c_7_1));
valve v_7_98 (.fluid_in(k_7_98), .fluid_out(k_6_49), .air_in(c_7_0));
valve v_7_99 (.fluid_in(k_7_99), .fluid_out(k_6_49), .air_in(c_7_1));
valve v_7_100 (.fluid_in(k_7_100), .fluid_out(k_6_50), .air_in(c_7_0));
valve v_7_101 (.fluid_in(k_7_101), .fluid_out(k_6_50), .air_in(c_7_1));
valve v_7_102 (.fluid_in(k_7_102), .fluid_out(k_6_51), .air_in(c_7_0));
valve v_7_103 (.fluid_in(k_7_103), .fluid_out(k_6_51), .air_in(c_7_1));
valve v_7_104 (.fluid_in(k_7_104), .fluid_out(k_6_52), .air_in(c_7_0));
valve v_7_105 (.fluid_in(k_7_105), .fluid_out(k_6_52), .air_in(c_7_1));
valve v_7_106 (.fluid_in(k_7_106), .fluid_out(k_6_53), .air_in(c_7_0));
valve v_7_107 (.fluid_in(k_7_107), .fluid_out(k_6_53), .air_in(c_7_1));
valve v_7_108 (.fluid_in(k_7_108), .fluid_out(k_6_54), .air_in(c_7_0));
valve v_7_109 (.fluid_in(k_7_109), .fluid_out(k_6_54), .air_in(c_7_1));
valve v_7_110 (.fluid_in(k_7_110), .fluid_out(k_6_55), .air_in(c_7_0));
valve v_7_111 (.fluid_in(k_7_111), .fluid_out(k_6_55), .air_in(c_7_1));
valve v_7_112 (.fluid_in(k_7_112), .fluid_out(k_6_56), .air_in(c_7_0));
valve v_7_113 (.fluid_in(k_7_113), .fluid_out(k_6_56), .air_in(c_7_1));
valve v_7_114 (.fluid_in(k_7_114), .fluid_out(k_6_57), .air_in(c_7_0));
valve v_7_115 (.fluid_in(k_7_115), .fluid_out(k_6_57), .air_in(c_7_1));
valve v_7_116 (.fluid_in(k_7_116), .fluid_out(k_6_58), .air_in(c_7_0));
valve v_7_117 (.fluid_in(k_7_117), .fluid_out(k_6_58), .air_in(c_7_1));
valve v_7_118 (.fluid_in(k_7_118), .fluid_out(k_6_59), .air_in(c_7_0));
valve v_7_119 (.fluid_in(k_7_119), .fluid_out(k_6_59), .air_in(c_7_1));
valve v_7_120 (.fluid_in(k_7_120), .fluid_out(k_6_60), .air_in(c_7_0));
valve v_7_121 (.fluid_in(k_7_121), .fluid_out(k_6_60), .air_in(c_7_1));
valve v_7_122 (.fluid_in(k_7_122), .fluid_out(k_6_61), .air_in(c_7_0));
valve v_7_123 (.fluid_in(k_7_123), .fluid_out(k_6_61), .air_in(c_7_1));
valve v_7_124 (.fluid_in(k_7_124), .fluid_out(k_6_62), .air_in(c_7_0));
valve v_7_125 (.fluid_in(k_7_125), .fluid_out(k_6_62), .air_in(c_7_1));
valve v_7_126 (.fluid_in(k_7_126), .fluid_out(k_6_63), .air_in(c_7_0));
valve v_7_127 (.fluid_in(k_7_127), .fluid_out(k_6_63), .air_in(c_7_1));
valve v_8_0 (.fluid_in(k_8_0), .fluid_out(k_7_0), .air_in(c_8_0));
valve v_8_1 (.fluid_in(k_8_1), .fluid_out(k_7_0), .air_in(c_8_1));
valve v_8_2 (.fluid_in(k_8_2), .fluid_out(k_7_1), .air_in(c_8_0));
valve v_8_3 (.fluid_in(k_8_3), .fluid_out(k_7_1), .air_in(c_8_1));
valve v_8_4 (.fluid_in(k_8_4), .fluid_out(k_7_2), .air_in(c_8_0));
valve v_8_5 (.fluid_in(k_8_5), .fluid_out(k_7_2), .air_in(c_8_1));
valve v_8_6 (.fluid_in(k_8_6), .fluid_out(k_7_3), .air_in(c_8_0));
valve v_8_7 (.fluid_in(k_8_7), .fluid_out(k_7_3), .air_in(c_8_1));
valve v_8_8 (.fluid_in(k_8_8), .fluid_out(k_7_4), .air_in(c_8_0));
valve v_8_9 (.fluid_in(k_8_9), .fluid_out(k_7_4), .air_in(c_8_1));
valve v_8_10 (.fluid_in(k_8_10), .fluid_out(k_7_5), .air_in(c_8_0));
valve v_8_11 (.fluid_in(k_8_11), .fluid_out(k_7_5), .air_in(c_8_1));
valve v_8_12 (.fluid_in(k_8_12), .fluid_out(k_7_6), .air_in(c_8_0));
valve v_8_13 (.fluid_in(k_8_13), .fluid_out(k_7_6), .air_in(c_8_1));
valve v_8_14 (.fluid_in(k_8_14), .fluid_out(k_7_7), .air_in(c_8_0));
valve v_8_15 (.fluid_in(k_8_15), .fluid_out(k_7_7), .air_in(c_8_1));
valve v_8_16 (.fluid_in(k_8_16), .fluid_out(k_7_8), .air_in(c_8_0));
valve v_8_17 (.fluid_in(k_8_17), .fluid_out(k_7_8), .air_in(c_8_1));
valve v_8_18 (.fluid_in(k_8_18), .fluid_out(k_7_9), .air_in(c_8_0));
valve v_8_19 (.fluid_in(k_8_19), .fluid_out(k_7_9), .air_in(c_8_1));
valve v_8_20 (.fluid_in(k_8_20), .fluid_out(k_7_10), .air_in(c_8_0));
valve v_8_21 (.fluid_in(k_8_21), .fluid_out(k_7_10), .air_in(c_8_1));
valve v_8_22 (.fluid_in(k_8_22), .fluid_out(k_7_11), .air_in(c_8_0));
valve v_8_23 (.fluid_in(k_8_23), .fluid_out(k_7_11), .air_in(c_8_1));
valve v_8_24 (.fluid_in(k_8_24), .fluid_out(k_7_12), .air_in(c_8_0));
valve v_8_25 (.fluid_in(k_8_25), .fluid_out(k_7_12), .air_in(c_8_1));
valve v_8_26 (.fluid_in(k_8_26), .fluid_out(k_7_13), .air_in(c_8_0));
valve v_8_27 (.fluid_in(k_8_27), .fluid_out(k_7_13), .air_in(c_8_1));
valve v_8_28 (.fluid_in(k_8_28), .fluid_out(k_7_14), .air_in(c_8_0));
valve v_8_29 (.fluid_in(k_8_29), .fluid_out(k_7_14), .air_in(c_8_1));
valve v_8_30 (.fluid_in(k_8_30), .fluid_out(k_7_15), .air_in(c_8_0));
valve v_8_31 (.fluid_in(k_8_31), .fluid_out(k_7_15), .air_in(c_8_1));
valve v_8_32 (.fluid_in(k_8_32), .fluid_out(k_7_16), .air_in(c_8_0));
valve v_8_33 (.fluid_in(k_8_33), .fluid_out(k_7_16), .air_in(c_8_1));
valve v_8_34 (.fluid_in(k_8_34), .fluid_out(k_7_17), .air_in(c_8_0));
valve v_8_35 (.fluid_in(k_8_35), .fluid_out(k_7_17), .air_in(c_8_1));
valve v_8_36 (.fluid_in(k_8_36), .fluid_out(k_7_18), .air_in(c_8_0));
valve v_8_37 (.fluid_in(k_8_37), .fluid_out(k_7_18), .air_in(c_8_1));
valve v_8_38 (.fluid_in(k_8_38), .fluid_out(k_7_19), .air_in(c_8_0));
valve v_8_39 (.fluid_in(k_8_39), .fluid_out(k_7_19), .air_in(c_8_1));
valve v_8_40 (.fluid_in(k_8_40), .fluid_out(k_7_20), .air_in(c_8_0));
valve v_8_41 (.fluid_in(k_8_41), .fluid_out(k_7_20), .air_in(c_8_1));
valve v_8_42 (.fluid_in(k_8_42), .fluid_out(k_7_21), .air_in(c_8_0));
valve v_8_43 (.fluid_in(k_8_43), .fluid_out(k_7_21), .air_in(c_8_1));
valve v_8_44 (.fluid_in(k_8_44), .fluid_out(k_7_22), .air_in(c_8_0));
valve v_8_45 (.fluid_in(k_8_45), .fluid_out(k_7_22), .air_in(c_8_1));
valve v_8_46 (.fluid_in(k_8_46), .fluid_out(k_7_23), .air_in(c_8_0));
valve v_8_47 (.fluid_in(k_8_47), .fluid_out(k_7_23), .air_in(c_8_1));
valve v_8_48 (.fluid_in(k_8_48), .fluid_out(k_7_24), .air_in(c_8_0));
valve v_8_49 (.fluid_in(k_8_49), .fluid_out(k_7_24), .air_in(c_8_1));
valve v_8_50 (.fluid_in(k_8_50), .fluid_out(k_7_25), .air_in(c_8_0));
valve v_8_51 (.fluid_in(k_8_51), .fluid_out(k_7_25), .air_in(c_8_1));
valve v_8_52 (.fluid_in(k_8_52), .fluid_out(k_7_26), .air_in(c_8_0));
valve v_8_53 (.fluid_in(k_8_53), .fluid_out(k_7_26), .air_in(c_8_1));
valve v_8_54 (.fluid_in(k_8_54), .fluid_out(k_7_27), .air_in(c_8_0));
valve v_8_55 (.fluid_in(k_8_55), .fluid_out(k_7_27), .air_in(c_8_1));
valve v_8_56 (.fluid_in(k_8_56), .fluid_out(k_7_28), .air_in(c_8_0));
valve v_8_57 (.fluid_in(k_8_57), .fluid_out(k_7_28), .air_in(c_8_1));
valve v_8_58 (.fluid_in(k_8_58), .fluid_out(k_7_29), .air_in(c_8_0));
valve v_8_59 (.fluid_in(k_8_59), .fluid_out(k_7_29), .air_in(c_8_1));
valve v_8_60 (.fluid_in(k_8_60), .fluid_out(k_7_30), .air_in(c_8_0));
valve v_8_61 (.fluid_in(k_8_61), .fluid_out(k_7_30), .air_in(c_8_1));
valve v_8_62 (.fluid_in(k_8_62), .fluid_out(k_7_31), .air_in(c_8_0));
valve v_8_63 (.fluid_in(k_8_63), .fluid_out(k_7_31), .air_in(c_8_1));
valve v_8_64 (.fluid_in(k_8_64), .fluid_out(k_7_32), .air_in(c_8_0));
valve v_8_65 (.fluid_in(k_8_65), .fluid_out(k_7_32), .air_in(c_8_1));
valve v_8_66 (.fluid_in(k_8_66), .fluid_out(k_7_33), .air_in(c_8_0));
valve v_8_67 (.fluid_in(k_8_67), .fluid_out(k_7_33), .air_in(c_8_1));
valve v_8_68 (.fluid_in(k_8_68), .fluid_out(k_7_34), .air_in(c_8_0));
valve v_8_69 (.fluid_in(k_8_69), .fluid_out(k_7_34), .air_in(c_8_1));
valve v_8_70 (.fluid_in(k_8_70), .fluid_out(k_7_35), .air_in(c_8_0));
valve v_8_71 (.fluid_in(k_8_71), .fluid_out(k_7_35), .air_in(c_8_1));
valve v_8_72 (.fluid_in(k_8_72), .fluid_out(k_7_36), .air_in(c_8_0));
valve v_8_73 (.fluid_in(k_8_73), .fluid_out(k_7_36), .air_in(c_8_1));
valve v_8_74 (.fluid_in(k_8_74), .fluid_out(k_7_37), .air_in(c_8_0));
valve v_8_75 (.fluid_in(k_8_75), .fluid_out(k_7_37), .air_in(c_8_1));
valve v_8_76 (.fluid_in(k_8_76), .fluid_out(k_7_38), .air_in(c_8_0));
valve v_8_77 (.fluid_in(k_8_77), .fluid_out(k_7_38), .air_in(c_8_1));
valve v_8_78 (.fluid_in(k_8_78), .fluid_out(k_7_39), .air_in(c_8_0));
valve v_8_79 (.fluid_in(k_8_79), .fluid_out(k_7_39), .air_in(c_8_1));
valve v_8_80 (.fluid_in(k_8_80), .fluid_out(k_7_40), .air_in(c_8_0));
valve v_8_81 (.fluid_in(k_8_81), .fluid_out(k_7_40), .air_in(c_8_1));
valve v_8_82 (.fluid_in(k_8_82), .fluid_out(k_7_41), .air_in(c_8_0));
valve v_8_83 (.fluid_in(k_8_83), .fluid_out(k_7_41), .air_in(c_8_1));
valve v_8_84 (.fluid_in(k_8_84), .fluid_out(k_7_42), .air_in(c_8_0));
valve v_8_85 (.fluid_in(k_8_85), .fluid_out(k_7_42), .air_in(c_8_1));
valve v_8_86 (.fluid_in(k_8_86), .fluid_out(k_7_43), .air_in(c_8_0));
valve v_8_87 (.fluid_in(k_8_87), .fluid_out(k_7_43), .air_in(c_8_1));
valve v_8_88 (.fluid_in(k_8_88), .fluid_out(k_7_44), .air_in(c_8_0));
valve v_8_89 (.fluid_in(k_8_89), .fluid_out(k_7_44), .air_in(c_8_1));
valve v_8_90 (.fluid_in(k_8_90), .fluid_out(k_7_45), .air_in(c_8_0));
valve v_8_91 (.fluid_in(k_8_91), .fluid_out(k_7_45), .air_in(c_8_1));
valve v_8_92 (.fluid_in(k_8_92), .fluid_out(k_7_46), .air_in(c_8_0));
valve v_8_93 (.fluid_in(k_8_93), .fluid_out(k_7_46), .air_in(c_8_1));
valve v_8_94 (.fluid_in(k_8_94), .fluid_out(k_7_47), .air_in(c_8_0));
valve v_8_95 (.fluid_in(k_8_95), .fluid_out(k_7_47), .air_in(c_8_1));
valve v_8_96 (.fluid_in(k_8_96), .fluid_out(k_7_48), .air_in(c_8_0));
valve v_8_97 (.fluid_in(k_8_97), .fluid_out(k_7_48), .air_in(c_8_1));
valve v_8_98 (.fluid_in(k_8_98), .fluid_out(k_7_49), .air_in(c_8_0));
valve v_8_99 (.fluid_in(k_8_99), .fluid_out(k_7_49), .air_in(c_8_1));
valve v_8_100 (.fluid_in(k_8_100), .fluid_out(k_7_50), .air_in(c_8_0));
valve v_8_101 (.fluid_in(k_8_101), .fluid_out(k_7_50), .air_in(c_8_1));
valve v_8_102 (.fluid_in(k_8_102), .fluid_out(k_7_51), .air_in(c_8_0));
valve v_8_103 (.fluid_in(k_8_103), .fluid_out(k_7_51), .air_in(c_8_1));
valve v_8_104 (.fluid_in(k_8_104), .fluid_out(k_7_52), .air_in(c_8_0));
valve v_8_105 (.fluid_in(k_8_105), .fluid_out(k_7_52), .air_in(c_8_1));
valve v_8_106 (.fluid_in(k_8_106), .fluid_out(k_7_53), .air_in(c_8_0));
valve v_8_107 (.fluid_in(k_8_107), .fluid_out(k_7_53), .air_in(c_8_1));
valve v_8_108 (.fluid_in(k_8_108), .fluid_out(k_7_54), .air_in(c_8_0));
valve v_8_109 (.fluid_in(k_8_109), .fluid_out(k_7_54), .air_in(c_8_1));
valve v_8_110 (.fluid_in(k_8_110), .fluid_out(k_7_55), .air_in(c_8_0));
valve v_8_111 (.fluid_in(k_8_111), .fluid_out(k_7_55), .air_in(c_8_1));
valve v_8_112 (.fluid_in(k_8_112), .fluid_out(k_7_56), .air_in(c_8_0));
valve v_8_113 (.fluid_in(k_8_113), .fluid_out(k_7_56), .air_in(c_8_1));
valve v_8_114 (.fluid_in(k_8_114), .fluid_out(k_7_57), .air_in(c_8_0));
valve v_8_115 (.fluid_in(k_8_115), .fluid_out(k_7_57), .air_in(c_8_1));
valve v_8_116 (.fluid_in(k_8_116), .fluid_out(k_7_58), .air_in(c_8_0));
valve v_8_117 (.fluid_in(k_8_117), .fluid_out(k_7_58), .air_in(c_8_1));
valve v_8_118 (.fluid_in(k_8_118), .fluid_out(k_7_59), .air_in(c_8_0));
valve v_8_119 (.fluid_in(k_8_119), .fluid_out(k_7_59), .air_in(c_8_1));
valve v_8_120 (.fluid_in(k_8_120), .fluid_out(k_7_60), .air_in(c_8_0));
valve v_8_121 (.fluid_in(k_8_121), .fluid_out(k_7_60), .air_in(c_8_1));
valve v_8_122 (.fluid_in(k_8_122), .fluid_out(k_7_61), .air_in(c_8_0));
valve v_8_123 (.fluid_in(k_8_123), .fluid_out(k_7_61), .air_in(c_8_1));
valve v_8_124 (.fluid_in(k_8_124), .fluid_out(k_7_62), .air_in(c_8_0));
valve v_8_125 (.fluid_in(k_8_125), .fluid_out(k_7_62), .air_in(c_8_1));
valve v_8_126 (.fluid_in(k_8_126), .fluid_out(k_7_63), .air_in(c_8_0));
valve v_8_127 (.fluid_in(k_8_127), .fluid_out(k_7_63), .air_in(c_8_1));
valve v_8_128 (.fluid_in(k_8_128), .fluid_out(k_7_64), .air_in(c_8_0));
valve v_8_129 (.fluid_in(k_8_129), .fluid_out(k_7_64), .air_in(c_8_1));
valve v_8_130 (.fluid_in(k_8_130), .fluid_out(k_7_65), .air_in(c_8_0));
valve v_8_131 (.fluid_in(k_8_131), .fluid_out(k_7_65), .air_in(c_8_1));
valve v_8_132 (.fluid_in(k_8_132), .fluid_out(k_7_66), .air_in(c_8_0));
valve v_8_133 (.fluid_in(k_8_133), .fluid_out(k_7_66), .air_in(c_8_1));
valve v_8_134 (.fluid_in(k_8_134), .fluid_out(k_7_67), .air_in(c_8_0));
valve v_8_135 (.fluid_in(k_8_135), .fluid_out(k_7_67), .air_in(c_8_1));
valve v_8_136 (.fluid_in(k_8_136), .fluid_out(k_7_68), .air_in(c_8_0));
valve v_8_137 (.fluid_in(k_8_137), .fluid_out(k_7_68), .air_in(c_8_1));
valve v_8_138 (.fluid_in(k_8_138), .fluid_out(k_7_69), .air_in(c_8_0));
valve v_8_139 (.fluid_in(k_8_139), .fluid_out(k_7_69), .air_in(c_8_1));
valve v_8_140 (.fluid_in(k_8_140), .fluid_out(k_7_70), .air_in(c_8_0));
valve v_8_141 (.fluid_in(k_8_141), .fluid_out(k_7_70), .air_in(c_8_1));
valve v_8_142 (.fluid_in(k_8_142), .fluid_out(k_7_71), .air_in(c_8_0));
valve v_8_143 (.fluid_in(k_8_143), .fluid_out(k_7_71), .air_in(c_8_1));
valve v_8_144 (.fluid_in(k_8_144), .fluid_out(k_7_72), .air_in(c_8_0));
valve v_8_145 (.fluid_in(k_8_145), .fluid_out(k_7_72), .air_in(c_8_1));
valve v_8_146 (.fluid_in(k_8_146), .fluid_out(k_7_73), .air_in(c_8_0));
valve v_8_147 (.fluid_in(k_8_147), .fluid_out(k_7_73), .air_in(c_8_1));
valve v_8_148 (.fluid_in(k_8_148), .fluid_out(k_7_74), .air_in(c_8_0));
valve v_8_149 (.fluid_in(k_8_149), .fluid_out(k_7_74), .air_in(c_8_1));
valve v_8_150 (.fluid_in(k_8_150), .fluid_out(k_7_75), .air_in(c_8_0));
valve v_8_151 (.fluid_in(k_8_151), .fluid_out(k_7_75), .air_in(c_8_1));
valve v_8_152 (.fluid_in(k_8_152), .fluid_out(k_7_76), .air_in(c_8_0));
valve v_8_153 (.fluid_in(k_8_153), .fluid_out(k_7_76), .air_in(c_8_1));
valve v_8_154 (.fluid_in(k_8_154), .fluid_out(k_7_77), .air_in(c_8_0));
valve v_8_155 (.fluid_in(k_8_155), .fluid_out(k_7_77), .air_in(c_8_1));
valve v_8_156 (.fluid_in(k_8_156), .fluid_out(k_7_78), .air_in(c_8_0));
valve v_8_157 (.fluid_in(k_8_157), .fluid_out(k_7_78), .air_in(c_8_1));
valve v_8_158 (.fluid_in(k_8_158), .fluid_out(k_7_79), .air_in(c_8_0));
valve v_8_159 (.fluid_in(k_8_159), .fluid_out(k_7_79), .air_in(c_8_1));
valve v_8_160 (.fluid_in(k_8_160), .fluid_out(k_7_80), .air_in(c_8_0));
valve v_8_161 (.fluid_in(k_8_161), .fluid_out(k_7_80), .air_in(c_8_1));
valve v_8_162 (.fluid_in(k_8_162), .fluid_out(k_7_81), .air_in(c_8_0));
valve v_8_163 (.fluid_in(k_8_163), .fluid_out(k_7_81), .air_in(c_8_1));
valve v_8_164 (.fluid_in(k_8_164), .fluid_out(k_7_82), .air_in(c_8_0));
valve v_8_165 (.fluid_in(k_8_165), .fluid_out(k_7_82), .air_in(c_8_1));
valve v_8_166 (.fluid_in(k_8_166), .fluid_out(k_7_83), .air_in(c_8_0));
valve v_8_167 (.fluid_in(k_8_167), .fluid_out(k_7_83), .air_in(c_8_1));
valve v_8_168 (.fluid_in(k_8_168), .fluid_out(k_7_84), .air_in(c_8_0));
valve v_8_169 (.fluid_in(k_8_169), .fluid_out(k_7_84), .air_in(c_8_1));
valve v_8_170 (.fluid_in(k_8_170), .fluid_out(k_7_85), .air_in(c_8_0));
valve v_8_171 (.fluid_in(k_8_171), .fluid_out(k_7_85), .air_in(c_8_1));
valve v_8_172 (.fluid_in(k_8_172), .fluid_out(k_7_86), .air_in(c_8_0));
valve v_8_173 (.fluid_in(k_8_173), .fluid_out(k_7_86), .air_in(c_8_1));
valve v_8_174 (.fluid_in(k_8_174), .fluid_out(k_7_87), .air_in(c_8_0));
valve v_8_175 (.fluid_in(k_8_175), .fluid_out(k_7_87), .air_in(c_8_1));
valve v_8_176 (.fluid_in(k_8_176), .fluid_out(k_7_88), .air_in(c_8_0));
valve v_8_177 (.fluid_in(k_8_177), .fluid_out(k_7_88), .air_in(c_8_1));
valve v_8_178 (.fluid_in(k_8_178), .fluid_out(k_7_89), .air_in(c_8_0));
valve v_8_179 (.fluid_in(k_8_179), .fluid_out(k_7_89), .air_in(c_8_1));
valve v_8_180 (.fluid_in(k_8_180), .fluid_out(k_7_90), .air_in(c_8_0));
valve v_8_181 (.fluid_in(k_8_181), .fluid_out(k_7_90), .air_in(c_8_1));
valve v_8_182 (.fluid_in(k_8_182), .fluid_out(k_7_91), .air_in(c_8_0));
valve v_8_183 (.fluid_in(k_8_183), .fluid_out(k_7_91), .air_in(c_8_1));
valve v_8_184 (.fluid_in(k_8_184), .fluid_out(k_7_92), .air_in(c_8_0));
valve v_8_185 (.fluid_in(k_8_185), .fluid_out(k_7_92), .air_in(c_8_1));
valve v_8_186 (.fluid_in(k_8_186), .fluid_out(k_7_93), .air_in(c_8_0));
valve v_8_187 (.fluid_in(k_8_187), .fluid_out(k_7_93), .air_in(c_8_1));
valve v_8_188 (.fluid_in(k_8_188), .fluid_out(k_7_94), .air_in(c_8_0));
valve v_8_189 (.fluid_in(k_8_189), .fluid_out(k_7_94), .air_in(c_8_1));
valve v_8_190 (.fluid_in(k_8_190), .fluid_out(k_7_95), .air_in(c_8_0));
valve v_8_191 (.fluid_in(k_8_191), .fluid_out(k_7_95), .air_in(c_8_1));
valve v_8_192 (.fluid_in(k_8_192), .fluid_out(k_7_96), .air_in(c_8_0));
valve v_8_193 (.fluid_in(k_8_193), .fluid_out(k_7_96), .air_in(c_8_1));
valve v_8_194 (.fluid_in(k_8_194), .fluid_out(k_7_97), .air_in(c_8_0));
valve v_8_195 (.fluid_in(k_8_195), .fluid_out(k_7_97), .air_in(c_8_1));
valve v_8_196 (.fluid_in(k_8_196), .fluid_out(k_7_98), .air_in(c_8_0));
valve v_8_197 (.fluid_in(k_8_197), .fluid_out(k_7_98), .air_in(c_8_1));
valve v_8_198 (.fluid_in(k_8_198), .fluid_out(k_7_99), .air_in(c_8_0));
valve v_8_199 (.fluid_in(k_8_199), .fluid_out(k_7_99), .air_in(c_8_1));
valve v_8_200 (.fluid_in(k_8_200), .fluid_out(k_7_100), .air_in(c_8_0));
valve v_8_201 (.fluid_in(k_8_201), .fluid_out(k_7_100), .air_in(c_8_1));
valve v_8_202 (.fluid_in(k_8_202), .fluid_out(k_7_101), .air_in(c_8_0));
valve v_8_203 (.fluid_in(k_8_203), .fluid_out(k_7_101), .air_in(c_8_1));
valve v_8_204 (.fluid_in(k_8_204), .fluid_out(k_7_102), .air_in(c_8_0));
valve v_8_205 (.fluid_in(k_8_205), .fluid_out(k_7_102), .air_in(c_8_1));
valve v_8_206 (.fluid_in(k_8_206), .fluid_out(k_7_103), .air_in(c_8_0));
valve v_8_207 (.fluid_in(k_8_207), .fluid_out(k_7_103), .air_in(c_8_1));
valve v_8_208 (.fluid_in(k_8_208), .fluid_out(k_7_104), .air_in(c_8_0));
valve v_8_209 (.fluid_in(k_8_209), .fluid_out(k_7_104), .air_in(c_8_1));
valve v_8_210 (.fluid_in(k_8_210), .fluid_out(k_7_105), .air_in(c_8_0));
valve v_8_211 (.fluid_in(k_8_211), .fluid_out(k_7_105), .air_in(c_8_1));
valve v_8_212 (.fluid_in(k_8_212), .fluid_out(k_7_106), .air_in(c_8_0));
valve v_8_213 (.fluid_in(k_8_213), .fluid_out(k_7_106), .air_in(c_8_1));
valve v_8_214 (.fluid_in(k_8_214), .fluid_out(k_7_107), .air_in(c_8_0));
valve v_8_215 (.fluid_in(k_8_215), .fluid_out(k_7_107), .air_in(c_8_1));
valve v_8_216 (.fluid_in(k_8_216), .fluid_out(k_7_108), .air_in(c_8_0));
valve v_8_217 (.fluid_in(k_8_217), .fluid_out(k_7_108), .air_in(c_8_1));
valve v_8_218 (.fluid_in(k_8_218), .fluid_out(k_7_109), .air_in(c_8_0));
valve v_8_219 (.fluid_in(k_8_219), .fluid_out(k_7_109), .air_in(c_8_1));
valve v_8_220 (.fluid_in(k_8_220), .fluid_out(k_7_110), .air_in(c_8_0));
valve v_8_221 (.fluid_in(k_8_221), .fluid_out(k_7_110), .air_in(c_8_1));
valve v_8_222 (.fluid_in(k_8_222), .fluid_out(k_7_111), .air_in(c_8_0));
valve v_8_223 (.fluid_in(k_8_223), .fluid_out(k_7_111), .air_in(c_8_1));
valve v_8_224 (.fluid_in(k_8_224), .fluid_out(k_7_112), .air_in(c_8_0));
valve v_8_225 (.fluid_in(k_8_225), .fluid_out(k_7_112), .air_in(c_8_1));
valve v_8_226 (.fluid_in(k_8_226), .fluid_out(k_7_113), .air_in(c_8_0));
valve v_8_227 (.fluid_in(k_8_227), .fluid_out(k_7_113), .air_in(c_8_1));
valve v_8_228 (.fluid_in(k_8_228), .fluid_out(k_7_114), .air_in(c_8_0));
valve v_8_229 (.fluid_in(k_8_229), .fluid_out(k_7_114), .air_in(c_8_1));
valve v_8_230 (.fluid_in(k_8_230), .fluid_out(k_7_115), .air_in(c_8_0));
valve v_8_231 (.fluid_in(k_8_231), .fluid_out(k_7_115), .air_in(c_8_1));
valve v_8_232 (.fluid_in(k_8_232), .fluid_out(k_7_116), .air_in(c_8_0));
valve v_8_233 (.fluid_in(k_8_233), .fluid_out(k_7_116), .air_in(c_8_1));
valve v_8_234 (.fluid_in(k_8_234), .fluid_out(k_7_117), .air_in(c_8_0));
valve v_8_235 (.fluid_in(k_8_235), .fluid_out(k_7_117), .air_in(c_8_1));
valve v_8_236 (.fluid_in(k_8_236), .fluid_out(k_7_118), .air_in(c_8_0));
valve v_8_237 (.fluid_in(k_8_237), .fluid_out(k_7_118), .air_in(c_8_1));
valve v_8_238 (.fluid_in(k_8_238), .fluid_out(k_7_119), .air_in(c_8_0));
valve v_8_239 (.fluid_in(k_8_239), .fluid_out(k_7_119), .air_in(c_8_1));
valve v_8_240 (.fluid_in(k_8_240), .fluid_out(k_7_120), .air_in(c_8_0));
valve v_8_241 (.fluid_in(k_8_241), .fluid_out(k_7_120), .air_in(c_8_1));
valve v_8_242 (.fluid_in(k_8_242), .fluid_out(k_7_121), .air_in(c_8_0));
valve v_8_243 (.fluid_in(k_8_243), .fluid_out(k_7_121), .air_in(c_8_1));
valve v_8_244 (.fluid_in(k_8_244), .fluid_out(k_7_122), .air_in(c_8_0));
valve v_8_245 (.fluid_in(k_8_245), .fluid_out(k_7_122), .air_in(c_8_1));
valve v_8_246 (.fluid_in(k_8_246), .fluid_out(k_7_123), .air_in(c_8_0));
valve v_8_247 (.fluid_in(k_8_247), .fluid_out(k_7_123), .air_in(c_8_1));
valve v_8_248 (.fluid_in(k_8_248), .fluid_out(k_7_124), .air_in(c_8_0));
valve v_8_249 (.fluid_in(k_8_249), .fluid_out(k_7_124), .air_in(c_8_1));
valve v_8_250 (.fluid_in(k_8_250), .fluid_out(k_7_125), .air_in(c_8_0));
valve v_8_251 (.fluid_in(k_8_251), .fluid_out(k_7_125), .air_in(c_8_1));
valve v_8_252 (.fluid_in(k_8_252), .fluid_out(k_7_126), .air_in(c_8_0));
valve v_8_253 (.fluid_in(k_8_253), .fluid_out(k_7_126), .air_in(c_8_1));
valve v_8_254 (.fluid_in(k_8_254), .fluid_out(k_7_127), .air_in(c_8_0));
valve v_8_255 (.fluid_in(k_8_255), .fluid_out(k_7_127), .air_in(c_8_1));
valve v_9_0 (.fluid_in(k_9_0), .fluid_out(k_8_0), .air_in(c_9_0));
valve v_9_1 (.fluid_in(k_9_1), .fluid_out(k_8_0), .air_in(c_9_1));
valve v_9_2 (.fluid_in(k_9_2), .fluid_out(k_8_1), .air_in(c_9_0));
valve v_9_3 (.fluid_in(k_9_3), .fluid_out(k_8_1), .air_in(c_9_1));
valve v_9_4 (.fluid_in(k_9_4), .fluid_out(k_8_2), .air_in(c_9_0));
valve v_9_5 (.fluid_in(k_9_5), .fluid_out(k_8_2), .air_in(c_9_1));
valve v_9_6 (.fluid_in(k_9_6), .fluid_out(k_8_3), .air_in(c_9_0));
valve v_9_7 (.fluid_in(k_9_7), .fluid_out(k_8_3), .air_in(c_9_1));
valve v_9_8 (.fluid_in(k_9_8), .fluid_out(k_8_4), .air_in(c_9_0));
valve v_9_9 (.fluid_in(k_9_9), .fluid_out(k_8_4), .air_in(c_9_1));
valve v_9_10 (.fluid_in(k_9_10), .fluid_out(k_8_5), .air_in(c_9_0));
valve v_9_11 (.fluid_in(k_9_11), .fluid_out(k_8_5), .air_in(c_9_1));
valve v_9_12 (.fluid_in(k_9_12), .fluid_out(k_8_6), .air_in(c_9_0));
valve v_9_13 (.fluid_in(k_9_13), .fluid_out(k_8_6), .air_in(c_9_1));
valve v_9_14 (.fluid_in(k_9_14), .fluid_out(k_8_7), .air_in(c_9_0));
valve v_9_15 (.fluid_in(k_9_15), .fluid_out(k_8_7), .air_in(c_9_1));
valve v_9_16 (.fluid_in(k_9_16), .fluid_out(k_8_8), .air_in(c_9_0));
valve v_9_17 (.fluid_in(k_9_17), .fluid_out(k_8_8), .air_in(c_9_1));
valve v_9_18 (.fluid_in(k_9_18), .fluid_out(k_8_9), .air_in(c_9_0));
valve v_9_19 (.fluid_in(k_9_19), .fluid_out(k_8_9), .air_in(c_9_1));
valve v_9_20 (.fluid_in(k_9_20), .fluid_out(k_8_10), .air_in(c_9_0));
valve v_9_21 (.fluid_in(k_9_21), .fluid_out(k_8_10), .air_in(c_9_1));
valve v_9_22 (.fluid_in(k_9_22), .fluid_out(k_8_11), .air_in(c_9_0));
valve v_9_23 (.fluid_in(k_9_23), .fluid_out(k_8_11), .air_in(c_9_1));
valve v_9_24 (.fluid_in(k_9_24), .fluid_out(k_8_12), .air_in(c_9_0));
valve v_9_25 (.fluid_in(k_9_25), .fluid_out(k_8_12), .air_in(c_9_1));
valve v_9_26 (.fluid_in(k_9_26), .fluid_out(k_8_13), .air_in(c_9_0));
valve v_9_27 (.fluid_in(k_9_27), .fluid_out(k_8_13), .air_in(c_9_1));
valve v_9_28 (.fluid_in(k_9_28), .fluid_out(k_8_14), .air_in(c_9_0));
valve v_9_29 (.fluid_in(k_9_29), .fluid_out(k_8_14), .air_in(c_9_1));
valve v_9_30 (.fluid_in(k_9_30), .fluid_out(k_8_15), .air_in(c_9_0));
valve v_9_31 (.fluid_in(k_9_31), .fluid_out(k_8_15), .air_in(c_9_1));
valve v_9_32 (.fluid_in(k_9_32), .fluid_out(k_8_16), .air_in(c_9_0));
valve v_9_33 (.fluid_in(k_9_33), .fluid_out(k_8_16), .air_in(c_9_1));
valve v_9_34 (.fluid_in(k_9_34), .fluid_out(k_8_17), .air_in(c_9_0));
valve v_9_35 (.fluid_in(k_9_35), .fluid_out(k_8_17), .air_in(c_9_1));
valve v_9_36 (.fluid_in(k_9_36), .fluid_out(k_8_18), .air_in(c_9_0));
valve v_9_37 (.fluid_in(k_9_37), .fluid_out(k_8_18), .air_in(c_9_1));
valve v_9_38 (.fluid_in(k_9_38), .fluid_out(k_8_19), .air_in(c_9_0));
valve v_9_39 (.fluid_in(k_9_39), .fluid_out(k_8_19), .air_in(c_9_1));
valve v_9_40 (.fluid_in(k_9_40), .fluid_out(k_8_20), .air_in(c_9_0));
valve v_9_41 (.fluid_in(k_9_41), .fluid_out(k_8_20), .air_in(c_9_1));
valve v_9_42 (.fluid_in(k_9_42), .fluid_out(k_8_21), .air_in(c_9_0));
valve v_9_43 (.fluid_in(k_9_43), .fluid_out(k_8_21), .air_in(c_9_1));
valve v_9_44 (.fluid_in(k_9_44), .fluid_out(k_8_22), .air_in(c_9_0));
valve v_9_45 (.fluid_in(k_9_45), .fluid_out(k_8_22), .air_in(c_9_1));
valve v_9_46 (.fluid_in(k_9_46), .fluid_out(k_8_23), .air_in(c_9_0));
valve v_9_47 (.fluid_in(k_9_47), .fluid_out(k_8_23), .air_in(c_9_1));
valve v_9_48 (.fluid_in(k_9_48), .fluid_out(k_8_24), .air_in(c_9_0));
valve v_9_49 (.fluid_in(k_9_49), .fluid_out(k_8_24), .air_in(c_9_1));
valve v_9_50 (.fluid_in(k_9_50), .fluid_out(k_8_25), .air_in(c_9_0));
valve v_9_51 (.fluid_in(k_9_51), .fluid_out(k_8_25), .air_in(c_9_1));
valve v_9_52 (.fluid_in(k_9_52), .fluid_out(k_8_26), .air_in(c_9_0));
valve v_9_53 (.fluid_in(k_9_53), .fluid_out(k_8_26), .air_in(c_9_1));
valve v_9_54 (.fluid_in(k_9_54), .fluid_out(k_8_27), .air_in(c_9_0));
valve v_9_55 (.fluid_in(k_9_55), .fluid_out(k_8_27), .air_in(c_9_1));
valve v_9_56 (.fluid_in(k_9_56), .fluid_out(k_8_28), .air_in(c_9_0));
valve v_9_57 (.fluid_in(k_9_57), .fluid_out(k_8_28), .air_in(c_9_1));
valve v_9_58 (.fluid_in(k_9_58), .fluid_out(k_8_29), .air_in(c_9_0));
valve v_9_59 (.fluid_in(k_9_59), .fluid_out(k_8_29), .air_in(c_9_1));
valve v_9_60 (.fluid_in(k_9_60), .fluid_out(k_8_30), .air_in(c_9_0));
valve v_9_61 (.fluid_in(k_9_61), .fluid_out(k_8_30), .air_in(c_9_1));
valve v_9_62 (.fluid_in(k_9_62), .fluid_out(k_8_31), .air_in(c_9_0));
valve v_9_63 (.fluid_in(k_9_63), .fluid_out(k_8_31), .air_in(c_9_1));
valve v_9_64 (.fluid_in(k_9_64), .fluid_out(k_8_32), .air_in(c_9_0));
valve v_9_65 (.fluid_in(k_9_65), .fluid_out(k_8_32), .air_in(c_9_1));
valve v_9_66 (.fluid_in(k_9_66), .fluid_out(k_8_33), .air_in(c_9_0));
valve v_9_67 (.fluid_in(k_9_67), .fluid_out(k_8_33), .air_in(c_9_1));
valve v_9_68 (.fluid_in(k_9_68), .fluid_out(k_8_34), .air_in(c_9_0));
valve v_9_69 (.fluid_in(k_9_69), .fluid_out(k_8_34), .air_in(c_9_1));
valve v_9_70 (.fluid_in(k_9_70), .fluid_out(k_8_35), .air_in(c_9_0));
valve v_9_71 (.fluid_in(k_9_71), .fluid_out(k_8_35), .air_in(c_9_1));
valve v_9_72 (.fluid_in(k_9_72), .fluid_out(k_8_36), .air_in(c_9_0));
valve v_9_73 (.fluid_in(k_9_73), .fluid_out(k_8_36), .air_in(c_9_1));
valve v_9_74 (.fluid_in(k_9_74), .fluid_out(k_8_37), .air_in(c_9_0));
valve v_9_75 (.fluid_in(k_9_75), .fluid_out(k_8_37), .air_in(c_9_1));
valve v_9_76 (.fluid_in(k_9_76), .fluid_out(k_8_38), .air_in(c_9_0));
valve v_9_77 (.fluid_in(k_9_77), .fluid_out(k_8_38), .air_in(c_9_1));
valve v_9_78 (.fluid_in(k_9_78), .fluid_out(k_8_39), .air_in(c_9_0));
valve v_9_79 (.fluid_in(k_9_79), .fluid_out(k_8_39), .air_in(c_9_1));
valve v_9_80 (.fluid_in(k_9_80), .fluid_out(k_8_40), .air_in(c_9_0));
valve v_9_81 (.fluid_in(k_9_81), .fluid_out(k_8_40), .air_in(c_9_1));
valve v_9_82 (.fluid_in(k_9_82), .fluid_out(k_8_41), .air_in(c_9_0));
valve v_9_83 (.fluid_in(k_9_83), .fluid_out(k_8_41), .air_in(c_9_1));
valve v_9_84 (.fluid_in(k_9_84), .fluid_out(k_8_42), .air_in(c_9_0));
valve v_9_85 (.fluid_in(k_9_85), .fluid_out(k_8_42), .air_in(c_9_1));
valve v_9_86 (.fluid_in(k_9_86), .fluid_out(k_8_43), .air_in(c_9_0));
valve v_9_87 (.fluid_in(k_9_87), .fluid_out(k_8_43), .air_in(c_9_1));
valve v_9_88 (.fluid_in(k_9_88), .fluid_out(k_8_44), .air_in(c_9_0));
valve v_9_89 (.fluid_in(k_9_89), .fluid_out(k_8_44), .air_in(c_9_1));
valve v_9_90 (.fluid_in(k_9_90), .fluid_out(k_8_45), .air_in(c_9_0));
valve v_9_91 (.fluid_in(k_9_91), .fluid_out(k_8_45), .air_in(c_9_1));
valve v_9_92 (.fluid_in(k_9_92), .fluid_out(k_8_46), .air_in(c_9_0));
valve v_9_93 (.fluid_in(k_9_93), .fluid_out(k_8_46), .air_in(c_9_1));
valve v_9_94 (.fluid_in(k_9_94), .fluid_out(k_8_47), .air_in(c_9_0));
valve v_9_95 (.fluid_in(k_9_95), .fluid_out(k_8_47), .air_in(c_9_1));
valve v_9_96 (.fluid_in(k_9_96), .fluid_out(k_8_48), .air_in(c_9_0));
valve v_9_97 (.fluid_in(k_9_97), .fluid_out(k_8_48), .air_in(c_9_1));
valve v_9_98 (.fluid_in(k_9_98), .fluid_out(k_8_49), .air_in(c_9_0));
valve v_9_99 (.fluid_in(k_9_99), .fluid_out(k_8_49), .air_in(c_9_1));
valve v_9_100 (.fluid_in(k_9_100), .fluid_out(k_8_50), .air_in(c_9_0));
valve v_9_101 (.fluid_in(k_9_101), .fluid_out(k_8_50), .air_in(c_9_1));
valve v_9_102 (.fluid_in(k_9_102), .fluid_out(k_8_51), .air_in(c_9_0));
valve v_9_103 (.fluid_in(k_9_103), .fluid_out(k_8_51), .air_in(c_9_1));
valve v_9_104 (.fluid_in(k_9_104), .fluid_out(k_8_52), .air_in(c_9_0));
valve v_9_105 (.fluid_in(k_9_105), .fluid_out(k_8_52), .air_in(c_9_1));
valve v_9_106 (.fluid_in(k_9_106), .fluid_out(k_8_53), .air_in(c_9_0));
valve v_9_107 (.fluid_in(k_9_107), .fluid_out(k_8_53), .air_in(c_9_1));
valve v_9_108 (.fluid_in(k_9_108), .fluid_out(k_8_54), .air_in(c_9_0));
valve v_9_109 (.fluid_in(k_9_109), .fluid_out(k_8_54), .air_in(c_9_1));
valve v_9_110 (.fluid_in(k_9_110), .fluid_out(k_8_55), .air_in(c_9_0));
valve v_9_111 (.fluid_in(k_9_111), .fluid_out(k_8_55), .air_in(c_9_1));
valve v_9_112 (.fluid_in(k_9_112), .fluid_out(k_8_56), .air_in(c_9_0));
valve v_9_113 (.fluid_in(k_9_113), .fluid_out(k_8_56), .air_in(c_9_1));
valve v_9_114 (.fluid_in(k_9_114), .fluid_out(k_8_57), .air_in(c_9_0));
valve v_9_115 (.fluid_in(k_9_115), .fluid_out(k_8_57), .air_in(c_9_1));
valve v_9_116 (.fluid_in(k_9_116), .fluid_out(k_8_58), .air_in(c_9_0));
valve v_9_117 (.fluid_in(k_9_117), .fluid_out(k_8_58), .air_in(c_9_1));
valve v_9_118 (.fluid_in(k_9_118), .fluid_out(k_8_59), .air_in(c_9_0));
valve v_9_119 (.fluid_in(k_9_119), .fluid_out(k_8_59), .air_in(c_9_1));
valve v_9_120 (.fluid_in(k_9_120), .fluid_out(k_8_60), .air_in(c_9_0));
valve v_9_121 (.fluid_in(k_9_121), .fluid_out(k_8_60), .air_in(c_9_1));
valve v_9_122 (.fluid_in(k_9_122), .fluid_out(k_8_61), .air_in(c_9_0));
valve v_9_123 (.fluid_in(k_9_123), .fluid_out(k_8_61), .air_in(c_9_1));
valve v_9_124 (.fluid_in(k_9_124), .fluid_out(k_8_62), .air_in(c_9_0));
valve v_9_125 (.fluid_in(k_9_125), .fluid_out(k_8_62), .air_in(c_9_1));
valve v_9_126 (.fluid_in(k_9_126), .fluid_out(k_8_63), .air_in(c_9_0));
valve v_9_127 (.fluid_in(k_9_127), .fluid_out(k_8_63), .air_in(c_9_1));
valve v_9_128 (.fluid_in(k_9_128), .fluid_out(k_8_64), .air_in(c_9_0));
valve v_9_129 (.fluid_in(k_9_129), .fluid_out(k_8_64), .air_in(c_9_1));
valve v_9_130 (.fluid_in(k_9_130), .fluid_out(k_8_65), .air_in(c_9_0));
valve v_9_131 (.fluid_in(k_9_131), .fluid_out(k_8_65), .air_in(c_9_1));
valve v_9_132 (.fluid_in(k_9_132), .fluid_out(k_8_66), .air_in(c_9_0));
valve v_9_133 (.fluid_in(k_9_133), .fluid_out(k_8_66), .air_in(c_9_1));
valve v_9_134 (.fluid_in(k_9_134), .fluid_out(k_8_67), .air_in(c_9_0));
valve v_9_135 (.fluid_in(k_9_135), .fluid_out(k_8_67), .air_in(c_9_1));
valve v_9_136 (.fluid_in(k_9_136), .fluid_out(k_8_68), .air_in(c_9_0));
valve v_9_137 (.fluid_in(k_9_137), .fluid_out(k_8_68), .air_in(c_9_1));
valve v_9_138 (.fluid_in(k_9_138), .fluid_out(k_8_69), .air_in(c_9_0));
valve v_9_139 (.fluid_in(k_9_139), .fluid_out(k_8_69), .air_in(c_9_1));
valve v_9_140 (.fluid_in(k_9_140), .fluid_out(k_8_70), .air_in(c_9_0));
valve v_9_141 (.fluid_in(k_9_141), .fluid_out(k_8_70), .air_in(c_9_1));
valve v_9_142 (.fluid_in(k_9_142), .fluid_out(k_8_71), .air_in(c_9_0));
valve v_9_143 (.fluid_in(k_9_143), .fluid_out(k_8_71), .air_in(c_9_1));
valve v_9_144 (.fluid_in(k_9_144), .fluid_out(k_8_72), .air_in(c_9_0));
valve v_9_145 (.fluid_in(k_9_145), .fluid_out(k_8_72), .air_in(c_9_1));
valve v_9_146 (.fluid_in(k_9_146), .fluid_out(k_8_73), .air_in(c_9_0));
valve v_9_147 (.fluid_in(k_9_147), .fluid_out(k_8_73), .air_in(c_9_1));
valve v_9_148 (.fluid_in(k_9_148), .fluid_out(k_8_74), .air_in(c_9_0));
valve v_9_149 (.fluid_in(k_9_149), .fluid_out(k_8_74), .air_in(c_9_1));
valve v_9_150 (.fluid_in(k_9_150), .fluid_out(k_8_75), .air_in(c_9_0));
valve v_9_151 (.fluid_in(k_9_151), .fluid_out(k_8_75), .air_in(c_9_1));
valve v_9_152 (.fluid_in(k_9_152), .fluid_out(k_8_76), .air_in(c_9_0));
valve v_9_153 (.fluid_in(k_9_153), .fluid_out(k_8_76), .air_in(c_9_1));
valve v_9_154 (.fluid_in(k_9_154), .fluid_out(k_8_77), .air_in(c_9_0));
valve v_9_155 (.fluid_in(k_9_155), .fluid_out(k_8_77), .air_in(c_9_1));
valve v_9_156 (.fluid_in(k_9_156), .fluid_out(k_8_78), .air_in(c_9_0));
valve v_9_157 (.fluid_in(k_9_157), .fluid_out(k_8_78), .air_in(c_9_1));
valve v_9_158 (.fluid_in(k_9_158), .fluid_out(k_8_79), .air_in(c_9_0));
valve v_9_159 (.fluid_in(k_9_159), .fluid_out(k_8_79), .air_in(c_9_1));
valve v_9_160 (.fluid_in(k_9_160), .fluid_out(k_8_80), .air_in(c_9_0));
valve v_9_161 (.fluid_in(k_9_161), .fluid_out(k_8_80), .air_in(c_9_1));
valve v_9_162 (.fluid_in(k_9_162), .fluid_out(k_8_81), .air_in(c_9_0));
valve v_9_163 (.fluid_in(k_9_163), .fluid_out(k_8_81), .air_in(c_9_1));
valve v_9_164 (.fluid_in(k_9_164), .fluid_out(k_8_82), .air_in(c_9_0));
valve v_9_165 (.fluid_in(k_9_165), .fluid_out(k_8_82), .air_in(c_9_1));
valve v_9_166 (.fluid_in(k_9_166), .fluid_out(k_8_83), .air_in(c_9_0));
valve v_9_167 (.fluid_in(k_9_167), .fluid_out(k_8_83), .air_in(c_9_1));
valve v_9_168 (.fluid_in(k_9_168), .fluid_out(k_8_84), .air_in(c_9_0));
valve v_9_169 (.fluid_in(k_9_169), .fluid_out(k_8_84), .air_in(c_9_1));
valve v_9_170 (.fluid_in(k_9_170), .fluid_out(k_8_85), .air_in(c_9_0));
valve v_9_171 (.fluid_in(k_9_171), .fluid_out(k_8_85), .air_in(c_9_1));
valve v_9_172 (.fluid_in(k_9_172), .fluid_out(k_8_86), .air_in(c_9_0));
valve v_9_173 (.fluid_in(k_9_173), .fluid_out(k_8_86), .air_in(c_9_1));
valve v_9_174 (.fluid_in(k_9_174), .fluid_out(k_8_87), .air_in(c_9_0));
valve v_9_175 (.fluid_in(k_9_175), .fluid_out(k_8_87), .air_in(c_9_1));
valve v_9_176 (.fluid_in(k_9_176), .fluid_out(k_8_88), .air_in(c_9_0));
valve v_9_177 (.fluid_in(k_9_177), .fluid_out(k_8_88), .air_in(c_9_1));
valve v_9_178 (.fluid_in(k_9_178), .fluid_out(k_8_89), .air_in(c_9_0));
valve v_9_179 (.fluid_in(k_9_179), .fluid_out(k_8_89), .air_in(c_9_1));
valve v_9_180 (.fluid_in(k_9_180), .fluid_out(k_8_90), .air_in(c_9_0));
valve v_9_181 (.fluid_in(k_9_181), .fluid_out(k_8_90), .air_in(c_9_1));
valve v_9_182 (.fluid_in(k_9_182), .fluid_out(k_8_91), .air_in(c_9_0));
valve v_9_183 (.fluid_in(k_9_183), .fluid_out(k_8_91), .air_in(c_9_1));
valve v_9_184 (.fluid_in(k_9_184), .fluid_out(k_8_92), .air_in(c_9_0));
valve v_9_185 (.fluid_in(k_9_185), .fluid_out(k_8_92), .air_in(c_9_1));
valve v_9_186 (.fluid_in(k_9_186), .fluid_out(k_8_93), .air_in(c_9_0));
valve v_9_187 (.fluid_in(k_9_187), .fluid_out(k_8_93), .air_in(c_9_1));
valve v_9_188 (.fluid_in(k_9_188), .fluid_out(k_8_94), .air_in(c_9_0));
valve v_9_189 (.fluid_in(k_9_189), .fluid_out(k_8_94), .air_in(c_9_1));
valve v_9_190 (.fluid_in(k_9_190), .fluid_out(k_8_95), .air_in(c_9_0));
valve v_9_191 (.fluid_in(k_9_191), .fluid_out(k_8_95), .air_in(c_9_1));
valve v_9_192 (.fluid_in(k_9_192), .fluid_out(k_8_96), .air_in(c_9_0));
valve v_9_193 (.fluid_in(k_9_193), .fluid_out(k_8_96), .air_in(c_9_1));
valve v_9_194 (.fluid_in(k_9_194), .fluid_out(k_8_97), .air_in(c_9_0));
valve v_9_195 (.fluid_in(k_9_195), .fluid_out(k_8_97), .air_in(c_9_1));
valve v_9_196 (.fluid_in(k_9_196), .fluid_out(k_8_98), .air_in(c_9_0));
valve v_9_197 (.fluid_in(k_9_197), .fluid_out(k_8_98), .air_in(c_9_1));
valve v_9_198 (.fluid_in(k_9_198), .fluid_out(k_8_99), .air_in(c_9_0));
valve v_9_199 (.fluid_in(k_9_199), .fluid_out(k_8_99), .air_in(c_9_1));
valve v_9_200 (.fluid_in(k_9_200), .fluid_out(k_8_100), .air_in(c_9_0));
valve v_9_201 (.fluid_in(k_9_201), .fluid_out(k_8_100), .air_in(c_9_1));
valve v_9_202 (.fluid_in(k_9_202), .fluid_out(k_8_101), .air_in(c_9_0));
valve v_9_203 (.fluid_in(k_9_203), .fluid_out(k_8_101), .air_in(c_9_1));
valve v_9_204 (.fluid_in(k_9_204), .fluid_out(k_8_102), .air_in(c_9_0));
valve v_9_205 (.fluid_in(k_9_205), .fluid_out(k_8_102), .air_in(c_9_1));
valve v_9_206 (.fluid_in(k_9_206), .fluid_out(k_8_103), .air_in(c_9_0));
valve v_9_207 (.fluid_in(k_9_207), .fluid_out(k_8_103), .air_in(c_9_1));
valve v_9_208 (.fluid_in(k_9_208), .fluid_out(k_8_104), .air_in(c_9_0));
valve v_9_209 (.fluid_in(k_9_209), .fluid_out(k_8_104), .air_in(c_9_1));
valve v_9_210 (.fluid_in(k_9_210), .fluid_out(k_8_105), .air_in(c_9_0));
valve v_9_211 (.fluid_in(k_9_211), .fluid_out(k_8_105), .air_in(c_9_1));
valve v_9_212 (.fluid_in(k_9_212), .fluid_out(k_8_106), .air_in(c_9_0));
valve v_9_213 (.fluid_in(k_9_213), .fluid_out(k_8_106), .air_in(c_9_1));
valve v_9_214 (.fluid_in(k_9_214), .fluid_out(k_8_107), .air_in(c_9_0));
valve v_9_215 (.fluid_in(k_9_215), .fluid_out(k_8_107), .air_in(c_9_1));
valve v_9_216 (.fluid_in(k_9_216), .fluid_out(k_8_108), .air_in(c_9_0));
valve v_9_217 (.fluid_in(k_9_217), .fluid_out(k_8_108), .air_in(c_9_1));
valve v_9_218 (.fluid_in(k_9_218), .fluid_out(k_8_109), .air_in(c_9_0));
valve v_9_219 (.fluid_in(k_9_219), .fluid_out(k_8_109), .air_in(c_9_1));
valve v_9_220 (.fluid_in(k_9_220), .fluid_out(k_8_110), .air_in(c_9_0));
valve v_9_221 (.fluid_in(k_9_221), .fluid_out(k_8_110), .air_in(c_9_1));
valve v_9_222 (.fluid_in(k_9_222), .fluid_out(k_8_111), .air_in(c_9_0));
valve v_9_223 (.fluid_in(k_9_223), .fluid_out(k_8_111), .air_in(c_9_1));
valve v_9_224 (.fluid_in(k_9_224), .fluid_out(k_8_112), .air_in(c_9_0));
valve v_9_225 (.fluid_in(k_9_225), .fluid_out(k_8_112), .air_in(c_9_1));
valve v_9_226 (.fluid_in(k_9_226), .fluid_out(k_8_113), .air_in(c_9_0));
valve v_9_227 (.fluid_in(k_9_227), .fluid_out(k_8_113), .air_in(c_9_1));
valve v_9_228 (.fluid_in(k_9_228), .fluid_out(k_8_114), .air_in(c_9_0));
valve v_9_229 (.fluid_in(k_9_229), .fluid_out(k_8_114), .air_in(c_9_1));
valve v_9_230 (.fluid_in(k_9_230), .fluid_out(k_8_115), .air_in(c_9_0));
valve v_9_231 (.fluid_in(k_9_231), .fluid_out(k_8_115), .air_in(c_9_1));
valve v_9_232 (.fluid_in(k_9_232), .fluid_out(k_8_116), .air_in(c_9_0));
valve v_9_233 (.fluid_in(k_9_233), .fluid_out(k_8_116), .air_in(c_9_1));
valve v_9_234 (.fluid_in(k_9_234), .fluid_out(k_8_117), .air_in(c_9_0));
valve v_9_235 (.fluid_in(k_9_235), .fluid_out(k_8_117), .air_in(c_9_1));
valve v_9_236 (.fluid_in(k_9_236), .fluid_out(k_8_118), .air_in(c_9_0));
valve v_9_237 (.fluid_in(k_9_237), .fluid_out(k_8_118), .air_in(c_9_1));
valve v_9_238 (.fluid_in(k_9_238), .fluid_out(k_8_119), .air_in(c_9_0));
valve v_9_239 (.fluid_in(k_9_239), .fluid_out(k_8_119), .air_in(c_9_1));
valve v_9_240 (.fluid_in(k_9_240), .fluid_out(k_8_120), .air_in(c_9_0));
valve v_9_241 (.fluid_in(k_9_241), .fluid_out(k_8_120), .air_in(c_9_1));
valve v_9_242 (.fluid_in(k_9_242), .fluid_out(k_8_121), .air_in(c_9_0));
valve v_9_243 (.fluid_in(k_9_243), .fluid_out(k_8_121), .air_in(c_9_1));
valve v_9_244 (.fluid_in(k_9_244), .fluid_out(k_8_122), .air_in(c_9_0));
valve v_9_245 (.fluid_in(k_9_245), .fluid_out(k_8_122), .air_in(c_9_1));
valve v_9_246 (.fluid_in(k_9_246), .fluid_out(k_8_123), .air_in(c_9_0));
valve v_9_247 (.fluid_in(k_9_247), .fluid_out(k_8_123), .air_in(c_9_1));
valve v_9_248 (.fluid_in(k_9_248), .fluid_out(k_8_124), .air_in(c_9_0));
valve v_9_249 (.fluid_in(k_9_249), .fluid_out(k_8_124), .air_in(c_9_1));
valve v_9_250 (.fluid_in(k_9_250), .fluid_out(k_8_125), .air_in(c_9_0));
valve v_9_251 (.fluid_in(k_9_251), .fluid_out(k_8_125), .air_in(c_9_1));
valve v_9_252 (.fluid_in(k_9_252), .fluid_out(k_8_126), .air_in(c_9_0));
valve v_9_253 (.fluid_in(k_9_253), .fluid_out(k_8_126), .air_in(c_9_1));
valve v_9_254 (.fluid_in(k_9_254), .fluid_out(k_8_127), .air_in(c_9_0));
valve v_9_255 (.fluid_in(k_9_255), .fluid_out(k_8_127), .air_in(c_9_1));
valve v_9_256 (.fluid_in(k_9_256), .fluid_out(k_8_128), .air_in(c_9_0));
valve v_9_257 (.fluid_in(k_9_257), .fluid_out(k_8_128), .air_in(c_9_1));
valve v_9_258 (.fluid_in(k_9_258), .fluid_out(k_8_129), .air_in(c_9_0));
valve v_9_259 (.fluid_in(k_9_259), .fluid_out(k_8_129), .air_in(c_9_1));
valve v_9_260 (.fluid_in(k_9_260), .fluid_out(k_8_130), .air_in(c_9_0));
valve v_9_261 (.fluid_in(k_9_261), .fluid_out(k_8_130), .air_in(c_9_1));
valve v_9_262 (.fluid_in(k_9_262), .fluid_out(k_8_131), .air_in(c_9_0));
valve v_9_263 (.fluid_in(k_9_263), .fluid_out(k_8_131), .air_in(c_9_1));
valve v_9_264 (.fluid_in(k_9_264), .fluid_out(k_8_132), .air_in(c_9_0));
valve v_9_265 (.fluid_in(k_9_265), .fluid_out(k_8_132), .air_in(c_9_1));
valve v_9_266 (.fluid_in(k_9_266), .fluid_out(k_8_133), .air_in(c_9_0));
valve v_9_267 (.fluid_in(k_9_267), .fluid_out(k_8_133), .air_in(c_9_1));
valve v_9_268 (.fluid_in(k_9_268), .fluid_out(k_8_134), .air_in(c_9_0));
valve v_9_269 (.fluid_in(k_9_269), .fluid_out(k_8_134), .air_in(c_9_1));
valve v_9_270 (.fluid_in(k_9_270), .fluid_out(k_8_135), .air_in(c_9_0));
valve v_9_271 (.fluid_in(k_9_271), .fluid_out(k_8_135), .air_in(c_9_1));
valve v_9_272 (.fluid_in(k_9_272), .fluid_out(k_8_136), .air_in(c_9_0));
valve v_9_273 (.fluid_in(k_9_273), .fluid_out(k_8_136), .air_in(c_9_1));
valve v_9_274 (.fluid_in(k_9_274), .fluid_out(k_8_137), .air_in(c_9_0));
valve v_9_275 (.fluid_in(k_9_275), .fluid_out(k_8_137), .air_in(c_9_1));
valve v_9_276 (.fluid_in(k_9_276), .fluid_out(k_8_138), .air_in(c_9_0));
valve v_9_277 (.fluid_in(k_9_277), .fluid_out(k_8_138), .air_in(c_9_1));
valve v_9_278 (.fluid_in(k_9_278), .fluid_out(k_8_139), .air_in(c_9_0));
valve v_9_279 (.fluid_in(k_9_279), .fluid_out(k_8_139), .air_in(c_9_1));
valve v_9_280 (.fluid_in(k_9_280), .fluid_out(k_8_140), .air_in(c_9_0));
valve v_9_281 (.fluid_in(k_9_281), .fluid_out(k_8_140), .air_in(c_9_1));
valve v_9_282 (.fluid_in(k_9_282), .fluid_out(k_8_141), .air_in(c_9_0));
valve v_9_283 (.fluid_in(k_9_283), .fluid_out(k_8_141), .air_in(c_9_1));
valve v_9_284 (.fluid_in(k_9_284), .fluid_out(k_8_142), .air_in(c_9_0));
valve v_9_285 (.fluid_in(k_9_285), .fluid_out(k_8_142), .air_in(c_9_1));
valve v_9_286 (.fluid_in(k_9_286), .fluid_out(k_8_143), .air_in(c_9_0));
valve v_9_287 (.fluid_in(k_9_287), .fluid_out(k_8_143), .air_in(c_9_1));
valve v_9_288 (.fluid_in(k_9_288), .fluid_out(k_8_144), .air_in(c_9_0));
valve v_9_289 (.fluid_in(k_9_289), .fluid_out(k_8_144), .air_in(c_9_1));
valve v_9_290 (.fluid_in(k_9_290), .fluid_out(k_8_145), .air_in(c_9_0));
valve v_9_291 (.fluid_in(k_9_291), .fluid_out(k_8_145), .air_in(c_9_1));
valve v_9_292 (.fluid_in(k_9_292), .fluid_out(k_8_146), .air_in(c_9_0));
valve v_9_293 (.fluid_in(k_9_293), .fluid_out(k_8_146), .air_in(c_9_1));
valve v_9_294 (.fluid_in(k_9_294), .fluid_out(k_8_147), .air_in(c_9_0));
valve v_9_295 (.fluid_in(k_9_295), .fluid_out(k_8_147), .air_in(c_9_1));
valve v_9_296 (.fluid_in(k_9_296), .fluid_out(k_8_148), .air_in(c_9_0));
valve v_9_297 (.fluid_in(k_9_297), .fluid_out(k_8_148), .air_in(c_9_1));
valve v_9_298 (.fluid_in(k_9_298), .fluid_out(k_8_149), .air_in(c_9_0));
valve v_9_299 (.fluid_in(k_9_299), .fluid_out(k_8_149), .air_in(c_9_1));
valve v_9_300 (.fluid_in(k_9_300), .fluid_out(k_8_150), .air_in(c_9_0));
valve v_9_301 (.fluid_in(k_9_301), .fluid_out(k_8_150), .air_in(c_9_1));
valve v_9_302 (.fluid_in(k_9_302), .fluid_out(k_8_151), .air_in(c_9_0));
valve v_9_303 (.fluid_in(k_9_303), .fluid_out(k_8_151), .air_in(c_9_1));
valve v_9_304 (.fluid_in(k_9_304), .fluid_out(k_8_152), .air_in(c_9_0));
valve v_9_305 (.fluid_in(k_9_305), .fluid_out(k_8_152), .air_in(c_9_1));
valve v_9_306 (.fluid_in(k_9_306), .fluid_out(k_8_153), .air_in(c_9_0));
valve v_9_307 (.fluid_in(k_9_307), .fluid_out(k_8_153), .air_in(c_9_1));
valve v_9_308 (.fluid_in(k_9_308), .fluid_out(k_8_154), .air_in(c_9_0));
valve v_9_309 (.fluid_in(k_9_309), .fluid_out(k_8_154), .air_in(c_9_1));
valve v_9_310 (.fluid_in(k_9_310), .fluid_out(k_8_155), .air_in(c_9_0));
valve v_9_311 (.fluid_in(k_9_311), .fluid_out(k_8_155), .air_in(c_9_1));
valve v_9_312 (.fluid_in(k_9_312), .fluid_out(k_8_156), .air_in(c_9_0));
valve v_9_313 (.fluid_in(k_9_313), .fluid_out(k_8_156), .air_in(c_9_1));
valve v_9_314 (.fluid_in(k_9_314), .fluid_out(k_8_157), .air_in(c_9_0));
valve v_9_315 (.fluid_in(k_9_315), .fluid_out(k_8_157), .air_in(c_9_1));
valve v_9_316 (.fluid_in(k_9_316), .fluid_out(k_8_158), .air_in(c_9_0));
valve v_9_317 (.fluid_in(k_9_317), .fluid_out(k_8_158), .air_in(c_9_1));
valve v_9_318 (.fluid_in(k_9_318), .fluid_out(k_8_159), .air_in(c_9_0));
valve v_9_319 (.fluid_in(k_9_319), .fluid_out(k_8_159), .air_in(c_9_1));
valve v_9_320 (.fluid_in(k_9_320), .fluid_out(k_8_160), .air_in(c_9_0));
valve v_9_321 (.fluid_in(k_9_321), .fluid_out(k_8_160), .air_in(c_9_1));
valve v_9_322 (.fluid_in(k_9_322), .fluid_out(k_8_161), .air_in(c_9_0));
valve v_9_323 (.fluid_in(k_9_323), .fluid_out(k_8_161), .air_in(c_9_1));
valve v_9_324 (.fluid_in(k_9_324), .fluid_out(k_8_162), .air_in(c_9_0));
valve v_9_325 (.fluid_in(k_9_325), .fluid_out(k_8_162), .air_in(c_9_1));
valve v_9_326 (.fluid_in(k_9_326), .fluid_out(k_8_163), .air_in(c_9_0));
valve v_9_327 (.fluid_in(k_9_327), .fluid_out(k_8_163), .air_in(c_9_1));
valve v_9_328 (.fluid_in(k_9_328), .fluid_out(k_8_164), .air_in(c_9_0));
valve v_9_329 (.fluid_in(k_9_329), .fluid_out(k_8_164), .air_in(c_9_1));
valve v_9_330 (.fluid_in(k_9_330), .fluid_out(k_8_165), .air_in(c_9_0));
valve v_9_331 (.fluid_in(k_9_331), .fluid_out(k_8_165), .air_in(c_9_1));
valve v_9_332 (.fluid_in(k_9_332), .fluid_out(k_8_166), .air_in(c_9_0));
valve v_9_333 (.fluid_in(k_9_333), .fluid_out(k_8_166), .air_in(c_9_1));
valve v_9_334 (.fluid_in(k_9_334), .fluid_out(k_8_167), .air_in(c_9_0));
valve v_9_335 (.fluid_in(k_9_335), .fluid_out(k_8_167), .air_in(c_9_1));
valve v_9_336 (.fluid_in(k_9_336), .fluid_out(k_8_168), .air_in(c_9_0));
valve v_9_337 (.fluid_in(k_9_337), .fluid_out(k_8_168), .air_in(c_9_1));
valve v_9_338 (.fluid_in(k_9_338), .fluid_out(k_8_169), .air_in(c_9_0));
valve v_9_339 (.fluid_in(k_9_339), .fluid_out(k_8_169), .air_in(c_9_1));
valve v_9_340 (.fluid_in(k_9_340), .fluid_out(k_8_170), .air_in(c_9_0));
valve v_9_341 (.fluid_in(k_9_341), .fluid_out(k_8_170), .air_in(c_9_1));
valve v_9_342 (.fluid_in(k_9_342), .fluid_out(k_8_171), .air_in(c_9_0));
valve v_9_343 (.fluid_in(k_9_343), .fluid_out(k_8_171), .air_in(c_9_1));
valve v_9_344 (.fluid_in(k_9_344), .fluid_out(k_8_172), .air_in(c_9_0));
valve v_9_345 (.fluid_in(k_9_345), .fluid_out(k_8_172), .air_in(c_9_1));
valve v_9_346 (.fluid_in(k_9_346), .fluid_out(k_8_173), .air_in(c_9_0));
valve v_9_347 (.fluid_in(k_9_347), .fluid_out(k_8_173), .air_in(c_9_1));
valve v_9_348 (.fluid_in(k_9_348), .fluid_out(k_8_174), .air_in(c_9_0));
valve v_9_349 (.fluid_in(k_9_349), .fluid_out(k_8_174), .air_in(c_9_1));
valve v_9_350 (.fluid_in(k_9_350), .fluid_out(k_8_175), .air_in(c_9_0));
valve v_9_351 (.fluid_in(k_9_351), .fluid_out(k_8_175), .air_in(c_9_1));
valve v_9_352 (.fluid_in(k_9_352), .fluid_out(k_8_176), .air_in(c_9_0));
valve v_9_353 (.fluid_in(k_9_353), .fluid_out(k_8_176), .air_in(c_9_1));
valve v_9_354 (.fluid_in(k_9_354), .fluid_out(k_8_177), .air_in(c_9_0));
valve v_9_355 (.fluid_in(k_9_355), .fluid_out(k_8_177), .air_in(c_9_1));
valve v_9_356 (.fluid_in(k_9_356), .fluid_out(k_8_178), .air_in(c_9_0));
valve v_9_357 (.fluid_in(k_9_357), .fluid_out(k_8_178), .air_in(c_9_1));
valve v_9_358 (.fluid_in(k_9_358), .fluid_out(k_8_179), .air_in(c_9_0));
valve v_9_359 (.fluid_in(k_9_359), .fluid_out(k_8_179), .air_in(c_9_1));
valve v_9_360 (.fluid_in(k_9_360), .fluid_out(k_8_180), .air_in(c_9_0));
valve v_9_361 (.fluid_in(k_9_361), .fluid_out(k_8_180), .air_in(c_9_1));
valve v_9_362 (.fluid_in(k_9_362), .fluid_out(k_8_181), .air_in(c_9_0));
valve v_9_363 (.fluid_in(k_9_363), .fluid_out(k_8_181), .air_in(c_9_1));
valve v_9_364 (.fluid_in(k_9_364), .fluid_out(k_8_182), .air_in(c_9_0));
valve v_9_365 (.fluid_in(k_9_365), .fluid_out(k_8_182), .air_in(c_9_1));
valve v_9_366 (.fluid_in(k_9_366), .fluid_out(k_8_183), .air_in(c_9_0));
valve v_9_367 (.fluid_in(k_9_367), .fluid_out(k_8_183), .air_in(c_9_1));
valve v_9_368 (.fluid_in(k_9_368), .fluid_out(k_8_184), .air_in(c_9_0));
valve v_9_369 (.fluid_in(k_9_369), .fluid_out(k_8_184), .air_in(c_9_1));
valve v_9_370 (.fluid_in(k_9_370), .fluid_out(k_8_185), .air_in(c_9_0));
valve v_9_371 (.fluid_in(k_9_371), .fluid_out(k_8_185), .air_in(c_9_1));
valve v_9_372 (.fluid_in(k_9_372), .fluid_out(k_8_186), .air_in(c_9_0));
valve v_9_373 (.fluid_in(k_9_373), .fluid_out(k_8_186), .air_in(c_9_1));
valve v_9_374 (.fluid_in(k_9_374), .fluid_out(k_8_187), .air_in(c_9_0));
valve v_9_375 (.fluid_in(k_9_375), .fluid_out(k_8_187), .air_in(c_9_1));
valve v_9_376 (.fluid_in(k_9_376), .fluid_out(k_8_188), .air_in(c_9_0));
valve v_9_377 (.fluid_in(k_9_377), .fluid_out(k_8_188), .air_in(c_9_1));
valve v_9_378 (.fluid_in(k_9_378), .fluid_out(k_8_189), .air_in(c_9_0));
valve v_9_379 (.fluid_in(k_9_379), .fluid_out(k_8_189), .air_in(c_9_1));
valve v_9_380 (.fluid_in(k_9_380), .fluid_out(k_8_190), .air_in(c_9_0));
valve v_9_381 (.fluid_in(k_9_381), .fluid_out(k_8_190), .air_in(c_9_1));
valve v_9_382 (.fluid_in(k_9_382), .fluid_out(k_8_191), .air_in(c_9_0));
valve v_9_383 (.fluid_in(k_9_383), .fluid_out(k_8_191), .air_in(c_9_1));
valve v_9_384 (.fluid_in(k_9_384), .fluid_out(k_8_192), .air_in(c_9_0));
valve v_9_385 (.fluid_in(k_9_385), .fluid_out(k_8_192), .air_in(c_9_1));
valve v_9_386 (.fluid_in(k_9_386), .fluid_out(k_8_193), .air_in(c_9_0));
valve v_9_387 (.fluid_in(k_9_387), .fluid_out(k_8_193), .air_in(c_9_1));
valve v_9_388 (.fluid_in(k_9_388), .fluid_out(k_8_194), .air_in(c_9_0));
valve v_9_389 (.fluid_in(k_9_389), .fluid_out(k_8_194), .air_in(c_9_1));
valve v_9_390 (.fluid_in(k_9_390), .fluid_out(k_8_195), .air_in(c_9_0));
valve v_9_391 (.fluid_in(k_9_391), .fluid_out(k_8_195), .air_in(c_9_1));
valve v_9_392 (.fluid_in(k_9_392), .fluid_out(k_8_196), .air_in(c_9_0));
valve v_9_393 (.fluid_in(k_9_393), .fluid_out(k_8_196), .air_in(c_9_1));
valve v_9_394 (.fluid_in(k_9_394), .fluid_out(k_8_197), .air_in(c_9_0));
valve v_9_395 (.fluid_in(k_9_395), .fluid_out(k_8_197), .air_in(c_9_1));
valve v_9_396 (.fluid_in(k_9_396), .fluid_out(k_8_198), .air_in(c_9_0));
valve v_9_397 (.fluid_in(k_9_397), .fluid_out(k_8_198), .air_in(c_9_1));
valve v_9_398 (.fluid_in(k_9_398), .fluid_out(k_8_199), .air_in(c_9_0));
valve v_9_399 (.fluid_in(k_9_399), .fluid_out(k_8_199), .air_in(c_9_1));
valve v_9_400 (.fluid_in(k_9_400), .fluid_out(k_8_200), .air_in(c_9_0));
valve v_9_401 (.fluid_in(k_9_401), .fluid_out(k_8_200), .air_in(c_9_1));
valve v_9_402 (.fluid_in(k_9_402), .fluid_out(k_8_201), .air_in(c_9_0));
valve v_9_403 (.fluid_in(k_9_403), .fluid_out(k_8_201), .air_in(c_9_1));
valve v_9_404 (.fluid_in(k_9_404), .fluid_out(k_8_202), .air_in(c_9_0));
valve v_9_405 (.fluid_in(k_9_405), .fluid_out(k_8_202), .air_in(c_9_1));
valve v_9_406 (.fluid_in(k_9_406), .fluid_out(k_8_203), .air_in(c_9_0));
valve v_9_407 (.fluid_in(k_9_407), .fluid_out(k_8_203), .air_in(c_9_1));
valve v_9_408 (.fluid_in(k_9_408), .fluid_out(k_8_204), .air_in(c_9_0));
valve v_9_409 (.fluid_in(k_9_409), .fluid_out(k_8_204), .air_in(c_9_1));
valve v_9_410 (.fluid_in(k_9_410), .fluid_out(k_8_205), .air_in(c_9_0));
valve v_9_411 (.fluid_in(k_9_411), .fluid_out(k_8_205), .air_in(c_9_1));
valve v_9_412 (.fluid_in(k_9_412), .fluid_out(k_8_206), .air_in(c_9_0));
valve v_9_413 (.fluid_in(k_9_413), .fluid_out(k_8_206), .air_in(c_9_1));
valve v_9_414 (.fluid_in(k_9_414), .fluid_out(k_8_207), .air_in(c_9_0));
valve v_9_415 (.fluid_in(k_9_415), .fluid_out(k_8_207), .air_in(c_9_1));
valve v_9_416 (.fluid_in(k_9_416), .fluid_out(k_8_208), .air_in(c_9_0));
valve v_9_417 (.fluid_in(k_9_417), .fluid_out(k_8_208), .air_in(c_9_1));
valve v_9_418 (.fluid_in(k_9_418), .fluid_out(k_8_209), .air_in(c_9_0));
valve v_9_419 (.fluid_in(k_9_419), .fluid_out(k_8_209), .air_in(c_9_1));
valve v_9_420 (.fluid_in(k_9_420), .fluid_out(k_8_210), .air_in(c_9_0));
valve v_9_421 (.fluid_in(k_9_421), .fluid_out(k_8_210), .air_in(c_9_1));
valve v_9_422 (.fluid_in(k_9_422), .fluid_out(k_8_211), .air_in(c_9_0));
valve v_9_423 (.fluid_in(k_9_423), .fluid_out(k_8_211), .air_in(c_9_1));
valve v_9_424 (.fluid_in(k_9_424), .fluid_out(k_8_212), .air_in(c_9_0));
valve v_9_425 (.fluid_in(k_9_425), .fluid_out(k_8_212), .air_in(c_9_1));
valve v_9_426 (.fluid_in(k_9_426), .fluid_out(k_8_213), .air_in(c_9_0));
valve v_9_427 (.fluid_in(k_9_427), .fluid_out(k_8_213), .air_in(c_9_1));
valve v_9_428 (.fluid_in(k_9_428), .fluid_out(k_8_214), .air_in(c_9_0));
valve v_9_429 (.fluid_in(k_9_429), .fluid_out(k_8_214), .air_in(c_9_1));
valve v_9_430 (.fluid_in(k_9_430), .fluid_out(k_8_215), .air_in(c_9_0));
valve v_9_431 (.fluid_in(k_9_431), .fluid_out(k_8_215), .air_in(c_9_1));
valve v_9_432 (.fluid_in(k_9_432), .fluid_out(k_8_216), .air_in(c_9_0));
valve v_9_433 (.fluid_in(k_9_433), .fluid_out(k_8_216), .air_in(c_9_1));
valve v_9_434 (.fluid_in(k_9_434), .fluid_out(k_8_217), .air_in(c_9_0));
valve v_9_435 (.fluid_in(k_9_435), .fluid_out(k_8_217), .air_in(c_9_1));
valve v_9_436 (.fluid_in(k_9_436), .fluid_out(k_8_218), .air_in(c_9_0));
valve v_9_437 (.fluid_in(k_9_437), .fluid_out(k_8_218), .air_in(c_9_1));
valve v_9_438 (.fluid_in(k_9_438), .fluid_out(k_8_219), .air_in(c_9_0));
valve v_9_439 (.fluid_in(k_9_439), .fluid_out(k_8_219), .air_in(c_9_1));
valve v_9_440 (.fluid_in(k_9_440), .fluid_out(k_8_220), .air_in(c_9_0));
valve v_9_441 (.fluid_in(k_9_441), .fluid_out(k_8_220), .air_in(c_9_1));
valve v_9_442 (.fluid_in(k_9_442), .fluid_out(k_8_221), .air_in(c_9_0));
valve v_9_443 (.fluid_in(k_9_443), .fluid_out(k_8_221), .air_in(c_9_1));
valve v_9_444 (.fluid_in(k_9_444), .fluid_out(k_8_222), .air_in(c_9_0));
valve v_9_445 (.fluid_in(k_9_445), .fluid_out(k_8_222), .air_in(c_9_1));
valve v_9_446 (.fluid_in(k_9_446), .fluid_out(k_8_223), .air_in(c_9_0));
valve v_9_447 (.fluid_in(k_9_447), .fluid_out(k_8_223), .air_in(c_9_1));
valve v_9_448 (.fluid_in(k_9_448), .fluid_out(k_8_224), .air_in(c_9_0));
valve v_9_449 (.fluid_in(k_9_449), .fluid_out(k_8_224), .air_in(c_9_1));
valve v_9_450 (.fluid_in(k_9_450), .fluid_out(k_8_225), .air_in(c_9_0));
valve v_9_451 (.fluid_in(k_9_451), .fluid_out(k_8_225), .air_in(c_9_1));
valve v_9_452 (.fluid_in(k_9_452), .fluid_out(k_8_226), .air_in(c_9_0));
valve v_9_453 (.fluid_in(k_9_453), .fluid_out(k_8_226), .air_in(c_9_1));
valve v_9_454 (.fluid_in(k_9_454), .fluid_out(k_8_227), .air_in(c_9_0));
valve v_9_455 (.fluid_in(k_9_455), .fluid_out(k_8_227), .air_in(c_9_1));
valve v_9_456 (.fluid_in(k_9_456), .fluid_out(k_8_228), .air_in(c_9_0));
valve v_9_457 (.fluid_in(k_9_457), .fluid_out(k_8_228), .air_in(c_9_1));
valve v_9_458 (.fluid_in(k_9_458), .fluid_out(k_8_229), .air_in(c_9_0));
valve v_9_459 (.fluid_in(k_9_459), .fluid_out(k_8_229), .air_in(c_9_1));
valve v_9_460 (.fluid_in(k_9_460), .fluid_out(k_8_230), .air_in(c_9_0));
valve v_9_461 (.fluid_in(k_9_461), .fluid_out(k_8_230), .air_in(c_9_1));
valve v_9_462 (.fluid_in(k_9_462), .fluid_out(k_8_231), .air_in(c_9_0));
valve v_9_463 (.fluid_in(k_9_463), .fluid_out(k_8_231), .air_in(c_9_1));
valve v_9_464 (.fluid_in(k_9_464), .fluid_out(k_8_232), .air_in(c_9_0));
valve v_9_465 (.fluid_in(k_9_465), .fluid_out(k_8_232), .air_in(c_9_1));
valve v_9_466 (.fluid_in(k_9_466), .fluid_out(k_8_233), .air_in(c_9_0));
valve v_9_467 (.fluid_in(k_9_467), .fluid_out(k_8_233), .air_in(c_9_1));
valve v_9_468 (.fluid_in(k_9_468), .fluid_out(k_8_234), .air_in(c_9_0));
valve v_9_469 (.fluid_in(k_9_469), .fluid_out(k_8_234), .air_in(c_9_1));
valve v_9_470 (.fluid_in(k_9_470), .fluid_out(k_8_235), .air_in(c_9_0));
valve v_9_471 (.fluid_in(k_9_471), .fluid_out(k_8_235), .air_in(c_9_1));
valve v_9_472 (.fluid_in(k_9_472), .fluid_out(k_8_236), .air_in(c_9_0));
valve v_9_473 (.fluid_in(k_9_473), .fluid_out(k_8_236), .air_in(c_9_1));
valve v_9_474 (.fluid_in(k_9_474), .fluid_out(k_8_237), .air_in(c_9_0));
valve v_9_475 (.fluid_in(k_9_475), .fluid_out(k_8_237), .air_in(c_9_1));
valve v_9_476 (.fluid_in(k_9_476), .fluid_out(k_8_238), .air_in(c_9_0));
valve v_9_477 (.fluid_in(k_9_477), .fluid_out(k_8_238), .air_in(c_9_1));
valve v_9_478 (.fluid_in(k_9_478), .fluid_out(k_8_239), .air_in(c_9_0));
valve v_9_479 (.fluid_in(k_9_479), .fluid_out(k_8_239), .air_in(c_9_1));
valve v_9_480 (.fluid_in(k_9_480), .fluid_out(k_8_240), .air_in(c_9_0));
valve v_9_481 (.fluid_in(k_9_481), .fluid_out(k_8_240), .air_in(c_9_1));
valve v_9_482 (.fluid_in(k_9_482), .fluid_out(k_8_241), .air_in(c_9_0));
valve v_9_483 (.fluid_in(k_9_483), .fluid_out(k_8_241), .air_in(c_9_1));
valve v_9_484 (.fluid_in(k_9_484), .fluid_out(k_8_242), .air_in(c_9_0));
valve v_9_485 (.fluid_in(k_9_485), .fluid_out(k_8_242), .air_in(c_9_1));
valve v_9_486 (.fluid_in(k_9_486), .fluid_out(k_8_243), .air_in(c_9_0));
valve v_9_487 (.fluid_in(k_9_487), .fluid_out(k_8_243), .air_in(c_9_1));
valve v_9_488 (.fluid_in(k_9_488), .fluid_out(k_8_244), .air_in(c_9_0));
valve v_9_489 (.fluid_in(k_9_489), .fluid_out(k_8_244), .air_in(c_9_1));
valve v_9_490 (.fluid_in(k_9_490), .fluid_out(k_8_245), .air_in(c_9_0));
valve v_9_491 (.fluid_in(k_9_491), .fluid_out(k_8_245), .air_in(c_9_1));
valve v_9_492 (.fluid_in(k_9_492), .fluid_out(k_8_246), .air_in(c_9_0));
valve v_9_493 (.fluid_in(k_9_493), .fluid_out(k_8_246), .air_in(c_9_1));
valve v_9_494 (.fluid_in(k_9_494), .fluid_out(k_8_247), .air_in(c_9_0));
valve v_9_495 (.fluid_in(k_9_495), .fluid_out(k_8_247), .air_in(c_9_1));
valve v_9_496 (.fluid_in(k_9_496), .fluid_out(k_8_248), .air_in(c_9_0));
valve v_9_497 (.fluid_in(k_9_497), .fluid_out(k_8_248), .air_in(c_9_1));
valve v_9_498 (.fluid_in(k_9_498), .fluid_out(k_8_249), .air_in(c_9_0));
valve v_9_499 (.fluid_in(k_9_499), .fluid_out(k_8_249), .air_in(c_9_1));
valve v_9_500 (.fluid_in(k_9_500), .fluid_out(k_8_250), .air_in(c_9_0));
valve v_9_501 (.fluid_in(k_9_501), .fluid_out(k_8_250), .air_in(c_9_1));
valve v_9_502 (.fluid_in(k_9_502), .fluid_out(k_8_251), .air_in(c_9_0));
valve v_9_503 (.fluid_in(k_9_503), .fluid_out(k_8_251), .air_in(c_9_1));
valve v_9_504 (.fluid_in(k_9_504), .fluid_out(k_8_252), .air_in(c_9_0));
valve v_9_505 (.fluid_in(k_9_505), .fluid_out(k_8_252), .air_in(c_9_1));
valve v_9_506 (.fluid_in(k_9_506), .fluid_out(k_8_253), .air_in(c_9_0));
valve v_9_507 (.fluid_in(k_9_507), .fluid_out(k_8_253), .air_in(c_9_1));
valve v_9_508 (.fluid_in(k_9_508), .fluid_out(k_8_254), .air_in(c_9_0));
valve v_9_509 (.fluid_in(k_9_509), .fluid_out(k_8_254), .air_in(c_9_1));
valve v_9_510 (.fluid_in(k_9_510), .fluid_out(k_8_255), .air_in(c_9_0));
valve v_9_511 (.fluid_in(k_9_511), .fluid_out(k_8_255), .air_in(c_9_1));
valve v_10_0 (.fluid_in(k_10_0), .fluid_out(k_9_0), .air_in(c_10_0));
valve v_10_1 (.fluid_in(k_10_1), .fluid_out(k_9_0), .air_in(c_10_1));
valve v_10_2 (.fluid_in(k_10_2), .fluid_out(k_9_1), .air_in(c_10_0));
valve v_10_3 (.fluid_in(k_10_3), .fluid_out(k_9_1), .air_in(c_10_1));
valve v_10_4 (.fluid_in(k_10_4), .fluid_out(k_9_2), .air_in(c_10_0));
valve v_10_5 (.fluid_in(k_10_5), .fluid_out(k_9_2), .air_in(c_10_1));
valve v_10_6 (.fluid_in(k_10_6), .fluid_out(k_9_3), .air_in(c_10_0));
valve v_10_7 (.fluid_in(k_10_7), .fluid_out(k_9_3), .air_in(c_10_1));
valve v_10_8 (.fluid_in(k_10_8), .fluid_out(k_9_4), .air_in(c_10_0));
valve v_10_9 (.fluid_in(k_10_9), .fluid_out(k_9_4), .air_in(c_10_1));
valve v_10_10 (.fluid_in(k_10_10), .fluid_out(k_9_5), .air_in(c_10_0));
valve v_10_11 (.fluid_in(k_10_11), .fluid_out(k_9_5), .air_in(c_10_1));
valve v_10_12 (.fluid_in(k_10_12), .fluid_out(k_9_6), .air_in(c_10_0));
valve v_10_13 (.fluid_in(k_10_13), .fluid_out(k_9_6), .air_in(c_10_1));
valve v_10_14 (.fluid_in(k_10_14), .fluid_out(k_9_7), .air_in(c_10_0));
valve v_10_15 (.fluid_in(k_10_15), .fluid_out(k_9_7), .air_in(c_10_1));
valve v_10_16 (.fluid_in(k_10_16), .fluid_out(k_9_8), .air_in(c_10_0));
valve v_10_17 (.fluid_in(k_10_17), .fluid_out(k_9_8), .air_in(c_10_1));
valve v_10_18 (.fluid_in(k_10_18), .fluid_out(k_9_9), .air_in(c_10_0));
valve v_10_19 (.fluid_in(k_10_19), .fluid_out(k_9_9), .air_in(c_10_1));
valve v_10_20 (.fluid_in(k_10_20), .fluid_out(k_9_10), .air_in(c_10_0));
valve v_10_21 (.fluid_in(k_10_21), .fluid_out(k_9_10), .air_in(c_10_1));
valve v_10_22 (.fluid_in(k_10_22), .fluid_out(k_9_11), .air_in(c_10_0));
valve v_10_23 (.fluid_in(k_10_23), .fluid_out(k_9_11), .air_in(c_10_1));
valve v_10_24 (.fluid_in(k_10_24), .fluid_out(k_9_12), .air_in(c_10_0));
valve v_10_25 (.fluid_in(k_10_25), .fluid_out(k_9_12), .air_in(c_10_1));
valve v_10_26 (.fluid_in(k_10_26), .fluid_out(k_9_13), .air_in(c_10_0));
valve v_10_27 (.fluid_in(k_10_27), .fluid_out(k_9_13), .air_in(c_10_1));
valve v_10_28 (.fluid_in(k_10_28), .fluid_out(k_9_14), .air_in(c_10_0));
valve v_10_29 (.fluid_in(k_10_29), .fluid_out(k_9_14), .air_in(c_10_1));
valve v_10_30 (.fluid_in(k_10_30), .fluid_out(k_9_15), .air_in(c_10_0));
valve v_10_31 (.fluid_in(k_10_31), .fluid_out(k_9_15), .air_in(c_10_1));
valve v_10_32 (.fluid_in(k_10_32), .fluid_out(k_9_16), .air_in(c_10_0));
valve v_10_33 (.fluid_in(k_10_33), .fluid_out(k_9_16), .air_in(c_10_1));
valve v_10_34 (.fluid_in(k_10_34), .fluid_out(k_9_17), .air_in(c_10_0));
valve v_10_35 (.fluid_in(k_10_35), .fluid_out(k_9_17), .air_in(c_10_1));
valve v_10_36 (.fluid_in(k_10_36), .fluid_out(k_9_18), .air_in(c_10_0));
valve v_10_37 (.fluid_in(k_10_37), .fluid_out(k_9_18), .air_in(c_10_1));
valve v_10_38 (.fluid_in(k_10_38), .fluid_out(k_9_19), .air_in(c_10_0));
valve v_10_39 (.fluid_in(k_10_39), .fluid_out(k_9_19), .air_in(c_10_1));
valve v_10_40 (.fluid_in(k_10_40), .fluid_out(k_9_20), .air_in(c_10_0));
valve v_10_41 (.fluid_in(k_10_41), .fluid_out(k_9_20), .air_in(c_10_1));
valve v_10_42 (.fluid_in(k_10_42), .fluid_out(k_9_21), .air_in(c_10_0));
valve v_10_43 (.fluid_in(k_10_43), .fluid_out(k_9_21), .air_in(c_10_1));
valve v_10_44 (.fluid_in(k_10_44), .fluid_out(k_9_22), .air_in(c_10_0));
valve v_10_45 (.fluid_in(k_10_45), .fluid_out(k_9_22), .air_in(c_10_1));
valve v_10_46 (.fluid_in(k_10_46), .fluid_out(k_9_23), .air_in(c_10_0));
valve v_10_47 (.fluid_in(k_10_47), .fluid_out(k_9_23), .air_in(c_10_1));
valve v_10_48 (.fluid_in(k_10_48), .fluid_out(k_9_24), .air_in(c_10_0));
valve v_10_49 (.fluid_in(k_10_49), .fluid_out(k_9_24), .air_in(c_10_1));
valve v_10_50 (.fluid_in(k_10_50), .fluid_out(k_9_25), .air_in(c_10_0));
valve v_10_51 (.fluid_in(k_10_51), .fluid_out(k_9_25), .air_in(c_10_1));
valve v_10_52 (.fluid_in(k_10_52), .fluid_out(k_9_26), .air_in(c_10_0));
valve v_10_53 (.fluid_in(k_10_53), .fluid_out(k_9_26), .air_in(c_10_1));
valve v_10_54 (.fluid_in(k_10_54), .fluid_out(k_9_27), .air_in(c_10_0));
valve v_10_55 (.fluid_in(k_10_55), .fluid_out(k_9_27), .air_in(c_10_1));
valve v_10_56 (.fluid_in(k_10_56), .fluid_out(k_9_28), .air_in(c_10_0));
valve v_10_57 (.fluid_in(k_10_57), .fluid_out(k_9_28), .air_in(c_10_1));
valve v_10_58 (.fluid_in(k_10_58), .fluid_out(k_9_29), .air_in(c_10_0));
valve v_10_59 (.fluid_in(k_10_59), .fluid_out(k_9_29), .air_in(c_10_1));
valve v_10_60 (.fluid_in(k_10_60), .fluid_out(k_9_30), .air_in(c_10_0));
valve v_10_61 (.fluid_in(k_10_61), .fluid_out(k_9_30), .air_in(c_10_1));
valve v_10_62 (.fluid_in(k_10_62), .fluid_out(k_9_31), .air_in(c_10_0));
valve v_10_63 (.fluid_in(k_10_63), .fluid_out(k_9_31), .air_in(c_10_1));
valve v_10_64 (.fluid_in(k_10_64), .fluid_out(k_9_32), .air_in(c_10_0));
valve v_10_65 (.fluid_in(k_10_65), .fluid_out(k_9_32), .air_in(c_10_1));
valve v_10_66 (.fluid_in(k_10_66), .fluid_out(k_9_33), .air_in(c_10_0));
valve v_10_67 (.fluid_in(k_10_67), .fluid_out(k_9_33), .air_in(c_10_1));
valve v_10_68 (.fluid_in(k_10_68), .fluid_out(k_9_34), .air_in(c_10_0));
valve v_10_69 (.fluid_in(k_10_69), .fluid_out(k_9_34), .air_in(c_10_1));
valve v_10_70 (.fluid_in(k_10_70), .fluid_out(k_9_35), .air_in(c_10_0));
valve v_10_71 (.fluid_in(k_10_71), .fluid_out(k_9_35), .air_in(c_10_1));
valve v_10_72 (.fluid_in(k_10_72), .fluid_out(k_9_36), .air_in(c_10_0));
valve v_10_73 (.fluid_in(k_10_73), .fluid_out(k_9_36), .air_in(c_10_1));
valve v_10_74 (.fluid_in(k_10_74), .fluid_out(k_9_37), .air_in(c_10_0));
valve v_10_75 (.fluid_in(k_10_75), .fluid_out(k_9_37), .air_in(c_10_1));
valve v_10_76 (.fluid_in(k_10_76), .fluid_out(k_9_38), .air_in(c_10_0));
valve v_10_77 (.fluid_in(k_10_77), .fluid_out(k_9_38), .air_in(c_10_1));
valve v_10_78 (.fluid_in(k_10_78), .fluid_out(k_9_39), .air_in(c_10_0));
valve v_10_79 (.fluid_in(k_10_79), .fluid_out(k_9_39), .air_in(c_10_1));
valve v_10_80 (.fluid_in(k_10_80), .fluid_out(k_9_40), .air_in(c_10_0));
valve v_10_81 (.fluid_in(k_10_81), .fluid_out(k_9_40), .air_in(c_10_1));
valve v_10_82 (.fluid_in(k_10_82), .fluid_out(k_9_41), .air_in(c_10_0));
valve v_10_83 (.fluid_in(k_10_83), .fluid_out(k_9_41), .air_in(c_10_1));
valve v_10_84 (.fluid_in(k_10_84), .fluid_out(k_9_42), .air_in(c_10_0));
valve v_10_85 (.fluid_in(k_10_85), .fluid_out(k_9_42), .air_in(c_10_1));
valve v_10_86 (.fluid_in(k_10_86), .fluid_out(k_9_43), .air_in(c_10_0));
valve v_10_87 (.fluid_in(k_10_87), .fluid_out(k_9_43), .air_in(c_10_1));
valve v_10_88 (.fluid_in(k_10_88), .fluid_out(k_9_44), .air_in(c_10_0));
valve v_10_89 (.fluid_in(k_10_89), .fluid_out(k_9_44), .air_in(c_10_1));
valve v_10_90 (.fluid_in(k_10_90), .fluid_out(k_9_45), .air_in(c_10_0));
valve v_10_91 (.fluid_in(k_10_91), .fluid_out(k_9_45), .air_in(c_10_1));
valve v_10_92 (.fluid_in(k_10_92), .fluid_out(k_9_46), .air_in(c_10_0));
valve v_10_93 (.fluid_in(k_10_93), .fluid_out(k_9_46), .air_in(c_10_1));
valve v_10_94 (.fluid_in(k_10_94), .fluid_out(k_9_47), .air_in(c_10_0));
valve v_10_95 (.fluid_in(k_10_95), .fluid_out(k_9_47), .air_in(c_10_1));
valve v_10_96 (.fluid_in(k_10_96), .fluid_out(k_9_48), .air_in(c_10_0));
valve v_10_97 (.fluid_in(k_10_97), .fluid_out(k_9_48), .air_in(c_10_1));
valve v_10_98 (.fluid_in(k_10_98), .fluid_out(k_9_49), .air_in(c_10_0));
valve v_10_99 (.fluid_in(k_10_99), .fluid_out(k_9_49), .air_in(c_10_1));
valve v_10_100 (.fluid_in(k_10_100), .fluid_out(k_9_50), .air_in(c_10_0));
valve v_10_101 (.fluid_in(k_10_101), .fluid_out(k_9_50), .air_in(c_10_1));
valve v_10_102 (.fluid_in(k_10_102), .fluid_out(k_9_51), .air_in(c_10_0));
valve v_10_103 (.fluid_in(k_10_103), .fluid_out(k_9_51), .air_in(c_10_1));
valve v_10_104 (.fluid_in(k_10_104), .fluid_out(k_9_52), .air_in(c_10_0));
valve v_10_105 (.fluid_in(k_10_105), .fluid_out(k_9_52), .air_in(c_10_1));
valve v_10_106 (.fluid_in(k_10_106), .fluid_out(k_9_53), .air_in(c_10_0));
valve v_10_107 (.fluid_in(k_10_107), .fluid_out(k_9_53), .air_in(c_10_1));
valve v_10_108 (.fluid_in(k_10_108), .fluid_out(k_9_54), .air_in(c_10_0));
valve v_10_109 (.fluid_in(k_10_109), .fluid_out(k_9_54), .air_in(c_10_1));
valve v_10_110 (.fluid_in(k_10_110), .fluid_out(k_9_55), .air_in(c_10_0));
valve v_10_111 (.fluid_in(k_10_111), .fluid_out(k_9_55), .air_in(c_10_1));
valve v_10_112 (.fluid_in(k_10_112), .fluid_out(k_9_56), .air_in(c_10_0));
valve v_10_113 (.fluid_in(k_10_113), .fluid_out(k_9_56), .air_in(c_10_1));
valve v_10_114 (.fluid_in(k_10_114), .fluid_out(k_9_57), .air_in(c_10_0));
valve v_10_115 (.fluid_in(k_10_115), .fluid_out(k_9_57), .air_in(c_10_1));
valve v_10_116 (.fluid_in(k_10_116), .fluid_out(k_9_58), .air_in(c_10_0));
valve v_10_117 (.fluid_in(k_10_117), .fluid_out(k_9_58), .air_in(c_10_1));
valve v_10_118 (.fluid_in(k_10_118), .fluid_out(k_9_59), .air_in(c_10_0));
valve v_10_119 (.fluid_in(k_10_119), .fluid_out(k_9_59), .air_in(c_10_1));
valve v_10_120 (.fluid_in(k_10_120), .fluid_out(k_9_60), .air_in(c_10_0));
valve v_10_121 (.fluid_in(k_10_121), .fluid_out(k_9_60), .air_in(c_10_1));
valve v_10_122 (.fluid_in(k_10_122), .fluid_out(k_9_61), .air_in(c_10_0));
valve v_10_123 (.fluid_in(k_10_123), .fluid_out(k_9_61), .air_in(c_10_1));
valve v_10_124 (.fluid_in(k_10_124), .fluid_out(k_9_62), .air_in(c_10_0));
valve v_10_125 (.fluid_in(k_10_125), .fluid_out(k_9_62), .air_in(c_10_1));
valve v_10_126 (.fluid_in(k_10_126), .fluid_out(k_9_63), .air_in(c_10_0));
valve v_10_127 (.fluid_in(k_10_127), .fluid_out(k_9_63), .air_in(c_10_1));
valve v_10_128 (.fluid_in(k_10_128), .fluid_out(k_9_64), .air_in(c_10_0));
valve v_10_129 (.fluid_in(k_10_129), .fluid_out(k_9_64), .air_in(c_10_1));
valve v_10_130 (.fluid_in(k_10_130), .fluid_out(k_9_65), .air_in(c_10_0));
valve v_10_131 (.fluid_in(k_10_131), .fluid_out(k_9_65), .air_in(c_10_1));
valve v_10_132 (.fluid_in(k_10_132), .fluid_out(k_9_66), .air_in(c_10_0));
valve v_10_133 (.fluid_in(k_10_133), .fluid_out(k_9_66), .air_in(c_10_1));
valve v_10_134 (.fluid_in(k_10_134), .fluid_out(k_9_67), .air_in(c_10_0));
valve v_10_135 (.fluid_in(k_10_135), .fluid_out(k_9_67), .air_in(c_10_1));
valve v_10_136 (.fluid_in(k_10_136), .fluid_out(k_9_68), .air_in(c_10_0));
valve v_10_137 (.fluid_in(k_10_137), .fluid_out(k_9_68), .air_in(c_10_1));
valve v_10_138 (.fluid_in(k_10_138), .fluid_out(k_9_69), .air_in(c_10_0));
valve v_10_139 (.fluid_in(k_10_139), .fluid_out(k_9_69), .air_in(c_10_1));
valve v_10_140 (.fluid_in(k_10_140), .fluid_out(k_9_70), .air_in(c_10_0));
valve v_10_141 (.fluid_in(k_10_141), .fluid_out(k_9_70), .air_in(c_10_1));
valve v_10_142 (.fluid_in(k_10_142), .fluid_out(k_9_71), .air_in(c_10_0));
valve v_10_143 (.fluid_in(k_10_143), .fluid_out(k_9_71), .air_in(c_10_1));
valve v_10_144 (.fluid_in(k_10_144), .fluid_out(k_9_72), .air_in(c_10_0));
valve v_10_145 (.fluid_in(k_10_145), .fluid_out(k_9_72), .air_in(c_10_1));
valve v_10_146 (.fluid_in(k_10_146), .fluid_out(k_9_73), .air_in(c_10_0));
valve v_10_147 (.fluid_in(k_10_147), .fluid_out(k_9_73), .air_in(c_10_1));
valve v_10_148 (.fluid_in(k_10_148), .fluid_out(k_9_74), .air_in(c_10_0));
valve v_10_149 (.fluid_in(k_10_149), .fluid_out(k_9_74), .air_in(c_10_1));
valve v_10_150 (.fluid_in(k_10_150), .fluid_out(k_9_75), .air_in(c_10_0));
valve v_10_151 (.fluid_in(k_10_151), .fluid_out(k_9_75), .air_in(c_10_1));
valve v_10_152 (.fluid_in(k_10_152), .fluid_out(k_9_76), .air_in(c_10_0));
valve v_10_153 (.fluid_in(k_10_153), .fluid_out(k_9_76), .air_in(c_10_1));
valve v_10_154 (.fluid_in(k_10_154), .fluid_out(k_9_77), .air_in(c_10_0));
valve v_10_155 (.fluid_in(k_10_155), .fluid_out(k_9_77), .air_in(c_10_1));
valve v_10_156 (.fluid_in(k_10_156), .fluid_out(k_9_78), .air_in(c_10_0));
valve v_10_157 (.fluid_in(k_10_157), .fluid_out(k_9_78), .air_in(c_10_1));
valve v_10_158 (.fluid_in(k_10_158), .fluid_out(k_9_79), .air_in(c_10_0));
valve v_10_159 (.fluid_in(k_10_159), .fluid_out(k_9_79), .air_in(c_10_1));
valve v_10_160 (.fluid_in(k_10_160), .fluid_out(k_9_80), .air_in(c_10_0));
valve v_10_161 (.fluid_in(k_10_161), .fluid_out(k_9_80), .air_in(c_10_1));
valve v_10_162 (.fluid_in(k_10_162), .fluid_out(k_9_81), .air_in(c_10_0));
valve v_10_163 (.fluid_in(k_10_163), .fluid_out(k_9_81), .air_in(c_10_1));
valve v_10_164 (.fluid_in(k_10_164), .fluid_out(k_9_82), .air_in(c_10_0));
valve v_10_165 (.fluid_in(k_10_165), .fluid_out(k_9_82), .air_in(c_10_1));
valve v_10_166 (.fluid_in(k_10_166), .fluid_out(k_9_83), .air_in(c_10_0));
valve v_10_167 (.fluid_in(k_10_167), .fluid_out(k_9_83), .air_in(c_10_1));
valve v_10_168 (.fluid_in(k_10_168), .fluid_out(k_9_84), .air_in(c_10_0));
valve v_10_169 (.fluid_in(k_10_169), .fluid_out(k_9_84), .air_in(c_10_1));
valve v_10_170 (.fluid_in(k_10_170), .fluid_out(k_9_85), .air_in(c_10_0));
valve v_10_171 (.fluid_in(k_10_171), .fluid_out(k_9_85), .air_in(c_10_1));
valve v_10_172 (.fluid_in(k_10_172), .fluid_out(k_9_86), .air_in(c_10_0));
valve v_10_173 (.fluid_in(k_10_173), .fluid_out(k_9_86), .air_in(c_10_1));
valve v_10_174 (.fluid_in(k_10_174), .fluid_out(k_9_87), .air_in(c_10_0));
valve v_10_175 (.fluid_in(k_10_175), .fluid_out(k_9_87), .air_in(c_10_1));
valve v_10_176 (.fluid_in(k_10_176), .fluid_out(k_9_88), .air_in(c_10_0));
valve v_10_177 (.fluid_in(k_10_177), .fluid_out(k_9_88), .air_in(c_10_1));
valve v_10_178 (.fluid_in(k_10_178), .fluid_out(k_9_89), .air_in(c_10_0));
valve v_10_179 (.fluid_in(k_10_179), .fluid_out(k_9_89), .air_in(c_10_1));
valve v_10_180 (.fluid_in(k_10_180), .fluid_out(k_9_90), .air_in(c_10_0));
valve v_10_181 (.fluid_in(k_10_181), .fluid_out(k_9_90), .air_in(c_10_1));
valve v_10_182 (.fluid_in(k_10_182), .fluid_out(k_9_91), .air_in(c_10_0));
valve v_10_183 (.fluid_in(k_10_183), .fluid_out(k_9_91), .air_in(c_10_1));
valve v_10_184 (.fluid_in(k_10_184), .fluid_out(k_9_92), .air_in(c_10_0));
valve v_10_185 (.fluid_in(k_10_185), .fluid_out(k_9_92), .air_in(c_10_1));
valve v_10_186 (.fluid_in(k_10_186), .fluid_out(k_9_93), .air_in(c_10_0));
valve v_10_187 (.fluid_in(k_10_187), .fluid_out(k_9_93), .air_in(c_10_1));
valve v_10_188 (.fluid_in(k_10_188), .fluid_out(k_9_94), .air_in(c_10_0));
valve v_10_189 (.fluid_in(k_10_189), .fluid_out(k_9_94), .air_in(c_10_1));
valve v_10_190 (.fluid_in(k_10_190), .fluid_out(k_9_95), .air_in(c_10_0));
valve v_10_191 (.fluid_in(k_10_191), .fluid_out(k_9_95), .air_in(c_10_1));
valve v_10_192 (.fluid_in(k_10_192), .fluid_out(k_9_96), .air_in(c_10_0));
valve v_10_193 (.fluid_in(k_10_193), .fluid_out(k_9_96), .air_in(c_10_1));
valve v_10_194 (.fluid_in(k_10_194), .fluid_out(k_9_97), .air_in(c_10_0));
valve v_10_195 (.fluid_in(k_10_195), .fluid_out(k_9_97), .air_in(c_10_1));
valve v_10_196 (.fluid_in(k_10_196), .fluid_out(k_9_98), .air_in(c_10_0));
valve v_10_197 (.fluid_in(k_10_197), .fluid_out(k_9_98), .air_in(c_10_1));
valve v_10_198 (.fluid_in(k_10_198), .fluid_out(k_9_99), .air_in(c_10_0));
valve v_10_199 (.fluid_in(k_10_199), .fluid_out(k_9_99), .air_in(c_10_1));
valve v_10_200 (.fluid_in(k_10_200), .fluid_out(k_9_100), .air_in(c_10_0));
valve v_10_201 (.fluid_in(k_10_201), .fluid_out(k_9_100), .air_in(c_10_1));
valve v_10_202 (.fluid_in(k_10_202), .fluid_out(k_9_101), .air_in(c_10_0));
valve v_10_203 (.fluid_in(k_10_203), .fluid_out(k_9_101), .air_in(c_10_1));
valve v_10_204 (.fluid_in(k_10_204), .fluid_out(k_9_102), .air_in(c_10_0));
valve v_10_205 (.fluid_in(k_10_205), .fluid_out(k_9_102), .air_in(c_10_1));
valve v_10_206 (.fluid_in(k_10_206), .fluid_out(k_9_103), .air_in(c_10_0));
valve v_10_207 (.fluid_in(k_10_207), .fluid_out(k_9_103), .air_in(c_10_1));
valve v_10_208 (.fluid_in(k_10_208), .fluid_out(k_9_104), .air_in(c_10_0));
valve v_10_209 (.fluid_in(k_10_209), .fluid_out(k_9_104), .air_in(c_10_1));
valve v_10_210 (.fluid_in(k_10_210), .fluid_out(k_9_105), .air_in(c_10_0));
valve v_10_211 (.fluid_in(k_10_211), .fluid_out(k_9_105), .air_in(c_10_1));
valve v_10_212 (.fluid_in(k_10_212), .fluid_out(k_9_106), .air_in(c_10_0));
valve v_10_213 (.fluid_in(k_10_213), .fluid_out(k_9_106), .air_in(c_10_1));
valve v_10_214 (.fluid_in(k_10_214), .fluid_out(k_9_107), .air_in(c_10_0));
valve v_10_215 (.fluid_in(k_10_215), .fluid_out(k_9_107), .air_in(c_10_1));
valve v_10_216 (.fluid_in(k_10_216), .fluid_out(k_9_108), .air_in(c_10_0));
valve v_10_217 (.fluid_in(k_10_217), .fluid_out(k_9_108), .air_in(c_10_1));
valve v_10_218 (.fluid_in(k_10_218), .fluid_out(k_9_109), .air_in(c_10_0));
valve v_10_219 (.fluid_in(k_10_219), .fluid_out(k_9_109), .air_in(c_10_1));
valve v_10_220 (.fluid_in(k_10_220), .fluid_out(k_9_110), .air_in(c_10_0));
valve v_10_221 (.fluid_in(k_10_221), .fluid_out(k_9_110), .air_in(c_10_1));
valve v_10_222 (.fluid_in(k_10_222), .fluid_out(k_9_111), .air_in(c_10_0));
valve v_10_223 (.fluid_in(k_10_223), .fluid_out(k_9_111), .air_in(c_10_1));
valve v_10_224 (.fluid_in(k_10_224), .fluid_out(k_9_112), .air_in(c_10_0));
valve v_10_225 (.fluid_in(k_10_225), .fluid_out(k_9_112), .air_in(c_10_1));
valve v_10_226 (.fluid_in(k_10_226), .fluid_out(k_9_113), .air_in(c_10_0));
valve v_10_227 (.fluid_in(k_10_227), .fluid_out(k_9_113), .air_in(c_10_1));
valve v_10_228 (.fluid_in(k_10_228), .fluid_out(k_9_114), .air_in(c_10_0));
valve v_10_229 (.fluid_in(k_10_229), .fluid_out(k_9_114), .air_in(c_10_1));
valve v_10_230 (.fluid_in(k_10_230), .fluid_out(k_9_115), .air_in(c_10_0));
valve v_10_231 (.fluid_in(k_10_231), .fluid_out(k_9_115), .air_in(c_10_1));
valve v_10_232 (.fluid_in(k_10_232), .fluid_out(k_9_116), .air_in(c_10_0));
valve v_10_233 (.fluid_in(k_10_233), .fluid_out(k_9_116), .air_in(c_10_1));
valve v_10_234 (.fluid_in(k_10_234), .fluid_out(k_9_117), .air_in(c_10_0));
valve v_10_235 (.fluid_in(k_10_235), .fluid_out(k_9_117), .air_in(c_10_1));
valve v_10_236 (.fluid_in(k_10_236), .fluid_out(k_9_118), .air_in(c_10_0));
valve v_10_237 (.fluid_in(k_10_237), .fluid_out(k_9_118), .air_in(c_10_1));
valve v_10_238 (.fluid_in(k_10_238), .fluid_out(k_9_119), .air_in(c_10_0));
valve v_10_239 (.fluid_in(k_10_239), .fluid_out(k_9_119), .air_in(c_10_1));
valve v_10_240 (.fluid_in(k_10_240), .fluid_out(k_9_120), .air_in(c_10_0));
valve v_10_241 (.fluid_in(k_10_241), .fluid_out(k_9_120), .air_in(c_10_1));
valve v_10_242 (.fluid_in(k_10_242), .fluid_out(k_9_121), .air_in(c_10_0));
valve v_10_243 (.fluid_in(k_10_243), .fluid_out(k_9_121), .air_in(c_10_1));
valve v_10_244 (.fluid_in(k_10_244), .fluid_out(k_9_122), .air_in(c_10_0));
valve v_10_245 (.fluid_in(k_10_245), .fluid_out(k_9_122), .air_in(c_10_1));
valve v_10_246 (.fluid_in(k_10_246), .fluid_out(k_9_123), .air_in(c_10_0));
valve v_10_247 (.fluid_in(k_10_247), .fluid_out(k_9_123), .air_in(c_10_1));
valve v_10_248 (.fluid_in(k_10_248), .fluid_out(k_9_124), .air_in(c_10_0));
valve v_10_249 (.fluid_in(k_10_249), .fluid_out(k_9_124), .air_in(c_10_1));
valve v_10_250 (.fluid_in(k_10_250), .fluid_out(k_9_125), .air_in(c_10_0));
valve v_10_251 (.fluid_in(k_10_251), .fluid_out(k_9_125), .air_in(c_10_1));
valve v_10_252 (.fluid_in(k_10_252), .fluid_out(k_9_126), .air_in(c_10_0));
valve v_10_253 (.fluid_in(k_10_253), .fluid_out(k_9_126), .air_in(c_10_1));
valve v_10_254 (.fluid_in(k_10_254), .fluid_out(k_9_127), .air_in(c_10_0));
valve v_10_255 (.fluid_in(k_10_255), .fluid_out(k_9_127), .air_in(c_10_1));
valve v_10_256 (.fluid_in(k_10_256), .fluid_out(k_9_128), .air_in(c_10_0));
valve v_10_257 (.fluid_in(k_10_257), .fluid_out(k_9_128), .air_in(c_10_1));
valve v_10_258 (.fluid_in(k_10_258), .fluid_out(k_9_129), .air_in(c_10_0));
valve v_10_259 (.fluid_in(k_10_259), .fluid_out(k_9_129), .air_in(c_10_1));
valve v_10_260 (.fluid_in(k_10_260), .fluid_out(k_9_130), .air_in(c_10_0));
valve v_10_261 (.fluid_in(k_10_261), .fluid_out(k_9_130), .air_in(c_10_1));
valve v_10_262 (.fluid_in(k_10_262), .fluid_out(k_9_131), .air_in(c_10_0));
valve v_10_263 (.fluid_in(k_10_263), .fluid_out(k_9_131), .air_in(c_10_1));
valve v_10_264 (.fluid_in(k_10_264), .fluid_out(k_9_132), .air_in(c_10_0));
valve v_10_265 (.fluid_in(k_10_265), .fluid_out(k_9_132), .air_in(c_10_1));
valve v_10_266 (.fluid_in(k_10_266), .fluid_out(k_9_133), .air_in(c_10_0));
valve v_10_267 (.fluid_in(k_10_267), .fluid_out(k_9_133), .air_in(c_10_1));
valve v_10_268 (.fluid_in(k_10_268), .fluid_out(k_9_134), .air_in(c_10_0));
valve v_10_269 (.fluid_in(k_10_269), .fluid_out(k_9_134), .air_in(c_10_1));
valve v_10_270 (.fluid_in(k_10_270), .fluid_out(k_9_135), .air_in(c_10_0));
valve v_10_271 (.fluid_in(k_10_271), .fluid_out(k_9_135), .air_in(c_10_1));
valve v_10_272 (.fluid_in(k_10_272), .fluid_out(k_9_136), .air_in(c_10_0));
valve v_10_273 (.fluid_in(k_10_273), .fluid_out(k_9_136), .air_in(c_10_1));
valve v_10_274 (.fluid_in(k_10_274), .fluid_out(k_9_137), .air_in(c_10_0));
valve v_10_275 (.fluid_in(k_10_275), .fluid_out(k_9_137), .air_in(c_10_1));
valve v_10_276 (.fluid_in(k_10_276), .fluid_out(k_9_138), .air_in(c_10_0));
valve v_10_277 (.fluid_in(k_10_277), .fluid_out(k_9_138), .air_in(c_10_1));
valve v_10_278 (.fluid_in(k_10_278), .fluid_out(k_9_139), .air_in(c_10_0));
valve v_10_279 (.fluid_in(k_10_279), .fluid_out(k_9_139), .air_in(c_10_1));
valve v_10_280 (.fluid_in(k_10_280), .fluid_out(k_9_140), .air_in(c_10_0));
valve v_10_281 (.fluid_in(k_10_281), .fluid_out(k_9_140), .air_in(c_10_1));
valve v_10_282 (.fluid_in(k_10_282), .fluid_out(k_9_141), .air_in(c_10_0));
valve v_10_283 (.fluid_in(k_10_283), .fluid_out(k_9_141), .air_in(c_10_1));
valve v_10_284 (.fluid_in(k_10_284), .fluid_out(k_9_142), .air_in(c_10_0));
valve v_10_285 (.fluid_in(k_10_285), .fluid_out(k_9_142), .air_in(c_10_1));
valve v_10_286 (.fluid_in(k_10_286), .fluid_out(k_9_143), .air_in(c_10_0));
valve v_10_287 (.fluid_in(k_10_287), .fluid_out(k_9_143), .air_in(c_10_1));
valve v_10_288 (.fluid_in(k_10_288), .fluid_out(k_9_144), .air_in(c_10_0));
valve v_10_289 (.fluid_in(k_10_289), .fluid_out(k_9_144), .air_in(c_10_1));
valve v_10_290 (.fluid_in(k_10_290), .fluid_out(k_9_145), .air_in(c_10_0));
valve v_10_291 (.fluid_in(k_10_291), .fluid_out(k_9_145), .air_in(c_10_1));
valve v_10_292 (.fluid_in(k_10_292), .fluid_out(k_9_146), .air_in(c_10_0));
valve v_10_293 (.fluid_in(k_10_293), .fluid_out(k_9_146), .air_in(c_10_1));
valve v_10_294 (.fluid_in(k_10_294), .fluid_out(k_9_147), .air_in(c_10_0));
valve v_10_295 (.fluid_in(k_10_295), .fluid_out(k_9_147), .air_in(c_10_1));
valve v_10_296 (.fluid_in(k_10_296), .fluid_out(k_9_148), .air_in(c_10_0));
valve v_10_297 (.fluid_in(k_10_297), .fluid_out(k_9_148), .air_in(c_10_1));
valve v_10_298 (.fluid_in(k_10_298), .fluid_out(k_9_149), .air_in(c_10_0));
valve v_10_299 (.fluid_in(k_10_299), .fluid_out(k_9_149), .air_in(c_10_1));
valve v_10_300 (.fluid_in(k_10_300), .fluid_out(k_9_150), .air_in(c_10_0));
valve v_10_301 (.fluid_in(k_10_301), .fluid_out(k_9_150), .air_in(c_10_1));
valve v_10_302 (.fluid_in(k_10_302), .fluid_out(k_9_151), .air_in(c_10_0));
valve v_10_303 (.fluid_in(k_10_303), .fluid_out(k_9_151), .air_in(c_10_1));
valve v_10_304 (.fluid_in(k_10_304), .fluid_out(k_9_152), .air_in(c_10_0));
valve v_10_305 (.fluid_in(k_10_305), .fluid_out(k_9_152), .air_in(c_10_1));
valve v_10_306 (.fluid_in(k_10_306), .fluid_out(k_9_153), .air_in(c_10_0));
valve v_10_307 (.fluid_in(k_10_307), .fluid_out(k_9_153), .air_in(c_10_1));
valve v_10_308 (.fluid_in(k_10_308), .fluid_out(k_9_154), .air_in(c_10_0));
valve v_10_309 (.fluid_in(k_10_309), .fluid_out(k_9_154), .air_in(c_10_1));
valve v_10_310 (.fluid_in(k_10_310), .fluid_out(k_9_155), .air_in(c_10_0));
valve v_10_311 (.fluid_in(k_10_311), .fluid_out(k_9_155), .air_in(c_10_1));
valve v_10_312 (.fluid_in(k_10_312), .fluid_out(k_9_156), .air_in(c_10_0));
valve v_10_313 (.fluid_in(k_10_313), .fluid_out(k_9_156), .air_in(c_10_1));
valve v_10_314 (.fluid_in(k_10_314), .fluid_out(k_9_157), .air_in(c_10_0));
valve v_10_315 (.fluid_in(k_10_315), .fluid_out(k_9_157), .air_in(c_10_1));
valve v_10_316 (.fluid_in(k_10_316), .fluid_out(k_9_158), .air_in(c_10_0));
valve v_10_317 (.fluid_in(k_10_317), .fluid_out(k_9_158), .air_in(c_10_1));
valve v_10_318 (.fluid_in(k_10_318), .fluid_out(k_9_159), .air_in(c_10_0));
valve v_10_319 (.fluid_in(k_10_319), .fluid_out(k_9_159), .air_in(c_10_1));
valve v_10_320 (.fluid_in(k_10_320), .fluid_out(k_9_160), .air_in(c_10_0));
valve v_10_321 (.fluid_in(k_10_321), .fluid_out(k_9_160), .air_in(c_10_1));
valve v_10_322 (.fluid_in(k_10_322), .fluid_out(k_9_161), .air_in(c_10_0));
valve v_10_323 (.fluid_in(k_10_323), .fluid_out(k_9_161), .air_in(c_10_1));
valve v_10_324 (.fluid_in(k_10_324), .fluid_out(k_9_162), .air_in(c_10_0));
valve v_10_325 (.fluid_in(k_10_325), .fluid_out(k_9_162), .air_in(c_10_1));
valve v_10_326 (.fluid_in(k_10_326), .fluid_out(k_9_163), .air_in(c_10_0));
valve v_10_327 (.fluid_in(k_10_327), .fluid_out(k_9_163), .air_in(c_10_1));
valve v_10_328 (.fluid_in(k_10_328), .fluid_out(k_9_164), .air_in(c_10_0));
valve v_10_329 (.fluid_in(k_10_329), .fluid_out(k_9_164), .air_in(c_10_1));
valve v_10_330 (.fluid_in(k_10_330), .fluid_out(k_9_165), .air_in(c_10_0));
valve v_10_331 (.fluid_in(k_10_331), .fluid_out(k_9_165), .air_in(c_10_1));
valve v_10_332 (.fluid_in(k_10_332), .fluid_out(k_9_166), .air_in(c_10_0));
valve v_10_333 (.fluid_in(k_10_333), .fluid_out(k_9_166), .air_in(c_10_1));
valve v_10_334 (.fluid_in(k_10_334), .fluid_out(k_9_167), .air_in(c_10_0));
valve v_10_335 (.fluid_in(k_10_335), .fluid_out(k_9_167), .air_in(c_10_1));
valve v_10_336 (.fluid_in(k_10_336), .fluid_out(k_9_168), .air_in(c_10_0));
valve v_10_337 (.fluid_in(k_10_337), .fluid_out(k_9_168), .air_in(c_10_1));
valve v_10_338 (.fluid_in(k_10_338), .fluid_out(k_9_169), .air_in(c_10_0));
valve v_10_339 (.fluid_in(k_10_339), .fluid_out(k_9_169), .air_in(c_10_1));
valve v_10_340 (.fluid_in(k_10_340), .fluid_out(k_9_170), .air_in(c_10_0));
valve v_10_341 (.fluid_in(k_10_341), .fluid_out(k_9_170), .air_in(c_10_1));
valve v_10_342 (.fluid_in(k_10_342), .fluid_out(k_9_171), .air_in(c_10_0));
valve v_10_343 (.fluid_in(k_10_343), .fluid_out(k_9_171), .air_in(c_10_1));
valve v_10_344 (.fluid_in(k_10_344), .fluid_out(k_9_172), .air_in(c_10_0));
valve v_10_345 (.fluid_in(k_10_345), .fluid_out(k_9_172), .air_in(c_10_1));
valve v_10_346 (.fluid_in(k_10_346), .fluid_out(k_9_173), .air_in(c_10_0));
valve v_10_347 (.fluid_in(k_10_347), .fluid_out(k_9_173), .air_in(c_10_1));
valve v_10_348 (.fluid_in(k_10_348), .fluid_out(k_9_174), .air_in(c_10_0));
valve v_10_349 (.fluid_in(k_10_349), .fluid_out(k_9_174), .air_in(c_10_1));
valve v_10_350 (.fluid_in(k_10_350), .fluid_out(k_9_175), .air_in(c_10_0));
valve v_10_351 (.fluid_in(k_10_351), .fluid_out(k_9_175), .air_in(c_10_1));
valve v_10_352 (.fluid_in(k_10_352), .fluid_out(k_9_176), .air_in(c_10_0));
valve v_10_353 (.fluid_in(k_10_353), .fluid_out(k_9_176), .air_in(c_10_1));
valve v_10_354 (.fluid_in(k_10_354), .fluid_out(k_9_177), .air_in(c_10_0));
valve v_10_355 (.fluid_in(k_10_355), .fluid_out(k_9_177), .air_in(c_10_1));
valve v_10_356 (.fluid_in(k_10_356), .fluid_out(k_9_178), .air_in(c_10_0));
valve v_10_357 (.fluid_in(k_10_357), .fluid_out(k_9_178), .air_in(c_10_1));
valve v_10_358 (.fluid_in(k_10_358), .fluid_out(k_9_179), .air_in(c_10_0));
valve v_10_359 (.fluid_in(k_10_359), .fluid_out(k_9_179), .air_in(c_10_1));
valve v_10_360 (.fluid_in(k_10_360), .fluid_out(k_9_180), .air_in(c_10_0));
valve v_10_361 (.fluid_in(k_10_361), .fluid_out(k_9_180), .air_in(c_10_1));
valve v_10_362 (.fluid_in(k_10_362), .fluid_out(k_9_181), .air_in(c_10_0));
valve v_10_363 (.fluid_in(k_10_363), .fluid_out(k_9_181), .air_in(c_10_1));
valve v_10_364 (.fluid_in(k_10_364), .fluid_out(k_9_182), .air_in(c_10_0));
valve v_10_365 (.fluid_in(k_10_365), .fluid_out(k_9_182), .air_in(c_10_1));
valve v_10_366 (.fluid_in(k_10_366), .fluid_out(k_9_183), .air_in(c_10_0));
valve v_10_367 (.fluid_in(k_10_367), .fluid_out(k_9_183), .air_in(c_10_1));
valve v_10_368 (.fluid_in(k_10_368), .fluid_out(k_9_184), .air_in(c_10_0));
valve v_10_369 (.fluid_in(k_10_369), .fluid_out(k_9_184), .air_in(c_10_1));
valve v_10_370 (.fluid_in(k_10_370), .fluid_out(k_9_185), .air_in(c_10_0));
valve v_10_371 (.fluid_in(k_10_371), .fluid_out(k_9_185), .air_in(c_10_1));
valve v_10_372 (.fluid_in(k_10_372), .fluid_out(k_9_186), .air_in(c_10_0));
valve v_10_373 (.fluid_in(k_10_373), .fluid_out(k_9_186), .air_in(c_10_1));
valve v_10_374 (.fluid_in(k_10_374), .fluid_out(k_9_187), .air_in(c_10_0));
valve v_10_375 (.fluid_in(k_10_375), .fluid_out(k_9_187), .air_in(c_10_1));
valve v_10_376 (.fluid_in(k_10_376), .fluid_out(k_9_188), .air_in(c_10_0));
valve v_10_377 (.fluid_in(k_10_377), .fluid_out(k_9_188), .air_in(c_10_1));
valve v_10_378 (.fluid_in(k_10_378), .fluid_out(k_9_189), .air_in(c_10_0));
valve v_10_379 (.fluid_in(k_10_379), .fluid_out(k_9_189), .air_in(c_10_1));
valve v_10_380 (.fluid_in(k_10_380), .fluid_out(k_9_190), .air_in(c_10_0));
valve v_10_381 (.fluid_in(k_10_381), .fluid_out(k_9_190), .air_in(c_10_1));
valve v_10_382 (.fluid_in(k_10_382), .fluid_out(k_9_191), .air_in(c_10_0));
valve v_10_383 (.fluid_in(k_10_383), .fluid_out(k_9_191), .air_in(c_10_1));
valve v_10_384 (.fluid_in(k_10_384), .fluid_out(k_9_192), .air_in(c_10_0));
valve v_10_385 (.fluid_in(k_10_385), .fluid_out(k_9_192), .air_in(c_10_1));
valve v_10_386 (.fluid_in(k_10_386), .fluid_out(k_9_193), .air_in(c_10_0));
valve v_10_387 (.fluid_in(k_10_387), .fluid_out(k_9_193), .air_in(c_10_1));
valve v_10_388 (.fluid_in(k_10_388), .fluid_out(k_9_194), .air_in(c_10_0));
valve v_10_389 (.fluid_in(k_10_389), .fluid_out(k_9_194), .air_in(c_10_1));
valve v_10_390 (.fluid_in(k_10_390), .fluid_out(k_9_195), .air_in(c_10_0));
valve v_10_391 (.fluid_in(k_10_391), .fluid_out(k_9_195), .air_in(c_10_1));
valve v_10_392 (.fluid_in(k_10_392), .fluid_out(k_9_196), .air_in(c_10_0));
valve v_10_393 (.fluid_in(k_10_393), .fluid_out(k_9_196), .air_in(c_10_1));
valve v_10_394 (.fluid_in(k_10_394), .fluid_out(k_9_197), .air_in(c_10_0));
valve v_10_395 (.fluid_in(k_10_395), .fluid_out(k_9_197), .air_in(c_10_1));
valve v_10_396 (.fluid_in(k_10_396), .fluid_out(k_9_198), .air_in(c_10_0));
valve v_10_397 (.fluid_in(k_10_397), .fluid_out(k_9_198), .air_in(c_10_1));
valve v_10_398 (.fluid_in(k_10_398), .fluid_out(k_9_199), .air_in(c_10_0));
valve v_10_399 (.fluid_in(k_10_399), .fluid_out(k_9_199), .air_in(c_10_1));
valve v_10_400 (.fluid_in(k_10_400), .fluid_out(k_9_200), .air_in(c_10_0));
valve v_10_401 (.fluid_in(k_10_401), .fluid_out(k_9_200), .air_in(c_10_1));
valve v_10_402 (.fluid_in(k_10_402), .fluid_out(k_9_201), .air_in(c_10_0));
valve v_10_403 (.fluid_in(k_10_403), .fluid_out(k_9_201), .air_in(c_10_1));
valve v_10_404 (.fluid_in(k_10_404), .fluid_out(k_9_202), .air_in(c_10_0));
valve v_10_405 (.fluid_in(k_10_405), .fluid_out(k_9_202), .air_in(c_10_1));
valve v_10_406 (.fluid_in(k_10_406), .fluid_out(k_9_203), .air_in(c_10_0));
valve v_10_407 (.fluid_in(k_10_407), .fluid_out(k_9_203), .air_in(c_10_1));
valve v_10_408 (.fluid_in(k_10_408), .fluid_out(k_9_204), .air_in(c_10_0));
valve v_10_409 (.fluid_in(k_10_409), .fluid_out(k_9_204), .air_in(c_10_1));
valve v_10_410 (.fluid_in(k_10_410), .fluid_out(k_9_205), .air_in(c_10_0));
valve v_10_411 (.fluid_in(k_10_411), .fluid_out(k_9_205), .air_in(c_10_1));
valve v_10_412 (.fluid_in(k_10_412), .fluid_out(k_9_206), .air_in(c_10_0));
valve v_10_413 (.fluid_in(k_10_413), .fluid_out(k_9_206), .air_in(c_10_1));
valve v_10_414 (.fluid_in(k_10_414), .fluid_out(k_9_207), .air_in(c_10_0));
valve v_10_415 (.fluid_in(k_10_415), .fluid_out(k_9_207), .air_in(c_10_1));
valve v_10_416 (.fluid_in(k_10_416), .fluid_out(k_9_208), .air_in(c_10_0));
valve v_10_417 (.fluid_in(k_10_417), .fluid_out(k_9_208), .air_in(c_10_1));
valve v_10_418 (.fluid_in(k_10_418), .fluid_out(k_9_209), .air_in(c_10_0));
valve v_10_419 (.fluid_in(k_10_419), .fluid_out(k_9_209), .air_in(c_10_1));
valve v_10_420 (.fluid_in(k_10_420), .fluid_out(k_9_210), .air_in(c_10_0));
valve v_10_421 (.fluid_in(k_10_421), .fluid_out(k_9_210), .air_in(c_10_1));
valve v_10_422 (.fluid_in(k_10_422), .fluid_out(k_9_211), .air_in(c_10_0));
valve v_10_423 (.fluid_in(k_10_423), .fluid_out(k_9_211), .air_in(c_10_1));
valve v_10_424 (.fluid_in(k_10_424), .fluid_out(k_9_212), .air_in(c_10_0));
valve v_10_425 (.fluid_in(k_10_425), .fluid_out(k_9_212), .air_in(c_10_1));
valve v_10_426 (.fluid_in(k_10_426), .fluid_out(k_9_213), .air_in(c_10_0));
valve v_10_427 (.fluid_in(k_10_427), .fluid_out(k_9_213), .air_in(c_10_1));
valve v_10_428 (.fluid_in(k_10_428), .fluid_out(k_9_214), .air_in(c_10_0));
valve v_10_429 (.fluid_in(k_10_429), .fluid_out(k_9_214), .air_in(c_10_1));
valve v_10_430 (.fluid_in(k_10_430), .fluid_out(k_9_215), .air_in(c_10_0));
valve v_10_431 (.fluid_in(k_10_431), .fluid_out(k_9_215), .air_in(c_10_1));
valve v_10_432 (.fluid_in(k_10_432), .fluid_out(k_9_216), .air_in(c_10_0));
valve v_10_433 (.fluid_in(k_10_433), .fluid_out(k_9_216), .air_in(c_10_1));
valve v_10_434 (.fluid_in(k_10_434), .fluid_out(k_9_217), .air_in(c_10_0));
valve v_10_435 (.fluid_in(k_10_435), .fluid_out(k_9_217), .air_in(c_10_1));
valve v_10_436 (.fluid_in(k_10_436), .fluid_out(k_9_218), .air_in(c_10_0));
valve v_10_437 (.fluid_in(k_10_437), .fluid_out(k_9_218), .air_in(c_10_1));
valve v_10_438 (.fluid_in(k_10_438), .fluid_out(k_9_219), .air_in(c_10_0));
valve v_10_439 (.fluid_in(k_10_439), .fluid_out(k_9_219), .air_in(c_10_1));
valve v_10_440 (.fluid_in(k_10_440), .fluid_out(k_9_220), .air_in(c_10_0));
valve v_10_441 (.fluid_in(k_10_441), .fluid_out(k_9_220), .air_in(c_10_1));
valve v_10_442 (.fluid_in(k_10_442), .fluid_out(k_9_221), .air_in(c_10_0));
valve v_10_443 (.fluid_in(k_10_443), .fluid_out(k_9_221), .air_in(c_10_1));
valve v_10_444 (.fluid_in(k_10_444), .fluid_out(k_9_222), .air_in(c_10_0));
valve v_10_445 (.fluid_in(k_10_445), .fluid_out(k_9_222), .air_in(c_10_1));
valve v_10_446 (.fluid_in(k_10_446), .fluid_out(k_9_223), .air_in(c_10_0));
valve v_10_447 (.fluid_in(k_10_447), .fluid_out(k_9_223), .air_in(c_10_1));
valve v_10_448 (.fluid_in(k_10_448), .fluid_out(k_9_224), .air_in(c_10_0));
valve v_10_449 (.fluid_in(k_10_449), .fluid_out(k_9_224), .air_in(c_10_1));
valve v_10_450 (.fluid_in(k_10_450), .fluid_out(k_9_225), .air_in(c_10_0));
valve v_10_451 (.fluid_in(k_10_451), .fluid_out(k_9_225), .air_in(c_10_1));
valve v_10_452 (.fluid_in(k_10_452), .fluid_out(k_9_226), .air_in(c_10_0));
valve v_10_453 (.fluid_in(k_10_453), .fluid_out(k_9_226), .air_in(c_10_1));
valve v_10_454 (.fluid_in(k_10_454), .fluid_out(k_9_227), .air_in(c_10_0));
valve v_10_455 (.fluid_in(k_10_455), .fluid_out(k_9_227), .air_in(c_10_1));
valve v_10_456 (.fluid_in(k_10_456), .fluid_out(k_9_228), .air_in(c_10_0));
valve v_10_457 (.fluid_in(k_10_457), .fluid_out(k_9_228), .air_in(c_10_1));
valve v_10_458 (.fluid_in(k_10_458), .fluid_out(k_9_229), .air_in(c_10_0));
valve v_10_459 (.fluid_in(k_10_459), .fluid_out(k_9_229), .air_in(c_10_1));
valve v_10_460 (.fluid_in(k_10_460), .fluid_out(k_9_230), .air_in(c_10_0));
valve v_10_461 (.fluid_in(k_10_461), .fluid_out(k_9_230), .air_in(c_10_1));
valve v_10_462 (.fluid_in(k_10_462), .fluid_out(k_9_231), .air_in(c_10_0));
valve v_10_463 (.fluid_in(k_10_463), .fluid_out(k_9_231), .air_in(c_10_1));
valve v_10_464 (.fluid_in(k_10_464), .fluid_out(k_9_232), .air_in(c_10_0));
valve v_10_465 (.fluid_in(k_10_465), .fluid_out(k_9_232), .air_in(c_10_1));
valve v_10_466 (.fluid_in(k_10_466), .fluid_out(k_9_233), .air_in(c_10_0));
valve v_10_467 (.fluid_in(k_10_467), .fluid_out(k_9_233), .air_in(c_10_1));
valve v_10_468 (.fluid_in(k_10_468), .fluid_out(k_9_234), .air_in(c_10_0));
valve v_10_469 (.fluid_in(k_10_469), .fluid_out(k_9_234), .air_in(c_10_1));
valve v_10_470 (.fluid_in(k_10_470), .fluid_out(k_9_235), .air_in(c_10_0));
valve v_10_471 (.fluid_in(k_10_471), .fluid_out(k_9_235), .air_in(c_10_1));
valve v_10_472 (.fluid_in(k_10_472), .fluid_out(k_9_236), .air_in(c_10_0));
valve v_10_473 (.fluid_in(k_10_473), .fluid_out(k_9_236), .air_in(c_10_1));
valve v_10_474 (.fluid_in(k_10_474), .fluid_out(k_9_237), .air_in(c_10_0));
valve v_10_475 (.fluid_in(k_10_475), .fluid_out(k_9_237), .air_in(c_10_1));
valve v_10_476 (.fluid_in(k_10_476), .fluid_out(k_9_238), .air_in(c_10_0));
valve v_10_477 (.fluid_in(k_10_477), .fluid_out(k_9_238), .air_in(c_10_1));
valve v_10_478 (.fluid_in(k_10_478), .fluid_out(k_9_239), .air_in(c_10_0));
valve v_10_479 (.fluid_in(k_10_479), .fluid_out(k_9_239), .air_in(c_10_1));
valve v_10_480 (.fluid_in(k_10_480), .fluid_out(k_9_240), .air_in(c_10_0));
valve v_10_481 (.fluid_in(k_10_481), .fluid_out(k_9_240), .air_in(c_10_1));
valve v_10_482 (.fluid_in(k_10_482), .fluid_out(k_9_241), .air_in(c_10_0));
valve v_10_483 (.fluid_in(k_10_483), .fluid_out(k_9_241), .air_in(c_10_1));
valve v_10_484 (.fluid_in(k_10_484), .fluid_out(k_9_242), .air_in(c_10_0));
valve v_10_485 (.fluid_in(k_10_485), .fluid_out(k_9_242), .air_in(c_10_1));
valve v_10_486 (.fluid_in(k_10_486), .fluid_out(k_9_243), .air_in(c_10_0));
valve v_10_487 (.fluid_in(k_10_487), .fluid_out(k_9_243), .air_in(c_10_1));
valve v_10_488 (.fluid_in(k_10_488), .fluid_out(k_9_244), .air_in(c_10_0));
valve v_10_489 (.fluid_in(k_10_489), .fluid_out(k_9_244), .air_in(c_10_1));
valve v_10_490 (.fluid_in(k_10_490), .fluid_out(k_9_245), .air_in(c_10_0));
valve v_10_491 (.fluid_in(k_10_491), .fluid_out(k_9_245), .air_in(c_10_1));
valve v_10_492 (.fluid_in(k_10_492), .fluid_out(k_9_246), .air_in(c_10_0));
valve v_10_493 (.fluid_in(k_10_493), .fluid_out(k_9_246), .air_in(c_10_1));
valve v_10_494 (.fluid_in(k_10_494), .fluid_out(k_9_247), .air_in(c_10_0));
valve v_10_495 (.fluid_in(k_10_495), .fluid_out(k_9_247), .air_in(c_10_1));
valve v_10_496 (.fluid_in(k_10_496), .fluid_out(k_9_248), .air_in(c_10_0));
valve v_10_497 (.fluid_in(k_10_497), .fluid_out(k_9_248), .air_in(c_10_1));
valve v_10_498 (.fluid_in(k_10_498), .fluid_out(k_9_249), .air_in(c_10_0));
valve v_10_499 (.fluid_in(k_10_499), .fluid_out(k_9_249), .air_in(c_10_1));
valve v_10_500 (.fluid_in(k_10_500), .fluid_out(k_9_250), .air_in(c_10_0));
valve v_10_501 (.fluid_in(k_10_501), .fluid_out(k_9_250), .air_in(c_10_1));
valve v_10_502 (.fluid_in(k_10_502), .fluid_out(k_9_251), .air_in(c_10_0));
valve v_10_503 (.fluid_in(k_10_503), .fluid_out(k_9_251), .air_in(c_10_1));
valve v_10_504 (.fluid_in(k_10_504), .fluid_out(k_9_252), .air_in(c_10_0));
valve v_10_505 (.fluid_in(k_10_505), .fluid_out(k_9_252), .air_in(c_10_1));
valve v_10_506 (.fluid_in(k_10_506), .fluid_out(k_9_253), .air_in(c_10_0));
valve v_10_507 (.fluid_in(k_10_507), .fluid_out(k_9_253), .air_in(c_10_1));
valve v_10_508 (.fluid_in(k_10_508), .fluid_out(k_9_254), .air_in(c_10_0));
valve v_10_509 (.fluid_in(k_10_509), .fluid_out(k_9_254), .air_in(c_10_1));
valve v_10_510 (.fluid_in(k_10_510), .fluid_out(k_9_255), .air_in(c_10_0));
valve v_10_511 (.fluid_in(k_10_511), .fluid_out(k_9_255), .air_in(c_10_1));
valve v_10_512 (.fluid_in(k_10_512), .fluid_out(k_9_256), .air_in(c_10_0));
valve v_10_513 (.fluid_in(k_10_513), .fluid_out(k_9_256), .air_in(c_10_1));
valve v_10_514 (.fluid_in(k_10_514), .fluid_out(k_9_257), .air_in(c_10_0));
valve v_10_515 (.fluid_in(k_10_515), .fluid_out(k_9_257), .air_in(c_10_1));
valve v_10_516 (.fluid_in(k_10_516), .fluid_out(k_9_258), .air_in(c_10_0));
valve v_10_517 (.fluid_in(k_10_517), .fluid_out(k_9_258), .air_in(c_10_1));
valve v_10_518 (.fluid_in(k_10_518), .fluid_out(k_9_259), .air_in(c_10_0));
valve v_10_519 (.fluid_in(k_10_519), .fluid_out(k_9_259), .air_in(c_10_1));
valve v_10_520 (.fluid_in(k_10_520), .fluid_out(k_9_260), .air_in(c_10_0));
valve v_10_521 (.fluid_in(k_10_521), .fluid_out(k_9_260), .air_in(c_10_1));
valve v_10_522 (.fluid_in(k_10_522), .fluid_out(k_9_261), .air_in(c_10_0));
valve v_10_523 (.fluid_in(k_10_523), .fluid_out(k_9_261), .air_in(c_10_1));
valve v_10_524 (.fluid_in(k_10_524), .fluid_out(k_9_262), .air_in(c_10_0));
valve v_10_525 (.fluid_in(k_10_525), .fluid_out(k_9_262), .air_in(c_10_1));
valve v_10_526 (.fluid_in(k_10_526), .fluid_out(k_9_263), .air_in(c_10_0));
valve v_10_527 (.fluid_in(k_10_527), .fluid_out(k_9_263), .air_in(c_10_1));
valve v_10_528 (.fluid_in(k_10_528), .fluid_out(k_9_264), .air_in(c_10_0));
valve v_10_529 (.fluid_in(k_10_529), .fluid_out(k_9_264), .air_in(c_10_1));
valve v_10_530 (.fluid_in(k_10_530), .fluid_out(k_9_265), .air_in(c_10_0));
valve v_10_531 (.fluid_in(k_10_531), .fluid_out(k_9_265), .air_in(c_10_1));
valve v_10_532 (.fluid_in(k_10_532), .fluid_out(k_9_266), .air_in(c_10_0));
valve v_10_533 (.fluid_in(k_10_533), .fluid_out(k_9_266), .air_in(c_10_1));
valve v_10_534 (.fluid_in(k_10_534), .fluid_out(k_9_267), .air_in(c_10_0));
valve v_10_535 (.fluid_in(k_10_535), .fluid_out(k_9_267), .air_in(c_10_1));
valve v_10_536 (.fluid_in(k_10_536), .fluid_out(k_9_268), .air_in(c_10_0));
valve v_10_537 (.fluid_in(k_10_537), .fluid_out(k_9_268), .air_in(c_10_1));
valve v_10_538 (.fluid_in(k_10_538), .fluid_out(k_9_269), .air_in(c_10_0));
valve v_10_539 (.fluid_in(k_10_539), .fluid_out(k_9_269), .air_in(c_10_1));
valve v_10_540 (.fluid_in(k_10_540), .fluid_out(k_9_270), .air_in(c_10_0));
valve v_10_541 (.fluid_in(k_10_541), .fluid_out(k_9_270), .air_in(c_10_1));
valve v_10_542 (.fluid_in(k_10_542), .fluid_out(k_9_271), .air_in(c_10_0));
valve v_10_543 (.fluid_in(k_10_543), .fluid_out(k_9_271), .air_in(c_10_1));
valve v_10_544 (.fluid_in(k_10_544), .fluid_out(k_9_272), .air_in(c_10_0));
valve v_10_545 (.fluid_in(k_10_545), .fluid_out(k_9_272), .air_in(c_10_1));
valve v_10_546 (.fluid_in(k_10_546), .fluid_out(k_9_273), .air_in(c_10_0));
valve v_10_547 (.fluid_in(k_10_547), .fluid_out(k_9_273), .air_in(c_10_1));
valve v_10_548 (.fluid_in(k_10_548), .fluid_out(k_9_274), .air_in(c_10_0));
valve v_10_549 (.fluid_in(k_10_549), .fluid_out(k_9_274), .air_in(c_10_1));
valve v_10_550 (.fluid_in(k_10_550), .fluid_out(k_9_275), .air_in(c_10_0));
valve v_10_551 (.fluid_in(k_10_551), .fluid_out(k_9_275), .air_in(c_10_1));
valve v_10_552 (.fluid_in(k_10_552), .fluid_out(k_9_276), .air_in(c_10_0));
valve v_10_553 (.fluid_in(k_10_553), .fluid_out(k_9_276), .air_in(c_10_1));
valve v_10_554 (.fluid_in(k_10_554), .fluid_out(k_9_277), .air_in(c_10_0));
valve v_10_555 (.fluid_in(k_10_555), .fluid_out(k_9_277), .air_in(c_10_1));
valve v_10_556 (.fluid_in(k_10_556), .fluid_out(k_9_278), .air_in(c_10_0));
valve v_10_557 (.fluid_in(k_10_557), .fluid_out(k_9_278), .air_in(c_10_1));
valve v_10_558 (.fluid_in(k_10_558), .fluid_out(k_9_279), .air_in(c_10_0));
valve v_10_559 (.fluid_in(k_10_559), .fluid_out(k_9_279), .air_in(c_10_1));
valve v_10_560 (.fluid_in(k_10_560), .fluid_out(k_9_280), .air_in(c_10_0));
valve v_10_561 (.fluid_in(k_10_561), .fluid_out(k_9_280), .air_in(c_10_1));
valve v_10_562 (.fluid_in(k_10_562), .fluid_out(k_9_281), .air_in(c_10_0));
valve v_10_563 (.fluid_in(k_10_563), .fluid_out(k_9_281), .air_in(c_10_1));
valve v_10_564 (.fluid_in(k_10_564), .fluid_out(k_9_282), .air_in(c_10_0));
valve v_10_565 (.fluid_in(k_10_565), .fluid_out(k_9_282), .air_in(c_10_1));
valve v_10_566 (.fluid_in(k_10_566), .fluid_out(k_9_283), .air_in(c_10_0));
valve v_10_567 (.fluid_in(k_10_567), .fluid_out(k_9_283), .air_in(c_10_1));
valve v_10_568 (.fluid_in(k_10_568), .fluid_out(k_9_284), .air_in(c_10_0));
valve v_10_569 (.fluid_in(k_10_569), .fluid_out(k_9_284), .air_in(c_10_1));
valve v_10_570 (.fluid_in(k_10_570), .fluid_out(k_9_285), .air_in(c_10_0));
valve v_10_571 (.fluid_in(k_10_571), .fluid_out(k_9_285), .air_in(c_10_1));
valve v_10_572 (.fluid_in(k_10_572), .fluid_out(k_9_286), .air_in(c_10_0));
valve v_10_573 (.fluid_in(k_10_573), .fluid_out(k_9_286), .air_in(c_10_1));
valve v_10_574 (.fluid_in(k_10_574), .fluid_out(k_9_287), .air_in(c_10_0));
valve v_10_575 (.fluid_in(k_10_575), .fluid_out(k_9_287), .air_in(c_10_1));
valve v_10_576 (.fluid_in(k_10_576), .fluid_out(k_9_288), .air_in(c_10_0));
valve v_10_577 (.fluid_in(k_10_577), .fluid_out(k_9_288), .air_in(c_10_1));
valve v_10_578 (.fluid_in(k_10_578), .fluid_out(k_9_289), .air_in(c_10_0));
valve v_10_579 (.fluid_in(k_10_579), .fluid_out(k_9_289), .air_in(c_10_1));
valve v_10_580 (.fluid_in(k_10_580), .fluid_out(k_9_290), .air_in(c_10_0));
valve v_10_581 (.fluid_in(k_10_581), .fluid_out(k_9_290), .air_in(c_10_1));
valve v_10_582 (.fluid_in(k_10_582), .fluid_out(k_9_291), .air_in(c_10_0));
valve v_10_583 (.fluid_in(k_10_583), .fluid_out(k_9_291), .air_in(c_10_1));
valve v_10_584 (.fluid_in(k_10_584), .fluid_out(k_9_292), .air_in(c_10_0));
valve v_10_585 (.fluid_in(k_10_585), .fluid_out(k_9_292), .air_in(c_10_1));
valve v_10_586 (.fluid_in(k_10_586), .fluid_out(k_9_293), .air_in(c_10_0));
valve v_10_587 (.fluid_in(k_10_587), .fluid_out(k_9_293), .air_in(c_10_1));
valve v_10_588 (.fluid_in(k_10_588), .fluid_out(k_9_294), .air_in(c_10_0));
valve v_10_589 (.fluid_in(k_10_589), .fluid_out(k_9_294), .air_in(c_10_1));
valve v_10_590 (.fluid_in(k_10_590), .fluid_out(k_9_295), .air_in(c_10_0));
valve v_10_591 (.fluid_in(k_10_591), .fluid_out(k_9_295), .air_in(c_10_1));
valve v_10_592 (.fluid_in(k_10_592), .fluid_out(k_9_296), .air_in(c_10_0));
valve v_10_593 (.fluid_in(k_10_593), .fluid_out(k_9_296), .air_in(c_10_1));
valve v_10_594 (.fluid_in(k_10_594), .fluid_out(k_9_297), .air_in(c_10_0));
valve v_10_595 (.fluid_in(k_10_595), .fluid_out(k_9_297), .air_in(c_10_1));
valve v_10_596 (.fluid_in(k_10_596), .fluid_out(k_9_298), .air_in(c_10_0));
valve v_10_597 (.fluid_in(k_10_597), .fluid_out(k_9_298), .air_in(c_10_1));
valve v_10_598 (.fluid_in(k_10_598), .fluid_out(k_9_299), .air_in(c_10_0));
valve v_10_599 (.fluid_in(k_10_599), .fluid_out(k_9_299), .air_in(c_10_1));
valve v_10_600 (.fluid_in(k_10_600), .fluid_out(k_9_300), .air_in(c_10_0));
valve v_10_601 (.fluid_in(k_10_601), .fluid_out(k_9_300), .air_in(c_10_1));
valve v_10_602 (.fluid_in(k_10_602), .fluid_out(k_9_301), .air_in(c_10_0));
valve v_10_603 (.fluid_in(k_10_603), .fluid_out(k_9_301), .air_in(c_10_1));
valve v_10_604 (.fluid_in(k_10_604), .fluid_out(k_9_302), .air_in(c_10_0));
valve v_10_605 (.fluid_in(k_10_605), .fluid_out(k_9_302), .air_in(c_10_1));
valve v_10_606 (.fluid_in(k_10_606), .fluid_out(k_9_303), .air_in(c_10_0));
valve v_10_607 (.fluid_in(k_10_607), .fluid_out(k_9_303), .air_in(c_10_1));
valve v_10_608 (.fluid_in(k_10_608), .fluid_out(k_9_304), .air_in(c_10_0));
valve v_10_609 (.fluid_in(k_10_609), .fluid_out(k_9_304), .air_in(c_10_1));
valve v_10_610 (.fluid_in(k_10_610), .fluid_out(k_9_305), .air_in(c_10_0));
valve v_10_611 (.fluid_in(k_10_611), .fluid_out(k_9_305), .air_in(c_10_1));
valve v_10_612 (.fluid_in(k_10_612), .fluid_out(k_9_306), .air_in(c_10_0));
valve v_10_613 (.fluid_in(k_10_613), .fluid_out(k_9_306), .air_in(c_10_1));
valve v_10_614 (.fluid_in(k_10_614), .fluid_out(k_9_307), .air_in(c_10_0));
valve v_10_615 (.fluid_in(k_10_615), .fluid_out(k_9_307), .air_in(c_10_1));
valve v_10_616 (.fluid_in(k_10_616), .fluid_out(k_9_308), .air_in(c_10_0));
valve v_10_617 (.fluid_in(k_10_617), .fluid_out(k_9_308), .air_in(c_10_1));
valve v_10_618 (.fluid_in(k_10_618), .fluid_out(k_9_309), .air_in(c_10_0));
valve v_10_619 (.fluid_in(k_10_619), .fluid_out(k_9_309), .air_in(c_10_1));
valve v_10_620 (.fluid_in(k_10_620), .fluid_out(k_9_310), .air_in(c_10_0));
valve v_10_621 (.fluid_in(k_10_621), .fluid_out(k_9_310), .air_in(c_10_1));
valve v_10_622 (.fluid_in(k_10_622), .fluid_out(k_9_311), .air_in(c_10_0));
valve v_10_623 (.fluid_in(k_10_623), .fluid_out(k_9_311), .air_in(c_10_1));
valve v_10_624 (.fluid_in(k_10_624), .fluid_out(k_9_312), .air_in(c_10_0));
valve v_10_625 (.fluid_in(k_10_625), .fluid_out(k_9_312), .air_in(c_10_1));
valve v_10_626 (.fluid_in(k_10_626), .fluid_out(k_9_313), .air_in(c_10_0));
valve v_10_627 (.fluid_in(k_10_627), .fluid_out(k_9_313), .air_in(c_10_1));
valve v_10_628 (.fluid_in(k_10_628), .fluid_out(k_9_314), .air_in(c_10_0));
valve v_10_629 (.fluid_in(k_10_629), .fluid_out(k_9_314), .air_in(c_10_1));
valve v_10_630 (.fluid_in(k_10_630), .fluid_out(k_9_315), .air_in(c_10_0));
valve v_10_631 (.fluid_in(k_10_631), .fluid_out(k_9_315), .air_in(c_10_1));
valve v_10_632 (.fluid_in(k_10_632), .fluid_out(k_9_316), .air_in(c_10_0));
valve v_10_633 (.fluid_in(k_10_633), .fluid_out(k_9_316), .air_in(c_10_1));
valve v_10_634 (.fluid_in(k_10_634), .fluid_out(k_9_317), .air_in(c_10_0));
valve v_10_635 (.fluid_in(k_10_635), .fluid_out(k_9_317), .air_in(c_10_1));
valve v_10_636 (.fluid_in(k_10_636), .fluid_out(k_9_318), .air_in(c_10_0));
valve v_10_637 (.fluid_in(k_10_637), .fluid_out(k_9_318), .air_in(c_10_1));
valve v_10_638 (.fluid_in(k_10_638), .fluid_out(k_9_319), .air_in(c_10_0));
valve v_10_639 (.fluid_in(k_10_639), .fluid_out(k_9_319), .air_in(c_10_1));
valve v_10_640 (.fluid_in(k_10_640), .fluid_out(k_9_320), .air_in(c_10_0));
valve v_10_641 (.fluid_in(k_10_641), .fluid_out(k_9_320), .air_in(c_10_1));
valve v_10_642 (.fluid_in(k_10_642), .fluid_out(k_9_321), .air_in(c_10_0));
valve v_10_643 (.fluid_in(k_10_643), .fluid_out(k_9_321), .air_in(c_10_1));
valve v_10_644 (.fluid_in(k_10_644), .fluid_out(k_9_322), .air_in(c_10_0));
valve v_10_645 (.fluid_in(k_10_645), .fluid_out(k_9_322), .air_in(c_10_1));
valve v_10_646 (.fluid_in(k_10_646), .fluid_out(k_9_323), .air_in(c_10_0));
valve v_10_647 (.fluid_in(k_10_647), .fluid_out(k_9_323), .air_in(c_10_1));
valve v_10_648 (.fluid_in(k_10_648), .fluid_out(k_9_324), .air_in(c_10_0));
valve v_10_649 (.fluid_in(k_10_649), .fluid_out(k_9_324), .air_in(c_10_1));
valve v_10_650 (.fluid_in(k_10_650), .fluid_out(k_9_325), .air_in(c_10_0));
valve v_10_651 (.fluid_in(k_10_651), .fluid_out(k_9_325), .air_in(c_10_1));
valve v_10_652 (.fluid_in(k_10_652), .fluid_out(k_9_326), .air_in(c_10_0));
valve v_10_653 (.fluid_in(k_10_653), .fluid_out(k_9_326), .air_in(c_10_1));
valve v_10_654 (.fluid_in(k_10_654), .fluid_out(k_9_327), .air_in(c_10_0));
valve v_10_655 (.fluid_in(k_10_655), .fluid_out(k_9_327), .air_in(c_10_1));
valve v_10_656 (.fluid_in(k_10_656), .fluid_out(k_9_328), .air_in(c_10_0));
valve v_10_657 (.fluid_in(k_10_657), .fluid_out(k_9_328), .air_in(c_10_1));
valve v_10_658 (.fluid_in(k_10_658), .fluid_out(k_9_329), .air_in(c_10_0));
valve v_10_659 (.fluid_in(k_10_659), .fluid_out(k_9_329), .air_in(c_10_1));
valve v_10_660 (.fluid_in(k_10_660), .fluid_out(k_9_330), .air_in(c_10_0));
valve v_10_661 (.fluid_in(k_10_661), .fluid_out(k_9_330), .air_in(c_10_1));
valve v_10_662 (.fluid_in(k_10_662), .fluid_out(k_9_331), .air_in(c_10_0));
valve v_10_663 (.fluid_in(k_10_663), .fluid_out(k_9_331), .air_in(c_10_1));
valve v_10_664 (.fluid_in(k_10_664), .fluid_out(k_9_332), .air_in(c_10_0));
valve v_10_665 (.fluid_in(k_10_665), .fluid_out(k_9_332), .air_in(c_10_1));
valve v_10_666 (.fluid_in(k_10_666), .fluid_out(k_9_333), .air_in(c_10_0));
valve v_10_667 (.fluid_in(k_10_667), .fluid_out(k_9_333), .air_in(c_10_1));
valve v_10_668 (.fluid_in(k_10_668), .fluid_out(k_9_334), .air_in(c_10_0));
valve v_10_669 (.fluid_in(k_10_669), .fluid_out(k_9_334), .air_in(c_10_1));
valve v_10_670 (.fluid_in(k_10_670), .fluid_out(k_9_335), .air_in(c_10_0));
valve v_10_671 (.fluid_in(k_10_671), .fluid_out(k_9_335), .air_in(c_10_1));
valve v_10_672 (.fluid_in(k_10_672), .fluid_out(k_9_336), .air_in(c_10_0));
valve v_10_673 (.fluid_in(k_10_673), .fluid_out(k_9_336), .air_in(c_10_1));
valve v_10_674 (.fluid_in(k_10_674), .fluid_out(k_9_337), .air_in(c_10_0));
valve v_10_675 (.fluid_in(k_10_675), .fluid_out(k_9_337), .air_in(c_10_1));
valve v_10_676 (.fluid_in(k_10_676), .fluid_out(k_9_338), .air_in(c_10_0));
valve v_10_677 (.fluid_in(k_10_677), .fluid_out(k_9_338), .air_in(c_10_1));
valve v_10_678 (.fluid_in(k_10_678), .fluid_out(k_9_339), .air_in(c_10_0));
valve v_10_679 (.fluid_in(k_10_679), .fluid_out(k_9_339), .air_in(c_10_1));
valve v_10_680 (.fluid_in(k_10_680), .fluid_out(k_9_340), .air_in(c_10_0));
valve v_10_681 (.fluid_in(k_10_681), .fluid_out(k_9_340), .air_in(c_10_1));
valve v_10_682 (.fluid_in(k_10_682), .fluid_out(k_9_341), .air_in(c_10_0));
valve v_10_683 (.fluid_in(k_10_683), .fluid_out(k_9_341), .air_in(c_10_1));
valve v_10_684 (.fluid_in(k_10_684), .fluid_out(k_9_342), .air_in(c_10_0));
valve v_10_685 (.fluid_in(k_10_685), .fluid_out(k_9_342), .air_in(c_10_1));
valve v_10_686 (.fluid_in(k_10_686), .fluid_out(k_9_343), .air_in(c_10_0));
valve v_10_687 (.fluid_in(k_10_687), .fluid_out(k_9_343), .air_in(c_10_1));
valve v_10_688 (.fluid_in(k_10_688), .fluid_out(k_9_344), .air_in(c_10_0));
valve v_10_689 (.fluid_in(k_10_689), .fluid_out(k_9_344), .air_in(c_10_1));
valve v_10_690 (.fluid_in(k_10_690), .fluid_out(k_9_345), .air_in(c_10_0));
valve v_10_691 (.fluid_in(k_10_691), .fluid_out(k_9_345), .air_in(c_10_1));
valve v_10_692 (.fluid_in(k_10_692), .fluid_out(k_9_346), .air_in(c_10_0));
valve v_10_693 (.fluid_in(k_10_693), .fluid_out(k_9_346), .air_in(c_10_1));
valve v_10_694 (.fluid_in(k_10_694), .fluid_out(k_9_347), .air_in(c_10_0));
valve v_10_695 (.fluid_in(k_10_695), .fluid_out(k_9_347), .air_in(c_10_1));
valve v_10_696 (.fluid_in(k_10_696), .fluid_out(k_9_348), .air_in(c_10_0));
valve v_10_697 (.fluid_in(k_10_697), .fluid_out(k_9_348), .air_in(c_10_1));
valve v_10_698 (.fluid_in(k_10_698), .fluid_out(k_9_349), .air_in(c_10_0));
valve v_10_699 (.fluid_in(k_10_699), .fluid_out(k_9_349), .air_in(c_10_1));
valve v_10_700 (.fluid_in(k_10_700), .fluid_out(k_9_350), .air_in(c_10_0));
valve v_10_701 (.fluid_in(k_10_701), .fluid_out(k_9_350), .air_in(c_10_1));
valve v_10_702 (.fluid_in(k_10_702), .fluid_out(k_9_351), .air_in(c_10_0));
valve v_10_703 (.fluid_in(k_10_703), .fluid_out(k_9_351), .air_in(c_10_1));
valve v_10_704 (.fluid_in(k_10_704), .fluid_out(k_9_352), .air_in(c_10_0));
valve v_10_705 (.fluid_in(k_10_705), .fluid_out(k_9_352), .air_in(c_10_1));
valve v_10_706 (.fluid_in(k_10_706), .fluid_out(k_9_353), .air_in(c_10_0));
valve v_10_707 (.fluid_in(k_10_707), .fluid_out(k_9_353), .air_in(c_10_1));
valve v_10_708 (.fluid_in(k_10_708), .fluid_out(k_9_354), .air_in(c_10_0));
valve v_10_709 (.fluid_in(k_10_709), .fluid_out(k_9_354), .air_in(c_10_1));
valve v_10_710 (.fluid_in(k_10_710), .fluid_out(k_9_355), .air_in(c_10_0));
valve v_10_711 (.fluid_in(k_10_711), .fluid_out(k_9_355), .air_in(c_10_1));
valve v_10_712 (.fluid_in(k_10_712), .fluid_out(k_9_356), .air_in(c_10_0));
valve v_10_713 (.fluid_in(k_10_713), .fluid_out(k_9_356), .air_in(c_10_1));
valve v_10_714 (.fluid_in(k_10_714), .fluid_out(k_9_357), .air_in(c_10_0));
valve v_10_715 (.fluid_in(k_10_715), .fluid_out(k_9_357), .air_in(c_10_1));
valve v_10_716 (.fluid_in(k_10_716), .fluid_out(k_9_358), .air_in(c_10_0));
valve v_10_717 (.fluid_in(k_10_717), .fluid_out(k_9_358), .air_in(c_10_1));
valve v_10_718 (.fluid_in(k_10_718), .fluid_out(k_9_359), .air_in(c_10_0));
valve v_10_719 (.fluid_in(k_10_719), .fluid_out(k_9_359), .air_in(c_10_1));
valve v_10_720 (.fluid_in(k_10_720), .fluid_out(k_9_360), .air_in(c_10_0));
valve v_10_721 (.fluid_in(k_10_721), .fluid_out(k_9_360), .air_in(c_10_1));
valve v_10_722 (.fluid_in(k_10_722), .fluid_out(k_9_361), .air_in(c_10_0));
valve v_10_723 (.fluid_in(k_10_723), .fluid_out(k_9_361), .air_in(c_10_1));
valve v_10_724 (.fluid_in(k_10_724), .fluid_out(k_9_362), .air_in(c_10_0));
valve v_10_725 (.fluid_in(k_10_725), .fluid_out(k_9_362), .air_in(c_10_1));
valve v_10_726 (.fluid_in(k_10_726), .fluid_out(k_9_363), .air_in(c_10_0));
valve v_10_727 (.fluid_in(k_10_727), .fluid_out(k_9_363), .air_in(c_10_1));
valve v_10_728 (.fluid_in(k_10_728), .fluid_out(k_9_364), .air_in(c_10_0));
valve v_10_729 (.fluid_in(k_10_729), .fluid_out(k_9_364), .air_in(c_10_1));
valve v_10_730 (.fluid_in(k_10_730), .fluid_out(k_9_365), .air_in(c_10_0));
valve v_10_731 (.fluid_in(k_10_731), .fluid_out(k_9_365), .air_in(c_10_1));
valve v_10_732 (.fluid_in(k_10_732), .fluid_out(k_9_366), .air_in(c_10_0));
valve v_10_733 (.fluid_in(k_10_733), .fluid_out(k_9_366), .air_in(c_10_1));
valve v_10_734 (.fluid_in(k_10_734), .fluid_out(k_9_367), .air_in(c_10_0));
valve v_10_735 (.fluid_in(k_10_735), .fluid_out(k_9_367), .air_in(c_10_1));
valve v_10_736 (.fluid_in(k_10_736), .fluid_out(k_9_368), .air_in(c_10_0));
valve v_10_737 (.fluid_in(k_10_737), .fluid_out(k_9_368), .air_in(c_10_1));
valve v_10_738 (.fluid_in(k_10_738), .fluid_out(k_9_369), .air_in(c_10_0));
valve v_10_739 (.fluid_in(k_10_739), .fluid_out(k_9_369), .air_in(c_10_1));
valve v_10_740 (.fluid_in(k_10_740), .fluid_out(k_9_370), .air_in(c_10_0));
valve v_10_741 (.fluid_in(k_10_741), .fluid_out(k_9_370), .air_in(c_10_1));
valve v_10_742 (.fluid_in(k_10_742), .fluid_out(k_9_371), .air_in(c_10_0));
valve v_10_743 (.fluid_in(k_10_743), .fluid_out(k_9_371), .air_in(c_10_1));
valve v_10_744 (.fluid_in(k_10_744), .fluid_out(k_9_372), .air_in(c_10_0));
valve v_10_745 (.fluid_in(k_10_745), .fluid_out(k_9_372), .air_in(c_10_1));
valve v_10_746 (.fluid_in(k_10_746), .fluid_out(k_9_373), .air_in(c_10_0));
valve v_10_747 (.fluid_in(k_10_747), .fluid_out(k_9_373), .air_in(c_10_1));
valve v_10_748 (.fluid_in(k_10_748), .fluid_out(k_9_374), .air_in(c_10_0));
valve v_10_749 (.fluid_in(k_10_749), .fluid_out(k_9_374), .air_in(c_10_1));
valve v_10_750 (.fluid_in(k_10_750), .fluid_out(k_9_375), .air_in(c_10_0));
valve v_10_751 (.fluid_in(k_10_751), .fluid_out(k_9_375), .air_in(c_10_1));
valve v_10_752 (.fluid_in(k_10_752), .fluid_out(k_9_376), .air_in(c_10_0));
valve v_10_753 (.fluid_in(k_10_753), .fluid_out(k_9_376), .air_in(c_10_1));
valve v_10_754 (.fluid_in(k_10_754), .fluid_out(k_9_377), .air_in(c_10_0));
valve v_10_755 (.fluid_in(k_10_755), .fluid_out(k_9_377), .air_in(c_10_1));
valve v_10_756 (.fluid_in(k_10_756), .fluid_out(k_9_378), .air_in(c_10_0));
valve v_10_757 (.fluid_in(k_10_757), .fluid_out(k_9_378), .air_in(c_10_1));
valve v_10_758 (.fluid_in(k_10_758), .fluid_out(k_9_379), .air_in(c_10_0));
valve v_10_759 (.fluid_in(k_10_759), .fluid_out(k_9_379), .air_in(c_10_1));
valve v_10_760 (.fluid_in(k_10_760), .fluid_out(k_9_380), .air_in(c_10_0));
valve v_10_761 (.fluid_in(k_10_761), .fluid_out(k_9_380), .air_in(c_10_1));
valve v_10_762 (.fluid_in(k_10_762), .fluid_out(k_9_381), .air_in(c_10_0));
valve v_10_763 (.fluid_in(k_10_763), .fluid_out(k_9_381), .air_in(c_10_1));
valve v_10_764 (.fluid_in(k_10_764), .fluid_out(k_9_382), .air_in(c_10_0));
valve v_10_765 (.fluid_in(k_10_765), .fluid_out(k_9_382), .air_in(c_10_1));
valve v_10_766 (.fluid_in(k_10_766), .fluid_out(k_9_383), .air_in(c_10_0));
valve v_10_767 (.fluid_in(k_10_767), .fluid_out(k_9_383), .air_in(c_10_1));
valve v_10_768 (.fluid_in(k_10_768), .fluid_out(k_9_384), .air_in(c_10_0));
valve v_10_769 (.fluid_in(k_10_769), .fluid_out(k_9_384), .air_in(c_10_1));
valve v_10_770 (.fluid_in(k_10_770), .fluid_out(k_9_385), .air_in(c_10_0));
valve v_10_771 (.fluid_in(k_10_771), .fluid_out(k_9_385), .air_in(c_10_1));
valve v_10_772 (.fluid_in(k_10_772), .fluid_out(k_9_386), .air_in(c_10_0));
valve v_10_773 (.fluid_in(k_10_773), .fluid_out(k_9_386), .air_in(c_10_1));
valve v_10_774 (.fluid_in(k_10_774), .fluid_out(k_9_387), .air_in(c_10_0));
valve v_10_775 (.fluid_in(k_10_775), .fluid_out(k_9_387), .air_in(c_10_1));
valve v_10_776 (.fluid_in(k_10_776), .fluid_out(k_9_388), .air_in(c_10_0));
valve v_10_777 (.fluid_in(k_10_777), .fluid_out(k_9_388), .air_in(c_10_1));
valve v_10_778 (.fluid_in(k_10_778), .fluid_out(k_9_389), .air_in(c_10_0));
valve v_10_779 (.fluid_in(k_10_779), .fluid_out(k_9_389), .air_in(c_10_1));
valve v_10_780 (.fluid_in(k_10_780), .fluid_out(k_9_390), .air_in(c_10_0));
valve v_10_781 (.fluid_in(k_10_781), .fluid_out(k_9_390), .air_in(c_10_1));
valve v_10_782 (.fluid_in(k_10_782), .fluid_out(k_9_391), .air_in(c_10_0));
valve v_10_783 (.fluid_in(k_10_783), .fluid_out(k_9_391), .air_in(c_10_1));
valve v_10_784 (.fluid_in(k_10_784), .fluid_out(k_9_392), .air_in(c_10_0));
valve v_10_785 (.fluid_in(k_10_785), .fluid_out(k_9_392), .air_in(c_10_1));
valve v_10_786 (.fluid_in(k_10_786), .fluid_out(k_9_393), .air_in(c_10_0));
valve v_10_787 (.fluid_in(k_10_787), .fluid_out(k_9_393), .air_in(c_10_1));
valve v_10_788 (.fluid_in(k_10_788), .fluid_out(k_9_394), .air_in(c_10_0));
valve v_10_789 (.fluid_in(k_10_789), .fluid_out(k_9_394), .air_in(c_10_1));
valve v_10_790 (.fluid_in(k_10_790), .fluid_out(k_9_395), .air_in(c_10_0));
valve v_10_791 (.fluid_in(k_10_791), .fluid_out(k_9_395), .air_in(c_10_1));
valve v_10_792 (.fluid_in(k_10_792), .fluid_out(k_9_396), .air_in(c_10_0));
valve v_10_793 (.fluid_in(k_10_793), .fluid_out(k_9_396), .air_in(c_10_1));
valve v_10_794 (.fluid_in(k_10_794), .fluid_out(k_9_397), .air_in(c_10_0));
valve v_10_795 (.fluid_in(k_10_795), .fluid_out(k_9_397), .air_in(c_10_1));
valve v_10_796 (.fluid_in(k_10_796), .fluid_out(k_9_398), .air_in(c_10_0));
valve v_10_797 (.fluid_in(k_10_797), .fluid_out(k_9_398), .air_in(c_10_1));
valve v_10_798 (.fluid_in(k_10_798), .fluid_out(k_9_399), .air_in(c_10_0));
valve v_10_799 (.fluid_in(k_10_799), .fluid_out(k_9_399), .air_in(c_10_1));
valve v_10_800 (.fluid_in(k_10_800), .fluid_out(k_9_400), .air_in(c_10_0));
valve v_10_801 (.fluid_in(k_10_801), .fluid_out(k_9_400), .air_in(c_10_1));
valve v_10_802 (.fluid_in(k_10_802), .fluid_out(k_9_401), .air_in(c_10_0));
valve v_10_803 (.fluid_in(k_10_803), .fluid_out(k_9_401), .air_in(c_10_1));
valve v_10_804 (.fluid_in(k_10_804), .fluid_out(k_9_402), .air_in(c_10_0));
valve v_10_805 (.fluid_in(k_10_805), .fluid_out(k_9_402), .air_in(c_10_1));
valve v_10_806 (.fluid_in(k_10_806), .fluid_out(k_9_403), .air_in(c_10_0));
valve v_10_807 (.fluid_in(k_10_807), .fluid_out(k_9_403), .air_in(c_10_1));
valve v_10_808 (.fluid_in(k_10_808), .fluid_out(k_9_404), .air_in(c_10_0));
valve v_10_809 (.fluid_in(k_10_809), .fluid_out(k_9_404), .air_in(c_10_1));
valve v_10_810 (.fluid_in(k_10_810), .fluid_out(k_9_405), .air_in(c_10_0));
valve v_10_811 (.fluid_in(k_10_811), .fluid_out(k_9_405), .air_in(c_10_1));
valve v_10_812 (.fluid_in(k_10_812), .fluid_out(k_9_406), .air_in(c_10_0));
valve v_10_813 (.fluid_in(k_10_813), .fluid_out(k_9_406), .air_in(c_10_1));
valve v_10_814 (.fluid_in(k_10_814), .fluid_out(k_9_407), .air_in(c_10_0));
valve v_10_815 (.fluid_in(k_10_815), .fluid_out(k_9_407), .air_in(c_10_1));
valve v_10_816 (.fluid_in(k_10_816), .fluid_out(k_9_408), .air_in(c_10_0));
valve v_10_817 (.fluid_in(k_10_817), .fluid_out(k_9_408), .air_in(c_10_1));
valve v_10_818 (.fluid_in(k_10_818), .fluid_out(k_9_409), .air_in(c_10_0));
valve v_10_819 (.fluid_in(k_10_819), .fluid_out(k_9_409), .air_in(c_10_1));
valve v_10_820 (.fluid_in(k_10_820), .fluid_out(k_9_410), .air_in(c_10_0));
valve v_10_821 (.fluid_in(k_10_821), .fluid_out(k_9_410), .air_in(c_10_1));
valve v_10_822 (.fluid_in(k_10_822), .fluid_out(k_9_411), .air_in(c_10_0));
valve v_10_823 (.fluid_in(k_10_823), .fluid_out(k_9_411), .air_in(c_10_1));
valve v_10_824 (.fluid_in(k_10_824), .fluid_out(k_9_412), .air_in(c_10_0));
valve v_10_825 (.fluid_in(k_10_825), .fluid_out(k_9_412), .air_in(c_10_1));
valve v_10_826 (.fluid_in(k_10_826), .fluid_out(k_9_413), .air_in(c_10_0));
valve v_10_827 (.fluid_in(k_10_827), .fluid_out(k_9_413), .air_in(c_10_1));
valve v_10_828 (.fluid_in(k_10_828), .fluid_out(k_9_414), .air_in(c_10_0));
valve v_10_829 (.fluid_in(k_10_829), .fluid_out(k_9_414), .air_in(c_10_1));
valve v_10_830 (.fluid_in(k_10_830), .fluid_out(k_9_415), .air_in(c_10_0));
valve v_10_831 (.fluid_in(k_10_831), .fluid_out(k_9_415), .air_in(c_10_1));
valve v_10_832 (.fluid_in(k_10_832), .fluid_out(k_9_416), .air_in(c_10_0));
valve v_10_833 (.fluid_in(k_10_833), .fluid_out(k_9_416), .air_in(c_10_1));
valve v_10_834 (.fluid_in(k_10_834), .fluid_out(k_9_417), .air_in(c_10_0));
valve v_10_835 (.fluid_in(k_10_835), .fluid_out(k_9_417), .air_in(c_10_1));
valve v_10_836 (.fluid_in(k_10_836), .fluid_out(k_9_418), .air_in(c_10_0));
valve v_10_837 (.fluid_in(k_10_837), .fluid_out(k_9_418), .air_in(c_10_1));
valve v_10_838 (.fluid_in(k_10_838), .fluid_out(k_9_419), .air_in(c_10_0));
valve v_10_839 (.fluid_in(k_10_839), .fluid_out(k_9_419), .air_in(c_10_1));
valve v_10_840 (.fluid_in(k_10_840), .fluid_out(k_9_420), .air_in(c_10_0));
valve v_10_841 (.fluid_in(k_10_841), .fluid_out(k_9_420), .air_in(c_10_1));
valve v_10_842 (.fluid_in(k_10_842), .fluid_out(k_9_421), .air_in(c_10_0));
valve v_10_843 (.fluid_in(k_10_843), .fluid_out(k_9_421), .air_in(c_10_1));
valve v_10_844 (.fluid_in(k_10_844), .fluid_out(k_9_422), .air_in(c_10_0));
valve v_10_845 (.fluid_in(k_10_845), .fluid_out(k_9_422), .air_in(c_10_1));
valve v_10_846 (.fluid_in(k_10_846), .fluid_out(k_9_423), .air_in(c_10_0));
valve v_10_847 (.fluid_in(k_10_847), .fluid_out(k_9_423), .air_in(c_10_1));
valve v_10_848 (.fluid_in(k_10_848), .fluid_out(k_9_424), .air_in(c_10_0));
valve v_10_849 (.fluid_in(k_10_849), .fluid_out(k_9_424), .air_in(c_10_1));
valve v_10_850 (.fluid_in(k_10_850), .fluid_out(k_9_425), .air_in(c_10_0));
valve v_10_851 (.fluid_in(k_10_851), .fluid_out(k_9_425), .air_in(c_10_1));
valve v_10_852 (.fluid_in(k_10_852), .fluid_out(k_9_426), .air_in(c_10_0));
valve v_10_853 (.fluid_in(k_10_853), .fluid_out(k_9_426), .air_in(c_10_1));
valve v_10_854 (.fluid_in(k_10_854), .fluid_out(k_9_427), .air_in(c_10_0));
valve v_10_855 (.fluid_in(k_10_855), .fluid_out(k_9_427), .air_in(c_10_1));
valve v_10_856 (.fluid_in(k_10_856), .fluid_out(k_9_428), .air_in(c_10_0));
valve v_10_857 (.fluid_in(k_10_857), .fluid_out(k_9_428), .air_in(c_10_1));
valve v_10_858 (.fluid_in(k_10_858), .fluid_out(k_9_429), .air_in(c_10_0));
valve v_10_859 (.fluid_in(k_10_859), .fluid_out(k_9_429), .air_in(c_10_1));
valve v_10_860 (.fluid_in(k_10_860), .fluid_out(k_9_430), .air_in(c_10_0));
valve v_10_861 (.fluid_in(k_10_861), .fluid_out(k_9_430), .air_in(c_10_1));
valve v_10_862 (.fluid_in(k_10_862), .fluid_out(k_9_431), .air_in(c_10_0));
valve v_10_863 (.fluid_in(k_10_863), .fluid_out(k_9_431), .air_in(c_10_1));
valve v_10_864 (.fluid_in(k_10_864), .fluid_out(k_9_432), .air_in(c_10_0));
valve v_10_865 (.fluid_in(k_10_865), .fluid_out(k_9_432), .air_in(c_10_1));
valve v_10_866 (.fluid_in(k_10_866), .fluid_out(k_9_433), .air_in(c_10_0));
valve v_10_867 (.fluid_in(k_10_867), .fluid_out(k_9_433), .air_in(c_10_1));
valve v_10_868 (.fluid_in(k_10_868), .fluid_out(k_9_434), .air_in(c_10_0));
valve v_10_869 (.fluid_in(k_10_869), .fluid_out(k_9_434), .air_in(c_10_1));
valve v_10_870 (.fluid_in(k_10_870), .fluid_out(k_9_435), .air_in(c_10_0));
valve v_10_871 (.fluid_in(k_10_871), .fluid_out(k_9_435), .air_in(c_10_1));
valve v_10_872 (.fluid_in(k_10_872), .fluid_out(k_9_436), .air_in(c_10_0));
valve v_10_873 (.fluid_in(k_10_873), .fluid_out(k_9_436), .air_in(c_10_1));
valve v_10_874 (.fluid_in(k_10_874), .fluid_out(k_9_437), .air_in(c_10_0));
valve v_10_875 (.fluid_in(k_10_875), .fluid_out(k_9_437), .air_in(c_10_1));
valve v_10_876 (.fluid_in(k_10_876), .fluid_out(k_9_438), .air_in(c_10_0));
valve v_10_877 (.fluid_in(k_10_877), .fluid_out(k_9_438), .air_in(c_10_1));
valve v_10_878 (.fluid_in(k_10_878), .fluid_out(k_9_439), .air_in(c_10_0));
valve v_10_879 (.fluid_in(k_10_879), .fluid_out(k_9_439), .air_in(c_10_1));
valve v_10_880 (.fluid_in(k_10_880), .fluid_out(k_9_440), .air_in(c_10_0));
valve v_10_881 (.fluid_in(k_10_881), .fluid_out(k_9_440), .air_in(c_10_1));
valve v_10_882 (.fluid_in(k_10_882), .fluid_out(k_9_441), .air_in(c_10_0));
valve v_10_883 (.fluid_in(k_10_883), .fluid_out(k_9_441), .air_in(c_10_1));
valve v_10_884 (.fluid_in(k_10_884), .fluid_out(k_9_442), .air_in(c_10_0));
valve v_10_885 (.fluid_in(k_10_885), .fluid_out(k_9_442), .air_in(c_10_1));
valve v_10_886 (.fluid_in(k_10_886), .fluid_out(k_9_443), .air_in(c_10_0));
valve v_10_887 (.fluid_in(k_10_887), .fluid_out(k_9_443), .air_in(c_10_1));
valve v_10_888 (.fluid_in(k_10_888), .fluid_out(k_9_444), .air_in(c_10_0));
valve v_10_889 (.fluid_in(k_10_889), .fluid_out(k_9_444), .air_in(c_10_1));
valve v_10_890 (.fluid_in(k_10_890), .fluid_out(k_9_445), .air_in(c_10_0));
valve v_10_891 (.fluid_in(k_10_891), .fluid_out(k_9_445), .air_in(c_10_1));
valve v_10_892 (.fluid_in(k_10_892), .fluid_out(k_9_446), .air_in(c_10_0));
valve v_10_893 (.fluid_in(k_10_893), .fluid_out(k_9_446), .air_in(c_10_1));
valve v_10_894 (.fluid_in(k_10_894), .fluid_out(k_9_447), .air_in(c_10_0));
valve v_10_895 (.fluid_in(k_10_895), .fluid_out(k_9_447), .air_in(c_10_1));
valve v_10_896 (.fluid_in(k_10_896), .fluid_out(k_9_448), .air_in(c_10_0));
valve v_10_897 (.fluid_in(k_10_897), .fluid_out(k_9_448), .air_in(c_10_1));
valve v_10_898 (.fluid_in(k_10_898), .fluid_out(k_9_449), .air_in(c_10_0));
valve v_10_899 (.fluid_in(k_10_899), .fluid_out(k_9_449), .air_in(c_10_1));
valve v_10_900 (.fluid_in(k_10_900), .fluid_out(k_9_450), .air_in(c_10_0));
valve v_10_901 (.fluid_in(k_10_901), .fluid_out(k_9_450), .air_in(c_10_1));
valve v_10_902 (.fluid_in(k_10_902), .fluid_out(k_9_451), .air_in(c_10_0));
valve v_10_903 (.fluid_in(k_10_903), .fluid_out(k_9_451), .air_in(c_10_1));
valve v_10_904 (.fluid_in(k_10_904), .fluid_out(k_9_452), .air_in(c_10_0));
valve v_10_905 (.fluid_in(k_10_905), .fluid_out(k_9_452), .air_in(c_10_1));
valve v_10_906 (.fluid_in(k_10_906), .fluid_out(k_9_453), .air_in(c_10_0));
valve v_10_907 (.fluid_in(k_10_907), .fluid_out(k_9_453), .air_in(c_10_1));
valve v_10_908 (.fluid_in(k_10_908), .fluid_out(k_9_454), .air_in(c_10_0));
valve v_10_909 (.fluid_in(k_10_909), .fluid_out(k_9_454), .air_in(c_10_1));
valve v_10_910 (.fluid_in(k_10_910), .fluid_out(k_9_455), .air_in(c_10_0));
valve v_10_911 (.fluid_in(k_10_911), .fluid_out(k_9_455), .air_in(c_10_1));
valve v_10_912 (.fluid_in(k_10_912), .fluid_out(k_9_456), .air_in(c_10_0));
valve v_10_913 (.fluid_in(k_10_913), .fluid_out(k_9_456), .air_in(c_10_1));
valve v_10_914 (.fluid_in(k_10_914), .fluid_out(k_9_457), .air_in(c_10_0));
valve v_10_915 (.fluid_in(k_10_915), .fluid_out(k_9_457), .air_in(c_10_1));
valve v_10_916 (.fluid_in(k_10_916), .fluid_out(k_9_458), .air_in(c_10_0));
valve v_10_917 (.fluid_in(k_10_917), .fluid_out(k_9_458), .air_in(c_10_1));
valve v_10_918 (.fluid_in(k_10_918), .fluid_out(k_9_459), .air_in(c_10_0));
valve v_10_919 (.fluid_in(k_10_919), .fluid_out(k_9_459), .air_in(c_10_1));
valve v_10_920 (.fluid_in(k_10_920), .fluid_out(k_9_460), .air_in(c_10_0));
valve v_10_921 (.fluid_in(k_10_921), .fluid_out(k_9_460), .air_in(c_10_1));
valve v_10_922 (.fluid_in(k_10_922), .fluid_out(k_9_461), .air_in(c_10_0));
valve v_10_923 (.fluid_in(k_10_923), .fluid_out(k_9_461), .air_in(c_10_1));
valve v_10_924 (.fluid_in(k_10_924), .fluid_out(k_9_462), .air_in(c_10_0));
valve v_10_925 (.fluid_in(k_10_925), .fluid_out(k_9_462), .air_in(c_10_1));
valve v_10_926 (.fluid_in(k_10_926), .fluid_out(k_9_463), .air_in(c_10_0));
valve v_10_927 (.fluid_in(k_10_927), .fluid_out(k_9_463), .air_in(c_10_1));
valve v_10_928 (.fluid_in(k_10_928), .fluid_out(k_9_464), .air_in(c_10_0));
valve v_10_929 (.fluid_in(k_10_929), .fluid_out(k_9_464), .air_in(c_10_1));
valve v_10_930 (.fluid_in(k_10_930), .fluid_out(k_9_465), .air_in(c_10_0));
valve v_10_931 (.fluid_in(k_10_931), .fluid_out(k_9_465), .air_in(c_10_1));
valve v_10_932 (.fluid_in(k_10_932), .fluid_out(k_9_466), .air_in(c_10_0));
valve v_10_933 (.fluid_in(k_10_933), .fluid_out(k_9_466), .air_in(c_10_1));
valve v_10_934 (.fluid_in(k_10_934), .fluid_out(k_9_467), .air_in(c_10_0));
valve v_10_935 (.fluid_in(k_10_935), .fluid_out(k_9_467), .air_in(c_10_1));
valve v_10_936 (.fluid_in(k_10_936), .fluid_out(k_9_468), .air_in(c_10_0));
valve v_10_937 (.fluid_in(k_10_937), .fluid_out(k_9_468), .air_in(c_10_1));
valve v_10_938 (.fluid_in(k_10_938), .fluid_out(k_9_469), .air_in(c_10_0));
valve v_10_939 (.fluid_in(k_10_939), .fluid_out(k_9_469), .air_in(c_10_1));
valve v_10_940 (.fluid_in(k_10_940), .fluid_out(k_9_470), .air_in(c_10_0));
valve v_10_941 (.fluid_in(k_10_941), .fluid_out(k_9_470), .air_in(c_10_1));
valve v_10_942 (.fluid_in(k_10_942), .fluid_out(k_9_471), .air_in(c_10_0));
valve v_10_943 (.fluid_in(k_10_943), .fluid_out(k_9_471), .air_in(c_10_1));
valve v_10_944 (.fluid_in(k_10_944), .fluid_out(k_9_472), .air_in(c_10_0));
valve v_10_945 (.fluid_in(k_10_945), .fluid_out(k_9_472), .air_in(c_10_1));
valve v_10_946 (.fluid_in(k_10_946), .fluid_out(k_9_473), .air_in(c_10_0));
valve v_10_947 (.fluid_in(k_10_947), .fluid_out(k_9_473), .air_in(c_10_1));
valve v_10_948 (.fluid_in(k_10_948), .fluid_out(k_9_474), .air_in(c_10_0));
valve v_10_949 (.fluid_in(k_10_949), .fluid_out(k_9_474), .air_in(c_10_1));
valve v_10_950 (.fluid_in(k_10_950), .fluid_out(k_9_475), .air_in(c_10_0));
valve v_10_951 (.fluid_in(k_10_951), .fluid_out(k_9_475), .air_in(c_10_1));
valve v_10_952 (.fluid_in(k_10_952), .fluid_out(k_9_476), .air_in(c_10_0));
valve v_10_953 (.fluid_in(k_10_953), .fluid_out(k_9_476), .air_in(c_10_1));
valve v_10_954 (.fluid_in(k_10_954), .fluid_out(k_9_477), .air_in(c_10_0));
valve v_10_955 (.fluid_in(k_10_955), .fluid_out(k_9_477), .air_in(c_10_1));
valve v_10_956 (.fluid_in(k_10_956), .fluid_out(k_9_478), .air_in(c_10_0));
valve v_10_957 (.fluid_in(k_10_957), .fluid_out(k_9_478), .air_in(c_10_1));
valve v_10_958 (.fluid_in(k_10_958), .fluid_out(k_9_479), .air_in(c_10_0));
valve v_10_959 (.fluid_in(k_10_959), .fluid_out(k_9_479), .air_in(c_10_1));
valve v_10_960 (.fluid_in(k_10_960), .fluid_out(k_9_480), .air_in(c_10_0));
valve v_10_961 (.fluid_in(k_10_961), .fluid_out(k_9_480), .air_in(c_10_1));
valve v_10_962 (.fluid_in(k_10_962), .fluid_out(k_9_481), .air_in(c_10_0));
valve v_10_963 (.fluid_in(k_10_963), .fluid_out(k_9_481), .air_in(c_10_1));
valve v_10_964 (.fluid_in(k_10_964), .fluid_out(k_9_482), .air_in(c_10_0));
valve v_10_965 (.fluid_in(k_10_965), .fluid_out(k_9_482), .air_in(c_10_1));
valve v_10_966 (.fluid_in(k_10_966), .fluid_out(k_9_483), .air_in(c_10_0));
valve v_10_967 (.fluid_in(k_10_967), .fluid_out(k_9_483), .air_in(c_10_1));
valve v_10_968 (.fluid_in(k_10_968), .fluid_out(k_9_484), .air_in(c_10_0));
valve v_10_969 (.fluid_in(k_10_969), .fluid_out(k_9_484), .air_in(c_10_1));
valve v_10_970 (.fluid_in(k_10_970), .fluid_out(k_9_485), .air_in(c_10_0));
valve v_10_971 (.fluid_in(k_10_971), .fluid_out(k_9_485), .air_in(c_10_1));
valve v_10_972 (.fluid_in(k_10_972), .fluid_out(k_9_486), .air_in(c_10_0));
valve v_10_973 (.fluid_in(k_10_973), .fluid_out(k_9_486), .air_in(c_10_1));
valve v_10_974 (.fluid_in(k_10_974), .fluid_out(k_9_487), .air_in(c_10_0));
valve v_10_975 (.fluid_in(k_10_975), .fluid_out(k_9_487), .air_in(c_10_1));
valve v_10_976 (.fluid_in(k_10_976), .fluid_out(k_9_488), .air_in(c_10_0));
valve v_10_977 (.fluid_in(k_10_977), .fluid_out(k_9_488), .air_in(c_10_1));
valve v_10_978 (.fluid_in(k_10_978), .fluid_out(k_9_489), .air_in(c_10_0));
valve v_10_979 (.fluid_in(k_10_979), .fluid_out(k_9_489), .air_in(c_10_1));
valve v_10_980 (.fluid_in(k_10_980), .fluid_out(k_9_490), .air_in(c_10_0));
valve v_10_981 (.fluid_in(k_10_981), .fluid_out(k_9_490), .air_in(c_10_1));
valve v_10_982 (.fluid_in(k_10_982), .fluid_out(k_9_491), .air_in(c_10_0));
valve v_10_983 (.fluid_in(k_10_983), .fluid_out(k_9_491), .air_in(c_10_1));
valve v_10_984 (.fluid_in(k_10_984), .fluid_out(k_9_492), .air_in(c_10_0));
valve v_10_985 (.fluid_in(k_10_985), .fluid_out(k_9_492), .air_in(c_10_1));
valve v_10_986 (.fluid_in(k_10_986), .fluid_out(k_9_493), .air_in(c_10_0));
valve v_10_987 (.fluid_in(k_10_987), .fluid_out(k_9_493), .air_in(c_10_1));
valve v_10_988 (.fluid_in(k_10_988), .fluid_out(k_9_494), .air_in(c_10_0));
valve v_10_989 (.fluid_in(k_10_989), .fluid_out(k_9_494), .air_in(c_10_1));
valve v_10_990 (.fluid_in(k_10_990), .fluid_out(k_9_495), .air_in(c_10_0));
valve v_10_991 (.fluid_in(k_10_991), .fluid_out(k_9_495), .air_in(c_10_1));
valve v_10_992 (.fluid_in(k_10_992), .fluid_out(k_9_496), .air_in(c_10_0));
valve v_10_993 (.fluid_in(k_10_993), .fluid_out(k_9_496), .air_in(c_10_1));
valve v_10_994 (.fluid_in(k_10_994), .fluid_out(k_9_497), .air_in(c_10_0));
valve v_10_995 (.fluid_in(k_10_995), .fluid_out(k_9_497), .air_in(c_10_1));
valve v_10_996 (.fluid_in(k_10_996), .fluid_out(k_9_498), .air_in(c_10_0));
valve v_10_997 (.fluid_in(k_10_997), .fluid_out(k_9_498), .air_in(c_10_1));
valve v_10_998 (.fluid_in(k_10_998), .fluid_out(k_9_499), .air_in(c_10_0));
valve v_10_999 (.fluid_in(k_10_999), .fluid_out(k_9_499), .air_in(c_10_1));
valve v_10_1000 (.fluid_in(k_10_1000), .fluid_out(k_9_500), .air_in(c_10_0));
valve v_10_1001 (.fluid_in(k_10_1001), .fluid_out(k_9_500), .air_in(c_10_1));
valve v_10_1002 (.fluid_in(k_10_1002), .fluid_out(k_9_501), .air_in(c_10_0));
valve v_10_1003 (.fluid_in(k_10_1003), .fluid_out(k_9_501), .air_in(c_10_1));
valve v_10_1004 (.fluid_in(k_10_1004), .fluid_out(k_9_502), .air_in(c_10_0));
valve v_10_1005 (.fluid_in(k_10_1005), .fluid_out(k_9_502), .air_in(c_10_1));
valve v_10_1006 (.fluid_in(k_10_1006), .fluid_out(k_9_503), .air_in(c_10_0));
valve v_10_1007 (.fluid_in(k_10_1007), .fluid_out(k_9_503), .air_in(c_10_1));
valve v_10_1008 (.fluid_in(k_10_1008), .fluid_out(k_9_504), .air_in(c_10_0));
valve v_10_1009 (.fluid_in(k_10_1009), .fluid_out(k_9_504), .air_in(c_10_1));
valve v_10_1010 (.fluid_in(k_10_1010), .fluid_out(k_9_505), .air_in(c_10_0));
valve v_10_1011 (.fluid_in(k_10_1011), .fluid_out(k_9_505), .air_in(c_10_1));
valve v_10_1012 (.fluid_in(k_10_1012), .fluid_out(k_9_506), .air_in(c_10_0));
valve v_10_1013 (.fluid_in(k_10_1013), .fluid_out(k_9_506), .air_in(c_10_1));
valve v_10_1014 (.fluid_in(k_10_1014), .fluid_out(k_9_507), .air_in(c_10_0));
valve v_10_1015 (.fluid_in(k_10_1015), .fluid_out(k_9_507), .air_in(c_10_1));
valve v_10_1016 (.fluid_in(k_10_1016), .fluid_out(k_9_508), .air_in(c_10_0));
valve v_10_1017 (.fluid_in(k_10_1017), .fluid_out(k_9_508), .air_in(c_10_1));
valve v_10_1018 (.fluid_in(k_10_1018), .fluid_out(k_9_509), .air_in(c_10_0));
valve v_10_1019 (.fluid_in(k_10_1019), .fluid_out(k_9_509), .air_in(c_10_1));
valve v_10_1020 (.fluid_in(k_10_1020), .fluid_out(k_9_510), .air_in(c_10_0));
valve v_10_1021 (.fluid_in(k_10_1021), .fluid_out(k_9_510), .air_in(c_10_1));
valve v_10_1022 (.fluid_in(k_10_1022), .fluid_out(k_9_511), .air_in(c_10_0));
valve v_10_1023 (.fluid_in(k_10_1023), .fluid_out(k_9_511), .air_in(c_10_1));
endmodule
