module fanout2_braid_4_8 (
output output_0,output output_1,output output_2,output output_3,input input_0,input input_1,input input_2,input input_3
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_1_3, output_1_0, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_0), .y(output_0_3));
wire output_2_3, output_2_0, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_0), .y(output_1_3));
wire output_3_3, output_3_0, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_0), .y(output_2_3));
wire output_4_3, output_4_0, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_0), .y(output_3_3));
wire output_1_4, output_1_1, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_1), .y(output_0_4));
wire output_2_4, output_2_1, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_1), .y(output_1_4));
wire output_3_4, output_3_1, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_1), .y(output_2_4));
wire output_4_4, output_4_1, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_1), .y(output_3_4));
wire output_1_5, output_1_2, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_2), .y(output_0_5));
wire output_2_5, output_2_2, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_2), .y(output_1_5));
wire output_3_5, output_3_2, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_2), .y(output_2_5));
wire output_4_5, output_4_2, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_2), .y(output_3_5));
wire output_1_6, output_1_3, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_3), .y(output_0_6));
wire output_2_6, output_2_3, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_3), .y(output_1_6));
wire output_3_6, output_3_3, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_3), .y(output_2_6));
wire output_4_6, output_4_3, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_3), .y(output_3_6));
wire output_1_7, output_1_0, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_0), .y(output_0_7));
wire output_2_7, output_2_0, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_0), .y(output_1_7));
wire output_3_7, output_3_0, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_0), .y(output_2_7));
wire output_4_7, output_4_0, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_0), .y(output_3_7));
assign output_0 = output_0_0;
wire output_0_8;
assign output_0_8 = input_0;
assign output_1 = output_1_0;
wire output_1_8;
assign output_1_8 = input_1;
assign output_2 = output_2_0;
wire output_2_8;
assign output_2_8 = input_2;
assign output_3 = output_3_0;
wire output_3_8;
assign output_3_8 = input_3;
endmodule
