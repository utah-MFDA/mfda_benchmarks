module multiplexer_8 (
inout k_0_0,k_8_0,k_8_1,k_8_2,k_8_3,k_8_4,k_8_5,k_8_6,k_8_7,k_8_8,k_8_9,k_8_10,k_8_11,k_8_12,k_8_13,k_8_14,k_8_15,k_8_16,k_8_17,k_8_18,k_8_19,k_8_20,k_8_21,k_8_22,k_8_23,k_8_24,k_8_25,k_8_26,k_8_27,k_8_28,k_8_29,k_8_30,k_8_31,k_8_32,k_8_33,k_8_34,k_8_35,k_8_36,k_8_37,k_8_38,k_8_39,k_8_40,k_8_41,k_8_42,k_8_43,k_8_44,k_8_45,k_8_46,k_8_47,k_8_48,k_8_49,k_8_50,k_8_51,k_8_52,k_8_53,k_8_54,k_8_55,k_8_56,k_8_57,k_8_58,k_8_59,k_8_60,k_8_61,k_8_62,k_8_63,k_8_64,k_8_65,k_8_66,k_8_67,k_8_68,k_8_69,k_8_70,k_8_71,k_8_72,k_8_73,k_8_74,k_8_75,k_8_76,k_8_77,k_8_78,k_8_79,k_8_80,k_8_81,k_8_82,k_8_83,k_8_84,k_8_85,k_8_86,k_8_87,k_8_88,k_8_89,k_8_90,k_8_91,k_8_92,k_8_93,k_8_94,k_8_95,k_8_96,k_8_97,k_8_98,k_8_99,k_8_100,k_8_101,k_8_102,k_8_103,k_8_104,k_8_105,k_8_106,k_8_107,k_8_108,k_8_109,k_8_110,k_8_111,k_8_112,k_8_113,k_8_114,k_8_115,k_8_116,k_8_117,k_8_118,k_8_119,k_8_120,k_8_121,k_8_122,k_8_123,k_8_124,k_8_125,k_8_126,k_8_127,k_8_128,k_8_129,k_8_130,k_8_131,k_8_132,k_8_133,k_8_134,k_8_135,k_8_136,k_8_137,k_8_138,k_8_139,k_8_140,k_8_141,k_8_142,k_8_143,k_8_144,k_8_145,k_8_146,k_8_147,k_8_148,k_8_149,k_8_150,k_8_151,k_8_152,k_8_153,k_8_154,k_8_155,k_8_156,k_8_157,k_8_158,k_8_159,k_8_160,k_8_161,k_8_162,k_8_163,k_8_164,k_8_165,k_8_166,k_8_167,k_8_168,k_8_169,k_8_170,k_8_171,k_8_172,k_8_173,k_8_174,k_8_175,k_8_176,k_8_177,k_8_178,k_8_179,k_8_180,k_8_181,k_8_182,k_8_183,k_8_184,k_8_185,k_8_186,k_8_187,k_8_188,k_8_189,k_8_190,k_8_191,k_8_192,k_8_193,k_8_194,k_8_195,k_8_196,k_8_197,k_8_198,k_8_199,k_8_200,k_8_201,k_8_202,k_8_203,k_8_204,k_8_205,k_8_206,k_8_207,k_8_208,k_8_209,k_8_210,k_8_211,k_8_212,k_8_213,k_8_214,k_8_215,k_8_216,k_8_217,k_8_218,k_8_219,k_8_220,k_8_221,k_8_222,k_8_223,k_8_224,k_8_225,k_8_226,k_8_227,k_8_228,k_8_229,k_8_230,k_8_231,k_8_232,k_8_233,k_8_234,k_8_235,k_8_236,k_8_237,k_8_238,k_8_239,k_8_240,k_8_241,k_8_242,k_8_243,k_8_244,k_8_245,k_8_246,k_8_247,k_8_248,k_8_249,k_8_250,k_8_251,k_8_252,k_8_253,k_8_254,k_8_255,
input c_0_0, c_0_1,
input c_1_0, c_1_1,
input c_2_0, c_2_1,
input c_3_0, c_3_1,
input c_4_0, c_4_1,
input c_5_0, c_5_1,
input c_6_0, c_6_1,
input c_7_0, c_7_1,
input c_8_0, c_8_1
);
wire k_1_0,k_1_1;
wire k_2_0,k_2_1,k_2_2,k_2_3;
wire k_3_0,k_3_1,k_3_2,k_3_3,k_3_4,k_3_5,k_3_6,k_3_7;
wire k_4_0,k_4_1,k_4_2,k_4_3,k_4_4,k_4_5,k_4_6,k_4_7,k_4_8,k_4_9,k_4_10,k_4_11,k_4_12,k_4_13,k_4_14,k_4_15;
wire k_5_0,k_5_1,k_5_2,k_5_3,k_5_4,k_5_5,k_5_6,k_5_7,k_5_8,k_5_9,k_5_10,k_5_11,k_5_12,k_5_13,k_5_14,k_5_15,k_5_16,k_5_17,k_5_18,k_5_19,k_5_20,k_5_21,k_5_22,k_5_23,k_5_24,k_5_25,k_5_26,k_5_27,k_5_28,k_5_29,k_5_30,k_5_31;
wire k_6_0,k_6_1,k_6_2,k_6_3,k_6_4,k_6_5,k_6_6,k_6_7,k_6_8,k_6_9,k_6_10,k_6_11,k_6_12,k_6_13,k_6_14,k_6_15,k_6_16,k_6_17,k_6_18,k_6_19,k_6_20,k_6_21,k_6_22,k_6_23,k_6_24,k_6_25,k_6_26,k_6_27,k_6_28,k_6_29,k_6_30,k_6_31,k_6_32,k_6_33,k_6_34,k_6_35,k_6_36,k_6_37,k_6_38,k_6_39,k_6_40,k_6_41,k_6_42,k_6_43,k_6_44,k_6_45,k_6_46,k_6_47,k_6_48,k_6_49,k_6_50,k_6_51,k_6_52,k_6_53,k_6_54,k_6_55,k_6_56,k_6_57,k_6_58,k_6_59,k_6_60,k_6_61,k_6_62,k_6_63;
wire k_7_0,k_7_1,k_7_2,k_7_3,k_7_4,k_7_5,k_7_6,k_7_7,k_7_8,k_7_9,k_7_10,k_7_11,k_7_12,k_7_13,k_7_14,k_7_15,k_7_16,k_7_17,k_7_18,k_7_19,k_7_20,k_7_21,k_7_22,k_7_23,k_7_24,k_7_25,k_7_26,k_7_27,k_7_28,k_7_29,k_7_30,k_7_31,k_7_32,k_7_33,k_7_34,k_7_35,k_7_36,k_7_37,k_7_38,k_7_39,k_7_40,k_7_41,k_7_42,k_7_43,k_7_44,k_7_45,k_7_46,k_7_47,k_7_48,k_7_49,k_7_50,k_7_51,k_7_52,k_7_53,k_7_54,k_7_55,k_7_56,k_7_57,k_7_58,k_7_59,k_7_60,k_7_61,k_7_62,k_7_63,k_7_64,k_7_65,k_7_66,k_7_67,k_7_68,k_7_69,k_7_70,k_7_71,k_7_72,k_7_73,k_7_74,k_7_75,k_7_76,k_7_77,k_7_78,k_7_79,k_7_80,k_7_81,k_7_82,k_7_83,k_7_84,k_7_85,k_7_86,k_7_87,k_7_88,k_7_89,k_7_90,k_7_91,k_7_92,k_7_93,k_7_94,k_7_95,k_7_96,k_7_97,k_7_98,k_7_99,k_7_100,k_7_101,k_7_102,k_7_103,k_7_104,k_7_105,k_7_106,k_7_107,k_7_108,k_7_109,k_7_110,k_7_111,k_7_112,k_7_113,k_7_114,k_7_115,k_7_116,k_7_117,k_7_118,k_7_119,k_7_120,k_7_121,k_7_122,k_7_123,k_7_124,k_7_125,k_7_126,k_7_127;
valve v_1_0 (.fluid_in(k_1_0), .fluid_out(k_0_0), .air_in(c_1_0));
valve v_1_1 (.fluid_in(k_1_1), .fluid_out(k_0_0), .air_in(c_1_1));
valve v_2_0 (.fluid_in(k_2_0), .fluid_out(k_1_0), .air_in(c_2_0));
valve v_2_1 (.fluid_in(k_2_1), .fluid_out(k_1_0), .air_in(c_2_1));
valve v_2_2 (.fluid_in(k_2_2), .fluid_out(k_1_1), .air_in(c_2_0));
valve v_2_3 (.fluid_in(k_2_3), .fluid_out(k_1_1), .air_in(c_2_1));
valve v_3_0 (.fluid_in(k_3_0), .fluid_out(k_2_0), .air_in(c_3_0));
valve v_3_1 (.fluid_in(k_3_1), .fluid_out(k_2_0), .air_in(c_3_1));
valve v_3_2 (.fluid_in(k_3_2), .fluid_out(k_2_1), .air_in(c_3_0));
valve v_3_3 (.fluid_in(k_3_3), .fluid_out(k_2_1), .air_in(c_3_1));
valve v_3_4 (.fluid_in(k_3_4), .fluid_out(k_2_2), .air_in(c_3_0));
valve v_3_5 (.fluid_in(k_3_5), .fluid_out(k_2_2), .air_in(c_3_1));
valve v_3_6 (.fluid_in(k_3_6), .fluid_out(k_2_3), .air_in(c_3_0));
valve v_3_7 (.fluid_in(k_3_7), .fluid_out(k_2_3), .air_in(c_3_1));
valve v_4_0 (.fluid_in(k_4_0), .fluid_out(k_3_0), .air_in(c_4_0));
valve v_4_1 (.fluid_in(k_4_1), .fluid_out(k_3_0), .air_in(c_4_1));
valve v_4_2 (.fluid_in(k_4_2), .fluid_out(k_3_1), .air_in(c_4_0));
valve v_4_3 (.fluid_in(k_4_3), .fluid_out(k_3_1), .air_in(c_4_1));
valve v_4_4 (.fluid_in(k_4_4), .fluid_out(k_3_2), .air_in(c_4_0));
valve v_4_5 (.fluid_in(k_4_5), .fluid_out(k_3_2), .air_in(c_4_1));
valve v_4_6 (.fluid_in(k_4_6), .fluid_out(k_3_3), .air_in(c_4_0));
valve v_4_7 (.fluid_in(k_4_7), .fluid_out(k_3_3), .air_in(c_4_1));
valve v_4_8 (.fluid_in(k_4_8), .fluid_out(k_3_4), .air_in(c_4_0));
valve v_4_9 (.fluid_in(k_4_9), .fluid_out(k_3_4), .air_in(c_4_1));
valve v_4_10 (.fluid_in(k_4_10), .fluid_out(k_3_5), .air_in(c_4_0));
valve v_4_11 (.fluid_in(k_4_11), .fluid_out(k_3_5), .air_in(c_4_1));
valve v_4_12 (.fluid_in(k_4_12), .fluid_out(k_3_6), .air_in(c_4_0));
valve v_4_13 (.fluid_in(k_4_13), .fluid_out(k_3_6), .air_in(c_4_1));
valve v_4_14 (.fluid_in(k_4_14), .fluid_out(k_3_7), .air_in(c_4_0));
valve v_4_15 (.fluid_in(k_4_15), .fluid_out(k_3_7), .air_in(c_4_1));
valve v_5_0 (.fluid_in(k_5_0), .fluid_out(k_4_0), .air_in(c_5_0));
valve v_5_1 (.fluid_in(k_5_1), .fluid_out(k_4_0), .air_in(c_5_1));
valve v_5_2 (.fluid_in(k_5_2), .fluid_out(k_4_1), .air_in(c_5_0));
valve v_5_3 (.fluid_in(k_5_3), .fluid_out(k_4_1), .air_in(c_5_1));
valve v_5_4 (.fluid_in(k_5_4), .fluid_out(k_4_2), .air_in(c_5_0));
valve v_5_5 (.fluid_in(k_5_5), .fluid_out(k_4_2), .air_in(c_5_1));
valve v_5_6 (.fluid_in(k_5_6), .fluid_out(k_4_3), .air_in(c_5_0));
valve v_5_7 (.fluid_in(k_5_7), .fluid_out(k_4_3), .air_in(c_5_1));
valve v_5_8 (.fluid_in(k_5_8), .fluid_out(k_4_4), .air_in(c_5_0));
valve v_5_9 (.fluid_in(k_5_9), .fluid_out(k_4_4), .air_in(c_5_1));
valve v_5_10 (.fluid_in(k_5_10), .fluid_out(k_4_5), .air_in(c_5_0));
valve v_5_11 (.fluid_in(k_5_11), .fluid_out(k_4_5), .air_in(c_5_1));
valve v_5_12 (.fluid_in(k_5_12), .fluid_out(k_4_6), .air_in(c_5_0));
valve v_5_13 (.fluid_in(k_5_13), .fluid_out(k_4_6), .air_in(c_5_1));
valve v_5_14 (.fluid_in(k_5_14), .fluid_out(k_4_7), .air_in(c_5_0));
valve v_5_15 (.fluid_in(k_5_15), .fluid_out(k_4_7), .air_in(c_5_1));
valve v_5_16 (.fluid_in(k_5_16), .fluid_out(k_4_8), .air_in(c_5_0));
valve v_5_17 (.fluid_in(k_5_17), .fluid_out(k_4_8), .air_in(c_5_1));
valve v_5_18 (.fluid_in(k_5_18), .fluid_out(k_4_9), .air_in(c_5_0));
valve v_5_19 (.fluid_in(k_5_19), .fluid_out(k_4_9), .air_in(c_5_1));
valve v_5_20 (.fluid_in(k_5_20), .fluid_out(k_4_10), .air_in(c_5_0));
valve v_5_21 (.fluid_in(k_5_21), .fluid_out(k_4_10), .air_in(c_5_1));
valve v_5_22 (.fluid_in(k_5_22), .fluid_out(k_4_11), .air_in(c_5_0));
valve v_5_23 (.fluid_in(k_5_23), .fluid_out(k_4_11), .air_in(c_5_1));
valve v_5_24 (.fluid_in(k_5_24), .fluid_out(k_4_12), .air_in(c_5_0));
valve v_5_25 (.fluid_in(k_5_25), .fluid_out(k_4_12), .air_in(c_5_1));
valve v_5_26 (.fluid_in(k_5_26), .fluid_out(k_4_13), .air_in(c_5_0));
valve v_5_27 (.fluid_in(k_5_27), .fluid_out(k_4_13), .air_in(c_5_1));
valve v_5_28 (.fluid_in(k_5_28), .fluid_out(k_4_14), .air_in(c_5_0));
valve v_5_29 (.fluid_in(k_5_29), .fluid_out(k_4_14), .air_in(c_5_1));
valve v_5_30 (.fluid_in(k_5_30), .fluid_out(k_4_15), .air_in(c_5_0));
valve v_5_31 (.fluid_in(k_5_31), .fluid_out(k_4_15), .air_in(c_5_1));
valve v_6_0 (.fluid_in(k_6_0), .fluid_out(k_5_0), .air_in(c_6_0));
valve v_6_1 (.fluid_in(k_6_1), .fluid_out(k_5_0), .air_in(c_6_1));
valve v_6_2 (.fluid_in(k_6_2), .fluid_out(k_5_1), .air_in(c_6_0));
valve v_6_3 (.fluid_in(k_6_3), .fluid_out(k_5_1), .air_in(c_6_1));
valve v_6_4 (.fluid_in(k_6_4), .fluid_out(k_5_2), .air_in(c_6_0));
valve v_6_5 (.fluid_in(k_6_5), .fluid_out(k_5_2), .air_in(c_6_1));
valve v_6_6 (.fluid_in(k_6_6), .fluid_out(k_5_3), .air_in(c_6_0));
valve v_6_7 (.fluid_in(k_6_7), .fluid_out(k_5_3), .air_in(c_6_1));
valve v_6_8 (.fluid_in(k_6_8), .fluid_out(k_5_4), .air_in(c_6_0));
valve v_6_9 (.fluid_in(k_6_9), .fluid_out(k_5_4), .air_in(c_6_1));
valve v_6_10 (.fluid_in(k_6_10), .fluid_out(k_5_5), .air_in(c_6_0));
valve v_6_11 (.fluid_in(k_6_11), .fluid_out(k_5_5), .air_in(c_6_1));
valve v_6_12 (.fluid_in(k_6_12), .fluid_out(k_5_6), .air_in(c_6_0));
valve v_6_13 (.fluid_in(k_6_13), .fluid_out(k_5_6), .air_in(c_6_1));
valve v_6_14 (.fluid_in(k_6_14), .fluid_out(k_5_7), .air_in(c_6_0));
valve v_6_15 (.fluid_in(k_6_15), .fluid_out(k_5_7), .air_in(c_6_1));
valve v_6_16 (.fluid_in(k_6_16), .fluid_out(k_5_8), .air_in(c_6_0));
valve v_6_17 (.fluid_in(k_6_17), .fluid_out(k_5_8), .air_in(c_6_1));
valve v_6_18 (.fluid_in(k_6_18), .fluid_out(k_5_9), .air_in(c_6_0));
valve v_6_19 (.fluid_in(k_6_19), .fluid_out(k_5_9), .air_in(c_6_1));
valve v_6_20 (.fluid_in(k_6_20), .fluid_out(k_5_10), .air_in(c_6_0));
valve v_6_21 (.fluid_in(k_6_21), .fluid_out(k_5_10), .air_in(c_6_1));
valve v_6_22 (.fluid_in(k_6_22), .fluid_out(k_5_11), .air_in(c_6_0));
valve v_6_23 (.fluid_in(k_6_23), .fluid_out(k_5_11), .air_in(c_6_1));
valve v_6_24 (.fluid_in(k_6_24), .fluid_out(k_5_12), .air_in(c_6_0));
valve v_6_25 (.fluid_in(k_6_25), .fluid_out(k_5_12), .air_in(c_6_1));
valve v_6_26 (.fluid_in(k_6_26), .fluid_out(k_5_13), .air_in(c_6_0));
valve v_6_27 (.fluid_in(k_6_27), .fluid_out(k_5_13), .air_in(c_6_1));
valve v_6_28 (.fluid_in(k_6_28), .fluid_out(k_5_14), .air_in(c_6_0));
valve v_6_29 (.fluid_in(k_6_29), .fluid_out(k_5_14), .air_in(c_6_1));
valve v_6_30 (.fluid_in(k_6_30), .fluid_out(k_5_15), .air_in(c_6_0));
valve v_6_31 (.fluid_in(k_6_31), .fluid_out(k_5_15), .air_in(c_6_1));
valve v_6_32 (.fluid_in(k_6_32), .fluid_out(k_5_16), .air_in(c_6_0));
valve v_6_33 (.fluid_in(k_6_33), .fluid_out(k_5_16), .air_in(c_6_1));
valve v_6_34 (.fluid_in(k_6_34), .fluid_out(k_5_17), .air_in(c_6_0));
valve v_6_35 (.fluid_in(k_6_35), .fluid_out(k_5_17), .air_in(c_6_1));
valve v_6_36 (.fluid_in(k_6_36), .fluid_out(k_5_18), .air_in(c_6_0));
valve v_6_37 (.fluid_in(k_6_37), .fluid_out(k_5_18), .air_in(c_6_1));
valve v_6_38 (.fluid_in(k_6_38), .fluid_out(k_5_19), .air_in(c_6_0));
valve v_6_39 (.fluid_in(k_6_39), .fluid_out(k_5_19), .air_in(c_6_1));
valve v_6_40 (.fluid_in(k_6_40), .fluid_out(k_5_20), .air_in(c_6_0));
valve v_6_41 (.fluid_in(k_6_41), .fluid_out(k_5_20), .air_in(c_6_1));
valve v_6_42 (.fluid_in(k_6_42), .fluid_out(k_5_21), .air_in(c_6_0));
valve v_6_43 (.fluid_in(k_6_43), .fluid_out(k_5_21), .air_in(c_6_1));
valve v_6_44 (.fluid_in(k_6_44), .fluid_out(k_5_22), .air_in(c_6_0));
valve v_6_45 (.fluid_in(k_6_45), .fluid_out(k_5_22), .air_in(c_6_1));
valve v_6_46 (.fluid_in(k_6_46), .fluid_out(k_5_23), .air_in(c_6_0));
valve v_6_47 (.fluid_in(k_6_47), .fluid_out(k_5_23), .air_in(c_6_1));
valve v_6_48 (.fluid_in(k_6_48), .fluid_out(k_5_24), .air_in(c_6_0));
valve v_6_49 (.fluid_in(k_6_49), .fluid_out(k_5_24), .air_in(c_6_1));
valve v_6_50 (.fluid_in(k_6_50), .fluid_out(k_5_25), .air_in(c_6_0));
valve v_6_51 (.fluid_in(k_6_51), .fluid_out(k_5_25), .air_in(c_6_1));
valve v_6_52 (.fluid_in(k_6_52), .fluid_out(k_5_26), .air_in(c_6_0));
valve v_6_53 (.fluid_in(k_6_53), .fluid_out(k_5_26), .air_in(c_6_1));
valve v_6_54 (.fluid_in(k_6_54), .fluid_out(k_5_27), .air_in(c_6_0));
valve v_6_55 (.fluid_in(k_6_55), .fluid_out(k_5_27), .air_in(c_6_1));
valve v_6_56 (.fluid_in(k_6_56), .fluid_out(k_5_28), .air_in(c_6_0));
valve v_6_57 (.fluid_in(k_6_57), .fluid_out(k_5_28), .air_in(c_6_1));
valve v_6_58 (.fluid_in(k_6_58), .fluid_out(k_5_29), .air_in(c_6_0));
valve v_6_59 (.fluid_in(k_6_59), .fluid_out(k_5_29), .air_in(c_6_1));
valve v_6_60 (.fluid_in(k_6_60), .fluid_out(k_5_30), .air_in(c_6_0));
valve v_6_61 (.fluid_in(k_6_61), .fluid_out(k_5_30), .air_in(c_6_1));
valve v_6_62 (.fluid_in(k_6_62), .fluid_out(k_5_31), .air_in(c_6_0));
valve v_6_63 (.fluid_in(k_6_63), .fluid_out(k_5_31), .air_in(c_6_1));
valve v_7_0 (.fluid_in(k_7_0), .fluid_out(k_6_0), .air_in(c_7_0));
valve v_7_1 (.fluid_in(k_7_1), .fluid_out(k_6_0), .air_in(c_7_1));
valve v_7_2 (.fluid_in(k_7_2), .fluid_out(k_6_1), .air_in(c_7_0));
valve v_7_3 (.fluid_in(k_7_3), .fluid_out(k_6_1), .air_in(c_7_1));
valve v_7_4 (.fluid_in(k_7_4), .fluid_out(k_6_2), .air_in(c_7_0));
valve v_7_5 (.fluid_in(k_7_5), .fluid_out(k_6_2), .air_in(c_7_1));
valve v_7_6 (.fluid_in(k_7_6), .fluid_out(k_6_3), .air_in(c_7_0));
valve v_7_7 (.fluid_in(k_7_7), .fluid_out(k_6_3), .air_in(c_7_1));
valve v_7_8 (.fluid_in(k_7_8), .fluid_out(k_6_4), .air_in(c_7_0));
valve v_7_9 (.fluid_in(k_7_9), .fluid_out(k_6_4), .air_in(c_7_1));
valve v_7_10 (.fluid_in(k_7_10), .fluid_out(k_6_5), .air_in(c_7_0));
valve v_7_11 (.fluid_in(k_7_11), .fluid_out(k_6_5), .air_in(c_7_1));
valve v_7_12 (.fluid_in(k_7_12), .fluid_out(k_6_6), .air_in(c_7_0));
valve v_7_13 (.fluid_in(k_7_13), .fluid_out(k_6_6), .air_in(c_7_1));
valve v_7_14 (.fluid_in(k_7_14), .fluid_out(k_6_7), .air_in(c_7_0));
valve v_7_15 (.fluid_in(k_7_15), .fluid_out(k_6_7), .air_in(c_7_1));
valve v_7_16 (.fluid_in(k_7_16), .fluid_out(k_6_8), .air_in(c_7_0));
valve v_7_17 (.fluid_in(k_7_17), .fluid_out(k_6_8), .air_in(c_7_1));
valve v_7_18 (.fluid_in(k_7_18), .fluid_out(k_6_9), .air_in(c_7_0));
valve v_7_19 (.fluid_in(k_7_19), .fluid_out(k_6_9), .air_in(c_7_1));
valve v_7_20 (.fluid_in(k_7_20), .fluid_out(k_6_10), .air_in(c_7_0));
valve v_7_21 (.fluid_in(k_7_21), .fluid_out(k_6_10), .air_in(c_7_1));
valve v_7_22 (.fluid_in(k_7_22), .fluid_out(k_6_11), .air_in(c_7_0));
valve v_7_23 (.fluid_in(k_7_23), .fluid_out(k_6_11), .air_in(c_7_1));
valve v_7_24 (.fluid_in(k_7_24), .fluid_out(k_6_12), .air_in(c_7_0));
valve v_7_25 (.fluid_in(k_7_25), .fluid_out(k_6_12), .air_in(c_7_1));
valve v_7_26 (.fluid_in(k_7_26), .fluid_out(k_6_13), .air_in(c_7_0));
valve v_7_27 (.fluid_in(k_7_27), .fluid_out(k_6_13), .air_in(c_7_1));
valve v_7_28 (.fluid_in(k_7_28), .fluid_out(k_6_14), .air_in(c_7_0));
valve v_7_29 (.fluid_in(k_7_29), .fluid_out(k_6_14), .air_in(c_7_1));
valve v_7_30 (.fluid_in(k_7_30), .fluid_out(k_6_15), .air_in(c_7_0));
valve v_7_31 (.fluid_in(k_7_31), .fluid_out(k_6_15), .air_in(c_7_1));
valve v_7_32 (.fluid_in(k_7_32), .fluid_out(k_6_16), .air_in(c_7_0));
valve v_7_33 (.fluid_in(k_7_33), .fluid_out(k_6_16), .air_in(c_7_1));
valve v_7_34 (.fluid_in(k_7_34), .fluid_out(k_6_17), .air_in(c_7_0));
valve v_7_35 (.fluid_in(k_7_35), .fluid_out(k_6_17), .air_in(c_7_1));
valve v_7_36 (.fluid_in(k_7_36), .fluid_out(k_6_18), .air_in(c_7_0));
valve v_7_37 (.fluid_in(k_7_37), .fluid_out(k_6_18), .air_in(c_7_1));
valve v_7_38 (.fluid_in(k_7_38), .fluid_out(k_6_19), .air_in(c_7_0));
valve v_7_39 (.fluid_in(k_7_39), .fluid_out(k_6_19), .air_in(c_7_1));
valve v_7_40 (.fluid_in(k_7_40), .fluid_out(k_6_20), .air_in(c_7_0));
valve v_7_41 (.fluid_in(k_7_41), .fluid_out(k_6_20), .air_in(c_7_1));
valve v_7_42 (.fluid_in(k_7_42), .fluid_out(k_6_21), .air_in(c_7_0));
valve v_7_43 (.fluid_in(k_7_43), .fluid_out(k_6_21), .air_in(c_7_1));
valve v_7_44 (.fluid_in(k_7_44), .fluid_out(k_6_22), .air_in(c_7_0));
valve v_7_45 (.fluid_in(k_7_45), .fluid_out(k_6_22), .air_in(c_7_1));
valve v_7_46 (.fluid_in(k_7_46), .fluid_out(k_6_23), .air_in(c_7_0));
valve v_7_47 (.fluid_in(k_7_47), .fluid_out(k_6_23), .air_in(c_7_1));
valve v_7_48 (.fluid_in(k_7_48), .fluid_out(k_6_24), .air_in(c_7_0));
valve v_7_49 (.fluid_in(k_7_49), .fluid_out(k_6_24), .air_in(c_7_1));
valve v_7_50 (.fluid_in(k_7_50), .fluid_out(k_6_25), .air_in(c_7_0));
valve v_7_51 (.fluid_in(k_7_51), .fluid_out(k_6_25), .air_in(c_7_1));
valve v_7_52 (.fluid_in(k_7_52), .fluid_out(k_6_26), .air_in(c_7_0));
valve v_7_53 (.fluid_in(k_7_53), .fluid_out(k_6_26), .air_in(c_7_1));
valve v_7_54 (.fluid_in(k_7_54), .fluid_out(k_6_27), .air_in(c_7_0));
valve v_7_55 (.fluid_in(k_7_55), .fluid_out(k_6_27), .air_in(c_7_1));
valve v_7_56 (.fluid_in(k_7_56), .fluid_out(k_6_28), .air_in(c_7_0));
valve v_7_57 (.fluid_in(k_7_57), .fluid_out(k_6_28), .air_in(c_7_1));
valve v_7_58 (.fluid_in(k_7_58), .fluid_out(k_6_29), .air_in(c_7_0));
valve v_7_59 (.fluid_in(k_7_59), .fluid_out(k_6_29), .air_in(c_7_1));
valve v_7_60 (.fluid_in(k_7_60), .fluid_out(k_6_30), .air_in(c_7_0));
valve v_7_61 (.fluid_in(k_7_61), .fluid_out(k_6_30), .air_in(c_7_1));
valve v_7_62 (.fluid_in(k_7_62), .fluid_out(k_6_31), .air_in(c_7_0));
valve v_7_63 (.fluid_in(k_7_63), .fluid_out(k_6_31), .air_in(c_7_1));
valve v_7_64 (.fluid_in(k_7_64), .fluid_out(k_6_32), .air_in(c_7_0));
valve v_7_65 (.fluid_in(k_7_65), .fluid_out(k_6_32), .air_in(c_7_1));
valve v_7_66 (.fluid_in(k_7_66), .fluid_out(k_6_33), .air_in(c_7_0));
valve v_7_67 (.fluid_in(k_7_67), .fluid_out(k_6_33), .air_in(c_7_1));
valve v_7_68 (.fluid_in(k_7_68), .fluid_out(k_6_34), .air_in(c_7_0));
valve v_7_69 (.fluid_in(k_7_69), .fluid_out(k_6_34), .air_in(c_7_1));
valve v_7_70 (.fluid_in(k_7_70), .fluid_out(k_6_35), .air_in(c_7_0));
valve v_7_71 (.fluid_in(k_7_71), .fluid_out(k_6_35), .air_in(c_7_1));
valve v_7_72 (.fluid_in(k_7_72), .fluid_out(k_6_36), .air_in(c_7_0));
valve v_7_73 (.fluid_in(k_7_73), .fluid_out(k_6_36), .air_in(c_7_1));
valve v_7_74 (.fluid_in(k_7_74), .fluid_out(k_6_37), .air_in(c_7_0));
valve v_7_75 (.fluid_in(k_7_75), .fluid_out(k_6_37), .air_in(c_7_1));
valve v_7_76 (.fluid_in(k_7_76), .fluid_out(k_6_38), .air_in(c_7_0));
valve v_7_77 (.fluid_in(k_7_77), .fluid_out(k_6_38), .air_in(c_7_1));
valve v_7_78 (.fluid_in(k_7_78), .fluid_out(k_6_39), .air_in(c_7_0));
valve v_7_79 (.fluid_in(k_7_79), .fluid_out(k_6_39), .air_in(c_7_1));
valve v_7_80 (.fluid_in(k_7_80), .fluid_out(k_6_40), .air_in(c_7_0));
valve v_7_81 (.fluid_in(k_7_81), .fluid_out(k_6_40), .air_in(c_7_1));
valve v_7_82 (.fluid_in(k_7_82), .fluid_out(k_6_41), .air_in(c_7_0));
valve v_7_83 (.fluid_in(k_7_83), .fluid_out(k_6_41), .air_in(c_7_1));
valve v_7_84 (.fluid_in(k_7_84), .fluid_out(k_6_42), .air_in(c_7_0));
valve v_7_85 (.fluid_in(k_7_85), .fluid_out(k_6_42), .air_in(c_7_1));
valve v_7_86 (.fluid_in(k_7_86), .fluid_out(k_6_43), .air_in(c_7_0));
valve v_7_87 (.fluid_in(k_7_87), .fluid_out(k_6_43), .air_in(c_7_1));
valve v_7_88 (.fluid_in(k_7_88), .fluid_out(k_6_44), .air_in(c_7_0));
valve v_7_89 (.fluid_in(k_7_89), .fluid_out(k_6_44), .air_in(c_7_1));
valve v_7_90 (.fluid_in(k_7_90), .fluid_out(k_6_45), .air_in(c_7_0));
valve v_7_91 (.fluid_in(k_7_91), .fluid_out(k_6_45), .air_in(c_7_1));
valve v_7_92 (.fluid_in(k_7_92), .fluid_out(k_6_46), .air_in(c_7_0));
valve v_7_93 (.fluid_in(k_7_93), .fluid_out(k_6_46), .air_in(c_7_1));
valve v_7_94 (.fluid_in(k_7_94), .fluid_out(k_6_47), .air_in(c_7_0));
valve v_7_95 (.fluid_in(k_7_95), .fluid_out(k_6_47), .air_in(c_7_1));
valve v_7_96 (.fluid_in(k_7_96), .fluid_out(k_6_48), .air_in(c_7_0));
valve v_7_97 (.fluid_in(k_7_97), .fluid_out(k_6_48), .air_in(c_7_1));
valve v_7_98 (.fluid_in(k_7_98), .fluid_out(k_6_49), .air_in(c_7_0));
valve v_7_99 (.fluid_in(k_7_99), .fluid_out(k_6_49), .air_in(c_7_1));
valve v_7_100 (.fluid_in(k_7_100), .fluid_out(k_6_50), .air_in(c_7_0));
valve v_7_101 (.fluid_in(k_7_101), .fluid_out(k_6_50), .air_in(c_7_1));
valve v_7_102 (.fluid_in(k_7_102), .fluid_out(k_6_51), .air_in(c_7_0));
valve v_7_103 (.fluid_in(k_7_103), .fluid_out(k_6_51), .air_in(c_7_1));
valve v_7_104 (.fluid_in(k_7_104), .fluid_out(k_6_52), .air_in(c_7_0));
valve v_7_105 (.fluid_in(k_7_105), .fluid_out(k_6_52), .air_in(c_7_1));
valve v_7_106 (.fluid_in(k_7_106), .fluid_out(k_6_53), .air_in(c_7_0));
valve v_7_107 (.fluid_in(k_7_107), .fluid_out(k_6_53), .air_in(c_7_1));
valve v_7_108 (.fluid_in(k_7_108), .fluid_out(k_6_54), .air_in(c_7_0));
valve v_7_109 (.fluid_in(k_7_109), .fluid_out(k_6_54), .air_in(c_7_1));
valve v_7_110 (.fluid_in(k_7_110), .fluid_out(k_6_55), .air_in(c_7_0));
valve v_7_111 (.fluid_in(k_7_111), .fluid_out(k_6_55), .air_in(c_7_1));
valve v_7_112 (.fluid_in(k_7_112), .fluid_out(k_6_56), .air_in(c_7_0));
valve v_7_113 (.fluid_in(k_7_113), .fluid_out(k_6_56), .air_in(c_7_1));
valve v_7_114 (.fluid_in(k_7_114), .fluid_out(k_6_57), .air_in(c_7_0));
valve v_7_115 (.fluid_in(k_7_115), .fluid_out(k_6_57), .air_in(c_7_1));
valve v_7_116 (.fluid_in(k_7_116), .fluid_out(k_6_58), .air_in(c_7_0));
valve v_7_117 (.fluid_in(k_7_117), .fluid_out(k_6_58), .air_in(c_7_1));
valve v_7_118 (.fluid_in(k_7_118), .fluid_out(k_6_59), .air_in(c_7_0));
valve v_7_119 (.fluid_in(k_7_119), .fluid_out(k_6_59), .air_in(c_7_1));
valve v_7_120 (.fluid_in(k_7_120), .fluid_out(k_6_60), .air_in(c_7_0));
valve v_7_121 (.fluid_in(k_7_121), .fluid_out(k_6_60), .air_in(c_7_1));
valve v_7_122 (.fluid_in(k_7_122), .fluid_out(k_6_61), .air_in(c_7_0));
valve v_7_123 (.fluid_in(k_7_123), .fluid_out(k_6_61), .air_in(c_7_1));
valve v_7_124 (.fluid_in(k_7_124), .fluid_out(k_6_62), .air_in(c_7_0));
valve v_7_125 (.fluid_in(k_7_125), .fluid_out(k_6_62), .air_in(c_7_1));
valve v_7_126 (.fluid_in(k_7_126), .fluid_out(k_6_63), .air_in(c_7_0));
valve v_7_127 (.fluid_in(k_7_127), .fluid_out(k_6_63), .air_in(c_7_1));
valve v_8_0 (.fluid_in(k_8_0), .fluid_out(k_7_0), .air_in(c_8_0));
valve v_8_1 (.fluid_in(k_8_1), .fluid_out(k_7_0), .air_in(c_8_1));
valve v_8_2 (.fluid_in(k_8_2), .fluid_out(k_7_1), .air_in(c_8_0));
valve v_8_3 (.fluid_in(k_8_3), .fluid_out(k_7_1), .air_in(c_8_1));
valve v_8_4 (.fluid_in(k_8_4), .fluid_out(k_7_2), .air_in(c_8_0));
valve v_8_5 (.fluid_in(k_8_5), .fluid_out(k_7_2), .air_in(c_8_1));
valve v_8_6 (.fluid_in(k_8_6), .fluid_out(k_7_3), .air_in(c_8_0));
valve v_8_7 (.fluid_in(k_8_7), .fluid_out(k_7_3), .air_in(c_8_1));
valve v_8_8 (.fluid_in(k_8_8), .fluid_out(k_7_4), .air_in(c_8_0));
valve v_8_9 (.fluid_in(k_8_9), .fluid_out(k_7_4), .air_in(c_8_1));
valve v_8_10 (.fluid_in(k_8_10), .fluid_out(k_7_5), .air_in(c_8_0));
valve v_8_11 (.fluid_in(k_8_11), .fluid_out(k_7_5), .air_in(c_8_1));
valve v_8_12 (.fluid_in(k_8_12), .fluid_out(k_7_6), .air_in(c_8_0));
valve v_8_13 (.fluid_in(k_8_13), .fluid_out(k_7_6), .air_in(c_8_1));
valve v_8_14 (.fluid_in(k_8_14), .fluid_out(k_7_7), .air_in(c_8_0));
valve v_8_15 (.fluid_in(k_8_15), .fluid_out(k_7_7), .air_in(c_8_1));
valve v_8_16 (.fluid_in(k_8_16), .fluid_out(k_7_8), .air_in(c_8_0));
valve v_8_17 (.fluid_in(k_8_17), .fluid_out(k_7_8), .air_in(c_8_1));
valve v_8_18 (.fluid_in(k_8_18), .fluid_out(k_7_9), .air_in(c_8_0));
valve v_8_19 (.fluid_in(k_8_19), .fluid_out(k_7_9), .air_in(c_8_1));
valve v_8_20 (.fluid_in(k_8_20), .fluid_out(k_7_10), .air_in(c_8_0));
valve v_8_21 (.fluid_in(k_8_21), .fluid_out(k_7_10), .air_in(c_8_1));
valve v_8_22 (.fluid_in(k_8_22), .fluid_out(k_7_11), .air_in(c_8_0));
valve v_8_23 (.fluid_in(k_8_23), .fluid_out(k_7_11), .air_in(c_8_1));
valve v_8_24 (.fluid_in(k_8_24), .fluid_out(k_7_12), .air_in(c_8_0));
valve v_8_25 (.fluid_in(k_8_25), .fluid_out(k_7_12), .air_in(c_8_1));
valve v_8_26 (.fluid_in(k_8_26), .fluid_out(k_7_13), .air_in(c_8_0));
valve v_8_27 (.fluid_in(k_8_27), .fluid_out(k_7_13), .air_in(c_8_1));
valve v_8_28 (.fluid_in(k_8_28), .fluid_out(k_7_14), .air_in(c_8_0));
valve v_8_29 (.fluid_in(k_8_29), .fluid_out(k_7_14), .air_in(c_8_1));
valve v_8_30 (.fluid_in(k_8_30), .fluid_out(k_7_15), .air_in(c_8_0));
valve v_8_31 (.fluid_in(k_8_31), .fluid_out(k_7_15), .air_in(c_8_1));
valve v_8_32 (.fluid_in(k_8_32), .fluid_out(k_7_16), .air_in(c_8_0));
valve v_8_33 (.fluid_in(k_8_33), .fluid_out(k_7_16), .air_in(c_8_1));
valve v_8_34 (.fluid_in(k_8_34), .fluid_out(k_7_17), .air_in(c_8_0));
valve v_8_35 (.fluid_in(k_8_35), .fluid_out(k_7_17), .air_in(c_8_1));
valve v_8_36 (.fluid_in(k_8_36), .fluid_out(k_7_18), .air_in(c_8_0));
valve v_8_37 (.fluid_in(k_8_37), .fluid_out(k_7_18), .air_in(c_8_1));
valve v_8_38 (.fluid_in(k_8_38), .fluid_out(k_7_19), .air_in(c_8_0));
valve v_8_39 (.fluid_in(k_8_39), .fluid_out(k_7_19), .air_in(c_8_1));
valve v_8_40 (.fluid_in(k_8_40), .fluid_out(k_7_20), .air_in(c_8_0));
valve v_8_41 (.fluid_in(k_8_41), .fluid_out(k_7_20), .air_in(c_8_1));
valve v_8_42 (.fluid_in(k_8_42), .fluid_out(k_7_21), .air_in(c_8_0));
valve v_8_43 (.fluid_in(k_8_43), .fluid_out(k_7_21), .air_in(c_8_1));
valve v_8_44 (.fluid_in(k_8_44), .fluid_out(k_7_22), .air_in(c_8_0));
valve v_8_45 (.fluid_in(k_8_45), .fluid_out(k_7_22), .air_in(c_8_1));
valve v_8_46 (.fluid_in(k_8_46), .fluid_out(k_7_23), .air_in(c_8_0));
valve v_8_47 (.fluid_in(k_8_47), .fluid_out(k_7_23), .air_in(c_8_1));
valve v_8_48 (.fluid_in(k_8_48), .fluid_out(k_7_24), .air_in(c_8_0));
valve v_8_49 (.fluid_in(k_8_49), .fluid_out(k_7_24), .air_in(c_8_1));
valve v_8_50 (.fluid_in(k_8_50), .fluid_out(k_7_25), .air_in(c_8_0));
valve v_8_51 (.fluid_in(k_8_51), .fluid_out(k_7_25), .air_in(c_8_1));
valve v_8_52 (.fluid_in(k_8_52), .fluid_out(k_7_26), .air_in(c_8_0));
valve v_8_53 (.fluid_in(k_8_53), .fluid_out(k_7_26), .air_in(c_8_1));
valve v_8_54 (.fluid_in(k_8_54), .fluid_out(k_7_27), .air_in(c_8_0));
valve v_8_55 (.fluid_in(k_8_55), .fluid_out(k_7_27), .air_in(c_8_1));
valve v_8_56 (.fluid_in(k_8_56), .fluid_out(k_7_28), .air_in(c_8_0));
valve v_8_57 (.fluid_in(k_8_57), .fluid_out(k_7_28), .air_in(c_8_1));
valve v_8_58 (.fluid_in(k_8_58), .fluid_out(k_7_29), .air_in(c_8_0));
valve v_8_59 (.fluid_in(k_8_59), .fluid_out(k_7_29), .air_in(c_8_1));
valve v_8_60 (.fluid_in(k_8_60), .fluid_out(k_7_30), .air_in(c_8_0));
valve v_8_61 (.fluid_in(k_8_61), .fluid_out(k_7_30), .air_in(c_8_1));
valve v_8_62 (.fluid_in(k_8_62), .fluid_out(k_7_31), .air_in(c_8_0));
valve v_8_63 (.fluid_in(k_8_63), .fluid_out(k_7_31), .air_in(c_8_1));
valve v_8_64 (.fluid_in(k_8_64), .fluid_out(k_7_32), .air_in(c_8_0));
valve v_8_65 (.fluid_in(k_8_65), .fluid_out(k_7_32), .air_in(c_8_1));
valve v_8_66 (.fluid_in(k_8_66), .fluid_out(k_7_33), .air_in(c_8_0));
valve v_8_67 (.fluid_in(k_8_67), .fluid_out(k_7_33), .air_in(c_8_1));
valve v_8_68 (.fluid_in(k_8_68), .fluid_out(k_7_34), .air_in(c_8_0));
valve v_8_69 (.fluid_in(k_8_69), .fluid_out(k_7_34), .air_in(c_8_1));
valve v_8_70 (.fluid_in(k_8_70), .fluid_out(k_7_35), .air_in(c_8_0));
valve v_8_71 (.fluid_in(k_8_71), .fluid_out(k_7_35), .air_in(c_8_1));
valve v_8_72 (.fluid_in(k_8_72), .fluid_out(k_7_36), .air_in(c_8_0));
valve v_8_73 (.fluid_in(k_8_73), .fluid_out(k_7_36), .air_in(c_8_1));
valve v_8_74 (.fluid_in(k_8_74), .fluid_out(k_7_37), .air_in(c_8_0));
valve v_8_75 (.fluid_in(k_8_75), .fluid_out(k_7_37), .air_in(c_8_1));
valve v_8_76 (.fluid_in(k_8_76), .fluid_out(k_7_38), .air_in(c_8_0));
valve v_8_77 (.fluid_in(k_8_77), .fluid_out(k_7_38), .air_in(c_8_1));
valve v_8_78 (.fluid_in(k_8_78), .fluid_out(k_7_39), .air_in(c_8_0));
valve v_8_79 (.fluid_in(k_8_79), .fluid_out(k_7_39), .air_in(c_8_1));
valve v_8_80 (.fluid_in(k_8_80), .fluid_out(k_7_40), .air_in(c_8_0));
valve v_8_81 (.fluid_in(k_8_81), .fluid_out(k_7_40), .air_in(c_8_1));
valve v_8_82 (.fluid_in(k_8_82), .fluid_out(k_7_41), .air_in(c_8_0));
valve v_8_83 (.fluid_in(k_8_83), .fluid_out(k_7_41), .air_in(c_8_1));
valve v_8_84 (.fluid_in(k_8_84), .fluid_out(k_7_42), .air_in(c_8_0));
valve v_8_85 (.fluid_in(k_8_85), .fluid_out(k_7_42), .air_in(c_8_1));
valve v_8_86 (.fluid_in(k_8_86), .fluid_out(k_7_43), .air_in(c_8_0));
valve v_8_87 (.fluid_in(k_8_87), .fluid_out(k_7_43), .air_in(c_8_1));
valve v_8_88 (.fluid_in(k_8_88), .fluid_out(k_7_44), .air_in(c_8_0));
valve v_8_89 (.fluid_in(k_8_89), .fluid_out(k_7_44), .air_in(c_8_1));
valve v_8_90 (.fluid_in(k_8_90), .fluid_out(k_7_45), .air_in(c_8_0));
valve v_8_91 (.fluid_in(k_8_91), .fluid_out(k_7_45), .air_in(c_8_1));
valve v_8_92 (.fluid_in(k_8_92), .fluid_out(k_7_46), .air_in(c_8_0));
valve v_8_93 (.fluid_in(k_8_93), .fluid_out(k_7_46), .air_in(c_8_1));
valve v_8_94 (.fluid_in(k_8_94), .fluid_out(k_7_47), .air_in(c_8_0));
valve v_8_95 (.fluid_in(k_8_95), .fluid_out(k_7_47), .air_in(c_8_1));
valve v_8_96 (.fluid_in(k_8_96), .fluid_out(k_7_48), .air_in(c_8_0));
valve v_8_97 (.fluid_in(k_8_97), .fluid_out(k_7_48), .air_in(c_8_1));
valve v_8_98 (.fluid_in(k_8_98), .fluid_out(k_7_49), .air_in(c_8_0));
valve v_8_99 (.fluid_in(k_8_99), .fluid_out(k_7_49), .air_in(c_8_1));
valve v_8_100 (.fluid_in(k_8_100), .fluid_out(k_7_50), .air_in(c_8_0));
valve v_8_101 (.fluid_in(k_8_101), .fluid_out(k_7_50), .air_in(c_8_1));
valve v_8_102 (.fluid_in(k_8_102), .fluid_out(k_7_51), .air_in(c_8_0));
valve v_8_103 (.fluid_in(k_8_103), .fluid_out(k_7_51), .air_in(c_8_1));
valve v_8_104 (.fluid_in(k_8_104), .fluid_out(k_7_52), .air_in(c_8_0));
valve v_8_105 (.fluid_in(k_8_105), .fluid_out(k_7_52), .air_in(c_8_1));
valve v_8_106 (.fluid_in(k_8_106), .fluid_out(k_7_53), .air_in(c_8_0));
valve v_8_107 (.fluid_in(k_8_107), .fluid_out(k_7_53), .air_in(c_8_1));
valve v_8_108 (.fluid_in(k_8_108), .fluid_out(k_7_54), .air_in(c_8_0));
valve v_8_109 (.fluid_in(k_8_109), .fluid_out(k_7_54), .air_in(c_8_1));
valve v_8_110 (.fluid_in(k_8_110), .fluid_out(k_7_55), .air_in(c_8_0));
valve v_8_111 (.fluid_in(k_8_111), .fluid_out(k_7_55), .air_in(c_8_1));
valve v_8_112 (.fluid_in(k_8_112), .fluid_out(k_7_56), .air_in(c_8_0));
valve v_8_113 (.fluid_in(k_8_113), .fluid_out(k_7_56), .air_in(c_8_1));
valve v_8_114 (.fluid_in(k_8_114), .fluid_out(k_7_57), .air_in(c_8_0));
valve v_8_115 (.fluid_in(k_8_115), .fluid_out(k_7_57), .air_in(c_8_1));
valve v_8_116 (.fluid_in(k_8_116), .fluid_out(k_7_58), .air_in(c_8_0));
valve v_8_117 (.fluid_in(k_8_117), .fluid_out(k_7_58), .air_in(c_8_1));
valve v_8_118 (.fluid_in(k_8_118), .fluid_out(k_7_59), .air_in(c_8_0));
valve v_8_119 (.fluid_in(k_8_119), .fluid_out(k_7_59), .air_in(c_8_1));
valve v_8_120 (.fluid_in(k_8_120), .fluid_out(k_7_60), .air_in(c_8_0));
valve v_8_121 (.fluid_in(k_8_121), .fluid_out(k_7_60), .air_in(c_8_1));
valve v_8_122 (.fluid_in(k_8_122), .fluid_out(k_7_61), .air_in(c_8_0));
valve v_8_123 (.fluid_in(k_8_123), .fluid_out(k_7_61), .air_in(c_8_1));
valve v_8_124 (.fluid_in(k_8_124), .fluid_out(k_7_62), .air_in(c_8_0));
valve v_8_125 (.fluid_in(k_8_125), .fluid_out(k_7_62), .air_in(c_8_1));
valve v_8_126 (.fluid_in(k_8_126), .fluid_out(k_7_63), .air_in(c_8_0));
valve v_8_127 (.fluid_in(k_8_127), .fluid_out(k_7_63), .air_in(c_8_1));
valve v_8_128 (.fluid_in(k_8_128), .fluid_out(k_7_64), .air_in(c_8_0));
valve v_8_129 (.fluid_in(k_8_129), .fluid_out(k_7_64), .air_in(c_8_1));
valve v_8_130 (.fluid_in(k_8_130), .fluid_out(k_7_65), .air_in(c_8_0));
valve v_8_131 (.fluid_in(k_8_131), .fluid_out(k_7_65), .air_in(c_8_1));
valve v_8_132 (.fluid_in(k_8_132), .fluid_out(k_7_66), .air_in(c_8_0));
valve v_8_133 (.fluid_in(k_8_133), .fluid_out(k_7_66), .air_in(c_8_1));
valve v_8_134 (.fluid_in(k_8_134), .fluid_out(k_7_67), .air_in(c_8_0));
valve v_8_135 (.fluid_in(k_8_135), .fluid_out(k_7_67), .air_in(c_8_1));
valve v_8_136 (.fluid_in(k_8_136), .fluid_out(k_7_68), .air_in(c_8_0));
valve v_8_137 (.fluid_in(k_8_137), .fluid_out(k_7_68), .air_in(c_8_1));
valve v_8_138 (.fluid_in(k_8_138), .fluid_out(k_7_69), .air_in(c_8_0));
valve v_8_139 (.fluid_in(k_8_139), .fluid_out(k_7_69), .air_in(c_8_1));
valve v_8_140 (.fluid_in(k_8_140), .fluid_out(k_7_70), .air_in(c_8_0));
valve v_8_141 (.fluid_in(k_8_141), .fluid_out(k_7_70), .air_in(c_8_1));
valve v_8_142 (.fluid_in(k_8_142), .fluid_out(k_7_71), .air_in(c_8_0));
valve v_8_143 (.fluid_in(k_8_143), .fluid_out(k_7_71), .air_in(c_8_1));
valve v_8_144 (.fluid_in(k_8_144), .fluid_out(k_7_72), .air_in(c_8_0));
valve v_8_145 (.fluid_in(k_8_145), .fluid_out(k_7_72), .air_in(c_8_1));
valve v_8_146 (.fluid_in(k_8_146), .fluid_out(k_7_73), .air_in(c_8_0));
valve v_8_147 (.fluid_in(k_8_147), .fluid_out(k_7_73), .air_in(c_8_1));
valve v_8_148 (.fluid_in(k_8_148), .fluid_out(k_7_74), .air_in(c_8_0));
valve v_8_149 (.fluid_in(k_8_149), .fluid_out(k_7_74), .air_in(c_8_1));
valve v_8_150 (.fluid_in(k_8_150), .fluid_out(k_7_75), .air_in(c_8_0));
valve v_8_151 (.fluid_in(k_8_151), .fluid_out(k_7_75), .air_in(c_8_1));
valve v_8_152 (.fluid_in(k_8_152), .fluid_out(k_7_76), .air_in(c_8_0));
valve v_8_153 (.fluid_in(k_8_153), .fluid_out(k_7_76), .air_in(c_8_1));
valve v_8_154 (.fluid_in(k_8_154), .fluid_out(k_7_77), .air_in(c_8_0));
valve v_8_155 (.fluid_in(k_8_155), .fluid_out(k_7_77), .air_in(c_8_1));
valve v_8_156 (.fluid_in(k_8_156), .fluid_out(k_7_78), .air_in(c_8_0));
valve v_8_157 (.fluid_in(k_8_157), .fluid_out(k_7_78), .air_in(c_8_1));
valve v_8_158 (.fluid_in(k_8_158), .fluid_out(k_7_79), .air_in(c_8_0));
valve v_8_159 (.fluid_in(k_8_159), .fluid_out(k_7_79), .air_in(c_8_1));
valve v_8_160 (.fluid_in(k_8_160), .fluid_out(k_7_80), .air_in(c_8_0));
valve v_8_161 (.fluid_in(k_8_161), .fluid_out(k_7_80), .air_in(c_8_1));
valve v_8_162 (.fluid_in(k_8_162), .fluid_out(k_7_81), .air_in(c_8_0));
valve v_8_163 (.fluid_in(k_8_163), .fluid_out(k_7_81), .air_in(c_8_1));
valve v_8_164 (.fluid_in(k_8_164), .fluid_out(k_7_82), .air_in(c_8_0));
valve v_8_165 (.fluid_in(k_8_165), .fluid_out(k_7_82), .air_in(c_8_1));
valve v_8_166 (.fluid_in(k_8_166), .fluid_out(k_7_83), .air_in(c_8_0));
valve v_8_167 (.fluid_in(k_8_167), .fluid_out(k_7_83), .air_in(c_8_1));
valve v_8_168 (.fluid_in(k_8_168), .fluid_out(k_7_84), .air_in(c_8_0));
valve v_8_169 (.fluid_in(k_8_169), .fluid_out(k_7_84), .air_in(c_8_1));
valve v_8_170 (.fluid_in(k_8_170), .fluid_out(k_7_85), .air_in(c_8_0));
valve v_8_171 (.fluid_in(k_8_171), .fluid_out(k_7_85), .air_in(c_8_1));
valve v_8_172 (.fluid_in(k_8_172), .fluid_out(k_7_86), .air_in(c_8_0));
valve v_8_173 (.fluid_in(k_8_173), .fluid_out(k_7_86), .air_in(c_8_1));
valve v_8_174 (.fluid_in(k_8_174), .fluid_out(k_7_87), .air_in(c_8_0));
valve v_8_175 (.fluid_in(k_8_175), .fluid_out(k_7_87), .air_in(c_8_1));
valve v_8_176 (.fluid_in(k_8_176), .fluid_out(k_7_88), .air_in(c_8_0));
valve v_8_177 (.fluid_in(k_8_177), .fluid_out(k_7_88), .air_in(c_8_1));
valve v_8_178 (.fluid_in(k_8_178), .fluid_out(k_7_89), .air_in(c_8_0));
valve v_8_179 (.fluid_in(k_8_179), .fluid_out(k_7_89), .air_in(c_8_1));
valve v_8_180 (.fluid_in(k_8_180), .fluid_out(k_7_90), .air_in(c_8_0));
valve v_8_181 (.fluid_in(k_8_181), .fluid_out(k_7_90), .air_in(c_8_1));
valve v_8_182 (.fluid_in(k_8_182), .fluid_out(k_7_91), .air_in(c_8_0));
valve v_8_183 (.fluid_in(k_8_183), .fluid_out(k_7_91), .air_in(c_8_1));
valve v_8_184 (.fluid_in(k_8_184), .fluid_out(k_7_92), .air_in(c_8_0));
valve v_8_185 (.fluid_in(k_8_185), .fluid_out(k_7_92), .air_in(c_8_1));
valve v_8_186 (.fluid_in(k_8_186), .fluid_out(k_7_93), .air_in(c_8_0));
valve v_8_187 (.fluid_in(k_8_187), .fluid_out(k_7_93), .air_in(c_8_1));
valve v_8_188 (.fluid_in(k_8_188), .fluid_out(k_7_94), .air_in(c_8_0));
valve v_8_189 (.fluid_in(k_8_189), .fluid_out(k_7_94), .air_in(c_8_1));
valve v_8_190 (.fluid_in(k_8_190), .fluid_out(k_7_95), .air_in(c_8_0));
valve v_8_191 (.fluid_in(k_8_191), .fluid_out(k_7_95), .air_in(c_8_1));
valve v_8_192 (.fluid_in(k_8_192), .fluid_out(k_7_96), .air_in(c_8_0));
valve v_8_193 (.fluid_in(k_8_193), .fluid_out(k_7_96), .air_in(c_8_1));
valve v_8_194 (.fluid_in(k_8_194), .fluid_out(k_7_97), .air_in(c_8_0));
valve v_8_195 (.fluid_in(k_8_195), .fluid_out(k_7_97), .air_in(c_8_1));
valve v_8_196 (.fluid_in(k_8_196), .fluid_out(k_7_98), .air_in(c_8_0));
valve v_8_197 (.fluid_in(k_8_197), .fluid_out(k_7_98), .air_in(c_8_1));
valve v_8_198 (.fluid_in(k_8_198), .fluid_out(k_7_99), .air_in(c_8_0));
valve v_8_199 (.fluid_in(k_8_199), .fluid_out(k_7_99), .air_in(c_8_1));
valve v_8_200 (.fluid_in(k_8_200), .fluid_out(k_7_100), .air_in(c_8_0));
valve v_8_201 (.fluid_in(k_8_201), .fluid_out(k_7_100), .air_in(c_8_1));
valve v_8_202 (.fluid_in(k_8_202), .fluid_out(k_7_101), .air_in(c_8_0));
valve v_8_203 (.fluid_in(k_8_203), .fluid_out(k_7_101), .air_in(c_8_1));
valve v_8_204 (.fluid_in(k_8_204), .fluid_out(k_7_102), .air_in(c_8_0));
valve v_8_205 (.fluid_in(k_8_205), .fluid_out(k_7_102), .air_in(c_8_1));
valve v_8_206 (.fluid_in(k_8_206), .fluid_out(k_7_103), .air_in(c_8_0));
valve v_8_207 (.fluid_in(k_8_207), .fluid_out(k_7_103), .air_in(c_8_1));
valve v_8_208 (.fluid_in(k_8_208), .fluid_out(k_7_104), .air_in(c_8_0));
valve v_8_209 (.fluid_in(k_8_209), .fluid_out(k_7_104), .air_in(c_8_1));
valve v_8_210 (.fluid_in(k_8_210), .fluid_out(k_7_105), .air_in(c_8_0));
valve v_8_211 (.fluid_in(k_8_211), .fluid_out(k_7_105), .air_in(c_8_1));
valve v_8_212 (.fluid_in(k_8_212), .fluid_out(k_7_106), .air_in(c_8_0));
valve v_8_213 (.fluid_in(k_8_213), .fluid_out(k_7_106), .air_in(c_8_1));
valve v_8_214 (.fluid_in(k_8_214), .fluid_out(k_7_107), .air_in(c_8_0));
valve v_8_215 (.fluid_in(k_8_215), .fluid_out(k_7_107), .air_in(c_8_1));
valve v_8_216 (.fluid_in(k_8_216), .fluid_out(k_7_108), .air_in(c_8_0));
valve v_8_217 (.fluid_in(k_8_217), .fluid_out(k_7_108), .air_in(c_8_1));
valve v_8_218 (.fluid_in(k_8_218), .fluid_out(k_7_109), .air_in(c_8_0));
valve v_8_219 (.fluid_in(k_8_219), .fluid_out(k_7_109), .air_in(c_8_1));
valve v_8_220 (.fluid_in(k_8_220), .fluid_out(k_7_110), .air_in(c_8_0));
valve v_8_221 (.fluid_in(k_8_221), .fluid_out(k_7_110), .air_in(c_8_1));
valve v_8_222 (.fluid_in(k_8_222), .fluid_out(k_7_111), .air_in(c_8_0));
valve v_8_223 (.fluid_in(k_8_223), .fluid_out(k_7_111), .air_in(c_8_1));
valve v_8_224 (.fluid_in(k_8_224), .fluid_out(k_7_112), .air_in(c_8_0));
valve v_8_225 (.fluid_in(k_8_225), .fluid_out(k_7_112), .air_in(c_8_1));
valve v_8_226 (.fluid_in(k_8_226), .fluid_out(k_7_113), .air_in(c_8_0));
valve v_8_227 (.fluid_in(k_8_227), .fluid_out(k_7_113), .air_in(c_8_1));
valve v_8_228 (.fluid_in(k_8_228), .fluid_out(k_7_114), .air_in(c_8_0));
valve v_8_229 (.fluid_in(k_8_229), .fluid_out(k_7_114), .air_in(c_8_1));
valve v_8_230 (.fluid_in(k_8_230), .fluid_out(k_7_115), .air_in(c_8_0));
valve v_8_231 (.fluid_in(k_8_231), .fluid_out(k_7_115), .air_in(c_8_1));
valve v_8_232 (.fluid_in(k_8_232), .fluid_out(k_7_116), .air_in(c_8_0));
valve v_8_233 (.fluid_in(k_8_233), .fluid_out(k_7_116), .air_in(c_8_1));
valve v_8_234 (.fluid_in(k_8_234), .fluid_out(k_7_117), .air_in(c_8_0));
valve v_8_235 (.fluid_in(k_8_235), .fluid_out(k_7_117), .air_in(c_8_1));
valve v_8_236 (.fluid_in(k_8_236), .fluid_out(k_7_118), .air_in(c_8_0));
valve v_8_237 (.fluid_in(k_8_237), .fluid_out(k_7_118), .air_in(c_8_1));
valve v_8_238 (.fluid_in(k_8_238), .fluid_out(k_7_119), .air_in(c_8_0));
valve v_8_239 (.fluid_in(k_8_239), .fluid_out(k_7_119), .air_in(c_8_1));
valve v_8_240 (.fluid_in(k_8_240), .fluid_out(k_7_120), .air_in(c_8_0));
valve v_8_241 (.fluid_in(k_8_241), .fluid_out(k_7_120), .air_in(c_8_1));
valve v_8_242 (.fluid_in(k_8_242), .fluid_out(k_7_121), .air_in(c_8_0));
valve v_8_243 (.fluid_in(k_8_243), .fluid_out(k_7_121), .air_in(c_8_1));
valve v_8_244 (.fluid_in(k_8_244), .fluid_out(k_7_122), .air_in(c_8_0));
valve v_8_245 (.fluid_in(k_8_245), .fluid_out(k_7_122), .air_in(c_8_1));
valve v_8_246 (.fluid_in(k_8_246), .fluid_out(k_7_123), .air_in(c_8_0));
valve v_8_247 (.fluid_in(k_8_247), .fluid_out(k_7_123), .air_in(c_8_1));
valve v_8_248 (.fluid_in(k_8_248), .fluid_out(k_7_124), .air_in(c_8_0));
valve v_8_249 (.fluid_in(k_8_249), .fluid_out(k_7_124), .air_in(c_8_1));
valve v_8_250 (.fluid_in(k_8_250), .fluid_out(k_7_125), .air_in(c_8_0));
valve v_8_251 (.fluid_in(k_8_251), .fluid_out(k_7_125), .air_in(c_8_1));
valve v_8_252 (.fluid_in(k_8_252), .fluid_out(k_7_126), .air_in(c_8_0));
valve v_8_253 (.fluid_in(k_8_253), .fluid_out(k_7_126), .air_in(c_8_1));
valve v_8_254 (.fluid_in(k_8_254), .fluid_out(k_7_127), .air_in(c_8_0));
valve v_8_255 (.fluid_in(k_8_255), .fluid_out(k_7_127), .air_in(c_8_1));
endmodule
