module complete_8 (
inout io_0,inout io_1,inout io_2,inout io_3,inout io_4,inout io_5,inout io_6,inout io_7
);
assign io_0 = input_0;
assign io_0 = input_1;
assign io_0 = input_2;
assign io_0 = input_3;
assign io_0 = input_4;
assign io_0 = input_5;
assign io_0 = input_6;
assign io_0 = input_7;
assign io_1 = input_1;
assign io_1 = input_2;
assign io_1 = input_3;
assign io_1 = input_4;
assign io_1 = input_5;
assign io_1 = input_6;
assign io_1 = input_7;
assign io_2 = input_2;
assign io_2 = input_3;
assign io_2 = input_4;
assign io_2 = input_5;
assign io_2 = input_6;
assign io_2 = input_7;
assign io_3 = input_3;
assign io_3 = input_4;
assign io_3 = input_5;
assign io_3 = input_6;
assign io_3 = input_7;
assign io_4 = input_4;
assign io_4 = input_5;
assign io_4 = input_6;
assign io_4 = input_7;
assign io_5 = input_5;
assign io_5 = input_6;
assign io_5 = input_7;
assign io_6 = input_6;
assign io_6 = input_7;
assign io_7 = input_7;
endmodule
