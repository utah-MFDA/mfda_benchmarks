module ljubljana();
	mixer m_0(.a(e_0_1), .b(e_0_2), .y(e_0_3));
	mixer m_1(.a(e_0_1), .b(e_1_108), .y(e_1_109));
	mixer m_2(.a(e_0_2), .b(e_2_106), .y(e_2_110));
	mixer m_3(.a(e_0_3), .b(e_3_107), .y(e_3_111));
	mixer m_4(.a(e_4_63), .b(e_4_64), .y(e_4_65));
	mixer m_5(.a(e_5_17), .b(e_5_48), .y(e_5_51));
	mixer m_6(.a(e_6_19), .b(e_6_49), .y(e_6_53));
	mixer m_7(.a(e_7_18), .b(e_7_50), .y(e_7_52));
	mixer m_8(.a(e_8_46), .b(e_8_51), .y(e_8_68));
	mixer m_9(.a(e_9_47), .b(e_9_53), .y(e_9_66));
	mixer m_10(.a(e_10_45), .b(e_10_52), .y(e_10_67));
	mixer m_11(.a(e_11_14), .b(e_11_45), .y(e_11_48));
	mixer m_12(.a(e_12_15), .b(e_12_47), .y(e_12_50));
	mixer m_13(.a(e_13_16), .b(e_13_46), .y(e_13_49));
	mixer m_14(.a(e_11_14), .b(e_14_28), .y(e_14_30));
	mixer m_15(.a(e_12_15), .b(e_15_27), .y(e_15_32));
	mixer m_16(.a(e_13_16), .b(e_16_29), .y(e_16_31));
	mixer m_17(.a(e_5_17), .b(e_17_22), .y(e_17_27));
	mixer m_18(.a(e_7_18), .b(e_18_23), .y(e_18_29));
	mixer m_19(.a(e_6_19), .b(e_19_21), .y(e_19_28));
	mixer m_20(.a(e_20_21), .b(e_20_22), .y(e_20_23));
	mixer m_21(.a(e_19_21), .b(e_20_21), .y(e_21_43));
	mixer m_22(.a(e_17_22), .b(e_20_22), .y(e_22_44));
	mixer m_23(.a(e_18_23), .b(e_20_23), .y(e_23_42));
	mixer m_24(.a(e_24_37), .b(e_24_54), .y(e_24_59));
	mixer m_25(.a(e_25_36), .b(e_25_56), .y(e_25_58));
	mixer m_26(.a(e_26_38), .b(e_26_55), .y(e_26_57));
	mixer m_27(.a(e_15_27), .b(e_17_27), .y(e_27_41));
	mixer m_28(.a(e_14_28), .b(e_19_28), .y(e_28_39));
	mixer m_29(.a(e_16_29), .b(e_18_29), .y(e_29_40));
	mixer m_30(.a(e_14_30), .b(e_30_40), .y(e_30_54));
	mixer m_31(.a(e_16_31), .b(e_31_41), .y(e_31_56));
	mixer m_32(.a(e_15_32), .b(e_32_39), .y(e_32_55));
	mixer m_33(.a(e_33_37), .b(e_33_44), .y(e_33_60));
	mixer m_34(.a(e_34_36), .b(e_34_43), .y(e_34_62));
	mixer m_35(.a(e_35_38), .b(e_35_42), .y(e_35_61));
	mixer m_36(.a(e_25_36), .b(e_34_36), .y(e_36_76));
	mixer m_37(.a(e_24_37), .b(e_33_37), .y(e_37_78));
	mixer m_38(.a(e_26_38), .b(e_35_38), .y(e_38_77));
	mixer m_39(.a(e_28_39), .b(e_32_39), .y(e_39_81));
	mixer m_40(.a(e_29_40), .b(e_30_40), .y(e_40_79));
	mixer m_41(.a(e_27_41), .b(e_31_41), .y(e_41_80));
	mixer m_42(.a(e_23_42), .b(e_35_42), .y(e_42_82));
	mixer m_43(.a(e_21_43), .b(e_34_43), .y(e_43_84));
	mixer m_44(.a(e_22_44), .b(e_33_44), .y(e_44_83));
	mixer m_45(.a(e_10_45), .b(e_11_45), .y(e_45_85));
	mixer m_46(.a(e_8_46), .b(e_13_46), .y(e_46_86));
	mixer m_47(.a(e_9_47), .b(e_12_47), .y(e_47_87));
	mixer m_48(.a(e_5_48), .b(e_11_48), .y(e_48_90));
	mixer m_49(.a(e_6_49), .b(e_13_49), .y(e_49_88));
	mixer m_50(.a(e_7_50), .b(e_12_50), .y(e_50_89));
	mixer m_51(.a(e_5_51), .b(e_8_51), .y(e_51_91));
	mixer m_52(.a(e_7_52), .b(e_10_52), .y(e_52_93));
	mixer m_53(.a(e_6_53), .b(e_9_53), .y(e_53_92));
	mixer m_54(.a(e_24_54), .b(e_30_54), .y(e_54_70));
	mixer m_55(.a(e_26_55), .b(e_32_55), .y(e_55_72));
	mixer m_56(.a(e_25_56), .b(e_31_56), .y(e_56_71));
	mixer m_57(.a(e_26_57), .b(e_57_75), .y(e_57_79));
	mixer m_58(.a(e_25_58), .b(e_58_74), .y(e_58_81));
	mixer m_59(.a(e_24_59), .b(e_59_73), .y(e_59_80));
	mixer m_60(.a(e_33_60), .b(e_60_76), .y(e_60_88));
	mixer m_61(.a(e_35_61), .b(e_61_78), .y(e_61_90));
	mixer m_62(.a(e_34_62), .b(e_62_77), .y(e_62_89));
	mixer m_63(.a(e_4_63), .b(e_63_82), .y(e_63_85));
	mixer m_64(.a(e_4_64), .b(e_64_84), .y(e_64_87));
	mixer m_65(.a(e_4_65), .b(e_65_83), .y(e_65_86));
	mixer m_66(.a(e_9_66), .b(e_66_74), .y(e_66_91));
	mixer m_67(.a(e_10_67), .b(e_67_75), .y(e_67_92));
	mixer m_68(.a(e_8_68), .b(e_68_73), .y(e_68_93));
	mixer m_69(.a(e_69_70), .b(e_69_71), .y(e_69_72));
	mixer m_70(.a(e_54_70), .b(e_69_70), .y(e_70_103));
	mixer m_71(.a(e_56_71), .b(e_69_71), .y(e_71_105));
	mixer m_72(.a(e_55_72), .b(e_69_72), .y(e_72_104));
	mixer m_73(.a(e_59_73), .b(e_68_73), .y(e_73_97));
	mixer m_74(.a(e_58_74), .b(e_66_74), .y(e_74_99));
	mixer m_75(.a(e_57_75), .b(e_67_75), .y(e_75_98));
	mixer m_76(.a(e_36_76), .b(e_60_76), .y(e_76_94));
	mixer m_77(.a(e_38_77), .b(e_62_77), .y(e_77_96));
	mixer m_78(.a(e_37_78), .b(e_61_78), .y(e_78_95));
	mixer m_79(.a(e_40_79), .b(e_57_79), .y(e_79_94));
	mixer m_80(.a(e_41_80), .b(e_59_80), .y(e_80_96));
	mixer m_81(.a(e_39_81), .b(e_58_81), .y(e_81_95));
	mixer m_82(.a(e_42_82), .b(e_63_82), .y(e_82_97));
	mixer m_83(.a(e_44_83), .b(e_65_83), .y(e_83_99));
	mixer m_84(.a(e_43_84), .b(e_64_84), .y(e_84_98));
	mixer m_85(.a(e_45_85), .b(e_63_85), .y(e_85_100));
	mixer m_86(.a(e_46_86), .b(e_65_86), .y(e_86_102));
	mixer m_87(.a(e_47_87), .b(e_64_87), .y(e_87_101));
	mixer m_88(.a(e_49_88), .b(e_60_88), .y(e_88_100));
	mixer m_89(.a(e_50_89), .b(e_62_89), .y(e_89_102));
	mixer m_90(.a(e_48_90), .b(e_61_90), .y(e_90_101));
	mixer m_91(.a(e_51_91), .b(e_66_91), .y(e_91_103));
	mixer m_92(.a(e_53_92), .b(e_67_92), .y(e_92_105));
	mixer m_93(.a(e_52_93), .b(e_68_93), .y(e_93_104));
	mixer m_94(.a(e_76_94), .b(e_79_94), .y(e_94_106));
	mixer m_95(.a(e_78_95), .b(e_81_95), .y(e_95_108));
	mixer m_96(.a(e_77_96), .b(e_80_96), .y(e_96_107));
	mixer m_97(.a(e_73_97), .b(e_82_97), .y(e_97_106));
	mixer m_98(.a(e_75_98), .b(e_84_98), .y(e_98_108));
	mixer m_99(.a(e_74_99), .b(e_83_99), .y(e_99_107));
	mixer m_100(.a(e_85_100), .b(e_88_100), .y(e_100_109));
	mixer m_101(.a(e_87_101), .b(e_90_101), .y(e_101_111));
	mixer m_102(.a(e_86_102), .b(e_89_102), .y(e_102_110));
	mixer m_103(.a(e_70_103), .b(e_91_103), .y(e_103_109));
	mixer m_104(.a(e_72_104), .b(e_93_104), .y(e_104_111));
	mixer m_105(.a(e_71_105), .b(e_92_105), .y(e_105_110));
	mixer m_106(.a(e_2_106), .b(e_94_106), .y(e_97_106));
	mixer m_107(.a(e_3_107), .b(e_96_107), .y(e_99_107));
	mixer m_108(.a(e_1_108), .b(e_95_108), .y(e_98_108));
	mixer m_109(.a(e_1_109), .b(e_100_109), .y(e_103_109));
	mixer m_110(.a(e_2_110), .b(e_102_110), .y(e_105_110));
	mixer m_111(.a(e_3_111), .b(e_101_111), .y(e_104_111));
wire e_0_1,
	e_0_2,
	e_0_3,
	e_1_108,
	e_1_109,
	e_2_106,
	e_2_110,
	e_3_107,
	e_3_111,
	e_4_63,
	e_4_64,
	e_4_65,
	e_5_17,
	e_5_48,
	e_5_51,
	e_6_19,
	e_6_49,
	e_6_53,
	e_7_18,
	e_7_50,
	e_7_52,
	e_8_46,
	e_8_51,
	e_8_68,
	e_9_47,
	e_9_53,
	e_9_66,
	e_10_45,
	e_10_52,
	e_10_67,
	e_11_14,
	e_11_45,
	e_11_48,
	e_12_15,
	e_12_47,
	e_12_50,
	e_13_16,
	e_13_46,
	e_13_49,
	e_14_28,
	e_14_30,
	e_15_27,
	e_15_32,
	e_16_29,
	e_16_31,
	e_17_22,
	e_17_27,
	e_18_23,
	e_18_29,
	e_19_21,
	e_19_28,
	e_20_21,
	e_20_22,
	e_20_23,
	e_21_43,
	e_22_44,
	e_23_42,
	e_24_37,
	e_24_54,
	e_24_59,
	e_25_36,
	e_25_56,
	e_25_58,
	e_26_38,
	e_26_55,
	e_26_57,
	e_27_41,
	e_28_39,
	e_29_40,
	e_30_40,
	e_30_54,
	e_31_41,
	e_31_56,
	e_32_39,
	e_32_55,
	e_33_37,
	e_33_44,
	e_33_60,
	e_34_36,
	e_34_43,
	e_34_62,
	e_35_38,
	e_35_42,
	e_35_61,
	e_36_76,
	e_37_78,
	e_38_77,
	e_39_81,
	e_40_79,
	e_41_80,
	e_42_82,
	e_43_84,
	e_44_83,
	e_45_85,
	e_46_86,
	e_47_87,
	e_48_90,
	e_49_88,
	e_50_89,
	e_51_91,
	e_52_93,
	e_53_92,
	e_54_70,
	e_55_72,
	e_56_71,
	e_57_75,
	e_57_79,
	e_58_74,
	e_58_81,
	e_59_73,
	e_59_80,
	e_60_76,
	e_60_88,
	e_61_78,
	e_61_90,
	e_62_77,
	e_62_89,
	e_63_82,
	e_63_85,
	e_64_84,
	e_64_87,
	e_65_83,
	e_65_86,
	e_66_74,
	e_66_91,
	e_67_75,
	e_67_92,
	e_68_73,
	e_68_93,
	e_69_70,
	e_69_71,
	e_69_72,
	e_70_103,
	e_71_105,
	e_72_104,
	e_73_97,
	e_74_99,
	e_75_98,
	e_76_94,
	e_77_96,
	e_78_95,
	e_79_94,
	e_80_96,
	e_81_95,
	e_82_97,
	e_83_99,
	e_84_98,
	e_85_100,
	e_86_102,
	e_87_101,
	e_88_100,
	e_89_102,
	e_90_101,
	e_91_103,
	e_92_105,
	e_93_104,
	e_94_106,
	e_95_108,
	e_96_107,
	e_97_106,
	e_98_108,
	e_99_107,
	e_100_109,
	e_101_111,
	e_102_110,
	e_103_109,
	e_104_111,
	e_105_110;
endmodule
