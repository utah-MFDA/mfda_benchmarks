module binary_tree_1_11 (
output out_0,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63,input input_64,input input_65,input input_66,input input_67,input input_68,input input_69,input input_70,input input_71,input input_72,input input_73,input input_74,input input_75,input input_76,input input_77,input input_78,input input_79,input input_80,input input_81,input input_82,input input_83,input input_84,input input_85,input input_86,input input_87,input input_88,input input_89,input input_90,input input_91,input input_92,input input_93,input input_94,input input_95,input input_96,input input_97,input input_98,input input_99,input input_100,input input_101,input input_102,input input_103,input input_104,input input_105,input input_106,input input_107,input input_108,input input_109,input input_110,input input_111,input input_112,input input_113,input input_114,input input_115,input input_116,input input_117,input input_118,input input_119,input input_120,input input_121,input input_122,input input_123,input input_124,input input_125,input input_126,input input_127,input input_128,input input_129,input input_130,input input_131,input input_132,input input_133,input input_134,input input_135,input input_136,input input_137,input input_138,input input_139,input input_140,input input_141,input input_142,input input_143,input input_144,input input_145,input input_146,input input_147,input input_148,input input_149,input input_150,input input_151,input input_152,input input_153,input input_154,input input_155,input input_156,input input_157,input input_158,input input_159,input input_160,input input_161,input input_162,input input_163,input input_164,input input_165,input input_166,input input_167,input input_168,input input_169,input input_170,input input_171,input input_172,input input_173,input input_174,input input_175,input input_176,input input_177,input input_178,input input_179,input input_180,input input_181,input input_182,input input_183,input input_184,input input_185,input input_186,input input_187,input input_188,input input_189,input input_190,input input_191,input input_192,input input_193,input input_194,input input_195,input input_196,input input_197,input input_198,input input_199,input input_200,input input_201,input input_202,input input_203,input input_204,input input_205,input input_206,input input_207,input input_208,input input_209,input input_210,input input_211,input input_212,input input_213,input input_214,input input_215,input input_216,input input_217,input input_218,input input_219,input input_220,input input_221,input input_222,input input_223,input input_224,input input_225,input input_226,input input_227,input input_228,input input_229,input input_230,input input_231,input input_232,input input_233,input input_234,input input_235,input input_236,input input_237,input input_238,input input_239,input input_240,input input_241,input input_242,input input_243,input input_244,input input_245,input input_246,input input_247,input input_248,input input_249,input input_250,input input_251,input input_252,input input_253,input input_254,input input_255,input input_256,input input_257,input input_258,input input_259,input input_260,input input_261,input input_262,input input_263,input input_264,input input_265,input input_266,input input_267,input input_268,input input_269,input input_270,input input_271,input input_272,input input_273,input input_274,input input_275,input input_276,input input_277,input input_278,input input_279,input input_280,input input_281,input input_282,input input_283,input input_284,input input_285,input input_286,input input_287,input input_288,input input_289,input input_290,input input_291,input input_292,input input_293,input input_294,input input_295,input input_296,input input_297,input input_298,input input_299,input input_300,input input_301,input input_302,input input_303,input input_304,input input_305,input input_306,input input_307,input input_308,input input_309,input input_310,input input_311,input input_312,input input_313,input input_314,input input_315,input input_316,input input_317,input input_318,input input_319,input input_320,input input_321,input input_322,input input_323,input input_324,input input_325,input input_326,input input_327,input input_328,input input_329,input input_330,input input_331,input input_332,input input_333,input input_334,input input_335,input input_336,input input_337,input input_338,input input_339,input input_340,input input_341,input input_342,input input_343,input input_344,input input_345,input input_346,input input_347,input input_348,input input_349,input input_350,input input_351,input input_352,input input_353,input input_354,input input_355,input input_356,input input_357,input input_358,input input_359,input input_360,input input_361,input input_362,input input_363,input input_364,input input_365,input input_366,input input_367,input input_368,input input_369,input input_370,input input_371,input input_372,input input_373,input input_374,input input_375,input input_376,input input_377,input input_378,input input_379,input input_380,input input_381,input input_382,input input_383,input input_384,input input_385,input input_386,input input_387,input input_388,input input_389,input input_390,input input_391,input input_392,input input_393,input input_394,input input_395,input input_396,input input_397,input input_398,input input_399,input input_400,input input_401,input input_402,input input_403,input input_404,input input_405,input input_406,input input_407,input input_408,input input_409,input input_410,input input_411,input input_412,input input_413,input input_414,input input_415,input input_416,input input_417,input input_418,input input_419,input input_420,input input_421,input input_422,input input_423,input input_424,input input_425,input input_426,input input_427,input input_428,input input_429,input input_430,input input_431,input input_432,input input_433,input input_434,input input_435,input input_436,input input_437,input input_438,input input_439,input input_440,input input_441,input input_442,input input_443,input input_444,input input_445,input input_446,input input_447,input input_448,input input_449,input input_450,input input_451,input input_452,input input_453,input input_454,input input_455,input input_456,input input_457,input input_458,input input_459,input input_460,input input_461,input input_462,input input_463,input input_464,input input_465,input input_466,input input_467,input input_468,input input_469,input input_470,input input_471,input input_472,input input_473,input input_474,input input_475,input input_476,input input_477,input input_478,input input_479,input input_480,input input_481,input input_482,input input_483,input input_484,input input_485,input input_486,input input_487,input input_488,input input_489,input input_490,input input_491,input input_492,input input_493,input input_494,input input_495,input input_496,input input_497,input input_498,input input_499,input input_500,input input_501,input input_502,input input_503,input input_504,input input_505,input input_506,input input_507,input input_508,input input_509,input input_510,input input_511,input input_512,input input_513,input input_514,input input_515,input input_516,input input_517,input input_518,input input_519,input input_520,input input_521,input input_522,input input_523,input input_524,input input_525,input input_526,input input_527,input input_528,input input_529,input input_530,input input_531,input input_532,input input_533,input input_534,input input_535,input input_536,input input_537,input input_538,input input_539,input input_540,input input_541,input input_542,input input_543,input input_544,input input_545,input input_546,input input_547,input input_548,input input_549,input input_550,input input_551,input input_552,input input_553,input input_554,input input_555,input input_556,input input_557,input input_558,input input_559,input input_560,input input_561,input input_562,input input_563,input input_564,input input_565,input input_566,input input_567,input input_568,input input_569,input input_570,input input_571,input input_572,input input_573,input input_574,input input_575,input input_576,input input_577,input input_578,input input_579,input input_580,input input_581,input input_582,input input_583,input input_584,input input_585,input input_586,input input_587,input input_588,input input_589,input input_590,input input_591,input input_592,input input_593,input input_594,input input_595,input input_596,input input_597,input input_598,input input_599,input input_600,input input_601,input input_602,input input_603,input input_604,input input_605,input input_606,input input_607,input input_608,input input_609,input input_610,input input_611,input input_612,input input_613,input input_614,input input_615,input input_616,input input_617,input input_618,input input_619,input input_620,input input_621,input input_622,input input_623,input input_624,input input_625,input input_626,input input_627,input input_628,input input_629,input input_630,input input_631,input input_632,input input_633,input input_634,input input_635,input input_636,input input_637,input input_638,input input_639,input input_640,input input_641,input input_642,input input_643,input input_644,input input_645,input input_646,input input_647,input input_648,input input_649,input input_650,input input_651,input input_652,input input_653,input input_654,input input_655,input input_656,input input_657,input input_658,input input_659,input input_660,input input_661,input input_662,input input_663,input input_664,input input_665,input input_666,input input_667,input input_668,input input_669,input input_670,input input_671,input input_672,input input_673,input input_674,input input_675,input input_676,input input_677,input input_678,input input_679,input input_680,input input_681,input input_682,input input_683,input input_684,input input_685,input input_686,input input_687,input input_688,input input_689,input input_690,input input_691,input input_692,input input_693,input input_694,input input_695,input input_696,input input_697,input input_698,input input_699,input input_700,input input_701,input input_702,input input_703,input input_704,input input_705,input input_706,input input_707,input input_708,input input_709,input input_710,input input_711,input input_712,input input_713,input input_714,input input_715,input input_716,input input_717,input input_718,input input_719,input input_720,input input_721,input input_722,input input_723,input input_724,input input_725,input input_726,input input_727,input input_728,input input_729,input input_730,input input_731,input input_732,input input_733,input input_734,input input_735,input input_736,input input_737,input input_738,input input_739,input input_740,input input_741,input input_742,input input_743,input input_744,input input_745,input input_746,input input_747,input input_748,input input_749,input input_750,input input_751,input input_752,input input_753,input input_754,input input_755,input input_756,input input_757,input input_758,input input_759,input input_760,input input_761,input input_762,input input_763,input input_764,input input_765,input input_766,input input_767,input input_768,input input_769,input input_770,input input_771,input input_772,input input_773,input input_774,input input_775,input input_776,input input_777,input input_778,input input_779,input input_780,input input_781,input input_782,input input_783,input input_784,input input_785,input input_786,input input_787,input input_788,input input_789,input input_790,input input_791,input input_792,input input_793,input input_794,input input_795,input input_796,input input_797,input input_798,input input_799,input input_800,input input_801,input input_802,input input_803,input input_804,input input_805,input input_806,input input_807,input input_808,input input_809,input input_810,input input_811,input input_812,input input_813,input input_814,input input_815,input input_816,input input_817,input input_818,input input_819,input input_820,input input_821,input input_822,input input_823,input input_824,input input_825,input input_826,input input_827,input input_828,input input_829,input input_830,input input_831,input input_832,input input_833,input input_834,input input_835,input input_836,input input_837,input input_838,input input_839,input input_840,input input_841,input input_842,input input_843,input input_844,input input_845,input input_846,input input_847,input input_848,input input_849,input input_850,input input_851,input input_852,input input_853,input input_854,input input_855,input input_856,input input_857,input input_858,input input_859,input input_860,input input_861,input input_862,input input_863,input input_864,input input_865,input input_866,input input_867,input input_868,input input_869,input input_870,input input_871,input input_872,input input_873,input input_874,input input_875,input input_876,input input_877,input input_878,input input_879,input input_880,input input_881,input input_882,input input_883,input input_884,input input_885,input input_886,input input_887,input input_888,input input_889,input input_890,input input_891,input input_892,input input_893,input input_894,input input_895,input input_896,input input_897,input input_898,input input_899,input input_900,input input_901,input input_902,input input_903,input input_904,input input_905,input input_906,input input_907,input input_908,input input_909,input input_910,input input_911,input input_912,input input_913,input input_914,input input_915,input input_916,input input_917,input input_918,input input_919,input input_920,input input_921,input input_922,input input_923,input input_924,input input_925,input input_926,input input_927,input input_928,input input_929,input input_930,input input_931,input input_932,input input_933,input input_934,input input_935,input input_936,input input_937,input input_938,input input_939,input input_940,input input_941,input input_942,input input_943,input input_944,input input_945,input input_946,input input_947,input input_948,input input_949,input input_950,input input_951,input input_952,input input_953,input input_954,input input_955,input input_956,input input_957,input input_958,input input_959,input input_960,input input_961,input input_962,input input_963,input input_964,input input_965,input input_966,input input_967,input input_968,input input_969,input input_970,input input_971,input input_972,input input_973,input input_974,input input_975,input input_976,input input_977,input input_978,input input_979,input input_980,input input_981,input input_982,input input_983,input input_984,input input_985,input input_986,input input_987,input input_988,input input_989,input input_990,input input_991,input input_992,input input_993,input input_994,input input_995,input input_996,input input_997,input input_998,input input_999,input input_1000,input input_1001,input input_1002,input input_1003,input input_1004,input input_1005,input input_1006,input input_1007,input input_1008,input input_1009,input input_1010,input input_1011,input input_1012,input input_1013,input input_1014,input input_1015,input input_1016,input input_1017,input input_1018,input input_1019,input input_1020,input input_1021,input input_1022,input input_1023,input input_1024,input input_1025,input input_1026,input input_1027,input input_1028,input input_1029,input input_1030,input input_1031,input input_1032,input input_1033,input input_1034,input input_1035,input input_1036,input input_1037,input input_1038,input input_1039,input input_1040,input input_1041,input input_1042,input input_1043,input input_1044,input input_1045,input input_1046,input input_1047,input input_1048,input input_1049,input input_1050,input input_1051,input input_1052,input input_1053,input input_1054,input input_1055,input input_1056,input input_1057,input input_1058,input input_1059,input input_1060,input input_1061,input input_1062,input input_1063,input input_1064,input input_1065,input input_1066,input input_1067,input input_1068,input input_1069,input input_1070,input input_1071,input input_1072,input input_1073,input input_1074,input input_1075,input input_1076,input input_1077,input input_1078,input input_1079,input input_1080,input input_1081,input input_1082,input input_1083,input input_1084,input input_1085,input input_1086,input input_1087,input input_1088,input input_1089,input input_1090,input input_1091,input input_1092,input input_1093,input input_1094,input input_1095,input input_1096,input input_1097,input input_1098,input input_1099,input input_1100,input input_1101,input input_1102,input input_1103,input input_1104,input input_1105,input input_1106,input input_1107,input input_1108,input input_1109,input input_1110,input input_1111,input input_1112,input input_1113,input input_1114,input input_1115,input input_1116,input input_1117,input input_1118,input input_1119,input input_1120,input input_1121,input input_1122,input input_1123,input input_1124,input input_1125,input input_1126,input input_1127,input input_1128,input input_1129,input input_1130,input input_1131,input input_1132,input input_1133,input input_1134,input input_1135,input input_1136,input input_1137,input input_1138,input input_1139,input input_1140,input input_1141,input input_1142,input input_1143,input input_1144,input input_1145,input input_1146,input input_1147,input input_1148,input input_1149,input input_1150,input input_1151,input input_1152,input input_1153,input input_1154,input input_1155,input input_1156,input input_1157,input input_1158,input input_1159,input input_1160,input input_1161,input input_1162,input input_1163,input input_1164,input input_1165,input input_1166,input input_1167,input input_1168,input input_1169,input input_1170,input input_1171,input input_1172,input input_1173,input input_1174,input input_1175,input input_1176,input input_1177,input input_1178,input input_1179,input input_1180,input input_1181,input input_1182,input input_1183,input input_1184,input input_1185,input input_1186,input input_1187,input input_1188,input input_1189,input input_1190,input input_1191,input input_1192,input input_1193,input input_1194,input input_1195,input input_1196,input input_1197,input input_1198,input input_1199,input input_1200,input input_1201,input input_1202,input input_1203,input input_1204,input input_1205,input input_1206,input input_1207,input input_1208,input input_1209,input input_1210,input input_1211,input input_1212,input input_1213,input input_1214,input input_1215,input input_1216,input input_1217,input input_1218,input input_1219,input input_1220,input input_1221,input input_1222,input input_1223,input input_1224,input input_1225,input input_1226,input input_1227,input input_1228,input input_1229,input input_1230,input input_1231,input input_1232,input input_1233,input input_1234,input input_1235,input input_1236,input input_1237,input input_1238,input input_1239,input input_1240,input input_1241,input input_1242,input input_1243,input input_1244,input input_1245,input input_1246,input input_1247,input input_1248,input input_1249,input input_1250,input input_1251,input input_1252,input input_1253,input input_1254,input input_1255,input input_1256,input input_1257,input input_1258,input input_1259,input input_1260,input input_1261,input input_1262,input input_1263,input input_1264,input input_1265,input input_1266,input input_1267,input input_1268,input input_1269,input input_1270,input input_1271,input input_1272,input input_1273,input input_1274,input input_1275,input input_1276,input input_1277,input input_1278,input input_1279,input input_1280,input input_1281,input input_1282,input input_1283,input input_1284,input input_1285,input input_1286,input input_1287,input input_1288,input input_1289,input input_1290,input input_1291,input input_1292,input input_1293,input input_1294,input input_1295,input input_1296,input input_1297,input input_1298,input input_1299,input input_1300,input input_1301,input input_1302,input input_1303,input input_1304,input input_1305,input input_1306,input input_1307,input input_1308,input input_1309,input input_1310,input input_1311,input input_1312,input input_1313,input input_1314,input input_1315,input input_1316,input input_1317,input input_1318,input input_1319,input input_1320,input input_1321,input input_1322,input input_1323,input input_1324,input input_1325,input input_1326,input input_1327,input input_1328,input input_1329,input input_1330,input input_1331,input input_1332,input input_1333,input input_1334,input input_1335,input input_1336,input input_1337,input input_1338,input input_1339,input input_1340,input input_1341,input input_1342,input input_1343,input input_1344,input input_1345,input input_1346,input input_1347,input input_1348,input input_1349,input input_1350,input input_1351,input input_1352,input input_1353,input input_1354,input input_1355,input input_1356,input input_1357,input input_1358,input input_1359,input input_1360,input input_1361,input input_1362,input input_1363,input input_1364,input input_1365,input input_1366,input input_1367,input input_1368,input input_1369,input input_1370,input input_1371,input input_1372,input input_1373,input input_1374,input input_1375,input input_1376,input input_1377,input input_1378,input input_1379,input input_1380,input input_1381,input input_1382,input input_1383,input input_1384,input input_1385,input input_1386,input input_1387,input input_1388,input input_1389,input input_1390,input input_1391,input input_1392,input input_1393,input input_1394,input input_1395,input input_1396,input input_1397,input input_1398,input input_1399,input input_1400,input input_1401,input input_1402,input input_1403,input input_1404,input input_1405,input input_1406,input input_1407,input input_1408,input input_1409,input input_1410,input input_1411,input input_1412,input input_1413,input input_1414,input input_1415,input input_1416,input input_1417,input input_1418,input input_1419,input input_1420,input input_1421,input input_1422,input input_1423,input input_1424,input input_1425,input input_1426,input input_1427,input input_1428,input input_1429,input input_1430,input input_1431,input input_1432,input input_1433,input input_1434,input input_1435,input input_1436,input input_1437,input input_1438,input input_1439,input input_1440,input input_1441,input input_1442,input input_1443,input input_1444,input input_1445,input input_1446,input input_1447,input input_1448,input input_1449,input input_1450,input input_1451,input input_1452,input input_1453,input input_1454,input input_1455,input input_1456,input input_1457,input input_1458,input input_1459,input input_1460,input input_1461,input input_1462,input input_1463,input input_1464,input input_1465,input input_1466,input input_1467,input input_1468,input input_1469,input input_1470,input input_1471,input input_1472,input input_1473,input input_1474,input input_1475,input input_1476,input input_1477,input input_1478,input input_1479,input input_1480,input input_1481,input input_1482,input input_1483,input input_1484,input input_1485,input input_1486,input input_1487,input input_1488,input input_1489,input input_1490,input input_1491,input input_1492,input input_1493,input input_1494,input input_1495,input input_1496,input input_1497,input input_1498,input input_1499,input input_1500,input input_1501,input input_1502,input input_1503,input input_1504,input input_1505,input input_1506,input input_1507,input input_1508,input input_1509,input input_1510,input input_1511,input input_1512,input input_1513,input input_1514,input input_1515,input input_1516,input input_1517,input input_1518,input input_1519,input input_1520,input input_1521,input input_1522,input input_1523,input input_1524,input input_1525,input input_1526,input input_1527,input input_1528,input input_1529,input input_1530,input input_1531,input input_1532,input input_1533,input input_1534,input input_1535,input input_1536,input input_1537,input input_1538,input input_1539,input input_1540,input input_1541,input input_1542,input input_1543,input input_1544,input input_1545,input input_1546,input input_1547,input input_1548,input input_1549,input input_1550,input input_1551,input input_1552,input input_1553,input input_1554,input input_1555,input input_1556,input input_1557,input input_1558,input input_1559,input input_1560,input input_1561,input input_1562,input input_1563,input input_1564,input input_1565,input input_1566,input input_1567,input input_1568,input input_1569,input input_1570,input input_1571,input input_1572,input input_1573,input input_1574,input input_1575,input input_1576,input input_1577,input input_1578,input input_1579,input input_1580,input input_1581,input input_1582,input input_1583,input input_1584,input input_1585,input input_1586,input input_1587,input input_1588,input input_1589,input input_1590,input input_1591,input input_1592,input input_1593,input input_1594,input input_1595,input input_1596,input input_1597,input input_1598,input input_1599,input input_1600,input input_1601,input input_1602,input input_1603,input input_1604,input input_1605,input input_1606,input input_1607,input input_1608,input input_1609,input input_1610,input input_1611,input input_1612,input input_1613,input input_1614,input input_1615,input input_1616,input input_1617,input input_1618,input input_1619,input input_1620,input input_1621,input input_1622,input input_1623,input input_1624,input input_1625,input input_1626,input input_1627,input input_1628,input input_1629,input input_1630,input input_1631,input input_1632,input input_1633,input input_1634,input input_1635,input input_1636,input input_1637,input input_1638,input input_1639,input input_1640,input input_1641,input input_1642,input input_1643,input input_1644,input input_1645,input input_1646,input input_1647,input input_1648,input input_1649,input input_1650,input input_1651,input input_1652,input input_1653,input input_1654,input input_1655,input input_1656,input input_1657,input input_1658,input input_1659,input input_1660,input input_1661,input input_1662,input input_1663,input input_1664,input input_1665,input input_1666,input input_1667,input input_1668,input input_1669,input input_1670,input input_1671,input input_1672,input input_1673,input input_1674,input input_1675,input input_1676,input input_1677,input input_1678,input input_1679,input input_1680,input input_1681,input input_1682,input input_1683,input input_1684,input input_1685,input input_1686,input input_1687,input input_1688,input input_1689,input input_1690,input input_1691,input input_1692,input input_1693,input input_1694,input input_1695,input input_1696,input input_1697,input input_1698,input input_1699,input input_1700,input input_1701,input input_1702,input input_1703,input input_1704,input input_1705,input input_1706,input input_1707,input input_1708,input input_1709,input input_1710,input input_1711,input input_1712,input input_1713,input input_1714,input input_1715,input input_1716,input input_1717,input input_1718,input input_1719,input input_1720,input input_1721,input input_1722,input input_1723,input input_1724,input input_1725,input input_1726,input input_1727,input input_1728,input input_1729,input input_1730,input input_1731,input input_1732,input input_1733,input input_1734,input input_1735,input input_1736,input input_1737,input input_1738,input input_1739,input input_1740,input input_1741,input input_1742,input input_1743,input input_1744,input input_1745,input input_1746,input input_1747,input input_1748,input input_1749,input input_1750,input input_1751,input input_1752,input input_1753,input input_1754,input input_1755,input input_1756,input input_1757,input input_1758,input input_1759,input input_1760,input input_1761,input input_1762,input input_1763,input input_1764,input input_1765,input input_1766,input input_1767,input input_1768,input input_1769,input input_1770,input input_1771,input input_1772,input input_1773,input input_1774,input input_1775,input input_1776,input input_1777,input input_1778,input input_1779,input input_1780,input input_1781,input input_1782,input input_1783,input input_1784,input input_1785,input input_1786,input input_1787,input input_1788,input input_1789,input input_1790,input input_1791,input input_1792,input input_1793,input input_1794,input input_1795,input input_1796,input input_1797,input input_1798,input input_1799,input input_1800,input input_1801,input input_1802,input input_1803,input input_1804,input input_1805,input input_1806,input input_1807,input input_1808,input input_1809,input input_1810,input input_1811,input input_1812,input input_1813,input input_1814,input input_1815,input input_1816,input input_1817,input input_1818,input input_1819,input input_1820,input input_1821,input input_1822,input input_1823,input input_1824,input input_1825,input input_1826,input input_1827,input input_1828,input input_1829,input input_1830,input input_1831,input input_1832,input input_1833,input input_1834,input input_1835,input input_1836,input input_1837,input input_1838,input input_1839,input input_1840,input input_1841,input input_1842,input input_1843,input input_1844,input input_1845,input input_1846,input input_1847,input input_1848,input input_1849,input input_1850,input input_1851,input input_1852,input input_1853,input input_1854,input input_1855,input input_1856,input input_1857,input input_1858,input input_1859,input input_1860,input input_1861,input input_1862,input input_1863,input input_1864,input input_1865,input input_1866,input input_1867,input input_1868,input input_1869,input input_1870,input input_1871,input input_1872,input input_1873,input input_1874,input input_1875,input input_1876,input input_1877,input input_1878,input input_1879,input input_1880,input input_1881,input input_1882,input input_1883,input input_1884,input input_1885,input input_1886,input input_1887,input input_1888,input input_1889,input input_1890,input input_1891,input input_1892,input input_1893,input input_1894,input input_1895,input input_1896,input input_1897,input input_1898,input input_1899,input input_1900,input input_1901,input input_1902,input input_1903,input input_1904,input input_1905,input input_1906,input input_1907,input input_1908,input input_1909,input input_1910,input input_1911,input input_1912,input input_1913,input input_1914,input input_1915,input input_1916,input input_1917,input input_1918,input input_1919,input input_1920,input input_1921,input input_1922,input input_1923,input input_1924,input input_1925,input input_1926,input input_1927,input input_1928,input input_1929,input input_1930,input input_1931,input input_1932,input input_1933,input input_1934,input input_1935,input input_1936,input input_1937,input input_1938,input input_1939,input input_1940,input input_1941,input input_1942,input input_1943,input input_1944,input input_1945,input input_1946,input input_1947,input input_1948,input input_1949,input input_1950,input input_1951,input input_1952,input input_1953,input input_1954,input input_1955,input input_1956,input input_1957,input input_1958,input input_1959,input input_1960,input input_1961,input input_1962,input input_1963,input input_1964,input input_1965,input input_1966,input input_1967,input input_1968,input input_1969,input input_1970,input input_1971,input input_1972,input input_1973,input input_1974,input input_1975,input input_1976,input input_1977,input input_1978,input input_1979,input input_1980,input input_1981,input input_1982,input input_1983,input input_1984,input input_1985,input input_1986,input input_1987,input input_1988,input input_1989,input input_1990,input input_1991,input input_1992,input input_1993,input input_1994,input input_1995,input input_1996,input input_1997,input input_1998,input input_1999,input input_2000,input input_2001,input input_2002,input input_2003,input input_2004,input input_2005,input input_2006,input input_2007,input input_2008,input input_2009,input input_2010,input input_2011,input input_2012,input input_2013,input input_2014,input input_2015,input input_2016,input input_2017,input input_2018,input input_2019,input input_2020,input input_2021,input input_2022,input input_2023,input input_2024,input input_2025,input input_2026,input input_2027,input input_2028,input input_2029,input input_2030,input input_2031,input input_2032,input input_2033,input input_2034,input input_2035,input input_2036,input input_2037,input input_2038,input input_2039,input input_2040,input input_2041,input input_2042,input input_2043,input input_2044,input input_2045,input input_2046,input input_2047
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_000000 (.a(t0_0000000), .b(t0_0000001), .y(t0_000000));
wire t0_0000000, t0_0000001;
mixer mix_t0_0000000 (.a(t0_00000000), .b(t0_00000001), .y(t0_0000000));
wire t0_00000000, t0_00000001;
mixer mix_t0_00000000 (.a(t0_000000000), .b(t0_000000001), .y(t0_00000000));
wire t0_000000000, t0_000000001;
mixer mix_t0_000000000 (.a(t0_0000000000), .b(t0_0000000001), .y(t0_000000000));
wire t0_0000000000, t0_0000000001;
mixer mix_t0_0000000000 (.a(t0_00000000000), .b(t0_00000000001), .y(t0_0000000000));
wire t0_00000000000, t0_00000000001;
mixer mix_t0_00000000000 (.a(t0_000000000000), .b(t0_000000000001), .y(t0_00000000000));
wire t0_000000000000, t0_000000000001;
mixer mix_t0_00000000001 (.a(t0_000000000010), .b(t0_000000000011), .y(t0_00000000001));
wire t0_000000000010, t0_000000000011;
mixer mix_t0_0000000001 (.a(t0_00000000010), .b(t0_00000000011), .y(t0_0000000001));
wire t0_00000000010, t0_00000000011;
mixer mix_t0_00000000010 (.a(t0_000000000100), .b(t0_000000000101), .y(t0_00000000010));
wire t0_000000000100, t0_000000000101;
mixer mix_t0_00000000011 (.a(t0_000000000110), .b(t0_000000000111), .y(t0_00000000011));
wire t0_000000000110, t0_000000000111;
mixer mix_t0_000000001 (.a(t0_0000000010), .b(t0_0000000011), .y(t0_000000001));
wire t0_0000000010, t0_0000000011;
mixer mix_t0_0000000010 (.a(t0_00000000100), .b(t0_00000000101), .y(t0_0000000010));
wire t0_00000000100, t0_00000000101;
mixer mix_t0_00000000100 (.a(t0_000000001000), .b(t0_000000001001), .y(t0_00000000100));
wire t0_000000001000, t0_000000001001;
mixer mix_t0_00000000101 (.a(t0_000000001010), .b(t0_000000001011), .y(t0_00000000101));
wire t0_000000001010, t0_000000001011;
mixer mix_t0_0000000011 (.a(t0_00000000110), .b(t0_00000000111), .y(t0_0000000011));
wire t0_00000000110, t0_00000000111;
mixer mix_t0_00000000110 (.a(t0_000000001100), .b(t0_000000001101), .y(t0_00000000110));
wire t0_000000001100, t0_000000001101;
mixer mix_t0_00000000111 (.a(t0_000000001110), .b(t0_000000001111), .y(t0_00000000111));
wire t0_000000001110, t0_000000001111;
mixer mix_t0_00000001 (.a(t0_000000010), .b(t0_000000011), .y(t0_00000001));
wire t0_000000010, t0_000000011;
mixer mix_t0_000000010 (.a(t0_0000000100), .b(t0_0000000101), .y(t0_000000010));
wire t0_0000000100, t0_0000000101;
mixer mix_t0_0000000100 (.a(t0_00000001000), .b(t0_00000001001), .y(t0_0000000100));
wire t0_00000001000, t0_00000001001;
mixer mix_t0_00000001000 (.a(t0_000000010000), .b(t0_000000010001), .y(t0_00000001000));
wire t0_000000010000, t0_000000010001;
mixer mix_t0_00000001001 (.a(t0_000000010010), .b(t0_000000010011), .y(t0_00000001001));
wire t0_000000010010, t0_000000010011;
mixer mix_t0_0000000101 (.a(t0_00000001010), .b(t0_00000001011), .y(t0_0000000101));
wire t0_00000001010, t0_00000001011;
mixer mix_t0_00000001010 (.a(t0_000000010100), .b(t0_000000010101), .y(t0_00000001010));
wire t0_000000010100, t0_000000010101;
mixer mix_t0_00000001011 (.a(t0_000000010110), .b(t0_000000010111), .y(t0_00000001011));
wire t0_000000010110, t0_000000010111;
mixer mix_t0_000000011 (.a(t0_0000000110), .b(t0_0000000111), .y(t0_000000011));
wire t0_0000000110, t0_0000000111;
mixer mix_t0_0000000110 (.a(t0_00000001100), .b(t0_00000001101), .y(t0_0000000110));
wire t0_00000001100, t0_00000001101;
mixer mix_t0_00000001100 (.a(t0_000000011000), .b(t0_000000011001), .y(t0_00000001100));
wire t0_000000011000, t0_000000011001;
mixer mix_t0_00000001101 (.a(t0_000000011010), .b(t0_000000011011), .y(t0_00000001101));
wire t0_000000011010, t0_000000011011;
mixer mix_t0_0000000111 (.a(t0_00000001110), .b(t0_00000001111), .y(t0_0000000111));
wire t0_00000001110, t0_00000001111;
mixer mix_t0_00000001110 (.a(t0_000000011100), .b(t0_000000011101), .y(t0_00000001110));
wire t0_000000011100, t0_000000011101;
mixer mix_t0_00000001111 (.a(t0_000000011110), .b(t0_000000011111), .y(t0_00000001111));
wire t0_000000011110, t0_000000011111;
mixer mix_t0_0000001 (.a(t0_00000010), .b(t0_00000011), .y(t0_0000001));
wire t0_00000010, t0_00000011;
mixer mix_t0_00000010 (.a(t0_000000100), .b(t0_000000101), .y(t0_00000010));
wire t0_000000100, t0_000000101;
mixer mix_t0_000000100 (.a(t0_0000001000), .b(t0_0000001001), .y(t0_000000100));
wire t0_0000001000, t0_0000001001;
mixer mix_t0_0000001000 (.a(t0_00000010000), .b(t0_00000010001), .y(t0_0000001000));
wire t0_00000010000, t0_00000010001;
mixer mix_t0_00000010000 (.a(t0_000000100000), .b(t0_000000100001), .y(t0_00000010000));
wire t0_000000100000, t0_000000100001;
mixer mix_t0_00000010001 (.a(t0_000000100010), .b(t0_000000100011), .y(t0_00000010001));
wire t0_000000100010, t0_000000100011;
mixer mix_t0_0000001001 (.a(t0_00000010010), .b(t0_00000010011), .y(t0_0000001001));
wire t0_00000010010, t0_00000010011;
mixer mix_t0_00000010010 (.a(t0_000000100100), .b(t0_000000100101), .y(t0_00000010010));
wire t0_000000100100, t0_000000100101;
mixer mix_t0_00000010011 (.a(t0_000000100110), .b(t0_000000100111), .y(t0_00000010011));
wire t0_000000100110, t0_000000100111;
mixer mix_t0_000000101 (.a(t0_0000001010), .b(t0_0000001011), .y(t0_000000101));
wire t0_0000001010, t0_0000001011;
mixer mix_t0_0000001010 (.a(t0_00000010100), .b(t0_00000010101), .y(t0_0000001010));
wire t0_00000010100, t0_00000010101;
mixer mix_t0_00000010100 (.a(t0_000000101000), .b(t0_000000101001), .y(t0_00000010100));
wire t0_000000101000, t0_000000101001;
mixer mix_t0_00000010101 (.a(t0_000000101010), .b(t0_000000101011), .y(t0_00000010101));
wire t0_000000101010, t0_000000101011;
mixer mix_t0_0000001011 (.a(t0_00000010110), .b(t0_00000010111), .y(t0_0000001011));
wire t0_00000010110, t0_00000010111;
mixer mix_t0_00000010110 (.a(t0_000000101100), .b(t0_000000101101), .y(t0_00000010110));
wire t0_000000101100, t0_000000101101;
mixer mix_t0_00000010111 (.a(t0_000000101110), .b(t0_000000101111), .y(t0_00000010111));
wire t0_000000101110, t0_000000101111;
mixer mix_t0_00000011 (.a(t0_000000110), .b(t0_000000111), .y(t0_00000011));
wire t0_000000110, t0_000000111;
mixer mix_t0_000000110 (.a(t0_0000001100), .b(t0_0000001101), .y(t0_000000110));
wire t0_0000001100, t0_0000001101;
mixer mix_t0_0000001100 (.a(t0_00000011000), .b(t0_00000011001), .y(t0_0000001100));
wire t0_00000011000, t0_00000011001;
mixer mix_t0_00000011000 (.a(t0_000000110000), .b(t0_000000110001), .y(t0_00000011000));
wire t0_000000110000, t0_000000110001;
mixer mix_t0_00000011001 (.a(t0_000000110010), .b(t0_000000110011), .y(t0_00000011001));
wire t0_000000110010, t0_000000110011;
mixer mix_t0_0000001101 (.a(t0_00000011010), .b(t0_00000011011), .y(t0_0000001101));
wire t0_00000011010, t0_00000011011;
mixer mix_t0_00000011010 (.a(t0_000000110100), .b(t0_000000110101), .y(t0_00000011010));
wire t0_000000110100, t0_000000110101;
mixer mix_t0_00000011011 (.a(t0_000000110110), .b(t0_000000110111), .y(t0_00000011011));
wire t0_000000110110, t0_000000110111;
mixer mix_t0_000000111 (.a(t0_0000001110), .b(t0_0000001111), .y(t0_000000111));
wire t0_0000001110, t0_0000001111;
mixer mix_t0_0000001110 (.a(t0_00000011100), .b(t0_00000011101), .y(t0_0000001110));
wire t0_00000011100, t0_00000011101;
mixer mix_t0_00000011100 (.a(t0_000000111000), .b(t0_000000111001), .y(t0_00000011100));
wire t0_000000111000, t0_000000111001;
mixer mix_t0_00000011101 (.a(t0_000000111010), .b(t0_000000111011), .y(t0_00000011101));
wire t0_000000111010, t0_000000111011;
mixer mix_t0_0000001111 (.a(t0_00000011110), .b(t0_00000011111), .y(t0_0000001111));
wire t0_00000011110, t0_00000011111;
mixer mix_t0_00000011110 (.a(t0_000000111100), .b(t0_000000111101), .y(t0_00000011110));
wire t0_000000111100, t0_000000111101;
mixer mix_t0_00000011111 (.a(t0_000000111110), .b(t0_000000111111), .y(t0_00000011111));
wire t0_000000111110, t0_000000111111;
mixer mix_t0_000001 (.a(t0_0000010), .b(t0_0000011), .y(t0_000001));
wire t0_0000010, t0_0000011;
mixer mix_t0_0000010 (.a(t0_00000100), .b(t0_00000101), .y(t0_0000010));
wire t0_00000100, t0_00000101;
mixer mix_t0_00000100 (.a(t0_000001000), .b(t0_000001001), .y(t0_00000100));
wire t0_000001000, t0_000001001;
mixer mix_t0_000001000 (.a(t0_0000010000), .b(t0_0000010001), .y(t0_000001000));
wire t0_0000010000, t0_0000010001;
mixer mix_t0_0000010000 (.a(t0_00000100000), .b(t0_00000100001), .y(t0_0000010000));
wire t0_00000100000, t0_00000100001;
mixer mix_t0_00000100000 (.a(t0_000001000000), .b(t0_000001000001), .y(t0_00000100000));
wire t0_000001000000, t0_000001000001;
mixer mix_t0_00000100001 (.a(t0_000001000010), .b(t0_000001000011), .y(t0_00000100001));
wire t0_000001000010, t0_000001000011;
mixer mix_t0_0000010001 (.a(t0_00000100010), .b(t0_00000100011), .y(t0_0000010001));
wire t0_00000100010, t0_00000100011;
mixer mix_t0_00000100010 (.a(t0_000001000100), .b(t0_000001000101), .y(t0_00000100010));
wire t0_000001000100, t0_000001000101;
mixer mix_t0_00000100011 (.a(t0_000001000110), .b(t0_000001000111), .y(t0_00000100011));
wire t0_000001000110, t0_000001000111;
mixer mix_t0_000001001 (.a(t0_0000010010), .b(t0_0000010011), .y(t0_000001001));
wire t0_0000010010, t0_0000010011;
mixer mix_t0_0000010010 (.a(t0_00000100100), .b(t0_00000100101), .y(t0_0000010010));
wire t0_00000100100, t0_00000100101;
mixer mix_t0_00000100100 (.a(t0_000001001000), .b(t0_000001001001), .y(t0_00000100100));
wire t0_000001001000, t0_000001001001;
mixer mix_t0_00000100101 (.a(t0_000001001010), .b(t0_000001001011), .y(t0_00000100101));
wire t0_000001001010, t0_000001001011;
mixer mix_t0_0000010011 (.a(t0_00000100110), .b(t0_00000100111), .y(t0_0000010011));
wire t0_00000100110, t0_00000100111;
mixer mix_t0_00000100110 (.a(t0_000001001100), .b(t0_000001001101), .y(t0_00000100110));
wire t0_000001001100, t0_000001001101;
mixer mix_t0_00000100111 (.a(t0_000001001110), .b(t0_000001001111), .y(t0_00000100111));
wire t0_000001001110, t0_000001001111;
mixer mix_t0_00000101 (.a(t0_000001010), .b(t0_000001011), .y(t0_00000101));
wire t0_000001010, t0_000001011;
mixer mix_t0_000001010 (.a(t0_0000010100), .b(t0_0000010101), .y(t0_000001010));
wire t0_0000010100, t0_0000010101;
mixer mix_t0_0000010100 (.a(t0_00000101000), .b(t0_00000101001), .y(t0_0000010100));
wire t0_00000101000, t0_00000101001;
mixer mix_t0_00000101000 (.a(t0_000001010000), .b(t0_000001010001), .y(t0_00000101000));
wire t0_000001010000, t0_000001010001;
mixer mix_t0_00000101001 (.a(t0_000001010010), .b(t0_000001010011), .y(t0_00000101001));
wire t0_000001010010, t0_000001010011;
mixer mix_t0_0000010101 (.a(t0_00000101010), .b(t0_00000101011), .y(t0_0000010101));
wire t0_00000101010, t0_00000101011;
mixer mix_t0_00000101010 (.a(t0_000001010100), .b(t0_000001010101), .y(t0_00000101010));
wire t0_000001010100, t0_000001010101;
mixer mix_t0_00000101011 (.a(t0_000001010110), .b(t0_000001010111), .y(t0_00000101011));
wire t0_000001010110, t0_000001010111;
mixer mix_t0_000001011 (.a(t0_0000010110), .b(t0_0000010111), .y(t0_000001011));
wire t0_0000010110, t0_0000010111;
mixer mix_t0_0000010110 (.a(t0_00000101100), .b(t0_00000101101), .y(t0_0000010110));
wire t0_00000101100, t0_00000101101;
mixer mix_t0_00000101100 (.a(t0_000001011000), .b(t0_000001011001), .y(t0_00000101100));
wire t0_000001011000, t0_000001011001;
mixer mix_t0_00000101101 (.a(t0_000001011010), .b(t0_000001011011), .y(t0_00000101101));
wire t0_000001011010, t0_000001011011;
mixer mix_t0_0000010111 (.a(t0_00000101110), .b(t0_00000101111), .y(t0_0000010111));
wire t0_00000101110, t0_00000101111;
mixer mix_t0_00000101110 (.a(t0_000001011100), .b(t0_000001011101), .y(t0_00000101110));
wire t0_000001011100, t0_000001011101;
mixer mix_t0_00000101111 (.a(t0_000001011110), .b(t0_000001011111), .y(t0_00000101111));
wire t0_000001011110, t0_000001011111;
mixer mix_t0_0000011 (.a(t0_00000110), .b(t0_00000111), .y(t0_0000011));
wire t0_00000110, t0_00000111;
mixer mix_t0_00000110 (.a(t0_000001100), .b(t0_000001101), .y(t0_00000110));
wire t0_000001100, t0_000001101;
mixer mix_t0_000001100 (.a(t0_0000011000), .b(t0_0000011001), .y(t0_000001100));
wire t0_0000011000, t0_0000011001;
mixer mix_t0_0000011000 (.a(t0_00000110000), .b(t0_00000110001), .y(t0_0000011000));
wire t0_00000110000, t0_00000110001;
mixer mix_t0_00000110000 (.a(t0_000001100000), .b(t0_000001100001), .y(t0_00000110000));
wire t0_000001100000, t0_000001100001;
mixer mix_t0_00000110001 (.a(t0_000001100010), .b(t0_000001100011), .y(t0_00000110001));
wire t0_000001100010, t0_000001100011;
mixer mix_t0_0000011001 (.a(t0_00000110010), .b(t0_00000110011), .y(t0_0000011001));
wire t0_00000110010, t0_00000110011;
mixer mix_t0_00000110010 (.a(t0_000001100100), .b(t0_000001100101), .y(t0_00000110010));
wire t0_000001100100, t0_000001100101;
mixer mix_t0_00000110011 (.a(t0_000001100110), .b(t0_000001100111), .y(t0_00000110011));
wire t0_000001100110, t0_000001100111;
mixer mix_t0_000001101 (.a(t0_0000011010), .b(t0_0000011011), .y(t0_000001101));
wire t0_0000011010, t0_0000011011;
mixer mix_t0_0000011010 (.a(t0_00000110100), .b(t0_00000110101), .y(t0_0000011010));
wire t0_00000110100, t0_00000110101;
mixer mix_t0_00000110100 (.a(t0_000001101000), .b(t0_000001101001), .y(t0_00000110100));
wire t0_000001101000, t0_000001101001;
mixer mix_t0_00000110101 (.a(t0_000001101010), .b(t0_000001101011), .y(t0_00000110101));
wire t0_000001101010, t0_000001101011;
mixer mix_t0_0000011011 (.a(t0_00000110110), .b(t0_00000110111), .y(t0_0000011011));
wire t0_00000110110, t0_00000110111;
mixer mix_t0_00000110110 (.a(t0_000001101100), .b(t0_000001101101), .y(t0_00000110110));
wire t0_000001101100, t0_000001101101;
mixer mix_t0_00000110111 (.a(t0_000001101110), .b(t0_000001101111), .y(t0_00000110111));
wire t0_000001101110, t0_000001101111;
mixer mix_t0_00000111 (.a(t0_000001110), .b(t0_000001111), .y(t0_00000111));
wire t0_000001110, t0_000001111;
mixer mix_t0_000001110 (.a(t0_0000011100), .b(t0_0000011101), .y(t0_000001110));
wire t0_0000011100, t0_0000011101;
mixer mix_t0_0000011100 (.a(t0_00000111000), .b(t0_00000111001), .y(t0_0000011100));
wire t0_00000111000, t0_00000111001;
mixer mix_t0_00000111000 (.a(t0_000001110000), .b(t0_000001110001), .y(t0_00000111000));
wire t0_000001110000, t0_000001110001;
mixer mix_t0_00000111001 (.a(t0_000001110010), .b(t0_000001110011), .y(t0_00000111001));
wire t0_000001110010, t0_000001110011;
mixer mix_t0_0000011101 (.a(t0_00000111010), .b(t0_00000111011), .y(t0_0000011101));
wire t0_00000111010, t0_00000111011;
mixer mix_t0_00000111010 (.a(t0_000001110100), .b(t0_000001110101), .y(t0_00000111010));
wire t0_000001110100, t0_000001110101;
mixer mix_t0_00000111011 (.a(t0_000001110110), .b(t0_000001110111), .y(t0_00000111011));
wire t0_000001110110, t0_000001110111;
mixer mix_t0_000001111 (.a(t0_0000011110), .b(t0_0000011111), .y(t0_000001111));
wire t0_0000011110, t0_0000011111;
mixer mix_t0_0000011110 (.a(t0_00000111100), .b(t0_00000111101), .y(t0_0000011110));
wire t0_00000111100, t0_00000111101;
mixer mix_t0_00000111100 (.a(t0_000001111000), .b(t0_000001111001), .y(t0_00000111100));
wire t0_000001111000, t0_000001111001;
mixer mix_t0_00000111101 (.a(t0_000001111010), .b(t0_000001111011), .y(t0_00000111101));
wire t0_000001111010, t0_000001111011;
mixer mix_t0_0000011111 (.a(t0_00000111110), .b(t0_00000111111), .y(t0_0000011111));
wire t0_00000111110, t0_00000111111;
mixer mix_t0_00000111110 (.a(t0_000001111100), .b(t0_000001111101), .y(t0_00000111110));
wire t0_000001111100, t0_000001111101;
mixer mix_t0_00000111111 (.a(t0_000001111110), .b(t0_000001111111), .y(t0_00000111111));
wire t0_000001111110, t0_000001111111;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_000010 (.a(t0_0000100), .b(t0_0000101), .y(t0_000010));
wire t0_0000100, t0_0000101;
mixer mix_t0_0000100 (.a(t0_00001000), .b(t0_00001001), .y(t0_0000100));
wire t0_00001000, t0_00001001;
mixer mix_t0_00001000 (.a(t0_000010000), .b(t0_000010001), .y(t0_00001000));
wire t0_000010000, t0_000010001;
mixer mix_t0_000010000 (.a(t0_0000100000), .b(t0_0000100001), .y(t0_000010000));
wire t0_0000100000, t0_0000100001;
mixer mix_t0_0000100000 (.a(t0_00001000000), .b(t0_00001000001), .y(t0_0000100000));
wire t0_00001000000, t0_00001000001;
mixer mix_t0_00001000000 (.a(t0_000010000000), .b(t0_000010000001), .y(t0_00001000000));
wire t0_000010000000, t0_000010000001;
mixer mix_t0_00001000001 (.a(t0_000010000010), .b(t0_000010000011), .y(t0_00001000001));
wire t0_000010000010, t0_000010000011;
mixer mix_t0_0000100001 (.a(t0_00001000010), .b(t0_00001000011), .y(t0_0000100001));
wire t0_00001000010, t0_00001000011;
mixer mix_t0_00001000010 (.a(t0_000010000100), .b(t0_000010000101), .y(t0_00001000010));
wire t0_000010000100, t0_000010000101;
mixer mix_t0_00001000011 (.a(t0_000010000110), .b(t0_000010000111), .y(t0_00001000011));
wire t0_000010000110, t0_000010000111;
mixer mix_t0_000010001 (.a(t0_0000100010), .b(t0_0000100011), .y(t0_000010001));
wire t0_0000100010, t0_0000100011;
mixer mix_t0_0000100010 (.a(t0_00001000100), .b(t0_00001000101), .y(t0_0000100010));
wire t0_00001000100, t0_00001000101;
mixer mix_t0_00001000100 (.a(t0_000010001000), .b(t0_000010001001), .y(t0_00001000100));
wire t0_000010001000, t0_000010001001;
mixer mix_t0_00001000101 (.a(t0_000010001010), .b(t0_000010001011), .y(t0_00001000101));
wire t0_000010001010, t0_000010001011;
mixer mix_t0_0000100011 (.a(t0_00001000110), .b(t0_00001000111), .y(t0_0000100011));
wire t0_00001000110, t0_00001000111;
mixer mix_t0_00001000110 (.a(t0_000010001100), .b(t0_000010001101), .y(t0_00001000110));
wire t0_000010001100, t0_000010001101;
mixer mix_t0_00001000111 (.a(t0_000010001110), .b(t0_000010001111), .y(t0_00001000111));
wire t0_000010001110, t0_000010001111;
mixer mix_t0_00001001 (.a(t0_000010010), .b(t0_000010011), .y(t0_00001001));
wire t0_000010010, t0_000010011;
mixer mix_t0_000010010 (.a(t0_0000100100), .b(t0_0000100101), .y(t0_000010010));
wire t0_0000100100, t0_0000100101;
mixer mix_t0_0000100100 (.a(t0_00001001000), .b(t0_00001001001), .y(t0_0000100100));
wire t0_00001001000, t0_00001001001;
mixer mix_t0_00001001000 (.a(t0_000010010000), .b(t0_000010010001), .y(t0_00001001000));
wire t0_000010010000, t0_000010010001;
mixer mix_t0_00001001001 (.a(t0_000010010010), .b(t0_000010010011), .y(t0_00001001001));
wire t0_000010010010, t0_000010010011;
mixer mix_t0_0000100101 (.a(t0_00001001010), .b(t0_00001001011), .y(t0_0000100101));
wire t0_00001001010, t0_00001001011;
mixer mix_t0_00001001010 (.a(t0_000010010100), .b(t0_000010010101), .y(t0_00001001010));
wire t0_000010010100, t0_000010010101;
mixer mix_t0_00001001011 (.a(t0_000010010110), .b(t0_000010010111), .y(t0_00001001011));
wire t0_000010010110, t0_000010010111;
mixer mix_t0_000010011 (.a(t0_0000100110), .b(t0_0000100111), .y(t0_000010011));
wire t0_0000100110, t0_0000100111;
mixer mix_t0_0000100110 (.a(t0_00001001100), .b(t0_00001001101), .y(t0_0000100110));
wire t0_00001001100, t0_00001001101;
mixer mix_t0_00001001100 (.a(t0_000010011000), .b(t0_000010011001), .y(t0_00001001100));
wire t0_000010011000, t0_000010011001;
mixer mix_t0_00001001101 (.a(t0_000010011010), .b(t0_000010011011), .y(t0_00001001101));
wire t0_000010011010, t0_000010011011;
mixer mix_t0_0000100111 (.a(t0_00001001110), .b(t0_00001001111), .y(t0_0000100111));
wire t0_00001001110, t0_00001001111;
mixer mix_t0_00001001110 (.a(t0_000010011100), .b(t0_000010011101), .y(t0_00001001110));
wire t0_000010011100, t0_000010011101;
mixer mix_t0_00001001111 (.a(t0_000010011110), .b(t0_000010011111), .y(t0_00001001111));
wire t0_000010011110, t0_000010011111;
mixer mix_t0_0000101 (.a(t0_00001010), .b(t0_00001011), .y(t0_0000101));
wire t0_00001010, t0_00001011;
mixer mix_t0_00001010 (.a(t0_000010100), .b(t0_000010101), .y(t0_00001010));
wire t0_000010100, t0_000010101;
mixer mix_t0_000010100 (.a(t0_0000101000), .b(t0_0000101001), .y(t0_000010100));
wire t0_0000101000, t0_0000101001;
mixer mix_t0_0000101000 (.a(t0_00001010000), .b(t0_00001010001), .y(t0_0000101000));
wire t0_00001010000, t0_00001010001;
mixer mix_t0_00001010000 (.a(t0_000010100000), .b(t0_000010100001), .y(t0_00001010000));
wire t0_000010100000, t0_000010100001;
mixer mix_t0_00001010001 (.a(t0_000010100010), .b(t0_000010100011), .y(t0_00001010001));
wire t0_000010100010, t0_000010100011;
mixer mix_t0_0000101001 (.a(t0_00001010010), .b(t0_00001010011), .y(t0_0000101001));
wire t0_00001010010, t0_00001010011;
mixer mix_t0_00001010010 (.a(t0_000010100100), .b(t0_000010100101), .y(t0_00001010010));
wire t0_000010100100, t0_000010100101;
mixer mix_t0_00001010011 (.a(t0_000010100110), .b(t0_000010100111), .y(t0_00001010011));
wire t0_000010100110, t0_000010100111;
mixer mix_t0_000010101 (.a(t0_0000101010), .b(t0_0000101011), .y(t0_000010101));
wire t0_0000101010, t0_0000101011;
mixer mix_t0_0000101010 (.a(t0_00001010100), .b(t0_00001010101), .y(t0_0000101010));
wire t0_00001010100, t0_00001010101;
mixer mix_t0_00001010100 (.a(t0_000010101000), .b(t0_000010101001), .y(t0_00001010100));
wire t0_000010101000, t0_000010101001;
mixer mix_t0_00001010101 (.a(t0_000010101010), .b(t0_000010101011), .y(t0_00001010101));
wire t0_000010101010, t0_000010101011;
mixer mix_t0_0000101011 (.a(t0_00001010110), .b(t0_00001010111), .y(t0_0000101011));
wire t0_00001010110, t0_00001010111;
mixer mix_t0_00001010110 (.a(t0_000010101100), .b(t0_000010101101), .y(t0_00001010110));
wire t0_000010101100, t0_000010101101;
mixer mix_t0_00001010111 (.a(t0_000010101110), .b(t0_000010101111), .y(t0_00001010111));
wire t0_000010101110, t0_000010101111;
mixer mix_t0_00001011 (.a(t0_000010110), .b(t0_000010111), .y(t0_00001011));
wire t0_000010110, t0_000010111;
mixer mix_t0_000010110 (.a(t0_0000101100), .b(t0_0000101101), .y(t0_000010110));
wire t0_0000101100, t0_0000101101;
mixer mix_t0_0000101100 (.a(t0_00001011000), .b(t0_00001011001), .y(t0_0000101100));
wire t0_00001011000, t0_00001011001;
mixer mix_t0_00001011000 (.a(t0_000010110000), .b(t0_000010110001), .y(t0_00001011000));
wire t0_000010110000, t0_000010110001;
mixer mix_t0_00001011001 (.a(t0_000010110010), .b(t0_000010110011), .y(t0_00001011001));
wire t0_000010110010, t0_000010110011;
mixer mix_t0_0000101101 (.a(t0_00001011010), .b(t0_00001011011), .y(t0_0000101101));
wire t0_00001011010, t0_00001011011;
mixer mix_t0_00001011010 (.a(t0_000010110100), .b(t0_000010110101), .y(t0_00001011010));
wire t0_000010110100, t0_000010110101;
mixer mix_t0_00001011011 (.a(t0_000010110110), .b(t0_000010110111), .y(t0_00001011011));
wire t0_000010110110, t0_000010110111;
mixer mix_t0_000010111 (.a(t0_0000101110), .b(t0_0000101111), .y(t0_000010111));
wire t0_0000101110, t0_0000101111;
mixer mix_t0_0000101110 (.a(t0_00001011100), .b(t0_00001011101), .y(t0_0000101110));
wire t0_00001011100, t0_00001011101;
mixer mix_t0_00001011100 (.a(t0_000010111000), .b(t0_000010111001), .y(t0_00001011100));
wire t0_000010111000, t0_000010111001;
mixer mix_t0_00001011101 (.a(t0_000010111010), .b(t0_000010111011), .y(t0_00001011101));
wire t0_000010111010, t0_000010111011;
mixer mix_t0_0000101111 (.a(t0_00001011110), .b(t0_00001011111), .y(t0_0000101111));
wire t0_00001011110, t0_00001011111;
mixer mix_t0_00001011110 (.a(t0_000010111100), .b(t0_000010111101), .y(t0_00001011110));
wire t0_000010111100, t0_000010111101;
mixer mix_t0_00001011111 (.a(t0_000010111110), .b(t0_000010111111), .y(t0_00001011111));
wire t0_000010111110, t0_000010111111;
mixer mix_t0_000011 (.a(t0_0000110), .b(t0_0000111), .y(t0_000011));
wire t0_0000110, t0_0000111;
mixer mix_t0_0000110 (.a(t0_00001100), .b(t0_00001101), .y(t0_0000110));
wire t0_00001100, t0_00001101;
mixer mix_t0_00001100 (.a(t0_000011000), .b(t0_000011001), .y(t0_00001100));
wire t0_000011000, t0_000011001;
mixer mix_t0_000011000 (.a(t0_0000110000), .b(t0_0000110001), .y(t0_000011000));
wire t0_0000110000, t0_0000110001;
mixer mix_t0_0000110000 (.a(t0_00001100000), .b(t0_00001100001), .y(t0_0000110000));
wire t0_00001100000, t0_00001100001;
mixer mix_t0_00001100000 (.a(t0_000011000000), .b(t0_000011000001), .y(t0_00001100000));
wire t0_000011000000, t0_000011000001;
mixer mix_t0_00001100001 (.a(t0_000011000010), .b(t0_000011000011), .y(t0_00001100001));
wire t0_000011000010, t0_000011000011;
mixer mix_t0_0000110001 (.a(t0_00001100010), .b(t0_00001100011), .y(t0_0000110001));
wire t0_00001100010, t0_00001100011;
mixer mix_t0_00001100010 (.a(t0_000011000100), .b(t0_000011000101), .y(t0_00001100010));
wire t0_000011000100, t0_000011000101;
mixer mix_t0_00001100011 (.a(t0_000011000110), .b(t0_000011000111), .y(t0_00001100011));
wire t0_000011000110, t0_000011000111;
mixer mix_t0_000011001 (.a(t0_0000110010), .b(t0_0000110011), .y(t0_000011001));
wire t0_0000110010, t0_0000110011;
mixer mix_t0_0000110010 (.a(t0_00001100100), .b(t0_00001100101), .y(t0_0000110010));
wire t0_00001100100, t0_00001100101;
mixer mix_t0_00001100100 (.a(t0_000011001000), .b(t0_000011001001), .y(t0_00001100100));
wire t0_000011001000, t0_000011001001;
mixer mix_t0_00001100101 (.a(t0_000011001010), .b(t0_000011001011), .y(t0_00001100101));
wire t0_000011001010, t0_000011001011;
mixer mix_t0_0000110011 (.a(t0_00001100110), .b(t0_00001100111), .y(t0_0000110011));
wire t0_00001100110, t0_00001100111;
mixer mix_t0_00001100110 (.a(t0_000011001100), .b(t0_000011001101), .y(t0_00001100110));
wire t0_000011001100, t0_000011001101;
mixer mix_t0_00001100111 (.a(t0_000011001110), .b(t0_000011001111), .y(t0_00001100111));
wire t0_000011001110, t0_000011001111;
mixer mix_t0_00001101 (.a(t0_000011010), .b(t0_000011011), .y(t0_00001101));
wire t0_000011010, t0_000011011;
mixer mix_t0_000011010 (.a(t0_0000110100), .b(t0_0000110101), .y(t0_000011010));
wire t0_0000110100, t0_0000110101;
mixer mix_t0_0000110100 (.a(t0_00001101000), .b(t0_00001101001), .y(t0_0000110100));
wire t0_00001101000, t0_00001101001;
mixer mix_t0_00001101000 (.a(t0_000011010000), .b(t0_000011010001), .y(t0_00001101000));
wire t0_000011010000, t0_000011010001;
mixer mix_t0_00001101001 (.a(t0_000011010010), .b(t0_000011010011), .y(t0_00001101001));
wire t0_000011010010, t0_000011010011;
mixer mix_t0_0000110101 (.a(t0_00001101010), .b(t0_00001101011), .y(t0_0000110101));
wire t0_00001101010, t0_00001101011;
mixer mix_t0_00001101010 (.a(t0_000011010100), .b(t0_000011010101), .y(t0_00001101010));
wire t0_000011010100, t0_000011010101;
mixer mix_t0_00001101011 (.a(t0_000011010110), .b(t0_000011010111), .y(t0_00001101011));
wire t0_000011010110, t0_000011010111;
mixer mix_t0_000011011 (.a(t0_0000110110), .b(t0_0000110111), .y(t0_000011011));
wire t0_0000110110, t0_0000110111;
mixer mix_t0_0000110110 (.a(t0_00001101100), .b(t0_00001101101), .y(t0_0000110110));
wire t0_00001101100, t0_00001101101;
mixer mix_t0_00001101100 (.a(t0_000011011000), .b(t0_000011011001), .y(t0_00001101100));
wire t0_000011011000, t0_000011011001;
mixer mix_t0_00001101101 (.a(t0_000011011010), .b(t0_000011011011), .y(t0_00001101101));
wire t0_000011011010, t0_000011011011;
mixer mix_t0_0000110111 (.a(t0_00001101110), .b(t0_00001101111), .y(t0_0000110111));
wire t0_00001101110, t0_00001101111;
mixer mix_t0_00001101110 (.a(t0_000011011100), .b(t0_000011011101), .y(t0_00001101110));
wire t0_000011011100, t0_000011011101;
mixer mix_t0_00001101111 (.a(t0_000011011110), .b(t0_000011011111), .y(t0_00001101111));
wire t0_000011011110, t0_000011011111;
mixer mix_t0_0000111 (.a(t0_00001110), .b(t0_00001111), .y(t0_0000111));
wire t0_00001110, t0_00001111;
mixer mix_t0_00001110 (.a(t0_000011100), .b(t0_000011101), .y(t0_00001110));
wire t0_000011100, t0_000011101;
mixer mix_t0_000011100 (.a(t0_0000111000), .b(t0_0000111001), .y(t0_000011100));
wire t0_0000111000, t0_0000111001;
mixer mix_t0_0000111000 (.a(t0_00001110000), .b(t0_00001110001), .y(t0_0000111000));
wire t0_00001110000, t0_00001110001;
mixer mix_t0_00001110000 (.a(t0_000011100000), .b(t0_000011100001), .y(t0_00001110000));
wire t0_000011100000, t0_000011100001;
mixer mix_t0_00001110001 (.a(t0_000011100010), .b(t0_000011100011), .y(t0_00001110001));
wire t0_000011100010, t0_000011100011;
mixer mix_t0_0000111001 (.a(t0_00001110010), .b(t0_00001110011), .y(t0_0000111001));
wire t0_00001110010, t0_00001110011;
mixer mix_t0_00001110010 (.a(t0_000011100100), .b(t0_000011100101), .y(t0_00001110010));
wire t0_000011100100, t0_000011100101;
mixer mix_t0_00001110011 (.a(t0_000011100110), .b(t0_000011100111), .y(t0_00001110011));
wire t0_000011100110, t0_000011100111;
mixer mix_t0_000011101 (.a(t0_0000111010), .b(t0_0000111011), .y(t0_000011101));
wire t0_0000111010, t0_0000111011;
mixer mix_t0_0000111010 (.a(t0_00001110100), .b(t0_00001110101), .y(t0_0000111010));
wire t0_00001110100, t0_00001110101;
mixer mix_t0_00001110100 (.a(t0_000011101000), .b(t0_000011101001), .y(t0_00001110100));
wire t0_000011101000, t0_000011101001;
mixer mix_t0_00001110101 (.a(t0_000011101010), .b(t0_000011101011), .y(t0_00001110101));
wire t0_000011101010, t0_000011101011;
mixer mix_t0_0000111011 (.a(t0_00001110110), .b(t0_00001110111), .y(t0_0000111011));
wire t0_00001110110, t0_00001110111;
mixer mix_t0_00001110110 (.a(t0_000011101100), .b(t0_000011101101), .y(t0_00001110110));
wire t0_000011101100, t0_000011101101;
mixer mix_t0_00001110111 (.a(t0_000011101110), .b(t0_000011101111), .y(t0_00001110111));
wire t0_000011101110, t0_000011101111;
mixer mix_t0_00001111 (.a(t0_000011110), .b(t0_000011111), .y(t0_00001111));
wire t0_000011110, t0_000011111;
mixer mix_t0_000011110 (.a(t0_0000111100), .b(t0_0000111101), .y(t0_000011110));
wire t0_0000111100, t0_0000111101;
mixer mix_t0_0000111100 (.a(t0_00001111000), .b(t0_00001111001), .y(t0_0000111100));
wire t0_00001111000, t0_00001111001;
mixer mix_t0_00001111000 (.a(t0_000011110000), .b(t0_000011110001), .y(t0_00001111000));
wire t0_000011110000, t0_000011110001;
mixer mix_t0_00001111001 (.a(t0_000011110010), .b(t0_000011110011), .y(t0_00001111001));
wire t0_000011110010, t0_000011110011;
mixer mix_t0_0000111101 (.a(t0_00001111010), .b(t0_00001111011), .y(t0_0000111101));
wire t0_00001111010, t0_00001111011;
mixer mix_t0_00001111010 (.a(t0_000011110100), .b(t0_000011110101), .y(t0_00001111010));
wire t0_000011110100, t0_000011110101;
mixer mix_t0_00001111011 (.a(t0_000011110110), .b(t0_000011110111), .y(t0_00001111011));
wire t0_000011110110, t0_000011110111;
mixer mix_t0_000011111 (.a(t0_0000111110), .b(t0_0000111111), .y(t0_000011111));
wire t0_0000111110, t0_0000111111;
mixer mix_t0_0000111110 (.a(t0_00001111100), .b(t0_00001111101), .y(t0_0000111110));
wire t0_00001111100, t0_00001111101;
mixer mix_t0_00001111100 (.a(t0_000011111000), .b(t0_000011111001), .y(t0_00001111100));
wire t0_000011111000, t0_000011111001;
mixer mix_t0_00001111101 (.a(t0_000011111010), .b(t0_000011111011), .y(t0_00001111101));
wire t0_000011111010, t0_000011111011;
mixer mix_t0_0000111111 (.a(t0_00001111110), .b(t0_00001111111), .y(t0_0000111111));
wire t0_00001111110, t0_00001111111;
mixer mix_t0_00001111110 (.a(t0_000011111100), .b(t0_000011111101), .y(t0_00001111110));
wire t0_000011111100, t0_000011111101;
mixer mix_t0_00001111111 (.a(t0_000011111110), .b(t0_000011111111), .y(t0_00001111111));
wire t0_000011111110, t0_000011111111;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_000100 (.a(t0_0001000), .b(t0_0001001), .y(t0_000100));
wire t0_0001000, t0_0001001;
mixer mix_t0_0001000 (.a(t0_00010000), .b(t0_00010001), .y(t0_0001000));
wire t0_00010000, t0_00010001;
mixer mix_t0_00010000 (.a(t0_000100000), .b(t0_000100001), .y(t0_00010000));
wire t0_000100000, t0_000100001;
mixer mix_t0_000100000 (.a(t0_0001000000), .b(t0_0001000001), .y(t0_000100000));
wire t0_0001000000, t0_0001000001;
mixer mix_t0_0001000000 (.a(t0_00010000000), .b(t0_00010000001), .y(t0_0001000000));
wire t0_00010000000, t0_00010000001;
mixer mix_t0_00010000000 (.a(t0_000100000000), .b(t0_000100000001), .y(t0_00010000000));
wire t0_000100000000, t0_000100000001;
mixer mix_t0_00010000001 (.a(t0_000100000010), .b(t0_000100000011), .y(t0_00010000001));
wire t0_000100000010, t0_000100000011;
mixer mix_t0_0001000001 (.a(t0_00010000010), .b(t0_00010000011), .y(t0_0001000001));
wire t0_00010000010, t0_00010000011;
mixer mix_t0_00010000010 (.a(t0_000100000100), .b(t0_000100000101), .y(t0_00010000010));
wire t0_000100000100, t0_000100000101;
mixer mix_t0_00010000011 (.a(t0_000100000110), .b(t0_000100000111), .y(t0_00010000011));
wire t0_000100000110, t0_000100000111;
mixer mix_t0_000100001 (.a(t0_0001000010), .b(t0_0001000011), .y(t0_000100001));
wire t0_0001000010, t0_0001000011;
mixer mix_t0_0001000010 (.a(t0_00010000100), .b(t0_00010000101), .y(t0_0001000010));
wire t0_00010000100, t0_00010000101;
mixer mix_t0_00010000100 (.a(t0_000100001000), .b(t0_000100001001), .y(t0_00010000100));
wire t0_000100001000, t0_000100001001;
mixer mix_t0_00010000101 (.a(t0_000100001010), .b(t0_000100001011), .y(t0_00010000101));
wire t0_000100001010, t0_000100001011;
mixer mix_t0_0001000011 (.a(t0_00010000110), .b(t0_00010000111), .y(t0_0001000011));
wire t0_00010000110, t0_00010000111;
mixer mix_t0_00010000110 (.a(t0_000100001100), .b(t0_000100001101), .y(t0_00010000110));
wire t0_000100001100, t0_000100001101;
mixer mix_t0_00010000111 (.a(t0_000100001110), .b(t0_000100001111), .y(t0_00010000111));
wire t0_000100001110, t0_000100001111;
mixer mix_t0_00010001 (.a(t0_000100010), .b(t0_000100011), .y(t0_00010001));
wire t0_000100010, t0_000100011;
mixer mix_t0_000100010 (.a(t0_0001000100), .b(t0_0001000101), .y(t0_000100010));
wire t0_0001000100, t0_0001000101;
mixer mix_t0_0001000100 (.a(t0_00010001000), .b(t0_00010001001), .y(t0_0001000100));
wire t0_00010001000, t0_00010001001;
mixer mix_t0_00010001000 (.a(t0_000100010000), .b(t0_000100010001), .y(t0_00010001000));
wire t0_000100010000, t0_000100010001;
mixer mix_t0_00010001001 (.a(t0_000100010010), .b(t0_000100010011), .y(t0_00010001001));
wire t0_000100010010, t0_000100010011;
mixer mix_t0_0001000101 (.a(t0_00010001010), .b(t0_00010001011), .y(t0_0001000101));
wire t0_00010001010, t0_00010001011;
mixer mix_t0_00010001010 (.a(t0_000100010100), .b(t0_000100010101), .y(t0_00010001010));
wire t0_000100010100, t0_000100010101;
mixer mix_t0_00010001011 (.a(t0_000100010110), .b(t0_000100010111), .y(t0_00010001011));
wire t0_000100010110, t0_000100010111;
mixer mix_t0_000100011 (.a(t0_0001000110), .b(t0_0001000111), .y(t0_000100011));
wire t0_0001000110, t0_0001000111;
mixer mix_t0_0001000110 (.a(t0_00010001100), .b(t0_00010001101), .y(t0_0001000110));
wire t0_00010001100, t0_00010001101;
mixer mix_t0_00010001100 (.a(t0_000100011000), .b(t0_000100011001), .y(t0_00010001100));
wire t0_000100011000, t0_000100011001;
mixer mix_t0_00010001101 (.a(t0_000100011010), .b(t0_000100011011), .y(t0_00010001101));
wire t0_000100011010, t0_000100011011;
mixer mix_t0_0001000111 (.a(t0_00010001110), .b(t0_00010001111), .y(t0_0001000111));
wire t0_00010001110, t0_00010001111;
mixer mix_t0_00010001110 (.a(t0_000100011100), .b(t0_000100011101), .y(t0_00010001110));
wire t0_000100011100, t0_000100011101;
mixer mix_t0_00010001111 (.a(t0_000100011110), .b(t0_000100011111), .y(t0_00010001111));
wire t0_000100011110, t0_000100011111;
mixer mix_t0_0001001 (.a(t0_00010010), .b(t0_00010011), .y(t0_0001001));
wire t0_00010010, t0_00010011;
mixer mix_t0_00010010 (.a(t0_000100100), .b(t0_000100101), .y(t0_00010010));
wire t0_000100100, t0_000100101;
mixer mix_t0_000100100 (.a(t0_0001001000), .b(t0_0001001001), .y(t0_000100100));
wire t0_0001001000, t0_0001001001;
mixer mix_t0_0001001000 (.a(t0_00010010000), .b(t0_00010010001), .y(t0_0001001000));
wire t0_00010010000, t0_00010010001;
mixer mix_t0_00010010000 (.a(t0_000100100000), .b(t0_000100100001), .y(t0_00010010000));
wire t0_000100100000, t0_000100100001;
mixer mix_t0_00010010001 (.a(t0_000100100010), .b(t0_000100100011), .y(t0_00010010001));
wire t0_000100100010, t0_000100100011;
mixer mix_t0_0001001001 (.a(t0_00010010010), .b(t0_00010010011), .y(t0_0001001001));
wire t0_00010010010, t0_00010010011;
mixer mix_t0_00010010010 (.a(t0_000100100100), .b(t0_000100100101), .y(t0_00010010010));
wire t0_000100100100, t0_000100100101;
mixer mix_t0_00010010011 (.a(t0_000100100110), .b(t0_000100100111), .y(t0_00010010011));
wire t0_000100100110, t0_000100100111;
mixer mix_t0_000100101 (.a(t0_0001001010), .b(t0_0001001011), .y(t0_000100101));
wire t0_0001001010, t0_0001001011;
mixer mix_t0_0001001010 (.a(t0_00010010100), .b(t0_00010010101), .y(t0_0001001010));
wire t0_00010010100, t0_00010010101;
mixer mix_t0_00010010100 (.a(t0_000100101000), .b(t0_000100101001), .y(t0_00010010100));
wire t0_000100101000, t0_000100101001;
mixer mix_t0_00010010101 (.a(t0_000100101010), .b(t0_000100101011), .y(t0_00010010101));
wire t0_000100101010, t0_000100101011;
mixer mix_t0_0001001011 (.a(t0_00010010110), .b(t0_00010010111), .y(t0_0001001011));
wire t0_00010010110, t0_00010010111;
mixer mix_t0_00010010110 (.a(t0_000100101100), .b(t0_000100101101), .y(t0_00010010110));
wire t0_000100101100, t0_000100101101;
mixer mix_t0_00010010111 (.a(t0_000100101110), .b(t0_000100101111), .y(t0_00010010111));
wire t0_000100101110, t0_000100101111;
mixer mix_t0_00010011 (.a(t0_000100110), .b(t0_000100111), .y(t0_00010011));
wire t0_000100110, t0_000100111;
mixer mix_t0_000100110 (.a(t0_0001001100), .b(t0_0001001101), .y(t0_000100110));
wire t0_0001001100, t0_0001001101;
mixer mix_t0_0001001100 (.a(t0_00010011000), .b(t0_00010011001), .y(t0_0001001100));
wire t0_00010011000, t0_00010011001;
mixer mix_t0_00010011000 (.a(t0_000100110000), .b(t0_000100110001), .y(t0_00010011000));
wire t0_000100110000, t0_000100110001;
mixer mix_t0_00010011001 (.a(t0_000100110010), .b(t0_000100110011), .y(t0_00010011001));
wire t0_000100110010, t0_000100110011;
mixer mix_t0_0001001101 (.a(t0_00010011010), .b(t0_00010011011), .y(t0_0001001101));
wire t0_00010011010, t0_00010011011;
mixer mix_t0_00010011010 (.a(t0_000100110100), .b(t0_000100110101), .y(t0_00010011010));
wire t0_000100110100, t0_000100110101;
mixer mix_t0_00010011011 (.a(t0_000100110110), .b(t0_000100110111), .y(t0_00010011011));
wire t0_000100110110, t0_000100110111;
mixer mix_t0_000100111 (.a(t0_0001001110), .b(t0_0001001111), .y(t0_000100111));
wire t0_0001001110, t0_0001001111;
mixer mix_t0_0001001110 (.a(t0_00010011100), .b(t0_00010011101), .y(t0_0001001110));
wire t0_00010011100, t0_00010011101;
mixer mix_t0_00010011100 (.a(t0_000100111000), .b(t0_000100111001), .y(t0_00010011100));
wire t0_000100111000, t0_000100111001;
mixer mix_t0_00010011101 (.a(t0_000100111010), .b(t0_000100111011), .y(t0_00010011101));
wire t0_000100111010, t0_000100111011;
mixer mix_t0_0001001111 (.a(t0_00010011110), .b(t0_00010011111), .y(t0_0001001111));
wire t0_00010011110, t0_00010011111;
mixer mix_t0_00010011110 (.a(t0_000100111100), .b(t0_000100111101), .y(t0_00010011110));
wire t0_000100111100, t0_000100111101;
mixer mix_t0_00010011111 (.a(t0_000100111110), .b(t0_000100111111), .y(t0_00010011111));
wire t0_000100111110, t0_000100111111;
mixer mix_t0_000101 (.a(t0_0001010), .b(t0_0001011), .y(t0_000101));
wire t0_0001010, t0_0001011;
mixer mix_t0_0001010 (.a(t0_00010100), .b(t0_00010101), .y(t0_0001010));
wire t0_00010100, t0_00010101;
mixer mix_t0_00010100 (.a(t0_000101000), .b(t0_000101001), .y(t0_00010100));
wire t0_000101000, t0_000101001;
mixer mix_t0_000101000 (.a(t0_0001010000), .b(t0_0001010001), .y(t0_000101000));
wire t0_0001010000, t0_0001010001;
mixer mix_t0_0001010000 (.a(t0_00010100000), .b(t0_00010100001), .y(t0_0001010000));
wire t0_00010100000, t0_00010100001;
mixer mix_t0_00010100000 (.a(t0_000101000000), .b(t0_000101000001), .y(t0_00010100000));
wire t0_000101000000, t0_000101000001;
mixer mix_t0_00010100001 (.a(t0_000101000010), .b(t0_000101000011), .y(t0_00010100001));
wire t0_000101000010, t0_000101000011;
mixer mix_t0_0001010001 (.a(t0_00010100010), .b(t0_00010100011), .y(t0_0001010001));
wire t0_00010100010, t0_00010100011;
mixer mix_t0_00010100010 (.a(t0_000101000100), .b(t0_000101000101), .y(t0_00010100010));
wire t0_000101000100, t0_000101000101;
mixer mix_t0_00010100011 (.a(t0_000101000110), .b(t0_000101000111), .y(t0_00010100011));
wire t0_000101000110, t0_000101000111;
mixer mix_t0_000101001 (.a(t0_0001010010), .b(t0_0001010011), .y(t0_000101001));
wire t0_0001010010, t0_0001010011;
mixer mix_t0_0001010010 (.a(t0_00010100100), .b(t0_00010100101), .y(t0_0001010010));
wire t0_00010100100, t0_00010100101;
mixer mix_t0_00010100100 (.a(t0_000101001000), .b(t0_000101001001), .y(t0_00010100100));
wire t0_000101001000, t0_000101001001;
mixer mix_t0_00010100101 (.a(t0_000101001010), .b(t0_000101001011), .y(t0_00010100101));
wire t0_000101001010, t0_000101001011;
mixer mix_t0_0001010011 (.a(t0_00010100110), .b(t0_00010100111), .y(t0_0001010011));
wire t0_00010100110, t0_00010100111;
mixer mix_t0_00010100110 (.a(t0_000101001100), .b(t0_000101001101), .y(t0_00010100110));
wire t0_000101001100, t0_000101001101;
mixer mix_t0_00010100111 (.a(t0_000101001110), .b(t0_000101001111), .y(t0_00010100111));
wire t0_000101001110, t0_000101001111;
mixer mix_t0_00010101 (.a(t0_000101010), .b(t0_000101011), .y(t0_00010101));
wire t0_000101010, t0_000101011;
mixer mix_t0_000101010 (.a(t0_0001010100), .b(t0_0001010101), .y(t0_000101010));
wire t0_0001010100, t0_0001010101;
mixer mix_t0_0001010100 (.a(t0_00010101000), .b(t0_00010101001), .y(t0_0001010100));
wire t0_00010101000, t0_00010101001;
mixer mix_t0_00010101000 (.a(t0_000101010000), .b(t0_000101010001), .y(t0_00010101000));
wire t0_000101010000, t0_000101010001;
mixer mix_t0_00010101001 (.a(t0_000101010010), .b(t0_000101010011), .y(t0_00010101001));
wire t0_000101010010, t0_000101010011;
mixer mix_t0_0001010101 (.a(t0_00010101010), .b(t0_00010101011), .y(t0_0001010101));
wire t0_00010101010, t0_00010101011;
mixer mix_t0_00010101010 (.a(t0_000101010100), .b(t0_000101010101), .y(t0_00010101010));
wire t0_000101010100, t0_000101010101;
mixer mix_t0_00010101011 (.a(t0_000101010110), .b(t0_000101010111), .y(t0_00010101011));
wire t0_000101010110, t0_000101010111;
mixer mix_t0_000101011 (.a(t0_0001010110), .b(t0_0001010111), .y(t0_000101011));
wire t0_0001010110, t0_0001010111;
mixer mix_t0_0001010110 (.a(t0_00010101100), .b(t0_00010101101), .y(t0_0001010110));
wire t0_00010101100, t0_00010101101;
mixer mix_t0_00010101100 (.a(t0_000101011000), .b(t0_000101011001), .y(t0_00010101100));
wire t0_000101011000, t0_000101011001;
mixer mix_t0_00010101101 (.a(t0_000101011010), .b(t0_000101011011), .y(t0_00010101101));
wire t0_000101011010, t0_000101011011;
mixer mix_t0_0001010111 (.a(t0_00010101110), .b(t0_00010101111), .y(t0_0001010111));
wire t0_00010101110, t0_00010101111;
mixer mix_t0_00010101110 (.a(t0_000101011100), .b(t0_000101011101), .y(t0_00010101110));
wire t0_000101011100, t0_000101011101;
mixer mix_t0_00010101111 (.a(t0_000101011110), .b(t0_000101011111), .y(t0_00010101111));
wire t0_000101011110, t0_000101011111;
mixer mix_t0_0001011 (.a(t0_00010110), .b(t0_00010111), .y(t0_0001011));
wire t0_00010110, t0_00010111;
mixer mix_t0_00010110 (.a(t0_000101100), .b(t0_000101101), .y(t0_00010110));
wire t0_000101100, t0_000101101;
mixer mix_t0_000101100 (.a(t0_0001011000), .b(t0_0001011001), .y(t0_000101100));
wire t0_0001011000, t0_0001011001;
mixer mix_t0_0001011000 (.a(t0_00010110000), .b(t0_00010110001), .y(t0_0001011000));
wire t0_00010110000, t0_00010110001;
mixer mix_t0_00010110000 (.a(t0_000101100000), .b(t0_000101100001), .y(t0_00010110000));
wire t0_000101100000, t0_000101100001;
mixer mix_t0_00010110001 (.a(t0_000101100010), .b(t0_000101100011), .y(t0_00010110001));
wire t0_000101100010, t0_000101100011;
mixer mix_t0_0001011001 (.a(t0_00010110010), .b(t0_00010110011), .y(t0_0001011001));
wire t0_00010110010, t0_00010110011;
mixer mix_t0_00010110010 (.a(t0_000101100100), .b(t0_000101100101), .y(t0_00010110010));
wire t0_000101100100, t0_000101100101;
mixer mix_t0_00010110011 (.a(t0_000101100110), .b(t0_000101100111), .y(t0_00010110011));
wire t0_000101100110, t0_000101100111;
mixer mix_t0_000101101 (.a(t0_0001011010), .b(t0_0001011011), .y(t0_000101101));
wire t0_0001011010, t0_0001011011;
mixer mix_t0_0001011010 (.a(t0_00010110100), .b(t0_00010110101), .y(t0_0001011010));
wire t0_00010110100, t0_00010110101;
mixer mix_t0_00010110100 (.a(t0_000101101000), .b(t0_000101101001), .y(t0_00010110100));
wire t0_000101101000, t0_000101101001;
mixer mix_t0_00010110101 (.a(t0_000101101010), .b(t0_000101101011), .y(t0_00010110101));
wire t0_000101101010, t0_000101101011;
mixer mix_t0_0001011011 (.a(t0_00010110110), .b(t0_00010110111), .y(t0_0001011011));
wire t0_00010110110, t0_00010110111;
mixer mix_t0_00010110110 (.a(t0_000101101100), .b(t0_000101101101), .y(t0_00010110110));
wire t0_000101101100, t0_000101101101;
mixer mix_t0_00010110111 (.a(t0_000101101110), .b(t0_000101101111), .y(t0_00010110111));
wire t0_000101101110, t0_000101101111;
mixer mix_t0_00010111 (.a(t0_000101110), .b(t0_000101111), .y(t0_00010111));
wire t0_000101110, t0_000101111;
mixer mix_t0_000101110 (.a(t0_0001011100), .b(t0_0001011101), .y(t0_000101110));
wire t0_0001011100, t0_0001011101;
mixer mix_t0_0001011100 (.a(t0_00010111000), .b(t0_00010111001), .y(t0_0001011100));
wire t0_00010111000, t0_00010111001;
mixer mix_t0_00010111000 (.a(t0_000101110000), .b(t0_000101110001), .y(t0_00010111000));
wire t0_000101110000, t0_000101110001;
mixer mix_t0_00010111001 (.a(t0_000101110010), .b(t0_000101110011), .y(t0_00010111001));
wire t0_000101110010, t0_000101110011;
mixer mix_t0_0001011101 (.a(t0_00010111010), .b(t0_00010111011), .y(t0_0001011101));
wire t0_00010111010, t0_00010111011;
mixer mix_t0_00010111010 (.a(t0_000101110100), .b(t0_000101110101), .y(t0_00010111010));
wire t0_000101110100, t0_000101110101;
mixer mix_t0_00010111011 (.a(t0_000101110110), .b(t0_000101110111), .y(t0_00010111011));
wire t0_000101110110, t0_000101110111;
mixer mix_t0_000101111 (.a(t0_0001011110), .b(t0_0001011111), .y(t0_000101111));
wire t0_0001011110, t0_0001011111;
mixer mix_t0_0001011110 (.a(t0_00010111100), .b(t0_00010111101), .y(t0_0001011110));
wire t0_00010111100, t0_00010111101;
mixer mix_t0_00010111100 (.a(t0_000101111000), .b(t0_000101111001), .y(t0_00010111100));
wire t0_000101111000, t0_000101111001;
mixer mix_t0_00010111101 (.a(t0_000101111010), .b(t0_000101111011), .y(t0_00010111101));
wire t0_000101111010, t0_000101111011;
mixer mix_t0_0001011111 (.a(t0_00010111110), .b(t0_00010111111), .y(t0_0001011111));
wire t0_00010111110, t0_00010111111;
mixer mix_t0_00010111110 (.a(t0_000101111100), .b(t0_000101111101), .y(t0_00010111110));
wire t0_000101111100, t0_000101111101;
mixer mix_t0_00010111111 (.a(t0_000101111110), .b(t0_000101111111), .y(t0_00010111111));
wire t0_000101111110, t0_000101111111;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_000110 (.a(t0_0001100), .b(t0_0001101), .y(t0_000110));
wire t0_0001100, t0_0001101;
mixer mix_t0_0001100 (.a(t0_00011000), .b(t0_00011001), .y(t0_0001100));
wire t0_00011000, t0_00011001;
mixer mix_t0_00011000 (.a(t0_000110000), .b(t0_000110001), .y(t0_00011000));
wire t0_000110000, t0_000110001;
mixer mix_t0_000110000 (.a(t0_0001100000), .b(t0_0001100001), .y(t0_000110000));
wire t0_0001100000, t0_0001100001;
mixer mix_t0_0001100000 (.a(t0_00011000000), .b(t0_00011000001), .y(t0_0001100000));
wire t0_00011000000, t0_00011000001;
mixer mix_t0_00011000000 (.a(t0_000110000000), .b(t0_000110000001), .y(t0_00011000000));
wire t0_000110000000, t0_000110000001;
mixer mix_t0_00011000001 (.a(t0_000110000010), .b(t0_000110000011), .y(t0_00011000001));
wire t0_000110000010, t0_000110000011;
mixer mix_t0_0001100001 (.a(t0_00011000010), .b(t0_00011000011), .y(t0_0001100001));
wire t0_00011000010, t0_00011000011;
mixer mix_t0_00011000010 (.a(t0_000110000100), .b(t0_000110000101), .y(t0_00011000010));
wire t0_000110000100, t0_000110000101;
mixer mix_t0_00011000011 (.a(t0_000110000110), .b(t0_000110000111), .y(t0_00011000011));
wire t0_000110000110, t0_000110000111;
mixer mix_t0_000110001 (.a(t0_0001100010), .b(t0_0001100011), .y(t0_000110001));
wire t0_0001100010, t0_0001100011;
mixer mix_t0_0001100010 (.a(t0_00011000100), .b(t0_00011000101), .y(t0_0001100010));
wire t0_00011000100, t0_00011000101;
mixer mix_t0_00011000100 (.a(t0_000110001000), .b(t0_000110001001), .y(t0_00011000100));
wire t0_000110001000, t0_000110001001;
mixer mix_t0_00011000101 (.a(t0_000110001010), .b(t0_000110001011), .y(t0_00011000101));
wire t0_000110001010, t0_000110001011;
mixer mix_t0_0001100011 (.a(t0_00011000110), .b(t0_00011000111), .y(t0_0001100011));
wire t0_00011000110, t0_00011000111;
mixer mix_t0_00011000110 (.a(t0_000110001100), .b(t0_000110001101), .y(t0_00011000110));
wire t0_000110001100, t0_000110001101;
mixer mix_t0_00011000111 (.a(t0_000110001110), .b(t0_000110001111), .y(t0_00011000111));
wire t0_000110001110, t0_000110001111;
mixer mix_t0_00011001 (.a(t0_000110010), .b(t0_000110011), .y(t0_00011001));
wire t0_000110010, t0_000110011;
mixer mix_t0_000110010 (.a(t0_0001100100), .b(t0_0001100101), .y(t0_000110010));
wire t0_0001100100, t0_0001100101;
mixer mix_t0_0001100100 (.a(t0_00011001000), .b(t0_00011001001), .y(t0_0001100100));
wire t0_00011001000, t0_00011001001;
mixer mix_t0_00011001000 (.a(t0_000110010000), .b(t0_000110010001), .y(t0_00011001000));
wire t0_000110010000, t0_000110010001;
mixer mix_t0_00011001001 (.a(t0_000110010010), .b(t0_000110010011), .y(t0_00011001001));
wire t0_000110010010, t0_000110010011;
mixer mix_t0_0001100101 (.a(t0_00011001010), .b(t0_00011001011), .y(t0_0001100101));
wire t0_00011001010, t0_00011001011;
mixer mix_t0_00011001010 (.a(t0_000110010100), .b(t0_000110010101), .y(t0_00011001010));
wire t0_000110010100, t0_000110010101;
mixer mix_t0_00011001011 (.a(t0_000110010110), .b(t0_000110010111), .y(t0_00011001011));
wire t0_000110010110, t0_000110010111;
mixer mix_t0_000110011 (.a(t0_0001100110), .b(t0_0001100111), .y(t0_000110011));
wire t0_0001100110, t0_0001100111;
mixer mix_t0_0001100110 (.a(t0_00011001100), .b(t0_00011001101), .y(t0_0001100110));
wire t0_00011001100, t0_00011001101;
mixer mix_t0_00011001100 (.a(t0_000110011000), .b(t0_000110011001), .y(t0_00011001100));
wire t0_000110011000, t0_000110011001;
mixer mix_t0_00011001101 (.a(t0_000110011010), .b(t0_000110011011), .y(t0_00011001101));
wire t0_000110011010, t0_000110011011;
mixer mix_t0_0001100111 (.a(t0_00011001110), .b(t0_00011001111), .y(t0_0001100111));
wire t0_00011001110, t0_00011001111;
mixer mix_t0_00011001110 (.a(t0_000110011100), .b(t0_000110011101), .y(t0_00011001110));
wire t0_000110011100, t0_000110011101;
mixer mix_t0_00011001111 (.a(t0_000110011110), .b(t0_000110011111), .y(t0_00011001111));
wire t0_000110011110, t0_000110011111;
mixer mix_t0_0001101 (.a(t0_00011010), .b(t0_00011011), .y(t0_0001101));
wire t0_00011010, t0_00011011;
mixer mix_t0_00011010 (.a(t0_000110100), .b(t0_000110101), .y(t0_00011010));
wire t0_000110100, t0_000110101;
mixer mix_t0_000110100 (.a(t0_0001101000), .b(t0_0001101001), .y(t0_000110100));
wire t0_0001101000, t0_0001101001;
mixer mix_t0_0001101000 (.a(t0_00011010000), .b(t0_00011010001), .y(t0_0001101000));
wire t0_00011010000, t0_00011010001;
mixer mix_t0_00011010000 (.a(t0_000110100000), .b(t0_000110100001), .y(t0_00011010000));
wire t0_000110100000, t0_000110100001;
mixer mix_t0_00011010001 (.a(t0_000110100010), .b(t0_000110100011), .y(t0_00011010001));
wire t0_000110100010, t0_000110100011;
mixer mix_t0_0001101001 (.a(t0_00011010010), .b(t0_00011010011), .y(t0_0001101001));
wire t0_00011010010, t0_00011010011;
mixer mix_t0_00011010010 (.a(t0_000110100100), .b(t0_000110100101), .y(t0_00011010010));
wire t0_000110100100, t0_000110100101;
mixer mix_t0_00011010011 (.a(t0_000110100110), .b(t0_000110100111), .y(t0_00011010011));
wire t0_000110100110, t0_000110100111;
mixer mix_t0_000110101 (.a(t0_0001101010), .b(t0_0001101011), .y(t0_000110101));
wire t0_0001101010, t0_0001101011;
mixer mix_t0_0001101010 (.a(t0_00011010100), .b(t0_00011010101), .y(t0_0001101010));
wire t0_00011010100, t0_00011010101;
mixer mix_t0_00011010100 (.a(t0_000110101000), .b(t0_000110101001), .y(t0_00011010100));
wire t0_000110101000, t0_000110101001;
mixer mix_t0_00011010101 (.a(t0_000110101010), .b(t0_000110101011), .y(t0_00011010101));
wire t0_000110101010, t0_000110101011;
mixer mix_t0_0001101011 (.a(t0_00011010110), .b(t0_00011010111), .y(t0_0001101011));
wire t0_00011010110, t0_00011010111;
mixer mix_t0_00011010110 (.a(t0_000110101100), .b(t0_000110101101), .y(t0_00011010110));
wire t0_000110101100, t0_000110101101;
mixer mix_t0_00011010111 (.a(t0_000110101110), .b(t0_000110101111), .y(t0_00011010111));
wire t0_000110101110, t0_000110101111;
mixer mix_t0_00011011 (.a(t0_000110110), .b(t0_000110111), .y(t0_00011011));
wire t0_000110110, t0_000110111;
mixer mix_t0_000110110 (.a(t0_0001101100), .b(t0_0001101101), .y(t0_000110110));
wire t0_0001101100, t0_0001101101;
mixer mix_t0_0001101100 (.a(t0_00011011000), .b(t0_00011011001), .y(t0_0001101100));
wire t0_00011011000, t0_00011011001;
mixer mix_t0_00011011000 (.a(t0_000110110000), .b(t0_000110110001), .y(t0_00011011000));
wire t0_000110110000, t0_000110110001;
mixer mix_t0_00011011001 (.a(t0_000110110010), .b(t0_000110110011), .y(t0_00011011001));
wire t0_000110110010, t0_000110110011;
mixer mix_t0_0001101101 (.a(t0_00011011010), .b(t0_00011011011), .y(t0_0001101101));
wire t0_00011011010, t0_00011011011;
mixer mix_t0_00011011010 (.a(t0_000110110100), .b(t0_000110110101), .y(t0_00011011010));
wire t0_000110110100, t0_000110110101;
mixer mix_t0_00011011011 (.a(t0_000110110110), .b(t0_000110110111), .y(t0_00011011011));
wire t0_000110110110, t0_000110110111;
mixer mix_t0_000110111 (.a(t0_0001101110), .b(t0_0001101111), .y(t0_000110111));
wire t0_0001101110, t0_0001101111;
mixer mix_t0_0001101110 (.a(t0_00011011100), .b(t0_00011011101), .y(t0_0001101110));
wire t0_00011011100, t0_00011011101;
mixer mix_t0_00011011100 (.a(t0_000110111000), .b(t0_000110111001), .y(t0_00011011100));
wire t0_000110111000, t0_000110111001;
mixer mix_t0_00011011101 (.a(t0_000110111010), .b(t0_000110111011), .y(t0_00011011101));
wire t0_000110111010, t0_000110111011;
mixer mix_t0_0001101111 (.a(t0_00011011110), .b(t0_00011011111), .y(t0_0001101111));
wire t0_00011011110, t0_00011011111;
mixer mix_t0_00011011110 (.a(t0_000110111100), .b(t0_000110111101), .y(t0_00011011110));
wire t0_000110111100, t0_000110111101;
mixer mix_t0_00011011111 (.a(t0_000110111110), .b(t0_000110111111), .y(t0_00011011111));
wire t0_000110111110, t0_000110111111;
mixer mix_t0_000111 (.a(t0_0001110), .b(t0_0001111), .y(t0_000111));
wire t0_0001110, t0_0001111;
mixer mix_t0_0001110 (.a(t0_00011100), .b(t0_00011101), .y(t0_0001110));
wire t0_00011100, t0_00011101;
mixer mix_t0_00011100 (.a(t0_000111000), .b(t0_000111001), .y(t0_00011100));
wire t0_000111000, t0_000111001;
mixer mix_t0_000111000 (.a(t0_0001110000), .b(t0_0001110001), .y(t0_000111000));
wire t0_0001110000, t0_0001110001;
mixer mix_t0_0001110000 (.a(t0_00011100000), .b(t0_00011100001), .y(t0_0001110000));
wire t0_00011100000, t0_00011100001;
mixer mix_t0_00011100000 (.a(t0_000111000000), .b(t0_000111000001), .y(t0_00011100000));
wire t0_000111000000, t0_000111000001;
mixer mix_t0_00011100001 (.a(t0_000111000010), .b(t0_000111000011), .y(t0_00011100001));
wire t0_000111000010, t0_000111000011;
mixer mix_t0_0001110001 (.a(t0_00011100010), .b(t0_00011100011), .y(t0_0001110001));
wire t0_00011100010, t0_00011100011;
mixer mix_t0_00011100010 (.a(t0_000111000100), .b(t0_000111000101), .y(t0_00011100010));
wire t0_000111000100, t0_000111000101;
mixer mix_t0_00011100011 (.a(t0_000111000110), .b(t0_000111000111), .y(t0_00011100011));
wire t0_000111000110, t0_000111000111;
mixer mix_t0_000111001 (.a(t0_0001110010), .b(t0_0001110011), .y(t0_000111001));
wire t0_0001110010, t0_0001110011;
mixer mix_t0_0001110010 (.a(t0_00011100100), .b(t0_00011100101), .y(t0_0001110010));
wire t0_00011100100, t0_00011100101;
mixer mix_t0_00011100100 (.a(t0_000111001000), .b(t0_000111001001), .y(t0_00011100100));
wire t0_000111001000, t0_000111001001;
mixer mix_t0_00011100101 (.a(t0_000111001010), .b(t0_000111001011), .y(t0_00011100101));
wire t0_000111001010, t0_000111001011;
mixer mix_t0_0001110011 (.a(t0_00011100110), .b(t0_00011100111), .y(t0_0001110011));
wire t0_00011100110, t0_00011100111;
mixer mix_t0_00011100110 (.a(t0_000111001100), .b(t0_000111001101), .y(t0_00011100110));
wire t0_000111001100, t0_000111001101;
mixer mix_t0_00011100111 (.a(t0_000111001110), .b(t0_000111001111), .y(t0_00011100111));
wire t0_000111001110, t0_000111001111;
mixer mix_t0_00011101 (.a(t0_000111010), .b(t0_000111011), .y(t0_00011101));
wire t0_000111010, t0_000111011;
mixer mix_t0_000111010 (.a(t0_0001110100), .b(t0_0001110101), .y(t0_000111010));
wire t0_0001110100, t0_0001110101;
mixer mix_t0_0001110100 (.a(t0_00011101000), .b(t0_00011101001), .y(t0_0001110100));
wire t0_00011101000, t0_00011101001;
mixer mix_t0_00011101000 (.a(t0_000111010000), .b(t0_000111010001), .y(t0_00011101000));
wire t0_000111010000, t0_000111010001;
mixer mix_t0_00011101001 (.a(t0_000111010010), .b(t0_000111010011), .y(t0_00011101001));
wire t0_000111010010, t0_000111010011;
mixer mix_t0_0001110101 (.a(t0_00011101010), .b(t0_00011101011), .y(t0_0001110101));
wire t0_00011101010, t0_00011101011;
mixer mix_t0_00011101010 (.a(t0_000111010100), .b(t0_000111010101), .y(t0_00011101010));
wire t0_000111010100, t0_000111010101;
mixer mix_t0_00011101011 (.a(t0_000111010110), .b(t0_000111010111), .y(t0_00011101011));
wire t0_000111010110, t0_000111010111;
mixer mix_t0_000111011 (.a(t0_0001110110), .b(t0_0001110111), .y(t0_000111011));
wire t0_0001110110, t0_0001110111;
mixer mix_t0_0001110110 (.a(t0_00011101100), .b(t0_00011101101), .y(t0_0001110110));
wire t0_00011101100, t0_00011101101;
mixer mix_t0_00011101100 (.a(t0_000111011000), .b(t0_000111011001), .y(t0_00011101100));
wire t0_000111011000, t0_000111011001;
mixer mix_t0_00011101101 (.a(t0_000111011010), .b(t0_000111011011), .y(t0_00011101101));
wire t0_000111011010, t0_000111011011;
mixer mix_t0_0001110111 (.a(t0_00011101110), .b(t0_00011101111), .y(t0_0001110111));
wire t0_00011101110, t0_00011101111;
mixer mix_t0_00011101110 (.a(t0_000111011100), .b(t0_000111011101), .y(t0_00011101110));
wire t0_000111011100, t0_000111011101;
mixer mix_t0_00011101111 (.a(t0_000111011110), .b(t0_000111011111), .y(t0_00011101111));
wire t0_000111011110, t0_000111011111;
mixer mix_t0_0001111 (.a(t0_00011110), .b(t0_00011111), .y(t0_0001111));
wire t0_00011110, t0_00011111;
mixer mix_t0_00011110 (.a(t0_000111100), .b(t0_000111101), .y(t0_00011110));
wire t0_000111100, t0_000111101;
mixer mix_t0_000111100 (.a(t0_0001111000), .b(t0_0001111001), .y(t0_000111100));
wire t0_0001111000, t0_0001111001;
mixer mix_t0_0001111000 (.a(t0_00011110000), .b(t0_00011110001), .y(t0_0001111000));
wire t0_00011110000, t0_00011110001;
mixer mix_t0_00011110000 (.a(t0_000111100000), .b(t0_000111100001), .y(t0_00011110000));
wire t0_000111100000, t0_000111100001;
mixer mix_t0_00011110001 (.a(t0_000111100010), .b(t0_000111100011), .y(t0_00011110001));
wire t0_000111100010, t0_000111100011;
mixer mix_t0_0001111001 (.a(t0_00011110010), .b(t0_00011110011), .y(t0_0001111001));
wire t0_00011110010, t0_00011110011;
mixer mix_t0_00011110010 (.a(t0_000111100100), .b(t0_000111100101), .y(t0_00011110010));
wire t0_000111100100, t0_000111100101;
mixer mix_t0_00011110011 (.a(t0_000111100110), .b(t0_000111100111), .y(t0_00011110011));
wire t0_000111100110, t0_000111100111;
mixer mix_t0_000111101 (.a(t0_0001111010), .b(t0_0001111011), .y(t0_000111101));
wire t0_0001111010, t0_0001111011;
mixer mix_t0_0001111010 (.a(t0_00011110100), .b(t0_00011110101), .y(t0_0001111010));
wire t0_00011110100, t0_00011110101;
mixer mix_t0_00011110100 (.a(t0_000111101000), .b(t0_000111101001), .y(t0_00011110100));
wire t0_000111101000, t0_000111101001;
mixer mix_t0_00011110101 (.a(t0_000111101010), .b(t0_000111101011), .y(t0_00011110101));
wire t0_000111101010, t0_000111101011;
mixer mix_t0_0001111011 (.a(t0_00011110110), .b(t0_00011110111), .y(t0_0001111011));
wire t0_00011110110, t0_00011110111;
mixer mix_t0_00011110110 (.a(t0_000111101100), .b(t0_000111101101), .y(t0_00011110110));
wire t0_000111101100, t0_000111101101;
mixer mix_t0_00011110111 (.a(t0_000111101110), .b(t0_000111101111), .y(t0_00011110111));
wire t0_000111101110, t0_000111101111;
mixer mix_t0_00011111 (.a(t0_000111110), .b(t0_000111111), .y(t0_00011111));
wire t0_000111110, t0_000111111;
mixer mix_t0_000111110 (.a(t0_0001111100), .b(t0_0001111101), .y(t0_000111110));
wire t0_0001111100, t0_0001111101;
mixer mix_t0_0001111100 (.a(t0_00011111000), .b(t0_00011111001), .y(t0_0001111100));
wire t0_00011111000, t0_00011111001;
mixer mix_t0_00011111000 (.a(t0_000111110000), .b(t0_000111110001), .y(t0_00011111000));
wire t0_000111110000, t0_000111110001;
mixer mix_t0_00011111001 (.a(t0_000111110010), .b(t0_000111110011), .y(t0_00011111001));
wire t0_000111110010, t0_000111110011;
mixer mix_t0_0001111101 (.a(t0_00011111010), .b(t0_00011111011), .y(t0_0001111101));
wire t0_00011111010, t0_00011111011;
mixer mix_t0_00011111010 (.a(t0_000111110100), .b(t0_000111110101), .y(t0_00011111010));
wire t0_000111110100, t0_000111110101;
mixer mix_t0_00011111011 (.a(t0_000111110110), .b(t0_000111110111), .y(t0_00011111011));
wire t0_000111110110, t0_000111110111;
mixer mix_t0_000111111 (.a(t0_0001111110), .b(t0_0001111111), .y(t0_000111111));
wire t0_0001111110, t0_0001111111;
mixer mix_t0_0001111110 (.a(t0_00011111100), .b(t0_00011111101), .y(t0_0001111110));
wire t0_00011111100, t0_00011111101;
mixer mix_t0_00011111100 (.a(t0_000111111000), .b(t0_000111111001), .y(t0_00011111100));
wire t0_000111111000, t0_000111111001;
mixer mix_t0_00011111101 (.a(t0_000111111010), .b(t0_000111111011), .y(t0_00011111101));
wire t0_000111111010, t0_000111111011;
mixer mix_t0_0001111111 (.a(t0_00011111110), .b(t0_00011111111), .y(t0_0001111111));
wire t0_00011111110, t0_00011111111;
mixer mix_t0_00011111110 (.a(t0_000111111100), .b(t0_000111111101), .y(t0_00011111110));
wire t0_000111111100, t0_000111111101;
mixer mix_t0_00011111111 (.a(t0_000111111110), .b(t0_000111111111), .y(t0_00011111111));
wire t0_000111111110, t0_000111111111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_001000 (.a(t0_0010000), .b(t0_0010001), .y(t0_001000));
wire t0_0010000, t0_0010001;
mixer mix_t0_0010000 (.a(t0_00100000), .b(t0_00100001), .y(t0_0010000));
wire t0_00100000, t0_00100001;
mixer mix_t0_00100000 (.a(t0_001000000), .b(t0_001000001), .y(t0_00100000));
wire t0_001000000, t0_001000001;
mixer mix_t0_001000000 (.a(t0_0010000000), .b(t0_0010000001), .y(t0_001000000));
wire t0_0010000000, t0_0010000001;
mixer mix_t0_0010000000 (.a(t0_00100000000), .b(t0_00100000001), .y(t0_0010000000));
wire t0_00100000000, t0_00100000001;
mixer mix_t0_00100000000 (.a(t0_001000000000), .b(t0_001000000001), .y(t0_00100000000));
wire t0_001000000000, t0_001000000001;
mixer mix_t0_00100000001 (.a(t0_001000000010), .b(t0_001000000011), .y(t0_00100000001));
wire t0_001000000010, t0_001000000011;
mixer mix_t0_0010000001 (.a(t0_00100000010), .b(t0_00100000011), .y(t0_0010000001));
wire t0_00100000010, t0_00100000011;
mixer mix_t0_00100000010 (.a(t0_001000000100), .b(t0_001000000101), .y(t0_00100000010));
wire t0_001000000100, t0_001000000101;
mixer mix_t0_00100000011 (.a(t0_001000000110), .b(t0_001000000111), .y(t0_00100000011));
wire t0_001000000110, t0_001000000111;
mixer mix_t0_001000001 (.a(t0_0010000010), .b(t0_0010000011), .y(t0_001000001));
wire t0_0010000010, t0_0010000011;
mixer mix_t0_0010000010 (.a(t0_00100000100), .b(t0_00100000101), .y(t0_0010000010));
wire t0_00100000100, t0_00100000101;
mixer mix_t0_00100000100 (.a(t0_001000001000), .b(t0_001000001001), .y(t0_00100000100));
wire t0_001000001000, t0_001000001001;
mixer mix_t0_00100000101 (.a(t0_001000001010), .b(t0_001000001011), .y(t0_00100000101));
wire t0_001000001010, t0_001000001011;
mixer mix_t0_0010000011 (.a(t0_00100000110), .b(t0_00100000111), .y(t0_0010000011));
wire t0_00100000110, t0_00100000111;
mixer mix_t0_00100000110 (.a(t0_001000001100), .b(t0_001000001101), .y(t0_00100000110));
wire t0_001000001100, t0_001000001101;
mixer mix_t0_00100000111 (.a(t0_001000001110), .b(t0_001000001111), .y(t0_00100000111));
wire t0_001000001110, t0_001000001111;
mixer mix_t0_00100001 (.a(t0_001000010), .b(t0_001000011), .y(t0_00100001));
wire t0_001000010, t0_001000011;
mixer mix_t0_001000010 (.a(t0_0010000100), .b(t0_0010000101), .y(t0_001000010));
wire t0_0010000100, t0_0010000101;
mixer mix_t0_0010000100 (.a(t0_00100001000), .b(t0_00100001001), .y(t0_0010000100));
wire t0_00100001000, t0_00100001001;
mixer mix_t0_00100001000 (.a(t0_001000010000), .b(t0_001000010001), .y(t0_00100001000));
wire t0_001000010000, t0_001000010001;
mixer mix_t0_00100001001 (.a(t0_001000010010), .b(t0_001000010011), .y(t0_00100001001));
wire t0_001000010010, t0_001000010011;
mixer mix_t0_0010000101 (.a(t0_00100001010), .b(t0_00100001011), .y(t0_0010000101));
wire t0_00100001010, t0_00100001011;
mixer mix_t0_00100001010 (.a(t0_001000010100), .b(t0_001000010101), .y(t0_00100001010));
wire t0_001000010100, t0_001000010101;
mixer mix_t0_00100001011 (.a(t0_001000010110), .b(t0_001000010111), .y(t0_00100001011));
wire t0_001000010110, t0_001000010111;
mixer mix_t0_001000011 (.a(t0_0010000110), .b(t0_0010000111), .y(t0_001000011));
wire t0_0010000110, t0_0010000111;
mixer mix_t0_0010000110 (.a(t0_00100001100), .b(t0_00100001101), .y(t0_0010000110));
wire t0_00100001100, t0_00100001101;
mixer mix_t0_00100001100 (.a(t0_001000011000), .b(t0_001000011001), .y(t0_00100001100));
wire t0_001000011000, t0_001000011001;
mixer mix_t0_00100001101 (.a(t0_001000011010), .b(t0_001000011011), .y(t0_00100001101));
wire t0_001000011010, t0_001000011011;
mixer mix_t0_0010000111 (.a(t0_00100001110), .b(t0_00100001111), .y(t0_0010000111));
wire t0_00100001110, t0_00100001111;
mixer mix_t0_00100001110 (.a(t0_001000011100), .b(t0_001000011101), .y(t0_00100001110));
wire t0_001000011100, t0_001000011101;
mixer mix_t0_00100001111 (.a(t0_001000011110), .b(t0_001000011111), .y(t0_00100001111));
wire t0_001000011110, t0_001000011111;
mixer mix_t0_0010001 (.a(t0_00100010), .b(t0_00100011), .y(t0_0010001));
wire t0_00100010, t0_00100011;
mixer mix_t0_00100010 (.a(t0_001000100), .b(t0_001000101), .y(t0_00100010));
wire t0_001000100, t0_001000101;
mixer mix_t0_001000100 (.a(t0_0010001000), .b(t0_0010001001), .y(t0_001000100));
wire t0_0010001000, t0_0010001001;
mixer mix_t0_0010001000 (.a(t0_00100010000), .b(t0_00100010001), .y(t0_0010001000));
wire t0_00100010000, t0_00100010001;
mixer mix_t0_00100010000 (.a(t0_001000100000), .b(t0_001000100001), .y(t0_00100010000));
wire t0_001000100000, t0_001000100001;
mixer mix_t0_00100010001 (.a(t0_001000100010), .b(t0_001000100011), .y(t0_00100010001));
wire t0_001000100010, t0_001000100011;
mixer mix_t0_0010001001 (.a(t0_00100010010), .b(t0_00100010011), .y(t0_0010001001));
wire t0_00100010010, t0_00100010011;
mixer mix_t0_00100010010 (.a(t0_001000100100), .b(t0_001000100101), .y(t0_00100010010));
wire t0_001000100100, t0_001000100101;
mixer mix_t0_00100010011 (.a(t0_001000100110), .b(t0_001000100111), .y(t0_00100010011));
wire t0_001000100110, t0_001000100111;
mixer mix_t0_001000101 (.a(t0_0010001010), .b(t0_0010001011), .y(t0_001000101));
wire t0_0010001010, t0_0010001011;
mixer mix_t0_0010001010 (.a(t0_00100010100), .b(t0_00100010101), .y(t0_0010001010));
wire t0_00100010100, t0_00100010101;
mixer mix_t0_00100010100 (.a(t0_001000101000), .b(t0_001000101001), .y(t0_00100010100));
wire t0_001000101000, t0_001000101001;
mixer mix_t0_00100010101 (.a(t0_001000101010), .b(t0_001000101011), .y(t0_00100010101));
wire t0_001000101010, t0_001000101011;
mixer mix_t0_0010001011 (.a(t0_00100010110), .b(t0_00100010111), .y(t0_0010001011));
wire t0_00100010110, t0_00100010111;
mixer mix_t0_00100010110 (.a(t0_001000101100), .b(t0_001000101101), .y(t0_00100010110));
wire t0_001000101100, t0_001000101101;
mixer mix_t0_00100010111 (.a(t0_001000101110), .b(t0_001000101111), .y(t0_00100010111));
wire t0_001000101110, t0_001000101111;
mixer mix_t0_00100011 (.a(t0_001000110), .b(t0_001000111), .y(t0_00100011));
wire t0_001000110, t0_001000111;
mixer mix_t0_001000110 (.a(t0_0010001100), .b(t0_0010001101), .y(t0_001000110));
wire t0_0010001100, t0_0010001101;
mixer mix_t0_0010001100 (.a(t0_00100011000), .b(t0_00100011001), .y(t0_0010001100));
wire t0_00100011000, t0_00100011001;
mixer mix_t0_00100011000 (.a(t0_001000110000), .b(t0_001000110001), .y(t0_00100011000));
wire t0_001000110000, t0_001000110001;
mixer mix_t0_00100011001 (.a(t0_001000110010), .b(t0_001000110011), .y(t0_00100011001));
wire t0_001000110010, t0_001000110011;
mixer mix_t0_0010001101 (.a(t0_00100011010), .b(t0_00100011011), .y(t0_0010001101));
wire t0_00100011010, t0_00100011011;
mixer mix_t0_00100011010 (.a(t0_001000110100), .b(t0_001000110101), .y(t0_00100011010));
wire t0_001000110100, t0_001000110101;
mixer mix_t0_00100011011 (.a(t0_001000110110), .b(t0_001000110111), .y(t0_00100011011));
wire t0_001000110110, t0_001000110111;
mixer mix_t0_001000111 (.a(t0_0010001110), .b(t0_0010001111), .y(t0_001000111));
wire t0_0010001110, t0_0010001111;
mixer mix_t0_0010001110 (.a(t0_00100011100), .b(t0_00100011101), .y(t0_0010001110));
wire t0_00100011100, t0_00100011101;
mixer mix_t0_00100011100 (.a(t0_001000111000), .b(t0_001000111001), .y(t0_00100011100));
wire t0_001000111000, t0_001000111001;
mixer mix_t0_00100011101 (.a(t0_001000111010), .b(t0_001000111011), .y(t0_00100011101));
wire t0_001000111010, t0_001000111011;
mixer mix_t0_0010001111 (.a(t0_00100011110), .b(t0_00100011111), .y(t0_0010001111));
wire t0_00100011110, t0_00100011111;
mixer mix_t0_00100011110 (.a(t0_001000111100), .b(t0_001000111101), .y(t0_00100011110));
wire t0_001000111100, t0_001000111101;
mixer mix_t0_00100011111 (.a(t0_001000111110), .b(t0_001000111111), .y(t0_00100011111));
wire t0_001000111110, t0_001000111111;
mixer mix_t0_001001 (.a(t0_0010010), .b(t0_0010011), .y(t0_001001));
wire t0_0010010, t0_0010011;
mixer mix_t0_0010010 (.a(t0_00100100), .b(t0_00100101), .y(t0_0010010));
wire t0_00100100, t0_00100101;
mixer mix_t0_00100100 (.a(t0_001001000), .b(t0_001001001), .y(t0_00100100));
wire t0_001001000, t0_001001001;
mixer mix_t0_001001000 (.a(t0_0010010000), .b(t0_0010010001), .y(t0_001001000));
wire t0_0010010000, t0_0010010001;
mixer mix_t0_0010010000 (.a(t0_00100100000), .b(t0_00100100001), .y(t0_0010010000));
wire t0_00100100000, t0_00100100001;
mixer mix_t0_00100100000 (.a(t0_001001000000), .b(t0_001001000001), .y(t0_00100100000));
wire t0_001001000000, t0_001001000001;
mixer mix_t0_00100100001 (.a(t0_001001000010), .b(t0_001001000011), .y(t0_00100100001));
wire t0_001001000010, t0_001001000011;
mixer mix_t0_0010010001 (.a(t0_00100100010), .b(t0_00100100011), .y(t0_0010010001));
wire t0_00100100010, t0_00100100011;
mixer mix_t0_00100100010 (.a(t0_001001000100), .b(t0_001001000101), .y(t0_00100100010));
wire t0_001001000100, t0_001001000101;
mixer mix_t0_00100100011 (.a(t0_001001000110), .b(t0_001001000111), .y(t0_00100100011));
wire t0_001001000110, t0_001001000111;
mixer mix_t0_001001001 (.a(t0_0010010010), .b(t0_0010010011), .y(t0_001001001));
wire t0_0010010010, t0_0010010011;
mixer mix_t0_0010010010 (.a(t0_00100100100), .b(t0_00100100101), .y(t0_0010010010));
wire t0_00100100100, t0_00100100101;
mixer mix_t0_00100100100 (.a(t0_001001001000), .b(t0_001001001001), .y(t0_00100100100));
wire t0_001001001000, t0_001001001001;
mixer mix_t0_00100100101 (.a(t0_001001001010), .b(t0_001001001011), .y(t0_00100100101));
wire t0_001001001010, t0_001001001011;
mixer mix_t0_0010010011 (.a(t0_00100100110), .b(t0_00100100111), .y(t0_0010010011));
wire t0_00100100110, t0_00100100111;
mixer mix_t0_00100100110 (.a(t0_001001001100), .b(t0_001001001101), .y(t0_00100100110));
wire t0_001001001100, t0_001001001101;
mixer mix_t0_00100100111 (.a(t0_001001001110), .b(t0_001001001111), .y(t0_00100100111));
wire t0_001001001110, t0_001001001111;
mixer mix_t0_00100101 (.a(t0_001001010), .b(t0_001001011), .y(t0_00100101));
wire t0_001001010, t0_001001011;
mixer mix_t0_001001010 (.a(t0_0010010100), .b(t0_0010010101), .y(t0_001001010));
wire t0_0010010100, t0_0010010101;
mixer mix_t0_0010010100 (.a(t0_00100101000), .b(t0_00100101001), .y(t0_0010010100));
wire t0_00100101000, t0_00100101001;
mixer mix_t0_00100101000 (.a(t0_001001010000), .b(t0_001001010001), .y(t0_00100101000));
wire t0_001001010000, t0_001001010001;
mixer mix_t0_00100101001 (.a(t0_001001010010), .b(t0_001001010011), .y(t0_00100101001));
wire t0_001001010010, t0_001001010011;
mixer mix_t0_0010010101 (.a(t0_00100101010), .b(t0_00100101011), .y(t0_0010010101));
wire t0_00100101010, t0_00100101011;
mixer mix_t0_00100101010 (.a(t0_001001010100), .b(t0_001001010101), .y(t0_00100101010));
wire t0_001001010100, t0_001001010101;
mixer mix_t0_00100101011 (.a(t0_001001010110), .b(t0_001001010111), .y(t0_00100101011));
wire t0_001001010110, t0_001001010111;
mixer mix_t0_001001011 (.a(t0_0010010110), .b(t0_0010010111), .y(t0_001001011));
wire t0_0010010110, t0_0010010111;
mixer mix_t0_0010010110 (.a(t0_00100101100), .b(t0_00100101101), .y(t0_0010010110));
wire t0_00100101100, t0_00100101101;
mixer mix_t0_00100101100 (.a(t0_001001011000), .b(t0_001001011001), .y(t0_00100101100));
wire t0_001001011000, t0_001001011001;
mixer mix_t0_00100101101 (.a(t0_001001011010), .b(t0_001001011011), .y(t0_00100101101));
wire t0_001001011010, t0_001001011011;
mixer mix_t0_0010010111 (.a(t0_00100101110), .b(t0_00100101111), .y(t0_0010010111));
wire t0_00100101110, t0_00100101111;
mixer mix_t0_00100101110 (.a(t0_001001011100), .b(t0_001001011101), .y(t0_00100101110));
wire t0_001001011100, t0_001001011101;
mixer mix_t0_00100101111 (.a(t0_001001011110), .b(t0_001001011111), .y(t0_00100101111));
wire t0_001001011110, t0_001001011111;
mixer mix_t0_0010011 (.a(t0_00100110), .b(t0_00100111), .y(t0_0010011));
wire t0_00100110, t0_00100111;
mixer mix_t0_00100110 (.a(t0_001001100), .b(t0_001001101), .y(t0_00100110));
wire t0_001001100, t0_001001101;
mixer mix_t0_001001100 (.a(t0_0010011000), .b(t0_0010011001), .y(t0_001001100));
wire t0_0010011000, t0_0010011001;
mixer mix_t0_0010011000 (.a(t0_00100110000), .b(t0_00100110001), .y(t0_0010011000));
wire t0_00100110000, t0_00100110001;
mixer mix_t0_00100110000 (.a(t0_001001100000), .b(t0_001001100001), .y(t0_00100110000));
wire t0_001001100000, t0_001001100001;
mixer mix_t0_00100110001 (.a(t0_001001100010), .b(t0_001001100011), .y(t0_00100110001));
wire t0_001001100010, t0_001001100011;
mixer mix_t0_0010011001 (.a(t0_00100110010), .b(t0_00100110011), .y(t0_0010011001));
wire t0_00100110010, t0_00100110011;
mixer mix_t0_00100110010 (.a(t0_001001100100), .b(t0_001001100101), .y(t0_00100110010));
wire t0_001001100100, t0_001001100101;
mixer mix_t0_00100110011 (.a(t0_001001100110), .b(t0_001001100111), .y(t0_00100110011));
wire t0_001001100110, t0_001001100111;
mixer mix_t0_001001101 (.a(t0_0010011010), .b(t0_0010011011), .y(t0_001001101));
wire t0_0010011010, t0_0010011011;
mixer mix_t0_0010011010 (.a(t0_00100110100), .b(t0_00100110101), .y(t0_0010011010));
wire t0_00100110100, t0_00100110101;
mixer mix_t0_00100110100 (.a(t0_001001101000), .b(t0_001001101001), .y(t0_00100110100));
wire t0_001001101000, t0_001001101001;
mixer mix_t0_00100110101 (.a(t0_001001101010), .b(t0_001001101011), .y(t0_00100110101));
wire t0_001001101010, t0_001001101011;
mixer mix_t0_0010011011 (.a(t0_00100110110), .b(t0_00100110111), .y(t0_0010011011));
wire t0_00100110110, t0_00100110111;
mixer mix_t0_00100110110 (.a(t0_001001101100), .b(t0_001001101101), .y(t0_00100110110));
wire t0_001001101100, t0_001001101101;
mixer mix_t0_00100110111 (.a(t0_001001101110), .b(t0_001001101111), .y(t0_00100110111));
wire t0_001001101110, t0_001001101111;
mixer mix_t0_00100111 (.a(t0_001001110), .b(t0_001001111), .y(t0_00100111));
wire t0_001001110, t0_001001111;
mixer mix_t0_001001110 (.a(t0_0010011100), .b(t0_0010011101), .y(t0_001001110));
wire t0_0010011100, t0_0010011101;
mixer mix_t0_0010011100 (.a(t0_00100111000), .b(t0_00100111001), .y(t0_0010011100));
wire t0_00100111000, t0_00100111001;
mixer mix_t0_00100111000 (.a(t0_001001110000), .b(t0_001001110001), .y(t0_00100111000));
wire t0_001001110000, t0_001001110001;
mixer mix_t0_00100111001 (.a(t0_001001110010), .b(t0_001001110011), .y(t0_00100111001));
wire t0_001001110010, t0_001001110011;
mixer mix_t0_0010011101 (.a(t0_00100111010), .b(t0_00100111011), .y(t0_0010011101));
wire t0_00100111010, t0_00100111011;
mixer mix_t0_00100111010 (.a(t0_001001110100), .b(t0_001001110101), .y(t0_00100111010));
wire t0_001001110100, t0_001001110101;
mixer mix_t0_00100111011 (.a(t0_001001110110), .b(t0_001001110111), .y(t0_00100111011));
wire t0_001001110110, t0_001001110111;
mixer mix_t0_001001111 (.a(t0_0010011110), .b(t0_0010011111), .y(t0_001001111));
wire t0_0010011110, t0_0010011111;
mixer mix_t0_0010011110 (.a(t0_00100111100), .b(t0_00100111101), .y(t0_0010011110));
wire t0_00100111100, t0_00100111101;
mixer mix_t0_00100111100 (.a(t0_001001111000), .b(t0_001001111001), .y(t0_00100111100));
wire t0_001001111000, t0_001001111001;
mixer mix_t0_00100111101 (.a(t0_001001111010), .b(t0_001001111011), .y(t0_00100111101));
wire t0_001001111010, t0_001001111011;
mixer mix_t0_0010011111 (.a(t0_00100111110), .b(t0_00100111111), .y(t0_0010011111));
wire t0_00100111110, t0_00100111111;
mixer mix_t0_00100111110 (.a(t0_001001111100), .b(t0_001001111101), .y(t0_00100111110));
wire t0_001001111100, t0_001001111101;
mixer mix_t0_00100111111 (.a(t0_001001111110), .b(t0_001001111111), .y(t0_00100111111));
wire t0_001001111110, t0_001001111111;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_001010 (.a(t0_0010100), .b(t0_0010101), .y(t0_001010));
wire t0_0010100, t0_0010101;
mixer mix_t0_0010100 (.a(t0_00101000), .b(t0_00101001), .y(t0_0010100));
wire t0_00101000, t0_00101001;
mixer mix_t0_00101000 (.a(t0_001010000), .b(t0_001010001), .y(t0_00101000));
wire t0_001010000, t0_001010001;
mixer mix_t0_001010000 (.a(t0_0010100000), .b(t0_0010100001), .y(t0_001010000));
wire t0_0010100000, t0_0010100001;
mixer mix_t0_0010100000 (.a(t0_00101000000), .b(t0_00101000001), .y(t0_0010100000));
wire t0_00101000000, t0_00101000001;
mixer mix_t0_00101000000 (.a(t0_001010000000), .b(t0_001010000001), .y(t0_00101000000));
wire t0_001010000000, t0_001010000001;
mixer mix_t0_00101000001 (.a(t0_001010000010), .b(t0_001010000011), .y(t0_00101000001));
wire t0_001010000010, t0_001010000011;
mixer mix_t0_0010100001 (.a(t0_00101000010), .b(t0_00101000011), .y(t0_0010100001));
wire t0_00101000010, t0_00101000011;
mixer mix_t0_00101000010 (.a(t0_001010000100), .b(t0_001010000101), .y(t0_00101000010));
wire t0_001010000100, t0_001010000101;
mixer mix_t0_00101000011 (.a(t0_001010000110), .b(t0_001010000111), .y(t0_00101000011));
wire t0_001010000110, t0_001010000111;
mixer mix_t0_001010001 (.a(t0_0010100010), .b(t0_0010100011), .y(t0_001010001));
wire t0_0010100010, t0_0010100011;
mixer mix_t0_0010100010 (.a(t0_00101000100), .b(t0_00101000101), .y(t0_0010100010));
wire t0_00101000100, t0_00101000101;
mixer mix_t0_00101000100 (.a(t0_001010001000), .b(t0_001010001001), .y(t0_00101000100));
wire t0_001010001000, t0_001010001001;
mixer mix_t0_00101000101 (.a(t0_001010001010), .b(t0_001010001011), .y(t0_00101000101));
wire t0_001010001010, t0_001010001011;
mixer mix_t0_0010100011 (.a(t0_00101000110), .b(t0_00101000111), .y(t0_0010100011));
wire t0_00101000110, t0_00101000111;
mixer mix_t0_00101000110 (.a(t0_001010001100), .b(t0_001010001101), .y(t0_00101000110));
wire t0_001010001100, t0_001010001101;
mixer mix_t0_00101000111 (.a(t0_001010001110), .b(t0_001010001111), .y(t0_00101000111));
wire t0_001010001110, t0_001010001111;
mixer mix_t0_00101001 (.a(t0_001010010), .b(t0_001010011), .y(t0_00101001));
wire t0_001010010, t0_001010011;
mixer mix_t0_001010010 (.a(t0_0010100100), .b(t0_0010100101), .y(t0_001010010));
wire t0_0010100100, t0_0010100101;
mixer mix_t0_0010100100 (.a(t0_00101001000), .b(t0_00101001001), .y(t0_0010100100));
wire t0_00101001000, t0_00101001001;
mixer mix_t0_00101001000 (.a(t0_001010010000), .b(t0_001010010001), .y(t0_00101001000));
wire t0_001010010000, t0_001010010001;
mixer mix_t0_00101001001 (.a(t0_001010010010), .b(t0_001010010011), .y(t0_00101001001));
wire t0_001010010010, t0_001010010011;
mixer mix_t0_0010100101 (.a(t0_00101001010), .b(t0_00101001011), .y(t0_0010100101));
wire t0_00101001010, t0_00101001011;
mixer mix_t0_00101001010 (.a(t0_001010010100), .b(t0_001010010101), .y(t0_00101001010));
wire t0_001010010100, t0_001010010101;
mixer mix_t0_00101001011 (.a(t0_001010010110), .b(t0_001010010111), .y(t0_00101001011));
wire t0_001010010110, t0_001010010111;
mixer mix_t0_001010011 (.a(t0_0010100110), .b(t0_0010100111), .y(t0_001010011));
wire t0_0010100110, t0_0010100111;
mixer mix_t0_0010100110 (.a(t0_00101001100), .b(t0_00101001101), .y(t0_0010100110));
wire t0_00101001100, t0_00101001101;
mixer mix_t0_00101001100 (.a(t0_001010011000), .b(t0_001010011001), .y(t0_00101001100));
wire t0_001010011000, t0_001010011001;
mixer mix_t0_00101001101 (.a(t0_001010011010), .b(t0_001010011011), .y(t0_00101001101));
wire t0_001010011010, t0_001010011011;
mixer mix_t0_0010100111 (.a(t0_00101001110), .b(t0_00101001111), .y(t0_0010100111));
wire t0_00101001110, t0_00101001111;
mixer mix_t0_00101001110 (.a(t0_001010011100), .b(t0_001010011101), .y(t0_00101001110));
wire t0_001010011100, t0_001010011101;
mixer mix_t0_00101001111 (.a(t0_001010011110), .b(t0_001010011111), .y(t0_00101001111));
wire t0_001010011110, t0_001010011111;
mixer mix_t0_0010101 (.a(t0_00101010), .b(t0_00101011), .y(t0_0010101));
wire t0_00101010, t0_00101011;
mixer mix_t0_00101010 (.a(t0_001010100), .b(t0_001010101), .y(t0_00101010));
wire t0_001010100, t0_001010101;
mixer mix_t0_001010100 (.a(t0_0010101000), .b(t0_0010101001), .y(t0_001010100));
wire t0_0010101000, t0_0010101001;
mixer mix_t0_0010101000 (.a(t0_00101010000), .b(t0_00101010001), .y(t0_0010101000));
wire t0_00101010000, t0_00101010001;
mixer mix_t0_00101010000 (.a(t0_001010100000), .b(t0_001010100001), .y(t0_00101010000));
wire t0_001010100000, t0_001010100001;
mixer mix_t0_00101010001 (.a(t0_001010100010), .b(t0_001010100011), .y(t0_00101010001));
wire t0_001010100010, t0_001010100011;
mixer mix_t0_0010101001 (.a(t0_00101010010), .b(t0_00101010011), .y(t0_0010101001));
wire t0_00101010010, t0_00101010011;
mixer mix_t0_00101010010 (.a(t0_001010100100), .b(t0_001010100101), .y(t0_00101010010));
wire t0_001010100100, t0_001010100101;
mixer mix_t0_00101010011 (.a(t0_001010100110), .b(t0_001010100111), .y(t0_00101010011));
wire t0_001010100110, t0_001010100111;
mixer mix_t0_001010101 (.a(t0_0010101010), .b(t0_0010101011), .y(t0_001010101));
wire t0_0010101010, t0_0010101011;
mixer mix_t0_0010101010 (.a(t0_00101010100), .b(t0_00101010101), .y(t0_0010101010));
wire t0_00101010100, t0_00101010101;
mixer mix_t0_00101010100 (.a(t0_001010101000), .b(t0_001010101001), .y(t0_00101010100));
wire t0_001010101000, t0_001010101001;
mixer mix_t0_00101010101 (.a(t0_001010101010), .b(t0_001010101011), .y(t0_00101010101));
wire t0_001010101010, t0_001010101011;
mixer mix_t0_0010101011 (.a(t0_00101010110), .b(t0_00101010111), .y(t0_0010101011));
wire t0_00101010110, t0_00101010111;
mixer mix_t0_00101010110 (.a(t0_001010101100), .b(t0_001010101101), .y(t0_00101010110));
wire t0_001010101100, t0_001010101101;
mixer mix_t0_00101010111 (.a(t0_001010101110), .b(t0_001010101111), .y(t0_00101010111));
wire t0_001010101110, t0_001010101111;
mixer mix_t0_00101011 (.a(t0_001010110), .b(t0_001010111), .y(t0_00101011));
wire t0_001010110, t0_001010111;
mixer mix_t0_001010110 (.a(t0_0010101100), .b(t0_0010101101), .y(t0_001010110));
wire t0_0010101100, t0_0010101101;
mixer mix_t0_0010101100 (.a(t0_00101011000), .b(t0_00101011001), .y(t0_0010101100));
wire t0_00101011000, t0_00101011001;
mixer mix_t0_00101011000 (.a(t0_001010110000), .b(t0_001010110001), .y(t0_00101011000));
wire t0_001010110000, t0_001010110001;
mixer mix_t0_00101011001 (.a(t0_001010110010), .b(t0_001010110011), .y(t0_00101011001));
wire t0_001010110010, t0_001010110011;
mixer mix_t0_0010101101 (.a(t0_00101011010), .b(t0_00101011011), .y(t0_0010101101));
wire t0_00101011010, t0_00101011011;
mixer mix_t0_00101011010 (.a(t0_001010110100), .b(t0_001010110101), .y(t0_00101011010));
wire t0_001010110100, t0_001010110101;
mixer mix_t0_00101011011 (.a(t0_001010110110), .b(t0_001010110111), .y(t0_00101011011));
wire t0_001010110110, t0_001010110111;
mixer mix_t0_001010111 (.a(t0_0010101110), .b(t0_0010101111), .y(t0_001010111));
wire t0_0010101110, t0_0010101111;
mixer mix_t0_0010101110 (.a(t0_00101011100), .b(t0_00101011101), .y(t0_0010101110));
wire t0_00101011100, t0_00101011101;
mixer mix_t0_00101011100 (.a(t0_001010111000), .b(t0_001010111001), .y(t0_00101011100));
wire t0_001010111000, t0_001010111001;
mixer mix_t0_00101011101 (.a(t0_001010111010), .b(t0_001010111011), .y(t0_00101011101));
wire t0_001010111010, t0_001010111011;
mixer mix_t0_0010101111 (.a(t0_00101011110), .b(t0_00101011111), .y(t0_0010101111));
wire t0_00101011110, t0_00101011111;
mixer mix_t0_00101011110 (.a(t0_001010111100), .b(t0_001010111101), .y(t0_00101011110));
wire t0_001010111100, t0_001010111101;
mixer mix_t0_00101011111 (.a(t0_001010111110), .b(t0_001010111111), .y(t0_00101011111));
wire t0_001010111110, t0_001010111111;
mixer mix_t0_001011 (.a(t0_0010110), .b(t0_0010111), .y(t0_001011));
wire t0_0010110, t0_0010111;
mixer mix_t0_0010110 (.a(t0_00101100), .b(t0_00101101), .y(t0_0010110));
wire t0_00101100, t0_00101101;
mixer mix_t0_00101100 (.a(t0_001011000), .b(t0_001011001), .y(t0_00101100));
wire t0_001011000, t0_001011001;
mixer mix_t0_001011000 (.a(t0_0010110000), .b(t0_0010110001), .y(t0_001011000));
wire t0_0010110000, t0_0010110001;
mixer mix_t0_0010110000 (.a(t0_00101100000), .b(t0_00101100001), .y(t0_0010110000));
wire t0_00101100000, t0_00101100001;
mixer mix_t0_00101100000 (.a(t0_001011000000), .b(t0_001011000001), .y(t0_00101100000));
wire t0_001011000000, t0_001011000001;
mixer mix_t0_00101100001 (.a(t0_001011000010), .b(t0_001011000011), .y(t0_00101100001));
wire t0_001011000010, t0_001011000011;
mixer mix_t0_0010110001 (.a(t0_00101100010), .b(t0_00101100011), .y(t0_0010110001));
wire t0_00101100010, t0_00101100011;
mixer mix_t0_00101100010 (.a(t0_001011000100), .b(t0_001011000101), .y(t0_00101100010));
wire t0_001011000100, t0_001011000101;
mixer mix_t0_00101100011 (.a(t0_001011000110), .b(t0_001011000111), .y(t0_00101100011));
wire t0_001011000110, t0_001011000111;
mixer mix_t0_001011001 (.a(t0_0010110010), .b(t0_0010110011), .y(t0_001011001));
wire t0_0010110010, t0_0010110011;
mixer mix_t0_0010110010 (.a(t0_00101100100), .b(t0_00101100101), .y(t0_0010110010));
wire t0_00101100100, t0_00101100101;
mixer mix_t0_00101100100 (.a(t0_001011001000), .b(t0_001011001001), .y(t0_00101100100));
wire t0_001011001000, t0_001011001001;
mixer mix_t0_00101100101 (.a(t0_001011001010), .b(t0_001011001011), .y(t0_00101100101));
wire t0_001011001010, t0_001011001011;
mixer mix_t0_0010110011 (.a(t0_00101100110), .b(t0_00101100111), .y(t0_0010110011));
wire t0_00101100110, t0_00101100111;
mixer mix_t0_00101100110 (.a(t0_001011001100), .b(t0_001011001101), .y(t0_00101100110));
wire t0_001011001100, t0_001011001101;
mixer mix_t0_00101100111 (.a(t0_001011001110), .b(t0_001011001111), .y(t0_00101100111));
wire t0_001011001110, t0_001011001111;
mixer mix_t0_00101101 (.a(t0_001011010), .b(t0_001011011), .y(t0_00101101));
wire t0_001011010, t0_001011011;
mixer mix_t0_001011010 (.a(t0_0010110100), .b(t0_0010110101), .y(t0_001011010));
wire t0_0010110100, t0_0010110101;
mixer mix_t0_0010110100 (.a(t0_00101101000), .b(t0_00101101001), .y(t0_0010110100));
wire t0_00101101000, t0_00101101001;
mixer mix_t0_00101101000 (.a(t0_001011010000), .b(t0_001011010001), .y(t0_00101101000));
wire t0_001011010000, t0_001011010001;
mixer mix_t0_00101101001 (.a(t0_001011010010), .b(t0_001011010011), .y(t0_00101101001));
wire t0_001011010010, t0_001011010011;
mixer mix_t0_0010110101 (.a(t0_00101101010), .b(t0_00101101011), .y(t0_0010110101));
wire t0_00101101010, t0_00101101011;
mixer mix_t0_00101101010 (.a(t0_001011010100), .b(t0_001011010101), .y(t0_00101101010));
wire t0_001011010100, t0_001011010101;
mixer mix_t0_00101101011 (.a(t0_001011010110), .b(t0_001011010111), .y(t0_00101101011));
wire t0_001011010110, t0_001011010111;
mixer mix_t0_001011011 (.a(t0_0010110110), .b(t0_0010110111), .y(t0_001011011));
wire t0_0010110110, t0_0010110111;
mixer mix_t0_0010110110 (.a(t0_00101101100), .b(t0_00101101101), .y(t0_0010110110));
wire t0_00101101100, t0_00101101101;
mixer mix_t0_00101101100 (.a(t0_001011011000), .b(t0_001011011001), .y(t0_00101101100));
wire t0_001011011000, t0_001011011001;
mixer mix_t0_00101101101 (.a(t0_001011011010), .b(t0_001011011011), .y(t0_00101101101));
wire t0_001011011010, t0_001011011011;
mixer mix_t0_0010110111 (.a(t0_00101101110), .b(t0_00101101111), .y(t0_0010110111));
wire t0_00101101110, t0_00101101111;
mixer mix_t0_00101101110 (.a(t0_001011011100), .b(t0_001011011101), .y(t0_00101101110));
wire t0_001011011100, t0_001011011101;
mixer mix_t0_00101101111 (.a(t0_001011011110), .b(t0_001011011111), .y(t0_00101101111));
wire t0_001011011110, t0_001011011111;
mixer mix_t0_0010111 (.a(t0_00101110), .b(t0_00101111), .y(t0_0010111));
wire t0_00101110, t0_00101111;
mixer mix_t0_00101110 (.a(t0_001011100), .b(t0_001011101), .y(t0_00101110));
wire t0_001011100, t0_001011101;
mixer mix_t0_001011100 (.a(t0_0010111000), .b(t0_0010111001), .y(t0_001011100));
wire t0_0010111000, t0_0010111001;
mixer mix_t0_0010111000 (.a(t0_00101110000), .b(t0_00101110001), .y(t0_0010111000));
wire t0_00101110000, t0_00101110001;
mixer mix_t0_00101110000 (.a(t0_001011100000), .b(t0_001011100001), .y(t0_00101110000));
wire t0_001011100000, t0_001011100001;
mixer mix_t0_00101110001 (.a(t0_001011100010), .b(t0_001011100011), .y(t0_00101110001));
wire t0_001011100010, t0_001011100011;
mixer mix_t0_0010111001 (.a(t0_00101110010), .b(t0_00101110011), .y(t0_0010111001));
wire t0_00101110010, t0_00101110011;
mixer mix_t0_00101110010 (.a(t0_001011100100), .b(t0_001011100101), .y(t0_00101110010));
wire t0_001011100100, t0_001011100101;
mixer mix_t0_00101110011 (.a(t0_001011100110), .b(t0_001011100111), .y(t0_00101110011));
wire t0_001011100110, t0_001011100111;
mixer mix_t0_001011101 (.a(t0_0010111010), .b(t0_0010111011), .y(t0_001011101));
wire t0_0010111010, t0_0010111011;
mixer mix_t0_0010111010 (.a(t0_00101110100), .b(t0_00101110101), .y(t0_0010111010));
wire t0_00101110100, t0_00101110101;
mixer mix_t0_00101110100 (.a(t0_001011101000), .b(t0_001011101001), .y(t0_00101110100));
wire t0_001011101000, t0_001011101001;
mixer mix_t0_00101110101 (.a(t0_001011101010), .b(t0_001011101011), .y(t0_00101110101));
wire t0_001011101010, t0_001011101011;
mixer mix_t0_0010111011 (.a(t0_00101110110), .b(t0_00101110111), .y(t0_0010111011));
wire t0_00101110110, t0_00101110111;
mixer mix_t0_00101110110 (.a(t0_001011101100), .b(t0_001011101101), .y(t0_00101110110));
wire t0_001011101100, t0_001011101101;
mixer mix_t0_00101110111 (.a(t0_001011101110), .b(t0_001011101111), .y(t0_00101110111));
wire t0_001011101110, t0_001011101111;
mixer mix_t0_00101111 (.a(t0_001011110), .b(t0_001011111), .y(t0_00101111));
wire t0_001011110, t0_001011111;
mixer mix_t0_001011110 (.a(t0_0010111100), .b(t0_0010111101), .y(t0_001011110));
wire t0_0010111100, t0_0010111101;
mixer mix_t0_0010111100 (.a(t0_00101111000), .b(t0_00101111001), .y(t0_0010111100));
wire t0_00101111000, t0_00101111001;
mixer mix_t0_00101111000 (.a(t0_001011110000), .b(t0_001011110001), .y(t0_00101111000));
wire t0_001011110000, t0_001011110001;
mixer mix_t0_00101111001 (.a(t0_001011110010), .b(t0_001011110011), .y(t0_00101111001));
wire t0_001011110010, t0_001011110011;
mixer mix_t0_0010111101 (.a(t0_00101111010), .b(t0_00101111011), .y(t0_0010111101));
wire t0_00101111010, t0_00101111011;
mixer mix_t0_00101111010 (.a(t0_001011110100), .b(t0_001011110101), .y(t0_00101111010));
wire t0_001011110100, t0_001011110101;
mixer mix_t0_00101111011 (.a(t0_001011110110), .b(t0_001011110111), .y(t0_00101111011));
wire t0_001011110110, t0_001011110111;
mixer mix_t0_001011111 (.a(t0_0010111110), .b(t0_0010111111), .y(t0_001011111));
wire t0_0010111110, t0_0010111111;
mixer mix_t0_0010111110 (.a(t0_00101111100), .b(t0_00101111101), .y(t0_0010111110));
wire t0_00101111100, t0_00101111101;
mixer mix_t0_00101111100 (.a(t0_001011111000), .b(t0_001011111001), .y(t0_00101111100));
wire t0_001011111000, t0_001011111001;
mixer mix_t0_00101111101 (.a(t0_001011111010), .b(t0_001011111011), .y(t0_00101111101));
wire t0_001011111010, t0_001011111011;
mixer mix_t0_0010111111 (.a(t0_00101111110), .b(t0_00101111111), .y(t0_0010111111));
wire t0_00101111110, t0_00101111111;
mixer mix_t0_00101111110 (.a(t0_001011111100), .b(t0_001011111101), .y(t0_00101111110));
wire t0_001011111100, t0_001011111101;
mixer mix_t0_00101111111 (.a(t0_001011111110), .b(t0_001011111111), .y(t0_00101111111));
wire t0_001011111110, t0_001011111111;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_001100 (.a(t0_0011000), .b(t0_0011001), .y(t0_001100));
wire t0_0011000, t0_0011001;
mixer mix_t0_0011000 (.a(t0_00110000), .b(t0_00110001), .y(t0_0011000));
wire t0_00110000, t0_00110001;
mixer mix_t0_00110000 (.a(t0_001100000), .b(t0_001100001), .y(t0_00110000));
wire t0_001100000, t0_001100001;
mixer mix_t0_001100000 (.a(t0_0011000000), .b(t0_0011000001), .y(t0_001100000));
wire t0_0011000000, t0_0011000001;
mixer mix_t0_0011000000 (.a(t0_00110000000), .b(t0_00110000001), .y(t0_0011000000));
wire t0_00110000000, t0_00110000001;
mixer mix_t0_00110000000 (.a(t0_001100000000), .b(t0_001100000001), .y(t0_00110000000));
wire t0_001100000000, t0_001100000001;
mixer mix_t0_00110000001 (.a(t0_001100000010), .b(t0_001100000011), .y(t0_00110000001));
wire t0_001100000010, t0_001100000011;
mixer mix_t0_0011000001 (.a(t0_00110000010), .b(t0_00110000011), .y(t0_0011000001));
wire t0_00110000010, t0_00110000011;
mixer mix_t0_00110000010 (.a(t0_001100000100), .b(t0_001100000101), .y(t0_00110000010));
wire t0_001100000100, t0_001100000101;
mixer mix_t0_00110000011 (.a(t0_001100000110), .b(t0_001100000111), .y(t0_00110000011));
wire t0_001100000110, t0_001100000111;
mixer mix_t0_001100001 (.a(t0_0011000010), .b(t0_0011000011), .y(t0_001100001));
wire t0_0011000010, t0_0011000011;
mixer mix_t0_0011000010 (.a(t0_00110000100), .b(t0_00110000101), .y(t0_0011000010));
wire t0_00110000100, t0_00110000101;
mixer mix_t0_00110000100 (.a(t0_001100001000), .b(t0_001100001001), .y(t0_00110000100));
wire t0_001100001000, t0_001100001001;
mixer mix_t0_00110000101 (.a(t0_001100001010), .b(t0_001100001011), .y(t0_00110000101));
wire t0_001100001010, t0_001100001011;
mixer mix_t0_0011000011 (.a(t0_00110000110), .b(t0_00110000111), .y(t0_0011000011));
wire t0_00110000110, t0_00110000111;
mixer mix_t0_00110000110 (.a(t0_001100001100), .b(t0_001100001101), .y(t0_00110000110));
wire t0_001100001100, t0_001100001101;
mixer mix_t0_00110000111 (.a(t0_001100001110), .b(t0_001100001111), .y(t0_00110000111));
wire t0_001100001110, t0_001100001111;
mixer mix_t0_00110001 (.a(t0_001100010), .b(t0_001100011), .y(t0_00110001));
wire t0_001100010, t0_001100011;
mixer mix_t0_001100010 (.a(t0_0011000100), .b(t0_0011000101), .y(t0_001100010));
wire t0_0011000100, t0_0011000101;
mixer mix_t0_0011000100 (.a(t0_00110001000), .b(t0_00110001001), .y(t0_0011000100));
wire t0_00110001000, t0_00110001001;
mixer mix_t0_00110001000 (.a(t0_001100010000), .b(t0_001100010001), .y(t0_00110001000));
wire t0_001100010000, t0_001100010001;
mixer mix_t0_00110001001 (.a(t0_001100010010), .b(t0_001100010011), .y(t0_00110001001));
wire t0_001100010010, t0_001100010011;
mixer mix_t0_0011000101 (.a(t0_00110001010), .b(t0_00110001011), .y(t0_0011000101));
wire t0_00110001010, t0_00110001011;
mixer mix_t0_00110001010 (.a(t0_001100010100), .b(t0_001100010101), .y(t0_00110001010));
wire t0_001100010100, t0_001100010101;
mixer mix_t0_00110001011 (.a(t0_001100010110), .b(t0_001100010111), .y(t0_00110001011));
wire t0_001100010110, t0_001100010111;
mixer mix_t0_001100011 (.a(t0_0011000110), .b(t0_0011000111), .y(t0_001100011));
wire t0_0011000110, t0_0011000111;
mixer mix_t0_0011000110 (.a(t0_00110001100), .b(t0_00110001101), .y(t0_0011000110));
wire t0_00110001100, t0_00110001101;
mixer mix_t0_00110001100 (.a(t0_001100011000), .b(t0_001100011001), .y(t0_00110001100));
wire t0_001100011000, t0_001100011001;
mixer mix_t0_00110001101 (.a(t0_001100011010), .b(t0_001100011011), .y(t0_00110001101));
wire t0_001100011010, t0_001100011011;
mixer mix_t0_0011000111 (.a(t0_00110001110), .b(t0_00110001111), .y(t0_0011000111));
wire t0_00110001110, t0_00110001111;
mixer mix_t0_00110001110 (.a(t0_001100011100), .b(t0_001100011101), .y(t0_00110001110));
wire t0_001100011100, t0_001100011101;
mixer mix_t0_00110001111 (.a(t0_001100011110), .b(t0_001100011111), .y(t0_00110001111));
wire t0_001100011110, t0_001100011111;
mixer mix_t0_0011001 (.a(t0_00110010), .b(t0_00110011), .y(t0_0011001));
wire t0_00110010, t0_00110011;
mixer mix_t0_00110010 (.a(t0_001100100), .b(t0_001100101), .y(t0_00110010));
wire t0_001100100, t0_001100101;
mixer mix_t0_001100100 (.a(t0_0011001000), .b(t0_0011001001), .y(t0_001100100));
wire t0_0011001000, t0_0011001001;
mixer mix_t0_0011001000 (.a(t0_00110010000), .b(t0_00110010001), .y(t0_0011001000));
wire t0_00110010000, t0_00110010001;
mixer mix_t0_00110010000 (.a(t0_001100100000), .b(t0_001100100001), .y(t0_00110010000));
wire t0_001100100000, t0_001100100001;
mixer mix_t0_00110010001 (.a(t0_001100100010), .b(t0_001100100011), .y(t0_00110010001));
wire t0_001100100010, t0_001100100011;
mixer mix_t0_0011001001 (.a(t0_00110010010), .b(t0_00110010011), .y(t0_0011001001));
wire t0_00110010010, t0_00110010011;
mixer mix_t0_00110010010 (.a(t0_001100100100), .b(t0_001100100101), .y(t0_00110010010));
wire t0_001100100100, t0_001100100101;
mixer mix_t0_00110010011 (.a(t0_001100100110), .b(t0_001100100111), .y(t0_00110010011));
wire t0_001100100110, t0_001100100111;
mixer mix_t0_001100101 (.a(t0_0011001010), .b(t0_0011001011), .y(t0_001100101));
wire t0_0011001010, t0_0011001011;
mixer mix_t0_0011001010 (.a(t0_00110010100), .b(t0_00110010101), .y(t0_0011001010));
wire t0_00110010100, t0_00110010101;
mixer mix_t0_00110010100 (.a(t0_001100101000), .b(t0_001100101001), .y(t0_00110010100));
wire t0_001100101000, t0_001100101001;
mixer mix_t0_00110010101 (.a(t0_001100101010), .b(t0_001100101011), .y(t0_00110010101));
wire t0_001100101010, t0_001100101011;
mixer mix_t0_0011001011 (.a(t0_00110010110), .b(t0_00110010111), .y(t0_0011001011));
wire t0_00110010110, t0_00110010111;
mixer mix_t0_00110010110 (.a(t0_001100101100), .b(t0_001100101101), .y(t0_00110010110));
wire t0_001100101100, t0_001100101101;
mixer mix_t0_00110010111 (.a(t0_001100101110), .b(t0_001100101111), .y(t0_00110010111));
wire t0_001100101110, t0_001100101111;
mixer mix_t0_00110011 (.a(t0_001100110), .b(t0_001100111), .y(t0_00110011));
wire t0_001100110, t0_001100111;
mixer mix_t0_001100110 (.a(t0_0011001100), .b(t0_0011001101), .y(t0_001100110));
wire t0_0011001100, t0_0011001101;
mixer mix_t0_0011001100 (.a(t0_00110011000), .b(t0_00110011001), .y(t0_0011001100));
wire t0_00110011000, t0_00110011001;
mixer mix_t0_00110011000 (.a(t0_001100110000), .b(t0_001100110001), .y(t0_00110011000));
wire t0_001100110000, t0_001100110001;
mixer mix_t0_00110011001 (.a(t0_001100110010), .b(t0_001100110011), .y(t0_00110011001));
wire t0_001100110010, t0_001100110011;
mixer mix_t0_0011001101 (.a(t0_00110011010), .b(t0_00110011011), .y(t0_0011001101));
wire t0_00110011010, t0_00110011011;
mixer mix_t0_00110011010 (.a(t0_001100110100), .b(t0_001100110101), .y(t0_00110011010));
wire t0_001100110100, t0_001100110101;
mixer mix_t0_00110011011 (.a(t0_001100110110), .b(t0_001100110111), .y(t0_00110011011));
wire t0_001100110110, t0_001100110111;
mixer mix_t0_001100111 (.a(t0_0011001110), .b(t0_0011001111), .y(t0_001100111));
wire t0_0011001110, t0_0011001111;
mixer mix_t0_0011001110 (.a(t0_00110011100), .b(t0_00110011101), .y(t0_0011001110));
wire t0_00110011100, t0_00110011101;
mixer mix_t0_00110011100 (.a(t0_001100111000), .b(t0_001100111001), .y(t0_00110011100));
wire t0_001100111000, t0_001100111001;
mixer mix_t0_00110011101 (.a(t0_001100111010), .b(t0_001100111011), .y(t0_00110011101));
wire t0_001100111010, t0_001100111011;
mixer mix_t0_0011001111 (.a(t0_00110011110), .b(t0_00110011111), .y(t0_0011001111));
wire t0_00110011110, t0_00110011111;
mixer mix_t0_00110011110 (.a(t0_001100111100), .b(t0_001100111101), .y(t0_00110011110));
wire t0_001100111100, t0_001100111101;
mixer mix_t0_00110011111 (.a(t0_001100111110), .b(t0_001100111111), .y(t0_00110011111));
wire t0_001100111110, t0_001100111111;
mixer mix_t0_001101 (.a(t0_0011010), .b(t0_0011011), .y(t0_001101));
wire t0_0011010, t0_0011011;
mixer mix_t0_0011010 (.a(t0_00110100), .b(t0_00110101), .y(t0_0011010));
wire t0_00110100, t0_00110101;
mixer mix_t0_00110100 (.a(t0_001101000), .b(t0_001101001), .y(t0_00110100));
wire t0_001101000, t0_001101001;
mixer mix_t0_001101000 (.a(t0_0011010000), .b(t0_0011010001), .y(t0_001101000));
wire t0_0011010000, t0_0011010001;
mixer mix_t0_0011010000 (.a(t0_00110100000), .b(t0_00110100001), .y(t0_0011010000));
wire t0_00110100000, t0_00110100001;
mixer mix_t0_00110100000 (.a(t0_001101000000), .b(t0_001101000001), .y(t0_00110100000));
wire t0_001101000000, t0_001101000001;
mixer mix_t0_00110100001 (.a(t0_001101000010), .b(t0_001101000011), .y(t0_00110100001));
wire t0_001101000010, t0_001101000011;
mixer mix_t0_0011010001 (.a(t0_00110100010), .b(t0_00110100011), .y(t0_0011010001));
wire t0_00110100010, t0_00110100011;
mixer mix_t0_00110100010 (.a(t0_001101000100), .b(t0_001101000101), .y(t0_00110100010));
wire t0_001101000100, t0_001101000101;
mixer mix_t0_00110100011 (.a(t0_001101000110), .b(t0_001101000111), .y(t0_00110100011));
wire t0_001101000110, t0_001101000111;
mixer mix_t0_001101001 (.a(t0_0011010010), .b(t0_0011010011), .y(t0_001101001));
wire t0_0011010010, t0_0011010011;
mixer mix_t0_0011010010 (.a(t0_00110100100), .b(t0_00110100101), .y(t0_0011010010));
wire t0_00110100100, t0_00110100101;
mixer mix_t0_00110100100 (.a(t0_001101001000), .b(t0_001101001001), .y(t0_00110100100));
wire t0_001101001000, t0_001101001001;
mixer mix_t0_00110100101 (.a(t0_001101001010), .b(t0_001101001011), .y(t0_00110100101));
wire t0_001101001010, t0_001101001011;
mixer mix_t0_0011010011 (.a(t0_00110100110), .b(t0_00110100111), .y(t0_0011010011));
wire t0_00110100110, t0_00110100111;
mixer mix_t0_00110100110 (.a(t0_001101001100), .b(t0_001101001101), .y(t0_00110100110));
wire t0_001101001100, t0_001101001101;
mixer mix_t0_00110100111 (.a(t0_001101001110), .b(t0_001101001111), .y(t0_00110100111));
wire t0_001101001110, t0_001101001111;
mixer mix_t0_00110101 (.a(t0_001101010), .b(t0_001101011), .y(t0_00110101));
wire t0_001101010, t0_001101011;
mixer mix_t0_001101010 (.a(t0_0011010100), .b(t0_0011010101), .y(t0_001101010));
wire t0_0011010100, t0_0011010101;
mixer mix_t0_0011010100 (.a(t0_00110101000), .b(t0_00110101001), .y(t0_0011010100));
wire t0_00110101000, t0_00110101001;
mixer mix_t0_00110101000 (.a(t0_001101010000), .b(t0_001101010001), .y(t0_00110101000));
wire t0_001101010000, t0_001101010001;
mixer mix_t0_00110101001 (.a(t0_001101010010), .b(t0_001101010011), .y(t0_00110101001));
wire t0_001101010010, t0_001101010011;
mixer mix_t0_0011010101 (.a(t0_00110101010), .b(t0_00110101011), .y(t0_0011010101));
wire t0_00110101010, t0_00110101011;
mixer mix_t0_00110101010 (.a(t0_001101010100), .b(t0_001101010101), .y(t0_00110101010));
wire t0_001101010100, t0_001101010101;
mixer mix_t0_00110101011 (.a(t0_001101010110), .b(t0_001101010111), .y(t0_00110101011));
wire t0_001101010110, t0_001101010111;
mixer mix_t0_001101011 (.a(t0_0011010110), .b(t0_0011010111), .y(t0_001101011));
wire t0_0011010110, t0_0011010111;
mixer mix_t0_0011010110 (.a(t0_00110101100), .b(t0_00110101101), .y(t0_0011010110));
wire t0_00110101100, t0_00110101101;
mixer mix_t0_00110101100 (.a(t0_001101011000), .b(t0_001101011001), .y(t0_00110101100));
wire t0_001101011000, t0_001101011001;
mixer mix_t0_00110101101 (.a(t0_001101011010), .b(t0_001101011011), .y(t0_00110101101));
wire t0_001101011010, t0_001101011011;
mixer mix_t0_0011010111 (.a(t0_00110101110), .b(t0_00110101111), .y(t0_0011010111));
wire t0_00110101110, t0_00110101111;
mixer mix_t0_00110101110 (.a(t0_001101011100), .b(t0_001101011101), .y(t0_00110101110));
wire t0_001101011100, t0_001101011101;
mixer mix_t0_00110101111 (.a(t0_001101011110), .b(t0_001101011111), .y(t0_00110101111));
wire t0_001101011110, t0_001101011111;
mixer mix_t0_0011011 (.a(t0_00110110), .b(t0_00110111), .y(t0_0011011));
wire t0_00110110, t0_00110111;
mixer mix_t0_00110110 (.a(t0_001101100), .b(t0_001101101), .y(t0_00110110));
wire t0_001101100, t0_001101101;
mixer mix_t0_001101100 (.a(t0_0011011000), .b(t0_0011011001), .y(t0_001101100));
wire t0_0011011000, t0_0011011001;
mixer mix_t0_0011011000 (.a(t0_00110110000), .b(t0_00110110001), .y(t0_0011011000));
wire t0_00110110000, t0_00110110001;
mixer mix_t0_00110110000 (.a(t0_001101100000), .b(t0_001101100001), .y(t0_00110110000));
wire t0_001101100000, t0_001101100001;
mixer mix_t0_00110110001 (.a(t0_001101100010), .b(t0_001101100011), .y(t0_00110110001));
wire t0_001101100010, t0_001101100011;
mixer mix_t0_0011011001 (.a(t0_00110110010), .b(t0_00110110011), .y(t0_0011011001));
wire t0_00110110010, t0_00110110011;
mixer mix_t0_00110110010 (.a(t0_001101100100), .b(t0_001101100101), .y(t0_00110110010));
wire t0_001101100100, t0_001101100101;
mixer mix_t0_00110110011 (.a(t0_001101100110), .b(t0_001101100111), .y(t0_00110110011));
wire t0_001101100110, t0_001101100111;
mixer mix_t0_001101101 (.a(t0_0011011010), .b(t0_0011011011), .y(t0_001101101));
wire t0_0011011010, t0_0011011011;
mixer mix_t0_0011011010 (.a(t0_00110110100), .b(t0_00110110101), .y(t0_0011011010));
wire t0_00110110100, t0_00110110101;
mixer mix_t0_00110110100 (.a(t0_001101101000), .b(t0_001101101001), .y(t0_00110110100));
wire t0_001101101000, t0_001101101001;
mixer mix_t0_00110110101 (.a(t0_001101101010), .b(t0_001101101011), .y(t0_00110110101));
wire t0_001101101010, t0_001101101011;
mixer mix_t0_0011011011 (.a(t0_00110110110), .b(t0_00110110111), .y(t0_0011011011));
wire t0_00110110110, t0_00110110111;
mixer mix_t0_00110110110 (.a(t0_001101101100), .b(t0_001101101101), .y(t0_00110110110));
wire t0_001101101100, t0_001101101101;
mixer mix_t0_00110110111 (.a(t0_001101101110), .b(t0_001101101111), .y(t0_00110110111));
wire t0_001101101110, t0_001101101111;
mixer mix_t0_00110111 (.a(t0_001101110), .b(t0_001101111), .y(t0_00110111));
wire t0_001101110, t0_001101111;
mixer mix_t0_001101110 (.a(t0_0011011100), .b(t0_0011011101), .y(t0_001101110));
wire t0_0011011100, t0_0011011101;
mixer mix_t0_0011011100 (.a(t0_00110111000), .b(t0_00110111001), .y(t0_0011011100));
wire t0_00110111000, t0_00110111001;
mixer mix_t0_00110111000 (.a(t0_001101110000), .b(t0_001101110001), .y(t0_00110111000));
wire t0_001101110000, t0_001101110001;
mixer mix_t0_00110111001 (.a(t0_001101110010), .b(t0_001101110011), .y(t0_00110111001));
wire t0_001101110010, t0_001101110011;
mixer mix_t0_0011011101 (.a(t0_00110111010), .b(t0_00110111011), .y(t0_0011011101));
wire t0_00110111010, t0_00110111011;
mixer mix_t0_00110111010 (.a(t0_001101110100), .b(t0_001101110101), .y(t0_00110111010));
wire t0_001101110100, t0_001101110101;
mixer mix_t0_00110111011 (.a(t0_001101110110), .b(t0_001101110111), .y(t0_00110111011));
wire t0_001101110110, t0_001101110111;
mixer mix_t0_001101111 (.a(t0_0011011110), .b(t0_0011011111), .y(t0_001101111));
wire t0_0011011110, t0_0011011111;
mixer mix_t0_0011011110 (.a(t0_00110111100), .b(t0_00110111101), .y(t0_0011011110));
wire t0_00110111100, t0_00110111101;
mixer mix_t0_00110111100 (.a(t0_001101111000), .b(t0_001101111001), .y(t0_00110111100));
wire t0_001101111000, t0_001101111001;
mixer mix_t0_00110111101 (.a(t0_001101111010), .b(t0_001101111011), .y(t0_00110111101));
wire t0_001101111010, t0_001101111011;
mixer mix_t0_0011011111 (.a(t0_00110111110), .b(t0_00110111111), .y(t0_0011011111));
wire t0_00110111110, t0_00110111111;
mixer mix_t0_00110111110 (.a(t0_001101111100), .b(t0_001101111101), .y(t0_00110111110));
wire t0_001101111100, t0_001101111101;
mixer mix_t0_00110111111 (.a(t0_001101111110), .b(t0_001101111111), .y(t0_00110111111));
wire t0_001101111110, t0_001101111111;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_001110 (.a(t0_0011100), .b(t0_0011101), .y(t0_001110));
wire t0_0011100, t0_0011101;
mixer mix_t0_0011100 (.a(t0_00111000), .b(t0_00111001), .y(t0_0011100));
wire t0_00111000, t0_00111001;
mixer mix_t0_00111000 (.a(t0_001110000), .b(t0_001110001), .y(t0_00111000));
wire t0_001110000, t0_001110001;
mixer mix_t0_001110000 (.a(t0_0011100000), .b(t0_0011100001), .y(t0_001110000));
wire t0_0011100000, t0_0011100001;
mixer mix_t0_0011100000 (.a(t0_00111000000), .b(t0_00111000001), .y(t0_0011100000));
wire t0_00111000000, t0_00111000001;
mixer mix_t0_00111000000 (.a(t0_001110000000), .b(t0_001110000001), .y(t0_00111000000));
wire t0_001110000000, t0_001110000001;
mixer mix_t0_00111000001 (.a(t0_001110000010), .b(t0_001110000011), .y(t0_00111000001));
wire t0_001110000010, t0_001110000011;
mixer mix_t0_0011100001 (.a(t0_00111000010), .b(t0_00111000011), .y(t0_0011100001));
wire t0_00111000010, t0_00111000011;
mixer mix_t0_00111000010 (.a(t0_001110000100), .b(t0_001110000101), .y(t0_00111000010));
wire t0_001110000100, t0_001110000101;
mixer mix_t0_00111000011 (.a(t0_001110000110), .b(t0_001110000111), .y(t0_00111000011));
wire t0_001110000110, t0_001110000111;
mixer mix_t0_001110001 (.a(t0_0011100010), .b(t0_0011100011), .y(t0_001110001));
wire t0_0011100010, t0_0011100011;
mixer mix_t0_0011100010 (.a(t0_00111000100), .b(t0_00111000101), .y(t0_0011100010));
wire t0_00111000100, t0_00111000101;
mixer mix_t0_00111000100 (.a(t0_001110001000), .b(t0_001110001001), .y(t0_00111000100));
wire t0_001110001000, t0_001110001001;
mixer mix_t0_00111000101 (.a(t0_001110001010), .b(t0_001110001011), .y(t0_00111000101));
wire t0_001110001010, t0_001110001011;
mixer mix_t0_0011100011 (.a(t0_00111000110), .b(t0_00111000111), .y(t0_0011100011));
wire t0_00111000110, t0_00111000111;
mixer mix_t0_00111000110 (.a(t0_001110001100), .b(t0_001110001101), .y(t0_00111000110));
wire t0_001110001100, t0_001110001101;
mixer mix_t0_00111000111 (.a(t0_001110001110), .b(t0_001110001111), .y(t0_00111000111));
wire t0_001110001110, t0_001110001111;
mixer mix_t0_00111001 (.a(t0_001110010), .b(t0_001110011), .y(t0_00111001));
wire t0_001110010, t0_001110011;
mixer mix_t0_001110010 (.a(t0_0011100100), .b(t0_0011100101), .y(t0_001110010));
wire t0_0011100100, t0_0011100101;
mixer mix_t0_0011100100 (.a(t0_00111001000), .b(t0_00111001001), .y(t0_0011100100));
wire t0_00111001000, t0_00111001001;
mixer mix_t0_00111001000 (.a(t0_001110010000), .b(t0_001110010001), .y(t0_00111001000));
wire t0_001110010000, t0_001110010001;
mixer mix_t0_00111001001 (.a(t0_001110010010), .b(t0_001110010011), .y(t0_00111001001));
wire t0_001110010010, t0_001110010011;
mixer mix_t0_0011100101 (.a(t0_00111001010), .b(t0_00111001011), .y(t0_0011100101));
wire t0_00111001010, t0_00111001011;
mixer mix_t0_00111001010 (.a(t0_001110010100), .b(t0_001110010101), .y(t0_00111001010));
wire t0_001110010100, t0_001110010101;
mixer mix_t0_00111001011 (.a(t0_001110010110), .b(t0_001110010111), .y(t0_00111001011));
wire t0_001110010110, t0_001110010111;
mixer mix_t0_001110011 (.a(t0_0011100110), .b(t0_0011100111), .y(t0_001110011));
wire t0_0011100110, t0_0011100111;
mixer mix_t0_0011100110 (.a(t0_00111001100), .b(t0_00111001101), .y(t0_0011100110));
wire t0_00111001100, t0_00111001101;
mixer mix_t0_00111001100 (.a(t0_001110011000), .b(t0_001110011001), .y(t0_00111001100));
wire t0_001110011000, t0_001110011001;
mixer mix_t0_00111001101 (.a(t0_001110011010), .b(t0_001110011011), .y(t0_00111001101));
wire t0_001110011010, t0_001110011011;
mixer mix_t0_0011100111 (.a(t0_00111001110), .b(t0_00111001111), .y(t0_0011100111));
wire t0_00111001110, t0_00111001111;
mixer mix_t0_00111001110 (.a(t0_001110011100), .b(t0_001110011101), .y(t0_00111001110));
wire t0_001110011100, t0_001110011101;
mixer mix_t0_00111001111 (.a(t0_001110011110), .b(t0_001110011111), .y(t0_00111001111));
wire t0_001110011110, t0_001110011111;
mixer mix_t0_0011101 (.a(t0_00111010), .b(t0_00111011), .y(t0_0011101));
wire t0_00111010, t0_00111011;
mixer mix_t0_00111010 (.a(t0_001110100), .b(t0_001110101), .y(t0_00111010));
wire t0_001110100, t0_001110101;
mixer mix_t0_001110100 (.a(t0_0011101000), .b(t0_0011101001), .y(t0_001110100));
wire t0_0011101000, t0_0011101001;
mixer mix_t0_0011101000 (.a(t0_00111010000), .b(t0_00111010001), .y(t0_0011101000));
wire t0_00111010000, t0_00111010001;
mixer mix_t0_00111010000 (.a(t0_001110100000), .b(t0_001110100001), .y(t0_00111010000));
wire t0_001110100000, t0_001110100001;
mixer mix_t0_00111010001 (.a(t0_001110100010), .b(t0_001110100011), .y(t0_00111010001));
wire t0_001110100010, t0_001110100011;
mixer mix_t0_0011101001 (.a(t0_00111010010), .b(t0_00111010011), .y(t0_0011101001));
wire t0_00111010010, t0_00111010011;
mixer mix_t0_00111010010 (.a(t0_001110100100), .b(t0_001110100101), .y(t0_00111010010));
wire t0_001110100100, t0_001110100101;
mixer mix_t0_00111010011 (.a(t0_001110100110), .b(t0_001110100111), .y(t0_00111010011));
wire t0_001110100110, t0_001110100111;
mixer mix_t0_001110101 (.a(t0_0011101010), .b(t0_0011101011), .y(t0_001110101));
wire t0_0011101010, t0_0011101011;
mixer mix_t0_0011101010 (.a(t0_00111010100), .b(t0_00111010101), .y(t0_0011101010));
wire t0_00111010100, t0_00111010101;
mixer mix_t0_00111010100 (.a(t0_001110101000), .b(t0_001110101001), .y(t0_00111010100));
wire t0_001110101000, t0_001110101001;
mixer mix_t0_00111010101 (.a(t0_001110101010), .b(t0_001110101011), .y(t0_00111010101));
wire t0_001110101010, t0_001110101011;
mixer mix_t0_0011101011 (.a(t0_00111010110), .b(t0_00111010111), .y(t0_0011101011));
wire t0_00111010110, t0_00111010111;
mixer mix_t0_00111010110 (.a(t0_001110101100), .b(t0_001110101101), .y(t0_00111010110));
wire t0_001110101100, t0_001110101101;
mixer mix_t0_00111010111 (.a(t0_001110101110), .b(t0_001110101111), .y(t0_00111010111));
wire t0_001110101110, t0_001110101111;
mixer mix_t0_00111011 (.a(t0_001110110), .b(t0_001110111), .y(t0_00111011));
wire t0_001110110, t0_001110111;
mixer mix_t0_001110110 (.a(t0_0011101100), .b(t0_0011101101), .y(t0_001110110));
wire t0_0011101100, t0_0011101101;
mixer mix_t0_0011101100 (.a(t0_00111011000), .b(t0_00111011001), .y(t0_0011101100));
wire t0_00111011000, t0_00111011001;
mixer mix_t0_00111011000 (.a(t0_001110110000), .b(t0_001110110001), .y(t0_00111011000));
wire t0_001110110000, t0_001110110001;
mixer mix_t0_00111011001 (.a(t0_001110110010), .b(t0_001110110011), .y(t0_00111011001));
wire t0_001110110010, t0_001110110011;
mixer mix_t0_0011101101 (.a(t0_00111011010), .b(t0_00111011011), .y(t0_0011101101));
wire t0_00111011010, t0_00111011011;
mixer mix_t0_00111011010 (.a(t0_001110110100), .b(t0_001110110101), .y(t0_00111011010));
wire t0_001110110100, t0_001110110101;
mixer mix_t0_00111011011 (.a(t0_001110110110), .b(t0_001110110111), .y(t0_00111011011));
wire t0_001110110110, t0_001110110111;
mixer mix_t0_001110111 (.a(t0_0011101110), .b(t0_0011101111), .y(t0_001110111));
wire t0_0011101110, t0_0011101111;
mixer mix_t0_0011101110 (.a(t0_00111011100), .b(t0_00111011101), .y(t0_0011101110));
wire t0_00111011100, t0_00111011101;
mixer mix_t0_00111011100 (.a(t0_001110111000), .b(t0_001110111001), .y(t0_00111011100));
wire t0_001110111000, t0_001110111001;
mixer mix_t0_00111011101 (.a(t0_001110111010), .b(t0_001110111011), .y(t0_00111011101));
wire t0_001110111010, t0_001110111011;
mixer mix_t0_0011101111 (.a(t0_00111011110), .b(t0_00111011111), .y(t0_0011101111));
wire t0_00111011110, t0_00111011111;
mixer mix_t0_00111011110 (.a(t0_001110111100), .b(t0_001110111101), .y(t0_00111011110));
wire t0_001110111100, t0_001110111101;
mixer mix_t0_00111011111 (.a(t0_001110111110), .b(t0_001110111111), .y(t0_00111011111));
wire t0_001110111110, t0_001110111111;
mixer mix_t0_001111 (.a(t0_0011110), .b(t0_0011111), .y(t0_001111));
wire t0_0011110, t0_0011111;
mixer mix_t0_0011110 (.a(t0_00111100), .b(t0_00111101), .y(t0_0011110));
wire t0_00111100, t0_00111101;
mixer mix_t0_00111100 (.a(t0_001111000), .b(t0_001111001), .y(t0_00111100));
wire t0_001111000, t0_001111001;
mixer mix_t0_001111000 (.a(t0_0011110000), .b(t0_0011110001), .y(t0_001111000));
wire t0_0011110000, t0_0011110001;
mixer mix_t0_0011110000 (.a(t0_00111100000), .b(t0_00111100001), .y(t0_0011110000));
wire t0_00111100000, t0_00111100001;
mixer mix_t0_00111100000 (.a(t0_001111000000), .b(t0_001111000001), .y(t0_00111100000));
wire t0_001111000000, t0_001111000001;
mixer mix_t0_00111100001 (.a(t0_001111000010), .b(t0_001111000011), .y(t0_00111100001));
wire t0_001111000010, t0_001111000011;
mixer mix_t0_0011110001 (.a(t0_00111100010), .b(t0_00111100011), .y(t0_0011110001));
wire t0_00111100010, t0_00111100011;
mixer mix_t0_00111100010 (.a(t0_001111000100), .b(t0_001111000101), .y(t0_00111100010));
wire t0_001111000100, t0_001111000101;
mixer mix_t0_00111100011 (.a(t0_001111000110), .b(t0_001111000111), .y(t0_00111100011));
wire t0_001111000110, t0_001111000111;
mixer mix_t0_001111001 (.a(t0_0011110010), .b(t0_0011110011), .y(t0_001111001));
wire t0_0011110010, t0_0011110011;
mixer mix_t0_0011110010 (.a(t0_00111100100), .b(t0_00111100101), .y(t0_0011110010));
wire t0_00111100100, t0_00111100101;
mixer mix_t0_00111100100 (.a(t0_001111001000), .b(t0_001111001001), .y(t0_00111100100));
wire t0_001111001000, t0_001111001001;
mixer mix_t0_00111100101 (.a(t0_001111001010), .b(t0_001111001011), .y(t0_00111100101));
wire t0_001111001010, t0_001111001011;
mixer mix_t0_0011110011 (.a(t0_00111100110), .b(t0_00111100111), .y(t0_0011110011));
wire t0_00111100110, t0_00111100111;
mixer mix_t0_00111100110 (.a(t0_001111001100), .b(t0_001111001101), .y(t0_00111100110));
wire t0_001111001100, t0_001111001101;
mixer mix_t0_00111100111 (.a(t0_001111001110), .b(t0_001111001111), .y(t0_00111100111));
wire t0_001111001110, t0_001111001111;
mixer mix_t0_00111101 (.a(t0_001111010), .b(t0_001111011), .y(t0_00111101));
wire t0_001111010, t0_001111011;
mixer mix_t0_001111010 (.a(t0_0011110100), .b(t0_0011110101), .y(t0_001111010));
wire t0_0011110100, t0_0011110101;
mixer mix_t0_0011110100 (.a(t0_00111101000), .b(t0_00111101001), .y(t0_0011110100));
wire t0_00111101000, t0_00111101001;
mixer mix_t0_00111101000 (.a(t0_001111010000), .b(t0_001111010001), .y(t0_00111101000));
wire t0_001111010000, t0_001111010001;
mixer mix_t0_00111101001 (.a(t0_001111010010), .b(t0_001111010011), .y(t0_00111101001));
wire t0_001111010010, t0_001111010011;
mixer mix_t0_0011110101 (.a(t0_00111101010), .b(t0_00111101011), .y(t0_0011110101));
wire t0_00111101010, t0_00111101011;
mixer mix_t0_00111101010 (.a(t0_001111010100), .b(t0_001111010101), .y(t0_00111101010));
wire t0_001111010100, t0_001111010101;
mixer mix_t0_00111101011 (.a(t0_001111010110), .b(t0_001111010111), .y(t0_00111101011));
wire t0_001111010110, t0_001111010111;
mixer mix_t0_001111011 (.a(t0_0011110110), .b(t0_0011110111), .y(t0_001111011));
wire t0_0011110110, t0_0011110111;
mixer mix_t0_0011110110 (.a(t0_00111101100), .b(t0_00111101101), .y(t0_0011110110));
wire t0_00111101100, t0_00111101101;
mixer mix_t0_00111101100 (.a(t0_001111011000), .b(t0_001111011001), .y(t0_00111101100));
wire t0_001111011000, t0_001111011001;
mixer mix_t0_00111101101 (.a(t0_001111011010), .b(t0_001111011011), .y(t0_00111101101));
wire t0_001111011010, t0_001111011011;
mixer mix_t0_0011110111 (.a(t0_00111101110), .b(t0_00111101111), .y(t0_0011110111));
wire t0_00111101110, t0_00111101111;
mixer mix_t0_00111101110 (.a(t0_001111011100), .b(t0_001111011101), .y(t0_00111101110));
wire t0_001111011100, t0_001111011101;
mixer mix_t0_00111101111 (.a(t0_001111011110), .b(t0_001111011111), .y(t0_00111101111));
wire t0_001111011110, t0_001111011111;
mixer mix_t0_0011111 (.a(t0_00111110), .b(t0_00111111), .y(t0_0011111));
wire t0_00111110, t0_00111111;
mixer mix_t0_00111110 (.a(t0_001111100), .b(t0_001111101), .y(t0_00111110));
wire t0_001111100, t0_001111101;
mixer mix_t0_001111100 (.a(t0_0011111000), .b(t0_0011111001), .y(t0_001111100));
wire t0_0011111000, t0_0011111001;
mixer mix_t0_0011111000 (.a(t0_00111110000), .b(t0_00111110001), .y(t0_0011111000));
wire t0_00111110000, t0_00111110001;
mixer mix_t0_00111110000 (.a(t0_001111100000), .b(t0_001111100001), .y(t0_00111110000));
wire t0_001111100000, t0_001111100001;
mixer mix_t0_00111110001 (.a(t0_001111100010), .b(t0_001111100011), .y(t0_00111110001));
wire t0_001111100010, t0_001111100011;
mixer mix_t0_0011111001 (.a(t0_00111110010), .b(t0_00111110011), .y(t0_0011111001));
wire t0_00111110010, t0_00111110011;
mixer mix_t0_00111110010 (.a(t0_001111100100), .b(t0_001111100101), .y(t0_00111110010));
wire t0_001111100100, t0_001111100101;
mixer mix_t0_00111110011 (.a(t0_001111100110), .b(t0_001111100111), .y(t0_00111110011));
wire t0_001111100110, t0_001111100111;
mixer mix_t0_001111101 (.a(t0_0011111010), .b(t0_0011111011), .y(t0_001111101));
wire t0_0011111010, t0_0011111011;
mixer mix_t0_0011111010 (.a(t0_00111110100), .b(t0_00111110101), .y(t0_0011111010));
wire t0_00111110100, t0_00111110101;
mixer mix_t0_00111110100 (.a(t0_001111101000), .b(t0_001111101001), .y(t0_00111110100));
wire t0_001111101000, t0_001111101001;
mixer mix_t0_00111110101 (.a(t0_001111101010), .b(t0_001111101011), .y(t0_00111110101));
wire t0_001111101010, t0_001111101011;
mixer mix_t0_0011111011 (.a(t0_00111110110), .b(t0_00111110111), .y(t0_0011111011));
wire t0_00111110110, t0_00111110111;
mixer mix_t0_00111110110 (.a(t0_001111101100), .b(t0_001111101101), .y(t0_00111110110));
wire t0_001111101100, t0_001111101101;
mixer mix_t0_00111110111 (.a(t0_001111101110), .b(t0_001111101111), .y(t0_00111110111));
wire t0_001111101110, t0_001111101111;
mixer mix_t0_00111111 (.a(t0_001111110), .b(t0_001111111), .y(t0_00111111));
wire t0_001111110, t0_001111111;
mixer mix_t0_001111110 (.a(t0_0011111100), .b(t0_0011111101), .y(t0_001111110));
wire t0_0011111100, t0_0011111101;
mixer mix_t0_0011111100 (.a(t0_00111111000), .b(t0_00111111001), .y(t0_0011111100));
wire t0_00111111000, t0_00111111001;
mixer mix_t0_00111111000 (.a(t0_001111110000), .b(t0_001111110001), .y(t0_00111111000));
wire t0_001111110000, t0_001111110001;
mixer mix_t0_00111111001 (.a(t0_001111110010), .b(t0_001111110011), .y(t0_00111111001));
wire t0_001111110010, t0_001111110011;
mixer mix_t0_0011111101 (.a(t0_00111111010), .b(t0_00111111011), .y(t0_0011111101));
wire t0_00111111010, t0_00111111011;
mixer mix_t0_00111111010 (.a(t0_001111110100), .b(t0_001111110101), .y(t0_00111111010));
wire t0_001111110100, t0_001111110101;
mixer mix_t0_00111111011 (.a(t0_001111110110), .b(t0_001111110111), .y(t0_00111111011));
wire t0_001111110110, t0_001111110111;
mixer mix_t0_001111111 (.a(t0_0011111110), .b(t0_0011111111), .y(t0_001111111));
wire t0_0011111110, t0_0011111111;
mixer mix_t0_0011111110 (.a(t0_00111111100), .b(t0_00111111101), .y(t0_0011111110));
wire t0_00111111100, t0_00111111101;
mixer mix_t0_00111111100 (.a(t0_001111111000), .b(t0_001111111001), .y(t0_00111111100));
wire t0_001111111000, t0_001111111001;
mixer mix_t0_00111111101 (.a(t0_001111111010), .b(t0_001111111011), .y(t0_00111111101));
wire t0_001111111010, t0_001111111011;
mixer mix_t0_0011111111 (.a(t0_00111111110), .b(t0_00111111111), .y(t0_0011111111));
wire t0_00111111110, t0_00111111111;
mixer mix_t0_00111111110 (.a(t0_001111111100), .b(t0_001111111101), .y(t0_00111111110));
wire t0_001111111100, t0_001111111101;
mixer mix_t0_00111111111 (.a(t0_001111111110), .b(t0_001111111111), .y(t0_00111111111));
wire t0_001111111110, t0_001111111111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_010000 (.a(t0_0100000), .b(t0_0100001), .y(t0_010000));
wire t0_0100000, t0_0100001;
mixer mix_t0_0100000 (.a(t0_01000000), .b(t0_01000001), .y(t0_0100000));
wire t0_01000000, t0_01000001;
mixer mix_t0_01000000 (.a(t0_010000000), .b(t0_010000001), .y(t0_01000000));
wire t0_010000000, t0_010000001;
mixer mix_t0_010000000 (.a(t0_0100000000), .b(t0_0100000001), .y(t0_010000000));
wire t0_0100000000, t0_0100000001;
mixer mix_t0_0100000000 (.a(t0_01000000000), .b(t0_01000000001), .y(t0_0100000000));
wire t0_01000000000, t0_01000000001;
mixer mix_t0_01000000000 (.a(t0_010000000000), .b(t0_010000000001), .y(t0_01000000000));
wire t0_010000000000, t0_010000000001;
mixer mix_t0_01000000001 (.a(t0_010000000010), .b(t0_010000000011), .y(t0_01000000001));
wire t0_010000000010, t0_010000000011;
mixer mix_t0_0100000001 (.a(t0_01000000010), .b(t0_01000000011), .y(t0_0100000001));
wire t0_01000000010, t0_01000000011;
mixer mix_t0_01000000010 (.a(t0_010000000100), .b(t0_010000000101), .y(t0_01000000010));
wire t0_010000000100, t0_010000000101;
mixer mix_t0_01000000011 (.a(t0_010000000110), .b(t0_010000000111), .y(t0_01000000011));
wire t0_010000000110, t0_010000000111;
mixer mix_t0_010000001 (.a(t0_0100000010), .b(t0_0100000011), .y(t0_010000001));
wire t0_0100000010, t0_0100000011;
mixer mix_t0_0100000010 (.a(t0_01000000100), .b(t0_01000000101), .y(t0_0100000010));
wire t0_01000000100, t0_01000000101;
mixer mix_t0_01000000100 (.a(t0_010000001000), .b(t0_010000001001), .y(t0_01000000100));
wire t0_010000001000, t0_010000001001;
mixer mix_t0_01000000101 (.a(t0_010000001010), .b(t0_010000001011), .y(t0_01000000101));
wire t0_010000001010, t0_010000001011;
mixer mix_t0_0100000011 (.a(t0_01000000110), .b(t0_01000000111), .y(t0_0100000011));
wire t0_01000000110, t0_01000000111;
mixer mix_t0_01000000110 (.a(t0_010000001100), .b(t0_010000001101), .y(t0_01000000110));
wire t0_010000001100, t0_010000001101;
mixer mix_t0_01000000111 (.a(t0_010000001110), .b(t0_010000001111), .y(t0_01000000111));
wire t0_010000001110, t0_010000001111;
mixer mix_t0_01000001 (.a(t0_010000010), .b(t0_010000011), .y(t0_01000001));
wire t0_010000010, t0_010000011;
mixer mix_t0_010000010 (.a(t0_0100000100), .b(t0_0100000101), .y(t0_010000010));
wire t0_0100000100, t0_0100000101;
mixer mix_t0_0100000100 (.a(t0_01000001000), .b(t0_01000001001), .y(t0_0100000100));
wire t0_01000001000, t0_01000001001;
mixer mix_t0_01000001000 (.a(t0_010000010000), .b(t0_010000010001), .y(t0_01000001000));
wire t0_010000010000, t0_010000010001;
mixer mix_t0_01000001001 (.a(t0_010000010010), .b(t0_010000010011), .y(t0_01000001001));
wire t0_010000010010, t0_010000010011;
mixer mix_t0_0100000101 (.a(t0_01000001010), .b(t0_01000001011), .y(t0_0100000101));
wire t0_01000001010, t0_01000001011;
mixer mix_t0_01000001010 (.a(t0_010000010100), .b(t0_010000010101), .y(t0_01000001010));
wire t0_010000010100, t0_010000010101;
mixer mix_t0_01000001011 (.a(t0_010000010110), .b(t0_010000010111), .y(t0_01000001011));
wire t0_010000010110, t0_010000010111;
mixer mix_t0_010000011 (.a(t0_0100000110), .b(t0_0100000111), .y(t0_010000011));
wire t0_0100000110, t0_0100000111;
mixer mix_t0_0100000110 (.a(t0_01000001100), .b(t0_01000001101), .y(t0_0100000110));
wire t0_01000001100, t0_01000001101;
mixer mix_t0_01000001100 (.a(t0_010000011000), .b(t0_010000011001), .y(t0_01000001100));
wire t0_010000011000, t0_010000011001;
mixer mix_t0_01000001101 (.a(t0_010000011010), .b(t0_010000011011), .y(t0_01000001101));
wire t0_010000011010, t0_010000011011;
mixer mix_t0_0100000111 (.a(t0_01000001110), .b(t0_01000001111), .y(t0_0100000111));
wire t0_01000001110, t0_01000001111;
mixer mix_t0_01000001110 (.a(t0_010000011100), .b(t0_010000011101), .y(t0_01000001110));
wire t0_010000011100, t0_010000011101;
mixer mix_t0_01000001111 (.a(t0_010000011110), .b(t0_010000011111), .y(t0_01000001111));
wire t0_010000011110, t0_010000011111;
mixer mix_t0_0100001 (.a(t0_01000010), .b(t0_01000011), .y(t0_0100001));
wire t0_01000010, t0_01000011;
mixer mix_t0_01000010 (.a(t0_010000100), .b(t0_010000101), .y(t0_01000010));
wire t0_010000100, t0_010000101;
mixer mix_t0_010000100 (.a(t0_0100001000), .b(t0_0100001001), .y(t0_010000100));
wire t0_0100001000, t0_0100001001;
mixer mix_t0_0100001000 (.a(t0_01000010000), .b(t0_01000010001), .y(t0_0100001000));
wire t0_01000010000, t0_01000010001;
mixer mix_t0_01000010000 (.a(t0_010000100000), .b(t0_010000100001), .y(t0_01000010000));
wire t0_010000100000, t0_010000100001;
mixer mix_t0_01000010001 (.a(t0_010000100010), .b(t0_010000100011), .y(t0_01000010001));
wire t0_010000100010, t0_010000100011;
mixer mix_t0_0100001001 (.a(t0_01000010010), .b(t0_01000010011), .y(t0_0100001001));
wire t0_01000010010, t0_01000010011;
mixer mix_t0_01000010010 (.a(t0_010000100100), .b(t0_010000100101), .y(t0_01000010010));
wire t0_010000100100, t0_010000100101;
mixer mix_t0_01000010011 (.a(t0_010000100110), .b(t0_010000100111), .y(t0_01000010011));
wire t0_010000100110, t0_010000100111;
mixer mix_t0_010000101 (.a(t0_0100001010), .b(t0_0100001011), .y(t0_010000101));
wire t0_0100001010, t0_0100001011;
mixer mix_t0_0100001010 (.a(t0_01000010100), .b(t0_01000010101), .y(t0_0100001010));
wire t0_01000010100, t0_01000010101;
mixer mix_t0_01000010100 (.a(t0_010000101000), .b(t0_010000101001), .y(t0_01000010100));
wire t0_010000101000, t0_010000101001;
mixer mix_t0_01000010101 (.a(t0_010000101010), .b(t0_010000101011), .y(t0_01000010101));
wire t0_010000101010, t0_010000101011;
mixer mix_t0_0100001011 (.a(t0_01000010110), .b(t0_01000010111), .y(t0_0100001011));
wire t0_01000010110, t0_01000010111;
mixer mix_t0_01000010110 (.a(t0_010000101100), .b(t0_010000101101), .y(t0_01000010110));
wire t0_010000101100, t0_010000101101;
mixer mix_t0_01000010111 (.a(t0_010000101110), .b(t0_010000101111), .y(t0_01000010111));
wire t0_010000101110, t0_010000101111;
mixer mix_t0_01000011 (.a(t0_010000110), .b(t0_010000111), .y(t0_01000011));
wire t0_010000110, t0_010000111;
mixer mix_t0_010000110 (.a(t0_0100001100), .b(t0_0100001101), .y(t0_010000110));
wire t0_0100001100, t0_0100001101;
mixer mix_t0_0100001100 (.a(t0_01000011000), .b(t0_01000011001), .y(t0_0100001100));
wire t0_01000011000, t0_01000011001;
mixer mix_t0_01000011000 (.a(t0_010000110000), .b(t0_010000110001), .y(t0_01000011000));
wire t0_010000110000, t0_010000110001;
mixer mix_t0_01000011001 (.a(t0_010000110010), .b(t0_010000110011), .y(t0_01000011001));
wire t0_010000110010, t0_010000110011;
mixer mix_t0_0100001101 (.a(t0_01000011010), .b(t0_01000011011), .y(t0_0100001101));
wire t0_01000011010, t0_01000011011;
mixer mix_t0_01000011010 (.a(t0_010000110100), .b(t0_010000110101), .y(t0_01000011010));
wire t0_010000110100, t0_010000110101;
mixer mix_t0_01000011011 (.a(t0_010000110110), .b(t0_010000110111), .y(t0_01000011011));
wire t0_010000110110, t0_010000110111;
mixer mix_t0_010000111 (.a(t0_0100001110), .b(t0_0100001111), .y(t0_010000111));
wire t0_0100001110, t0_0100001111;
mixer mix_t0_0100001110 (.a(t0_01000011100), .b(t0_01000011101), .y(t0_0100001110));
wire t0_01000011100, t0_01000011101;
mixer mix_t0_01000011100 (.a(t0_010000111000), .b(t0_010000111001), .y(t0_01000011100));
wire t0_010000111000, t0_010000111001;
mixer mix_t0_01000011101 (.a(t0_010000111010), .b(t0_010000111011), .y(t0_01000011101));
wire t0_010000111010, t0_010000111011;
mixer mix_t0_0100001111 (.a(t0_01000011110), .b(t0_01000011111), .y(t0_0100001111));
wire t0_01000011110, t0_01000011111;
mixer mix_t0_01000011110 (.a(t0_010000111100), .b(t0_010000111101), .y(t0_01000011110));
wire t0_010000111100, t0_010000111101;
mixer mix_t0_01000011111 (.a(t0_010000111110), .b(t0_010000111111), .y(t0_01000011111));
wire t0_010000111110, t0_010000111111;
mixer mix_t0_010001 (.a(t0_0100010), .b(t0_0100011), .y(t0_010001));
wire t0_0100010, t0_0100011;
mixer mix_t0_0100010 (.a(t0_01000100), .b(t0_01000101), .y(t0_0100010));
wire t0_01000100, t0_01000101;
mixer mix_t0_01000100 (.a(t0_010001000), .b(t0_010001001), .y(t0_01000100));
wire t0_010001000, t0_010001001;
mixer mix_t0_010001000 (.a(t0_0100010000), .b(t0_0100010001), .y(t0_010001000));
wire t0_0100010000, t0_0100010001;
mixer mix_t0_0100010000 (.a(t0_01000100000), .b(t0_01000100001), .y(t0_0100010000));
wire t0_01000100000, t0_01000100001;
mixer mix_t0_01000100000 (.a(t0_010001000000), .b(t0_010001000001), .y(t0_01000100000));
wire t0_010001000000, t0_010001000001;
mixer mix_t0_01000100001 (.a(t0_010001000010), .b(t0_010001000011), .y(t0_01000100001));
wire t0_010001000010, t0_010001000011;
mixer mix_t0_0100010001 (.a(t0_01000100010), .b(t0_01000100011), .y(t0_0100010001));
wire t0_01000100010, t0_01000100011;
mixer mix_t0_01000100010 (.a(t0_010001000100), .b(t0_010001000101), .y(t0_01000100010));
wire t0_010001000100, t0_010001000101;
mixer mix_t0_01000100011 (.a(t0_010001000110), .b(t0_010001000111), .y(t0_01000100011));
wire t0_010001000110, t0_010001000111;
mixer mix_t0_010001001 (.a(t0_0100010010), .b(t0_0100010011), .y(t0_010001001));
wire t0_0100010010, t0_0100010011;
mixer mix_t0_0100010010 (.a(t0_01000100100), .b(t0_01000100101), .y(t0_0100010010));
wire t0_01000100100, t0_01000100101;
mixer mix_t0_01000100100 (.a(t0_010001001000), .b(t0_010001001001), .y(t0_01000100100));
wire t0_010001001000, t0_010001001001;
mixer mix_t0_01000100101 (.a(t0_010001001010), .b(t0_010001001011), .y(t0_01000100101));
wire t0_010001001010, t0_010001001011;
mixer mix_t0_0100010011 (.a(t0_01000100110), .b(t0_01000100111), .y(t0_0100010011));
wire t0_01000100110, t0_01000100111;
mixer mix_t0_01000100110 (.a(t0_010001001100), .b(t0_010001001101), .y(t0_01000100110));
wire t0_010001001100, t0_010001001101;
mixer mix_t0_01000100111 (.a(t0_010001001110), .b(t0_010001001111), .y(t0_01000100111));
wire t0_010001001110, t0_010001001111;
mixer mix_t0_01000101 (.a(t0_010001010), .b(t0_010001011), .y(t0_01000101));
wire t0_010001010, t0_010001011;
mixer mix_t0_010001010 (.a(t0_0100010100), .b(t0_0100010101), .y(t0_010001010));
wire t0_0100010100, t0_0100010101;
mixer mix_t0_0100010100 (.a(t0_01000101000), .b(t0_01000101001), .y(t0_0100010100));
wire t0_01000101000, t0_01000101001;
mixer mix_t0_01000101000 (.a(t0_010001010000), .b(t0_010001010001), .y(t0_01000101000));
wire t0_010001010000, t0_010001010001;
mixer mix_t0_01000101001 (.a(t0_010001010010), .b(t0_010001010011), .y(t0_01000101001));
wire t0_010001010010, t0_010001010011;
mixer mix_t0_0100010101 (.a(t0_01000101010), .b(t0_01000101011), .y(t0_0100010101));
wire t0_01000101010, t0_01000101011;
mixer mix_t0_01000101010 (.a(t0_010001010100), .b(t0_010001010101), .y(t0_01000101010));
wire t0_010001010100, t0_010001010101;
mixer mix_t0_01000101011 (.a(t0_010001010110), .b(t0_010001010111), .y(t0_01000101011));
wire t0_010001010110, t0_010001010111;
mixer mix_t0_010001011 (.a(t0_0100010110), .b(t0_0100010111), .y(t0_010001011));
wire t0_0100010110, t0_0100010111;
mixer mix_t0_0100010110 (.a(t0_01000101100), .b(t0_01000101101), .y(t0_0100010110));
wire t0_01000101100, t0_01000101101;
mixer mix_t0_01000101100 (.a(t0_010001011000), .b(t0_010001011001), .y(t0_01000101100));
wire t0_010001011000, t0_010001011001;
mixer mix_t0_01000101101 (.a(t0_010001011010), .b(t0_010001011011), .y(t0_01000101101));
wire t0_010001011010, t0_010001011011;
mixer mix_t0_0100010111 (.a(t0_01000101110), .b(t0_01000101111), .y(t0_0100010111));
wire t0_01000101110, t0_01000101111;
mixer mix_t0_01000101110 (.a(t0_010001011100), .b(t0_010001011101), .y(t0_01000101110));
wire t0_010001011100, t0_010001011101;
mixer mix_t0_01000101111 (.a(t0_010001011110), .b(t0_010001011111), .y(t0_01000101111));
wire t0_010001011110, t0_010001011111;
mixer mix_t0_0100011 (.a(t0_01000110), .b(t0_01000111), .y(t0_0100011));
wire t0_01000110, t0_01000111;
mixer mix_t0_01000110 (.a(t0_010001100), .b(t0_010001101), .y(t0_01000110));
wire t0_010001100, t0_010001101;
mixer mix_t0_010001100 (.a(t0_0100011000), .b(t0_0100011001), .y(t0_010001100));
wire t0_0100011000, t0_0100011001;
mixer mix_t0_0100011000 (.a(t0_01000110000), .b(t0_01000110001), .y(t0_0100011000));
wire t0_01000110000, t0_01000110001;
mixer mix_t0_01000110000 (.a(t0_010001100000), .b(t0_010001100001), .y(t0_01000110000));
wire t0_010001100000, t0_010001100001;
mixer mix_t0_01000110001 (.a(t0_010001100010), .b(t0_010001100011), .y(t0_01000110001));
wire t0_010001100010, t0_010001100011;
mixer mix_t0_0100011001 (.a(t0_01000110010), .b(t0_01000110011), .y(t0_0100011001));
wire t0_01000110010, t0_01000110011;
mixer mix_t0_01000110010 (.a(t0_010001100100), .b(t0_010001100101), .y(t0_01000110010));
wire t0_010001100100, t0_010001100101;
mixer mix_t0_01000110011 (.a(t0_010001100110), .b(t0_010001100111), .y(t0_01000110011));
wire t0_010001100110, t0_010001100111;
mixer mix_t0_010001101 (.a(t0_0100011010), .b(t0_0100011011), .y(t0_010001101));
wire t0_0100011010, t0_0100011011;
mixer mix_t0_0100011010 (.a(t0_01000110100), .b(t0_01000110101), .y(t0_0100011010));
wire t0_01000110100, t0_01000110101;
mixer mix_t0_01000110100 (.a(t0_010001101000), .b(t0_010001101001), .y(t0_01000110100));
wire t0_010001101000, t0_010001101001;
mixer mix_t0_01000110101 (.a(t0_010001101010), .b(t0_010001101011), .y(t0_01000110101));
wire t0_010001101010, t0_010001101011;
mixer mix_t0_0100011011 (.a(t0_01000110110), .b(t0_01000110111), .y(t0_0100011011));
wire t0_01000110110, t0_01000110111;
mixer mix_t0_01000110110 (.a(t0_010001101100), .b(t0_010001101101), .y(t0_01000110110));
wire t0_010001101100, t0_010001101101;
mixer mix_t0_01000110111 (.a(t0_010001101110), .b(t0_010001101111), .y(t0_01000110111));
wire t0_010001101110, t0_010001101111;
mixer mix_t0_01000111 (.a(t0_010001110), .b(t0_010001111), .y(t0_01000111));
wire t0_010001110, t0_010001111;
mixer mix_t0_010001110 (.a(t0_0100011100), .b(t0_0100011101), .y(t0_010001110));
wire t0_0100011100, t0_0100011101;
mixer mix_t0_0100011100 (.a(t0_01000111000), .b(t0_01000111001), .y(t0_0100011100));
wire t0_01000111000, t0_01000111001;
mixer mix_t0_01000111000 (.a(t0_010001110000), .b(t0_010001110001), .y(t0_01000111000));
wire t0_010001110000, t0_010001110001;
mixer mix_t0_01000111001 (.a(t0_010001110010), .b(t0_010001110011), .y(t0_01000111001));
wire t0_010001110010, t0_010001110011;
mixer mix_t0_0100011101 (.a(t0_01000111010), .b(t0_01000111011), .y(t0_0100011101));
wire t0_01000111010, t0_01000111011;
mixer mix_t0_01000111010 (.a(t0_010001110100), .b(t0_010001110101), .y(t0_01000111010));
wire t0_010001110100, t0_010001110101;
mixer mix_t0_01000111011 (.a(t0_010001110110), .b(t0_010001110111), .y(t0_01000111011));
wire t0_010001110110, t0_010001110111;
mixer mix_t0_010001111 (.a(t0_0100011110), .b(t0_0100011111), .y(t0_010001111));
wire t0_0100011110, t0_0100011111;
mixer mix_t0_0100011110 (.a(t0_01000111100), .b(t0_01000111101), .y(t0_0100011110));
wire t0_01000111100, t0_01000111101;
mixer mix_t0_01000111100 (.a(t0_010001111000), .b(t0_010001111001), .y(t0_01000111100));
wire t0_010001111000, t0_010001111001;
mixer mix_t0_01000111101 (.a(t0_010001111010), .b(t0_010001111011), .y(t0_01000111101));
wire t0_010001111010, t0_010001111011;
mixer mix_t0_0100011111 (.a(t0_01000111110), .b(t0_01000111111), .y(t0_0100011111));
wire t0_01000111110, t0_01000111111;
mixer mix_t0_01000111110 (.a(t0_010001111100), .b(t0_010001111101), .y(t0_01000111110));
wire t0_010001111100, t0_010001111101;
mixer mix_t0_01000111111 (.a(t0_010001111110), .b(t0_010001111111), .y(t0_01000111111));
wire t0_010001111110, t0_010001111111;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_010010 (.a(t0_0100100), .b(t0_0100101), .y(t0_010010));
wire t0_0100100, t0_0100101;
mixer mix_t0_0100100 (.a(t0_01001000), .b(t0_01001001), .y(t0_0100100));
wire t0_01001000, t0_01001001;
mixer mix_t0_01001000 (.a(t0_010010000), .b(t0_010010001), .y(t0_01001000));
wire t0_010010000, t0_010010001;
mixer mix_t0_010010000 (.a(t0_0100100000), .b(t0_0100100001), .y(t0_010010000));
wire t0_0100100000, t0_0100100001;
mixer mix_t0_0100100000 (.a(t0_01001000000), .b(t0_01001000001), .y(t0_0100100000));
wire t0_01001000000, t0_01001000001;
mixer mix_t0_01001000000 (.a(t0_010010000000), .b(t0_010010000001), .y(t0_01001000000));
wire t0_010010000000, t0_010010000001;
mixer mix_t0_01001000001 (.a(t0_010010000010), .b(t0_010010000011), .y(t0_01001000001));
wire t0_010010000010, t0_010010000011;
mixer mix_t0_0100100001 (.a(t0_01001000010), .b(t0_01001000011), .y(t0_0100100001));
wire t0_01001000010, t0_01001000011;
mixer mix_t0_01001000010 (.a(t0_010010000100), .b(t0_010010000101), .y(t0_01001000010));
wire t0_010010000100, t0_010010000101;
mixer mix_t0_01001000011 (.a(t0_010010000110), .b(t0_010010000111), .y(t0_01001000011));
wire t0_010010000110, t0_010010000111;
mixer mix_t0_010010001 (.a(t0_0100100010), .b(t0_0100100011), .y(t0_010010001));
wire t0_0100100010, t0_0100100011;
mixer mix_t0_0100100010 (.a(t0_01001000100), .b(t0_01001000101), .y(t0_0100100010));
wire t0_01001000100, t0_01001000101;
mixer mix_t0_01001000100 (.a(t0_010010001000), .b(t0_010010001001), .y(t0_01001000100));
wire t0_010010001000, t0_010010001001;
mixer mix_t0_01001000101 (.a(t0_010010001010), .b(t0_010010001011), .y(t0_01001000101));
wire t0_010010001010, t0_010010001011;
mixer mix_t0_0100100011 (.a(t0_01001000110), .b(t0_01001000111), .y(t0_0100100011));
wire t0_01001000110, t0_01001000111;
mixer mix_t0_01001000110 (.a(t0_010010001100), .b(t0_010010001101), .y(t0_01001000110));
wire t0_010010001100, t0_010010001101;
mixer mix_t0_01001000111 (.a(t0_010010001110), .b(t0_010010001111), .y(t0_01001000111));
wire t0_010010001110, t0_010010001111;
mixer mix_t0_01001001 (.a(t0_010010010), .b(t0_010010011), .y(t0_01001001));
wire t0_010010010, t0_010010011;
mixer mix_t0_010010010 (.a(t0_0100100100), .b(t0_0100100101), .y(t0_010010010));
wire t0_0100100100, t0_0100100101;
mixer mix_t0_0100100100 (.a(t0_01001001000), .b(t0_01001001001), .y(t0_0100100100));
wire t0_01001001000, t0_01001001001;
mixer mix_t0_01001001000 (.a(t0_010010010000), .b(t0_010010010001), .y(t0_01001001000));
wire t0_010010010000, t0_010010010001;
mixer mix_t0_01001001001 (.a(t0_010010010010), .b(t0_010010010011), .y(t0_01001001001));
wire t0_010010010010, t0_010010010011;
mixer mix_t0_0100100101 (.a(t0_01001001010), .b(t0_01001001011), .y(t0_0100100101));
wire t0_01001001010, t0_01001001011;
mixer mix_t0_01001001010 (.a(t0_010010010100), .b(t0_010010010101), .y(t0_01001001010));
wire t0_010010010100, t0_010010010101;
mixer mix_t0_01001001011 (.a(t0_010010010110), .b(t0_010010010111), .y(t0_01001001011));
wire t0_010010010110, t0_010010010111;
mixer mix_t0_010010011 (.a(t0_0100100110), .b(t0_0100100111), .y(t0_010010011));
wire t0_0100100110, t0_0100100111;
mixer mix_t0_0100100110 (.a(t0_01001001100), .b(t0_01001001101), .y(t0_0100100110));
wire t0_01001001100, t0_01001001101;
mixer mix_t0_01001001100 (.a(t0_010010011000), .b(t0_010010011001), .y(t0_01001001100));
wire t0_010010011000, t0_010010011001;
mixer mix_t0_01001001101 (.a(t0_010010011010), .b(t0_010010011011), .y(t0_01001001101));
wire t0_010010011010, t0_010010011011;
mixer mix_t0_0100100111 (.a(t0_01001001110), .b(t0_01001001111), .y(t0_0100100111));
wire t0_01001001110, t0_01001001111;
mixer mix_t0_01001001110 (.a(t0_010010011100), .b(t0_010010011101), .y(t0_01001001110));
wire t0_010010011100, t0_010010011101;
mixer mix_t0_01001001111 (.a(t0_010010011110), .b(t0_010010011111), .y(t0_01001001111));
wire t0_010010011110, t0_010010011111;
mixer mix_t0_0100101 (.a(t0_01001010), .b(t0_01001011), .y(t0_0100101));
wire t0_01001010, t0_01001011;
mixer mix_t0_01001010 (.a(t0_010010100), .b(t0_010010101), .y(t0_01001010));
wire t0_010010100, t0_010010101;
mixer mix_t0_010010100 (.a(t0_0100101000), .b(t0_0100101001), .y(t0_010010100));
wire t0_0100101000, t0_0100101001;
mixer mix_t0_0100101000 (.a(t0_01001010000), .b(t0_01001010001), .y(t0_0100101000));
wire t0_01001010000, t0_01001010001;
mixer mix_t0_01001010000 (.a(t0_010010100000), .b(t0_010010100001), .y(t0_01001010000));
wire t0_010010100000, t0_010010100001;
mixer mix_t0_01001010001 (.a(t0_010010100010), .b(t0_010010100011), .y(t0_01001010001));
wire t0_010010100010, t0_010010100011;
mixer mix_t0_0100101001 (.a(t0_01001010010), .b(t0_01001010011), .y(t0_0100101001));
wire t0_01001010010, t0_01001010011;
mixer mix_t0_01001010010 (.a(t0_010010100100), .b(t0_010010100101), .y(t0_01001010010));
wire t0_010010100100, t0_010010100101;
mixer mix_t0_01001010011 (.a(t0_010010100110), .b(t0_010010100111), .y(t0_01001010011));
wire t0_010010100110, t0_010010100111;
mixer mix_t0_010010101 (.a(t0_0100101010), .b(t0_0100101011), .y(t0_010010101));
wire t0_0100101010, t0_0100101011;
mixer mix_t0_0100101010 (.a(t0_01001010100), .b(t0_01001010101), .y(t0_0100101010));
wire t0_01001010100, t0_01001010101;
mixer mix_t0_01001010100 (.a(t0_010010101000), .b(t0_010010101001), .y(t0_01001010100));
wire t0_010010101000, t0_010010101001;
mixer mix_t0_01001010101 (.a(t0_010010101010), .b(t0_010010101011), .y(t0_01001010101));
wire t0_010010101010, t0_010010101011;
mixer mix_t0_0100101011 (.a(t0_01001010110), .b(t0_01001010111), .y(t0_0100101011));
wire t0_01001010110, t0_01001010111;
mixer mix_t0_01001010110 (.a(t0_010010101100), .b(t0_010010101101), .y(t0_01001010110));
wire t0_010010101100, t0_010010101101;
mixer mix_t0_01001010111 (.a(t0_010010101110), .b(t0_010010101111), .y(t0_01001010111));
wire t0_010010101110, t0_010010101111;
mixer mix_t0_01001011 (.a(t0_010010110), .b(t0_010010111), .y(t0_01001011));
wire t0_010010110, t0_010010111;
mixer mix_t0_010010110 (.a(t0_0100101100), .b(t0_0100101101), .y(t0_010010110));
wire t0_0100101100, t0_0100101101;
mixer mix_t0_0100101100 (.a(t0_01001011000), .b(t0_01001011001), .y(t0_0100101100));
wire t0_01001011000, t0_01001011001;
mixer mix_t0_01001011000 (.a(t0_010010110000), .b(t0_010010110001), .y(t0_01001011000));
wire t0_010010110000, t0_010010110001;
mixer mix_t0_01001011001 (.a(t0_010010110010), .b(t0_010010110011), .y(t0_01001011001));
wire t0_010010110010, t0_010010110011;
mixer mix_t0_0100101101 (.a(t0_01001011010), .b(t0_01001011011), .y(t0_0100101101));
wire t0_01001011010, t0_01001011011;
mixer mix_t0_01001011010 (.a(t0_010010110100), .b(t0_010010110101), .y(t0_01001011010));
wire t0_010010110100, t0_010010110101;
mixer mix_t0_01001011011 (.a(t0_010010110110), .b(t0_010010110111), .y(t0_01001011011));
wire t0_010010110110, t0_010010110111;
mixer mix_t0_010010111 (.a(t0_0100101110), .b(t0_0100101111), .y(t0_010010111));
wire t0_0100101110, t0_0100101111;
mixer mix_t0_0100101110 (.a(t0_01001011100), .b(t0_01001011101), .y(t0_0100101110));
wire t0_01001011100, t0_01001011101;
mixer mix_t0_01001011100 (.a(t0_010010111000), .b(t0_010010111001), .y(t0_01001011100));
wire t0_010010111000, t0_010010111001;
mixer mix_t0_01001011101 (.a(t0_010010111010), .b(t0_010010111011), .y(t0_01001011101));
wire t0_010010111010, t0_010010111011;
mixer mix_t0_0100101111 (.a(t0_01001011110), .b(t0_01001011111), .y(t0_0100101111));
wire t0_01001011110, t0_01001011111;
mixer mix_t0_01001011110 (.a(t0_010010111100), .b(t0_010010111101), .y(t0_01001011110));
wire t0_010010111100, t0_010010111101;
mixer mix_t0_01001011111 (.a(t0_010010111110), .b(t0_010010111111), .y(t0_01001011111));
wire t0_010010111110, t0_010010111111;
mixer mix_t0_010011 (.a(t0_0100110), .b(t0_0100111), .y(t0_010011));
wire t0_0100110, t0_0100111;
mixer mix_t0_0100110 (.a(t0_01001100), .b(t0_01001101), .y(t0_0100110));
wire t0_01001100, t0_01001101;
mixer mix_t0_01001100 (.a(t0_010011000), .b(t0_010011001), .y(t0_01001100));
wire t0_010011000, t0_010011001;
mixer mix_t0_010011000 (.a(t0_0100110000), .b(t0_0100110001), .y(t0_010011000));
wire t0_0100110000, t0_0100110001;
mixer mix_t0_0100110000 (.a(t0_01001100000), .b(t0_01001100001), .y(t0_0100110000));
wire t0_01001100000, t0_01001100001;
mixer mix_t0_01001100000 (.a(t0_010011000000), .b(t0_010011000001), .y(t0_01001100000));
wire t0_010011000000, t0_010011000001;
mixer mix_t0_01001100001 (.a(t0_010011000010), .b(t0_010011000011), .y(t0_01001100001));
wire t0_010011000010, t0_010011000011;
mixer mix_t0_0100110001 (.a(t0_01001100010), .b(t0_01001100011), .y(t0_0100110001));
wire t0_01001100010, t0_01001100011;
mixer mix_t0_01001100010 (.a(t0_010011000100), .b(t0_010011000101), .y(t0_01001100010));
wire t0_010011000100, t0_010011000101;
mixer mix_t0_01001100011 (.a(t0_010011000110), .b(t0_010011000111), .y(t0_01001100011));
wire t0_010011000110, t0_010011000111;
mixer mix_t0_010011001 (.a(t0_0100110010), .b(t0_0100110011), .y(t0_010011001));
wire t0_0100110010, t0_0100110011;
mixer mix_t0_0100110010 (.a(t0_01001100100), .b(t0_01001100101), .y(t0_0100110010));
wire t0_01001100100, t0_01001100101;
mixer mix_t0_01001100100 (.a(t0_010011001000), .b(t0_010011001001), .y(t0_01001100100));
wire t0_010011001000, t0_010011001001;
mixer mix_t0_01001100101 (.a(t0_010011001010), .b(t0_010011001011), .y(t0_01001100101));
wire t0_010011001010, t0_010011001011;
mixer mix_t0_0100110011 (.a(t0_01001100110), .b(t0_01001100111), .y(t0_0100110011));
wire t0_01001100110, t0_01001100111;
mixer mix_t0_01001100110 (.a(t0_010011001100), .b(t0_010011001101), .y(t0_01001100110));
wire t0_010011001100, t0_010011001101;
mixer mix_t0_01001100111 (.a(t0_010011001110), .b(t0_010011001111), .y(t0_01001100111));
wire t0_010011001110, t0_010011001111;
mixer mix_t0_01001101 (.a(t0_010011010), .b(t0_010011011), .y(t0_01001101));
wire t0_010011010, t0_010011011;
mixer mix_t0_010011010 (.a(t0_0100110100), .b(t0_0100110101), .y(t0_010011010));
wire t0_0100110100, t0_0100110101;
mixer mix_t0_0100110100 (.a(t0_01001101000), .b(t0_01001101001), .y(t0_0100110100));
wire t0_01001101000, t0_01001101001;
mixer mix_t0_01001101000 (.a(t0_010011010000), .b(t0_010011010001), .y(t0_01001101000));
wire t0_010011010000, t0_010011010001;
mixer mix_t0_01001101001 (.a(t0_010011010010), .b(t0_010011010011), .y(t0_01001101001));
wire t0_010011010010, t0_010011010011;
mixer mix_t0_0100110101 (.a(t0_01001101010), .b(t0_01001101011), .y(t0_0100110101));
wire t0_01001101010, t0_01001101011;
mixer mix_t0_01001101010 (.a(t0_010011010100), .b(t0_010011010101), .y(t0_01001101010));
wire t0_010011010100, t0_010011010101;
mixer mix_t0_01001101011 (.a(t0_010011010110), .b(t0_010011010111), .y(t0_01001101011));
wire t0_010011010110, t0_010011010111;
mixer mix_t0_010011011 (.a(t0_0100110110), .b(t0_0100110111), .y(t0_010011011));
wire t0_0100110110, t0_0100110111;
mixer mix_t0_0100110110 (.a(t0_01001101100), .b(t0_01001101101), .y(t0_0100110110));
wire t0_01001101100, t0_01001101101;
mixer mix_t0_01001101100 (.a(t0_010011011000), .b(t0_010011011001), .y(t0_01001101100));
wire t0_010011011000, t0_010011011001;
mixer mix_t0_01001101101 (.a(t0_010011011010), .b(t0_010011011011), .y(t0_01001101101));
wire t0_010011011010, t0_010011011011;
mixer mix_t0_0100110111 (.a(t0_01001101110), .b(t0_01001101111), .y(t0_0100110111));
wire t0_01001101110, t0_01001101111;
mixer mix_t0_01001101110 (.a(t0_010011011100), .b(t0_010011011101), .y(t0_01001101110));
wire t0_010011011100, t0_010011011101;
mixer mix_t0_01001101111 (.a(t0_010011011110), .b(t0_010011011111), .y(t0_01001101111));
wire t0_010011011110, t0_010011011111;
mixer mix_t0_0100111 (.a(t0_01001110), .b(t0_01001111), .y(t0_0100111));
wire t0_01001110, t0_01001111;
mixer mix_t0_01001110 (.a(t0_010011100), .b(t0_010011101), .y(t0_01001110));
wire t0_010011100, t0_010011101;
mixer mix_t0_010011100 (.a(t0_0100111000), .b(t0_0100111001), .y(t0_010011100));
wire t0_0100111000, t0_0100111001;
mixer mix_t0_0100111000 (.a(t0_01001110000), .b(t0_01001110001), .y(t0_0100111000));
wire t0_01001110000, t0_01001110001;
mixer mix_t0_01001110000 (.a(t0_010011100000), .b(t0_010011100001), .y(t0_01001110000));
wire t0_010011100000, t0_010011100001;
mixer mix_t0_01001110001 (.a(t0_010011100010), .b(t0_010011100011), .y(t0_01001110001));
wire t0_010011100010, t0_010011100011;
mixer mix_t0_0100111001 (.a(t0_01001110010), .b(t0_01001110011), .y(t0_0100111001));
wire t0_01001110010, t0_01001110011;
mixer mix_t0_01001110010 (.a(t0_010011100100), .b(t0_010011100101), .y(t0_01001110010));
wire t0_010011100100, t0_010011100101;
mixer mix_t0_01001110011 (.a(t0_010011100110), .b(t0_010011100111), .y(t0_01001110011));
wire t0_010011100110, t0_010011100111;
mixer mix_t0_010011101 (.a(t0_0100111010), .b(t0_0100111011), .y(t0_010011101));
wire t0_0100111010, t0_0100111011;
mixer mix_t0_0100111010 (.a(t0_01001110100), .b(t0_01001110101), .y(t0_0100111010));
wire t0_01001110100, t0_01001110101;
mixer mix_t0_01001110100 (.a(t0_010011101000), .b(t0_010011101001), .y(t0_01001110100));
wire t0_010011101000, t0_010011101001;
mixer mix_t0_01001110101 (.a(t0_010011101010), .b(t0_010011101011), .y(t0_01001110101));
wire t0_010011101010, t0_010011101011;
mixer mix_t0_0100111011 (.a(t0_01001110110), .b(t0_01001110111), .y(t0_0100111011));
wire t0_01001110110, t0_01001110111;
mixer mix_t0_01001110110 (.a(t0_010011101100), .b(t0_010011101101), .y(t0_01001110110));
wire t0_010011101100, t0_010011101101;
mixer mix_t0_01001110111 (.a(t0_010011101110), .b(t0_010011101111), .y(t0_01001110111));
wire t0_010011101110, t0_010011101111;
mixer mix_t0_01001111 (.a(t0_010011110), .b(t0_010011111), .y(t0_01001111));
wire t0_010011110, t0_010011111;
mixer mix_t0_010011110 (.a(t0_0100111100), .b(t0_0100111101), .y(t0_010011110));
wire t0_0100111100, t0_0100111101;
mixer mix_t0_0100111100 (.a(t0_01001111000), .b(t0_01001111001), .y(t0_0100111100));
wire t0_01001111000, t0_01001111001;
mixer mix_t0_01001111000 (.a(t0_010011110000), .b(t0_010011110001), .y(t0_01001111000));
wire t0_010011110000, t0_010011110001;
mixer mix_t0_01001111001 (.a(t0_010011110010), .b(t0_010011110011), .y(t0_01001111001));
wire t0_010011110010, t0_010011110011;
mixer mix_t0_0100111101 (.a(t0_01001111010), .b(t0_01001111011), .y(t0_0100111101));
wire t0_01001111010, t0_01001111011;
mixer mix_t0_01001111010 (.a(t0_010011110100), .b(t0_010011110101), .y(t0_01001111010));
wire t0_010011110100, t0_010011110101;
mixer mix_t0_01001111011 (.a(t0_010011110110), .b(t0_010011110111), .y(t0_01001111011));
wire t0_010011110110, t0_010011110111;
mixer mix_t0_010011111 (.a(t0_0100111110), .b(t0_0100111111), .y(t0_010011111));
wire t0_0100111110, t0_0100111111;
mixer mix_t0_0100111110 (.a(t0_01001111100), .b(t0_01001111101), .y(t0_0100111110));
wire t0_01001111100, t0_01001111101;
mixer mix_t0_01001111100 (.a(t0_010011111000), .b(t0_010011111001), .y(t0_01001111100));
wire t0_010011111000, t0_010011111001;
mixer mix_t0_01001111101 (.a(t0_010011111010), .b(t0_010011111011), .y(t0_01001111101));
wire t0_010011111010, t0_010011111011;
mixer mix_t0_0100111111 (.a(t0_01001111110), .b(t0_01001111111), .y(t0_0100111111));
wire t0_01001111110, t0_01001111111;
mixer mix_t0_01001111110 (.a(t0_010011111100), .b(t0_010011111101), .y(t0_01001111110));
wire t0_010011111100, t0_010011111101;
mixer mix_t0_01001111111 (.a(t0_010011111110), .b(t0_010011111111), .y(t0_01001111111));
wire t0_010011111110, t0_010011111111;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_010100 (.a(t0_0101000), .b(t0_0101001), .y(t0_010100));
wire t0_0101000, t0_0101001;
mixer mix_t0_0101000 (.a(t0_01010000), .b(t0_01010001), .y(t0_0101000));
wire t0_01010000, t0_01010001;
mixer mix_t0_01010000 (.a(t0_010100000), .b(t0_010100001), .y(t0_01010000));
wire t0_010100000, t0_010100001;
mixer mix_t0_010100000 (.a(t0_0101000000), .b(t0_0101000001), .y(t0_010100000));
wire t0_0101000000, t0_0101000001;
mixer mix_t0_0101000000 (.a(t0_01010000000), .b(t0_01010000001), .y(t0_0101000000));
wire t0_01010000000, t0_01010000001;
mixer mix_t0_01010000000 (.a(t0_010100000000), .b(t0_010100000001), .y(t0_01010000000));
wire t0_010100000000, t0_010100000001;
mixer mix_t0_01010000001 (.a(t0_010100000010), .b(t0_010100000011), .y(t0_01010000001));
wire t0_010100000010, t0_010100000011;
mixer mix_t0_0101000001 (.a(t0_01010000010), .b(t0_01010000011), .y(t0_0101000001));
wire t0_01010000010, t0_01010000011;
mixer mix_t0_01010000010 (.a(t0_010100000100), .b(t0_010100000101), .y(t0_01010000010));
wire t0_010100000100, t0_010100000101;
mixer mix_t0_01010000011 (.a(t0_010100000110), .b(t0_010100000111), .y(t0_01010000011));
wire t0_010100000110, t0_010100000111;
mixer mix_t0_010100001 (.a(t0_0101000010), .b(t0_0101000011), .y(t0_010100001));
wire t0_0101000010, t0_0101000011;
mixer mix_t0_0101000010 (.a(t0_01010000100), .b(t0_01010000101), .y(t0_0101000010));
wire t0_01010000100, t0_01010000101;
mixer mix_t0_01010000100 (.a(t0_010100001000), .b(t0_010100001001), .y(t0_01010000100));
wire t0_010100001000, t0_010100001001;
mixer mix_t0_01010000101 (.a(t0_010100001010), .b(t0_010100001011), .y(t0_01010000101));
wire t0_010100001010, t0_010100001011;
mixer mix_t0_0101000011 (.a(t0_01010000110), .b(t0_01010000111), .y(t0_0101000011));
wire t0_01010000110, t0_01010000111;
mixer mix_t0_01010000110 (.a(t0_010100001100), .b(t0_010100001101), .y(t0_01010000110));
wire t0_010100001100, t0_010100001101;
mixer mix_t0_01010000111 (.a(t0_010100001110), .b(t0_010100001111), .y(t0_01010000111));
wire t0_010100001110, t0_010100001111;
mixer mix_t0_01010001 (.a(t0_010100010), .b(t0_010100011), .y(t0_01010001));
wire t0_010100010, t0_010100011;
mixer mix_t0_010100010 (.a(t0_0101000100), .b(t0_0101000101), .y(t0_010100010));
wire t0_0101000100, t0_0101000101;
mixer mix_t0_0101000100 (.a(t0_01010001000), .b(t0_01010001001), .y(t0_0101000100));
wire t0_01010001000, t0_01010001001;
mixer mix_t0_01010001000 (.a(t0_010100010000), .b(t0_010100010001), .y(t0_01010001000));
wire t0_010100010000, t0_010100010001;
mixer mix_t0_01010001001 (.a(t0_010100010010), .b(t0_010100010011), .y(t0_01010001001));
wire t0_010100010010, t0_010100010011;
mixer mix_t0_0101000101 (.a(t0_01010001010), .b(t0_01010001011), .y(t0_0101000101));
wire t0_01010001010, t0_01010001011;
mixer mix_t0_01010001010 (.a(t0_010100010100), .b(t0_010100010101), .y(t0_01010001010));
wire t0_010100010100, t0_010100010101;
mixer mix_t0_01010001011 (.a(t0_010100010110), .b(t0_010100010111), .y(t0_01010001011));
wire t0_010100010110, t0_010100010111;
mixer mix_t0_010100011 (.a(t0_0101000110), .b(t0_0101000111), .y(t0_010100011));
wire t0_0101000110, t0_0101000111;
mixer mix_t0_0101000110 (.a(t0_01010001100), .b(t0_01010001101), .y(t0_0101000110));
wire t0_01010001100, t0_01010001101;
mixer mix_t0_01010001100 (.a(t0_010100011000), .b(t0_010100011001), .y(t0_01010001100));
wire t0_010100011000, t0_010100011001;
mixer mix_t0_01010001101 (.a(t0_010100011010), .b(t0_010100011011), .y(t0_01010001101));
wire t0_010100011010, t0_010100011011;
mixer mix_t0_0101000111 (.a(t0_01010001110), .b(t0_01010001111), .y(t0_0101000111));
wire t0_01010001110, t0_01010001111;
mixer mix_t0_01010001110 (.a(t0_010100011100), .b(t0_010100011101), .y(t0_01010001110));
wire t0_010100011100, t0_010100011101;
mixer mix_t0_01010001111 (.a(t0_010100011110), .b(t0_010100011111), .y(t0_01010001111));
wire t0_010100011110, t0_010100011111;
mixer mix_t0_0101001 (.a(t0_01010010), .b(t0_01010011), .y(t0_0101001));
wire t0_01010010, t0_01010011;
mixer mix_t0_01010010 (.a(t0_010100100), .b(t0_010100101), .y(t0_01010010));
wire t0_010100100, t0_010100101;
mixer mix_t0_010100100 (.a(t0_0101001000), .b(t0_0101001001), .y(t0_010100100));
wire t0_0101001000, t0_0101001001;
mixer mix_t0_0101001000 (.a(t0_01010010000), .b(t0_01010010001), .y(t0_0101001000));
wire t0_01010010000, t0_01010010001;
mixer mix_t0_01010010000 (.a(t0_010100100000), .b(t0_010100100001), .y(t0_01010010000));
wire t0_010100100000, t0_010100100001;
mixer mix_t0_01010010001 (.a(t0_010100100010), .b(t0_010100100011), .y(t0_01010010001));
wire t0_010100100010, t0_010100100011;
mixer mix_t0_0101001001 (.a(t0_01010010010), .b(t0_01010010011), .y(t0_0101001001));
wire t0_01010010010, t0_01010010011;
mixer mix_t0_01010010010 (.a(t0_010100100100), .b(t0_010100100101), .y(t0_01010010010));
wire t0_010100100100, t0_010100100101;
mixer mix_t0_01010010011 (.a(t0_010100100110), .b(t0_010100100111), .y(t0_01010010011));
wire t0_010100100110, t0_010100100111;
mixer mix_t0_010100101 (.a(t0_0101001010), .b(t0_0101001011), .y(t0_010100101));
wire t0_0101001010, t0_0101001011;
mixer mix_t0_0101001010 (.a(t0_01010010100), .b(t0_01010010101), .y(t0_0101001010));
wire t0_01010010100, t0_01010010101;
mixer mix_t0_01010010100 (.a(t0_010100101000), .b(t0_010100101001), .y(t0_01010010100));
wire t0_010100101000, t0_010100101001;
mixer mix_t0_01010010101 (.a(t0_010100101010), .b(t0_010100101011), .y(t0_01010010101));
wire t0_010100101010, t0_010100101011;
mixer mix_t0_0101001011 (.a(t0_01010010110), .b(t0_01010010111), .y(t0_0101001011));
wire t0_01010010110, t0_01010010111;
mixer mix_t0_01010010110 (.a(t0_010100101100), .b(t0_010100101101), .y(t0_01010010110));
wire t0_010100101100, t0_010100101101;
mixer mix_t0_01010010111 (.a(t0_010100101110), .b(t0_010100101111), .y(t0_01010010111));
wire t0_010100101110, t0_010100101111;
mixer mix_t0_01010011 (.a(t0_010100110), .b(t0_010100111), .y(t0_01010011));
wire t0_010100110, t0_010100111;
mixer mix_t0_010100110 (.a(t0_0101001100), .b(t0_0101001101), .y(t0_010100110));
wire t0_0101001100, t0_0101001101;
mixer mix_t0_0101001100 (.a(t0_01010011000), .b(t0_01010011001), .y(t0_0101001100));
wire t0_01010011000, t0_01010011001;
mixer mix_t0_01010011000 (.a(t0_010100110000), .b(t0_010100110001), .y(t0_01010011000));
wire t0_010100110000, t0_010100110001;
mixer mix_t0_01010011001 (.a(t0_010100110010), .b(t0_010100110011), .y(t0_01010011001));
wire t0_010100110010, t0_010100110011;
mixer mix_t0_0101001101 (.a(t0_01010011010), .b(t0_01010011011), .y(t0_0101001101));
wire t0_01010011010, t0_01010011011;
mixer mix_t0_01010011010 (.a(t0_010100110100), .b(t0_010100110101), .y(t0_01010011010));
wire t0_010100110100, t0_010100110101;
mixer mix_t0_01010011011 (.a(t0_010100110110), .b(t0_010100110111), .y(t0_01010011011));
wire t0_010100110110, t0_010100110111;
mixer mix_t0_010100111 (.a(t0_0101001110), .b(t0_0101001111), .y(t0_010100111));
wire t0_0101001110, t0_0101001111;
mixer mix_t0_0101001110 (.a(t0_01010011100), .b(t0_01010011101), .y(t0_0101001110));
wire t0_01010011100, t0_01010011101;
mixer mix_t0_01010011100 (.a(t0_010100111000), .b(t0_010100111001), .y(t0_01010011100));
wire t0_010100111000, t0_010100111001;
mixer mix_t0_01010011101 (.a(t0_010100111010), .b(t0_010100111011), .y(t0_01010011101));
wire t0_010100111010, t0_010100111011;
mixer mix_t0_0101001111 (.a(t0_01010011110), .b(t0_01010011111), .y(t0_0101001111));
wire t0_01010011110, t0_01010011111;
mixer mix_t0_01010011110 (.a(t0_010100111100), .b(t0_010100111101), .y(t0_01010011110));
wire t0_010100111100, t0_010100111101;
mixer mix_t0_01010011111 (.a(t0_010100111110), .b(t0_010100111111), .y(t0_01010011111));
wire t0_010100111110, t0_010100111111;
mixer mix_t0_010101 (.a(t0_0101010), .b(t0_0101011), .y(t0_010101));
wire t0_0101010, t0_0101011;
mixer mix_t0_0101010 (.a(t0_01010100), .b(t0_01010101), .y(t0_0101010));
wire t0_01010100, t0_01010101;
mixer mix_t0_01010100 (.a(t0_010101000), .b(t0_010101001), .y(t0_01010100));
wire t0_010101000, t0_010101001;
mixer mix_t0_010101000 (.a(t0_0101010000), .b(t0_0101010001), .y(t0_010101000));
wire t0_0101010000, t0_0101010001;
mixer mix_t0_0101010000 (.a(t0_01010100000), .b(t0_01010100001), .y(t0_0101010000));
wire t0_01010100000, t0_01010100001;
mixer mix_t0_01010100000 (.a(t0_010101000000), .b(t0_010101000001), .y(t0_01010100000));
wire t0_010101000000, t0_010101000001;
mixer mix_t0_01010100001 (.a(t0_010101000010), .b(t0_010101000011), .y(t0_01010100001));
wire t0_010101000010, t0_010101000011;
mixer mix_t0_0101010001 (.a(t0_01010100010), .b(t0_01010100011), .y(t0_0101010001));
wire t0_01010100010, t0_01010100011;
mixer mix_t0_01010100010 (.a(t0_010101000100), .b(t0_010101000101), .y(t0_01010100010));
wire t0_010101000100, t0_010101000101;
mixer mix_t0_01010100011 (.a(t0_010101000110), .b(t0_010101000111), .y(t0_01010100011));
wire t0_010101000110, t0_010101000111;
mixer mix_t0_010101001 (.a(t0_0101010010), .b(t0_0101010011), .y(t0_010101001));
wire t0_0101010010, t0_0101010011;
mixer mix_t0_0101010010 (.a(t0_01010100100), .b(t0_01010100101), .y(t0_0101010010));
wire t0_01010100100, t0_01010100101;
mixer mix_t0_01010100100 (.a(t0_010101001000), .b(t0_010101001001), .y(t0_01010100100));
wire t0_010101001000, t0_010101001001;
mixer mix_t0_01010100101 (.a(t0_010101001010), .b(t0_010101001011), .y(t0_01010100101));
wire t0_010101001010, t0_010101001011;
mixer mix_t0_0101010011 (.a(t0_01010100110), .b(t0_01010100111), .y(t0_0101010011));
wire t0_01010100110, t0_01010100111;
mixer mix_t0_01010100110 (.a(t0_010101001100), .b(t0_010101001101), .y(t0_01010100110));
wire t0_010101001100, t0_010101001101;
mixer mix_t0_01010100111 (.a(t0_010101001110), .b(t0_010101001111), .y(t0_01010100111));
wire t0_010101001110, t0_010101001111;
mixer mix_t0_01010101 (.a(t0_010101010), .b(t0_010101011), .y(t0_01010101));
wire t0_010101010, t0_010101011;
mixer mix_t0_010101010 (.a(t0_0101010100), .b(t0_0101010101), .y(t0_010101010));
wire t0_0101010100, t0_0101010101;
mixer mix_t0_0101010100 (.a(t0_01010101000), .b(t0_01010101001), .y(t0_0101010100));
wire t0_01010101000, t0_01010101001;
mixer mix_t0_01010101000 (.a(t0_010101010000), .b(t0_010101010001), .y(t0_01010101000));
wire t0_010101010000, t0_010101010001;
mixer mix_t0_01010101001 (.a(t0_010101010010), .b(t0_010101010011), .y(t0_01010101001));
wire t0_010101010010, t0_010101010011;
mixer mix_t0_0101010101 (.a(t0_01010101010), .b(t0_01010101011), .y(t0_0101010101));
wire t0_01010101010, t0_01010101011;
mixer mix_t0_01010101010 (.a(t0_010101010100), .b(t0_010101010101), .y(t0_01010101010));
wire t0_010101010100, t0_010101010101;
mixer mix_t0_01010101011 (.a(t0_010101010110), .b(t0_010101010111), .y(t0_01010101011));
wire t0_010101010110, t0_010101010111;
mixer mix_t0_010101011 (.a(t0_0101010110), .b(t0_0101010111), .y(t0_010101011));
wire t0_0101010110, t0_0101010111;
mixer mix_t0_0101010110 (.a(t0_01010101100), .b(t0_01010101101), .y(t0_0101010110));
wire t0_01010101100, t0_01010101101;
mixer mix_t0_01010101100 (.a(t0_010101011000), .b(t0_010101011001), .y(t0_01010101100));
wire t0_010101011000, t0_010101011001;
mixer mix_t0_01010101101 (.a(t0_010101011010), .b(t0_010101011011), .y(t0_01010101101));
wire t0_010101011010, t0_010101011011;
mixer mix_t0_0101010111 (.a(t0_01010101110), .b(t0_01010101111), .y(t0_0101010111));
wire t0_01010101110, t0_01010101111;
mixer mix_t0_01010101110 (.a(t0_010101011100), .b(t0_010101011101), .y(t0_01010101110));
wire t0_010101011100, t0_010101011101;
mixer mix_t0_01010101111 (.a(t0_010101011110), .b(t0_010101011111), .y(t0_01010101111));
wire t0_010101011110, t0_010101011111;
mixer mix_t0_0101011 (.a(t0_01010110), .b(t0_01010111), .y(t0_0101011));
wire t0_01010110, t0_01010111;
mixer mix_t0_01010110 (.a(t0_010101100), .b(t0_010101101), .y(t0_01010110));
wire t0_010101100, t0_010101101;
mixer mix_t0_010101100 (.a(t0_0101011000), .b(t0_0101011001), .y(t0_010101100));
wire t0_0101011000, t0_0101011001;
mixer mix_t0_0101011000 (.a(t0_01010110000), .b(t0_01010110001), .y(t0_0101011000));
wire t0_01010110000, t0_01010110001;
mixer mix_t0_01010110000 (.a(t0_010101100000), .b(t0_010101100001), .y(t0_01010110000));
wire t0_010101100000, t0_010101100001;
mixer mix_t0_01010110001 (.a(t0_010101100010), .b(t0_010101100011), .y(t0_01010110001));
wire t0_010101100010, t0_010101100011;
mixer mix_t0_0101011001 (.a(t0_01010110010), .b(t0_01010110011), .y(t0_0101011001));
wire t0_01010110010, t0_01010110011;
mixer mix_t0_01010110010 (.a(t0_010101100100), .b(t0_010101100101), .y(t0_01010110010));
wire t0_010101100100, t0_010101100101;
mixer mix_t0_01010110011 (.a(t0_010101100110), .b(t0_010101100111), .y(t0_01010110011));
wire t0_010101100110, t0_010101100111;
mixer mix_t0_010101101 (.a(t0_0101011010), .b(t0_0101011011), .y(t0_010101101));
wire t0_0101011010, t0_0101011011;
mixer mix_t0_0101011010 (.a(t0_01010110100), .b(t0_01010110101), .y(t0_0101011010));
wire t0_01010110100, t0_01010110101;
mixer mix_t0_01010110100 (.a(t0_010101101000), .b(t0_010101101001), .y(t0_01010110100));
wire t0_010101101000, t0_010101101001;
mixer mix_t0_01010110101 (.a(t0_010101101010), .b(t0_010101101011), .y(t0_01010110101));
wire t0_010101101010, t0_010101101011;
mixer mix_t0_0101011011 (.a(t0_01010110110), .b(t0_01010110111), .y(t0_0101011011));
wire t0_01010110110, t0_01010110111;
mixer mix_t0_01010110110 (.a(t0_010101101100), .b(t0_010101101101), .y(t0_01010110110));
wire t0_010101101100, t0_010101101101;
mixer mix_t0_01010110111 (.a(t0_010101101110), .b(t0_010101101111), .y(t0_01010110111));
wire t0_010101101110, t0_010101101111;
mixer mix_t0_01010111 (.a(t0_010101110), .b(t0_010101111), .y(t0_01010111));
wire t0_010101110, t0_010101111;
mixer mix_t0_010101110 (.a(t0_0101011100), .b(t0_0101011101), .y(t0_010101110));
wire t0_0101011100, t0_0101011101;
mixer mix_t0_0101011100 (.a(t0_01010111000), .b(t0_01010111001), .y(t0_0101011100));
wire t0_01010111000, t0_01010111001;
mixer mix_t0_01010111000 (.a(t0_010101110000), .b(t0_010101110001), .y(t0_01010111000));
wire t0_010101110000, t0_010101110001;
mixer mix_t0_01010111001 (.a(t0_010101110010), .b(t0_010101110011), .y(t0_01010111001));
wire t0_010101110010, t0_010101110011;
mixer mix_t0_0101011101 (.a(t0_01010111010), .b(t0_01010111011), .y(t0_0101011101));
wire t0_01010111010, t0_01010111011;
mixer mix_t0_01010111010 (.a(t0_010101110100), .b(t0_010101110101), .y(t0_01010111010));
wire t0_010101110100, t0_010101110101;
mixer mix_t0_01010111011 (.a(t0_010101110110), .b(t0_010101110111), .y(t0_01010111011));
wire t0_010101110110, t0_010101110111;
mixer mix_t0_010101111 (.a(t0_0101011110), .b(t0_0101011111), .y(t0_010101111));
wire t0_0101011110, t0_0101011111;
mixer mix_t0_0101011110 (.a(t0_01010111100), .b(t0_01010111101), .y(t0_0101011110));
wire t0_01010111100, t0_01010111101;
mixer mix_t0_01010111100 (.a(t0_010101111000), .b(t0_010101111001), .y(t0_01010111100));
wire t0_010101111000, t0_010101111001;
mixer mix_t0_01010111101 (.a(t0_010101111010), .b(t0_010101111011), .y(t0_01010111101));
wire t0_010101111010, t0_010101111011;
mixer mix_t0_0101011111 (.a(t0_01010111110), .b(t0_01010111111), .y(t0_0101011111));
wire t0_01010111110, t0_01010111111;
mixer mix_t0_01010111110 (.a(t0_010101111100), .b(t0_010101111101), .y(t0_01010111110));
wire t0_010101111100, t0_010101111101;
mixer mix_t0_01010111111 (.a(t0_010101111110), .b(t0_010101111111), .y(t0_01010111111));
wire t0_010101111110, t0_010101111111;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_010110 (.a(t0_0101100), .b(t0_0101101), .y(t0_010110));
wire t0_0101100, t0_0101101;
mixer mix_t0_0101100 (.a(t0_01011000), .b(t0_01011001), .y(t0_0101100));
wire t0_01011000, t0_01011001;
mixer mix_t0_01011000 (.a(t0_010110000), .b(t0_010110001), .y(t0_01011000));
wire t0_010110000, t0_010110001;
mixer mix_t0_010110000 (.a(t0_0101100000), .b(t0_0101100001), .y(t0_010110000));
wire t0_0101100000, t0_0101100001;
mixer mix_t0_0101100000 (.a(t0_01011000000), .b(t0_01011000001), .y(t0_0101100000));
wire t0_01011000000, t0_01011000001;
mixer mix_t0_01011000000 (.a(t0_010110000000), .b(t0_010110000001), .y(t0_01011000000));
wire t0_010110000000, t0_010110000001;
mixer mix_t0_01011000001 (.a(t0_010110000010), .b(t0_010110000011), .y(t0_01011000001));
wire t0_010110000010, t0_010110000011;
mixer mix_t0_0101100001 (.a(t0_01011000010), .b(t0_01011000011), .y(t0_0101100001));
wire t0_01011000010, t0_01011000011;
mixer mix_t0_01011000010 (.a(t0_010110000100), .b(t0_010110000101), .y(t0_01011000010));
wire t0_010110000100, t0_010110000101;
mixer mix_t0_01011000011 (.a(t0_010110000110), .b(t0_010110000111), .y(t0_01011000011));
wire t0_010110000110, t0_010110000111;
mixer mix_t0_010110001 (.a(t0_0101100010), .b(t0_0101100011), .y(t0_010110001));
wire t0_0101100010, t0_0101100011;
mixer mix_t0_0101100010 (.a(t0_01011000100), .b(t0_01011000101), .y(t0_0101100010));
wire t0_01011000100, t0_01011000101;
mixer mix_t0_01011000100 (.a(t0_010110001000), .b(t0_010110001001), .y(t0_01011000100));
wire t0_010110001000, t0_010110001001;
mixer mix_t0_01011000101 (.a(t0_010110001010), .b(t0_010110001011), .y(t0_01011000101));
wire t0_010110001010, t0_010110001011;
mixer mix_t0_0101100011 (.a(t0_01011000110), .b(t0_01011000111), .y(t0_0101100011));
wire t0_01011000110, t0_01011000111;
mixer mix_t0_01011000110 (.a(t0_010110001100), .b(t0_010110001101), .y(t0_01011000110));
wire t0_010110001100, t0_010110001101;
mixer mix_t0_01011000111 (.a(t0_010110001110), .b(t0_010110001111), .y(t0_01011000111));
wire t0_010110001110, t0_010110001111;
mixer mix_t0_01011001 (.a(t0_010110010), .b(t0_010110011), .y(t0_01011001));
wire t0_010110010, t0_010110011;
mixer mix_t0_010110010 (.a(t0_0101100100), .b(t0_0101100101), .y(t0_010110010));
wire t0_0101100100, t0_0101100101;
mixer mix_t0_0101100100 (.a(t0_01011001000), .b(t0_01011001001), .y(t0_0101100100));
wire t0_01011001000, t0_01011001001;
mixer mix_t0_01011001000 (.a(t0_010110010000), .b(t0_010110010001), .y(t0_01011001000));
wire t0_010110010000, t0_010110010001;
mixer mix_t0_01011001001 (.a(t0_010110010010), .b(t0_010110010011), .y(t0_01011001001));
wire t0_010110010010, t0_010110010011;
mixer mix_t0_0101100101 (.a(t0_01011001010), .b(t0_01011001011), .y(t0_0101100101));
wire t0_01011001010, t0_01011001011;
mixer mix_t0_01011001010 (.a(t0_010110010100), .b(t0_010110010101), .y(t0_01011001010));
wire t0_010110010100, t0_010110010101;
mixer mix_t0_01011001011 (.a(t0_010110010110), .b(t0_010110010111), .y(t0_01011001011));
wire t0_010110010110, t0_010110010111;
mixer mix_t0_010110011 (.a(t0_0101100110), .b(t0_0101100111), .y(t0_010110011));
wire t0_0101100110, t0_0101100111;
mixer mix_t0_0101100110 (.a(t0_01011001100), .b(t0_01011001101), .y(t0_0101100110));
wire t0_01011001100, t0_01011001101;
mixer mix_t0_01011001100 (.a(t0_010110011000), .b(t0_010110011001), .y(t0_01011001100));
wire t0_010110011000, t0_010110011001;
mixer mix_t0_01011001101 (.a(t0_010110011010), .b(t0_010110011011), .y(t0_01011001101));
wire t0_010110011010, t0_010110011011;
mixer mix_t0_0101100111 (.a(t0_01011001110), .b(t0_01011001111), .y(t0_0101100111));
wire t0_01011001110, t0_01011001111;
mixer mix_t0_01011001110 (.a(t0_010110011100), .b(t0_010110011101), .y(t0_01011001110));
wire t0_010110011100, t0_010110011101;
mixer mix_t0_01011001111 (.a(t0_010110011110), .b(t0_010110011111), .y(t0_01011001111));
wire t0_010110011110, t0_010110011111;
mixer mix_t0_0101101 (.a(t0_01011010), .b(t0_01011011), .y(t0_0101101));
wire t0_01011010, t0_01011011;
mixer mix_t0_01011010 (.a(t0_010110100), .b(t0_010110101), .y(t0_01011010));
wire t0_010110100, t0_010110101;
mixer mix_t0_010110100 (.a(t0_0101101000), .b(t0_0101101001), .y(t0_010110100));
wire t0_0101101000, t0_0101101001;
mixer mix_t0_0101101000 (.a(t0_01011010000), .b(t0_01011010001), .y(t0_0101101000));
wire t0_01011010000, t0_01011010001;
mixer mix_t0_01011010000 (.a(t0_010110100000), .b(t0_010110100001), .y(t0_01011010000));
wire t0_010110100000, t0_010110100001;
mixer mix_t0_01011010001 (.a(t0_010110100010), .b(t0_010110100011), .y(t0_01011010001));
wire t0_010110100010, t0_010110100011;
mixer mix_t0_0101101001 (.a(t0_01011010010), .b(t0_01011010011), .y(t0_0101101001));
wire t0_01011010010, t0_01011010011;
mixer mix_t0_01011010010 (.a(t0_010110100100), .b(t0_010110100101), .y(t0_01011010010));
wire t0_010110100100, t0_010110100101;
mixer mix_t0_01011010011 (.a(t0_010110100110), .b(t0_010110100111), .y(t0_01011010011));
wire t0_010110100110, t0_010110100111;
mixer mix_t0_010110101 (.a(t0_0101101010), .b(t0_0101101011), .y(t0_010110101));
wire t0_0101101010, t0_0101101011;
mixer mix_t0_0101101010 (.a(t0_01011010100), .b(t0_01011010101), .y(t0_0101101010));
wire t0_01011010100, t0_01011010101;
mixer mix_t0_01011010100 (.a(t0_010110101000), .b(t0_010110101001), .y(t0_01011010100));
wire t0_010110101000, t0_010110101001;
mixer mix_t0_01011010101 (.a(t0_010110101010), .b(t0_010110101011), .y(t0_01011010101));
wire t0_010110101010, t0_010110101011;
mixer mix_t0_0101101011 (.a(t0_01011010110), .b(t0_01011010111), .y(t0_0101101011));
wire t0_01011010110, t0_01011010111;
mixer mix_t0_01011010110 (.a(t0_010110101100), .b(t0_010110101101), .y(t0_01011010110));
wire t0_010110101100, t0_010110101101;
mixer mix_t0_01011010111 (.a(t0_010110101110), .b(t0_010110101111), .y(t0_01011010111));
wire t0_010110101110, t0_010110101111;
mixer mix_t0_01011011 (.a(t0_010110110), .b(t0_010110111), .y(t0_01011011));
wire t0_010110110, t0_010110111;
mixer mix_t0_010110110 (.a(t0_0101101100), .b(t0_0101101101), .y(t0_010110110));
wire t0_0101101100, t0_0101101101;
mixer mix_t0_0101101100 (.a(t0_01011011000), .b(t0_01011011001), .y(t0_0101101100));
wire t0_01011011000, t0_01011011001;
mixer mix_t0_01011011000 (.a(t0_010110110000), .b(t0_010110110001), .y(t0_01011011000));
wire t0_010110110000, t0_010110110001;
mixer mix_t0_01011011001 (.a(t0_010110110010), .b(t0_010110110011), .y(t0_01011011001));
wire t0_010110110010, t0_010110110011;
mixer mix_t0_0101101101 (.a(t0_01011011010), .b(t0_01011011011), .y(t0_0101101101));
wire t0_01011011010, t0_01011011011;
mixer mix_t0_01011011010 (.a(t0_010110110100), .b(t0_010110110101), .y(t0_01011011010));
wire t0_010110110100, t0_010110110101;
mixer mix_t0_01011011011 (.a(t0_010110110110), .b(t0_010110110111), .y(t0_01011011011));
wire t0_010110110110, t0_010110110111;
mixer mix_t0_010110111 (.a(t0_0101101110), .b(t0_0101101111), .y(t0_010110111));
wire t0_0101101110, t0_0101101111;
mixer mix_t0_0101101110 (.a(t0_01011011100), .b(t0_01011011101), .y(t0_0101101110));
wire t0_01011011100, t0_01011011101;
mixer mix_t0_01011011100 (.a(t0_010110111000), .b(t0_010110111001), .y(t0_01011011100));
wire t0_010110111000, t0_010110111001;
mixer mix_t0_01011011101 (.a(t0_010110111010), .b(t0_010110111011), .y(t0_01011011101));
wire t0_010110111010, t0_010110111011;
mixer mix_t0_0101101111 (.a(t0_01011011110), .b(t0_01011011111), .y(t0_0101101111));
wire t0_01011011110, t0_01011011111;
mixer mix_t0_01011011110 (.a(t0_010110111100), .b(t0_010110111101), .y(t0_01011011110));
wire t0_010110111100, t0_010110111101;
mixer mix_t0_01011011111 (.a(t0_010110111110), .b(t0_010110111111), .y(t0_01011011111));
wire t0_010110111110, t0_010110111111;
mixer mix_t0_010111 (.a(t0_0101110), .b(t0_0101111), .y(t0_010111));
wire t0_0101110, t0_0101111;
mixer mix_t0_0101110 (.a(t0_01011100), .b(t0_01011101), .y(t0_0101110));
wire t0_01011100, t0_01011101;
mixer mix_t0_01011100 (.a(t0_010111000), .b(t0_010111001), .y(t0_01011100));
wire t0_010111000, t0_010111001;
mixer mix_t0_010111000 (.a(t0_0101110000), .b(t0_0101110001), .y(t0_010111000));
wire t0_0101110000, t0_0101110001;
mixer mix_t0_0101110000 (.a(t0_01011100000), .b(t0_01011100001), .y(t0_0101110000));
wire t0_01011100000, t0_01011100001;
mixer mix_t0_01011100000 (.a(t0_010111000000), .b(t0_010111000001), .y(t0_01011100000));
wire t0_010111000000, t0_010111000001;
mixer mix_t0_01011100001 (.a(t0_010111000010), .b(t0_010111000011), .y(t0_01011100001));
wire t0_010111000010, t0_010111000011;
mixer mix_t0_0101110001 (.a(t0_01011100010), .b(t0_01011100011), .y(t0_0101110001));
wire t0_01011100010, t0_01011100011;
mixer mix_t0_01011100010 (.a(t0_010111000100), .b(t0_010111000101), .y(t0_01011100010));
wire t0_010111000100, t0_010111000101;
mixer mix_t0_01011100011 (.a(t0_010111000110), .b(t0_010111000111), .y(t0_01011100011));
wire t0_010111000110, t0_010111000111;
mixer mix_t0_010111001 (.a(t0_0101110010), .b(t0_0101110011), .y(t0_010111001));
wire t0_0101110010, t0_0101110011;
mixer mix_t0_0101110010 (.a(t0_01011100100), .b(t0_01011100101), .y(t0_0101110010));
wire t0_01011100100, t0_01011100101;
mixer mix_t0_01011100100 (.a(t0_010111001000), .b(t0_010111001001), .y(t0_01011100100));
wire t0_010111001000, t0_010111001001;
mixer mix_t0_01011100101 (.a(t0_010111001010), .b(t0_010111001011), .y(t0_01011100101));
wire t0_010111001010, t0_010111001011;
mixer mix_t0_0101110011 (.a(t0_01011100110), .b(t0_01011100111), .y(t0_0101110011));
wire t0_01011100110, t0_01011100111;
mixer mix_t0_01011100110 (.a(t0_010111001100), .b(t0_010111001101), .y(t0_01011100110));
wire t0_010111001100, t0_010111001101;
mixer mix_t0_01011100111 (.a(t0_010111001110), .b(t0_010111001111), .y(t0_01011100111));
wire t0_010111001110, t0_010111001111;
mixer mix_t0_01011101 (.a(t0_010111010), .b(t0_010111011), .y(t0_01011101));
wire t0_010111010, t0_010111011;
mixer mix_t0_010111010 (.a(t0_0101110100), .b(t0_0101110101), .y(t0_010111010));
wire t0_0101110100, t0_0101110101;
mixer mix_t0_0101110100 (.a(t0_01011101000), .b(t0_01011101001), .y(t0_0101110100));
wire t0_01011101000, t0_01011101001;
mixer mix_t0_01011101000 (.a(t0_010111010000), .b(t0_010111010001), .y(t0_01011101000));
wire t0_010111010000, t0_010111010001;
mixer mix_t0_01011101001 (.a(t0_010111010010), .b(t0_010111010011), .y(t0_01011101001));
wire t0_010111010010, t0_010111010011;
mixer mix_t0_0101110101 (.a(t0_01011101010), .b(t0_01011101011), .y(t0_0101110101));
wire t0_01011101010, t0_01011101011;
mixer mix_t0_01011101010 (.a(t0_010111010100), .b(t0_010111010101), .y(t0_01011101010));
wire t0_010111010100, t0_010111010101;
mixer mix_t0_01011101011 (.a(t0_010111010110), .b(t0_010111010111), .y(t0_01011101011));
wire t0_010111010110, t0_010111010111;
mixer mix_t0_010111011 (.a(t0_0101110110), .b(t0_0101110111), .y(t0_010111011));
wire t0_0101110110, t0_0101110111;
mixer mix_t0_0101110110 (.a(t0_01011101100), .b(t0_01011101101), .y(t0_0101110110));
wire t0_01011101100, t0_01011101101;
mixer mix_t0_01011101100 (.a(t0_010111011000), .b(t0_010111011001), .y(t0_01011101100));
wire t0_010111011000, t0_010111011001;
mixer mix_t0_01011101101 (.a(t0_010111011010), .b(t0_010111011011), .y(t0_01011101101));
wire t0_010111011010, t0_010111011011;
mixer mix_t0_0101110111 (.a(t0_01011101110), .b(t0_01011101111), .y(t0_0101110111));
wire t0_01011101110, t0_01011101111;
mixer mix_t0_01011101110 (.a(t0_010111011100), .b(t0_010111011101), .y(t0_01011101110));
wire t0_010111011100, t0_010111011101;
mixer mix_t0_01011101111 (.a(t0_010111011110), .b(t0_010111011111), .y(t0_01011101111));
wire t0_010111011110, t0_010111011111;
mixer mix_t0_0101111 (.a(t0_01011110), .b(t0_01011111), .y(t0_0101111));
wire t0_01011110, t0_01011111;
mixer mix_t0_01011110 (.a(t0_010111100), .b(t0_010111101), .y(t0_01011110));
wire t0_010111100, t0_010111101;
mixer mix_t0_010111100 (.a(t0_0101111000), .b(t0_0101111001), .y(t0_010111100));
wire t0_0101111000, t0_0101111001;
mixer mix_t0_0101111000 (.a(t0_01011110000), .b(t0_01011110001), .y(t0_0101111000));
wire t0_01011110000, t0_01011110001;
mixer mix_t0_01011110000 (.a(t0_010111100000), .b(t0_010111100001), .y(t0_01011110000));
wire t0_010111100000, t0_010111100001;
mixer mix_t0_01011110001 (.a(t0_010111100010), .b(t0_010111100011), .y(t0_01011110001));
wire t0_010111100010, t0_010111100011;
mixer mix_t0_0101111001 (.a(t0_01011110010), .b(t0_01011110011), .y(t0_0101111001));
wire t0_01011110010, t0_01011110011;
mixer mix_t0_01011110010 (.a(t0_010111100100), .b(t0_010111100101), .y(t0_01011110010));
wire t0_010111100100, t0_010111100101;
mixer mix_t0_01011110011 (.a(t0_010111100110), .b(t0_010111100111), .y(t0_01011110011));
wire t0_010111100110, t0_010111100111;
mixer mix_t0_010111101 (.a(t0_0101111010), .b(t0_0101111011), .y(t0_010111101));
wire t0_0101111010, t0_0101111011;
mixer mix_t0_0101111010 (.a(t0_01011110100), .b(t0_01011110101), .y(t0_0101111010));
wire t0_01011110100, t0_01011110101;
mixer mix_t0_01011110100 (.a(t0_010111101000), .b(t0_010111101001), .y(t0_01011110100));
wire t0_010111101000, t0_010111101001;
mixer mix_t0_01011110101 (.a(t0_010111101010), .b(t0_010111101011), .y(t0_01011110101));
wire t0_010111101010, t0_010111101011;
mixer mix_t0_0101111011 (.a(t0_01011110110), .b(t0_01011110111), .y(t0_0101111011));
wire t0_01011110110, t0_01011110111;
mixer mix_t0_01011110110 (.a(t0_010111101100), .b(t0_010111101101), .y(t0_01011110110));
wire t0_010111101100, t0_010111101101;
mixer mix_t0_01011110111 (.a(t0_010111101110), .b(t0_010111101111), .y(t0_01011110111));
wire t0_010111101110, t0_010111101111;
mixer mix_t0_01011111 (.a(t0_010111110), .b(t0_010111111), .y(t0_01011111));
wire t0_010111110, t0_010111111;
mixer mix_t0_010111110 (.a(t0_0101111100), .b(t0_0101111101), .y(t0_010111110));
wire t0_0101111100, t0_0101111101;
mixer mix_t0_0101111100 (.a(t0_01011111000), .b(t0_01011111001), .y(t0_0101111100));
wire t0_01011111000, t0_01011111001;
mixer mix_t0_01011111000 (.a(t0_010111110000), .b(t0_010111110001), .y(t0_01011111000));
wire t0_010111110000, t0_010111110001;
mixer mix_t0_01011111001 (.a(t0_010111110010), .b(t0_010111110011), .y(t0_01011111001));
wire t0_010111110010, t0_010111110011;
mixer mix_t0_0101111101 (.a(t0_01011111010), .b(t0_01011111011), .y(t0_0101111101));
wire t0_01011111010, t0_01011111011;
mixer mix_t0_01011111010 (.a(t0_010111110100), .b(t0_010111110101), .y(t0_01011111010));
wire t0_010111110100, t0_010111110101;
mixer mix_t0_01011111011 (.a(t0_010111110110), .b(t0_010111110111), .y(t0_01011111011));
wire t0_010111110110, t0_010111110111;
mixer mix_t0_010111111 (.a(t0_0101111110), .b(t0_0101111111), .y(t0_010111111));
wire t0_0101111110, t0_0101111111;
mixer mix_t0_0101111110 (.a(t0_01011111100), .b(t0_01011111101), .y(t0_0101111110));
wire t0_01011111100, t0_01011111101;
mixer mix_t0_01011111100 (.a(t0_010111111000), .b(t0_010111111001), .y(t0_01011111100));
wire t0_010111111000, t0_010111111001;
mixer mix_t0_01011111101 (.a(t0_010111111010), .b(t0_010111111011), .y(t0_01011111101));
wire t0_010111111010, t0_010111111011;
mixer mix_t0_0101111111 (.a(t0_01011111110), .b(t0_01011111111), .y(t0_0101111111));
wire t0_01011111110, t0_01011111111;
mixer mix_t0_01011111110 (.a(t0_010111111100), .b(t0_010111111101), .y(t0_01011111110));
wire t0_010111111100, t0_010111111101;
mixer mix_t0_01011111111 (.a(t0_010111111110), .b(t0_010111111111), .y(t0_01011111111));
wire t0_010111111110, t0_010111111111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_011000 (.a(t0_0110000), .b(t0_0110001), .y(t0_011000));
wire t0_0110000, t0_0110001;
mixer mix_t0_0110000 (.a(t0_01100000), .b(t0_01100001), .y(t0_0110000));
wire t0_01100000, t0_01100001;
mixer mix_t0_01100000 (.a(t0_011000000), .b(t0_011000001), .y(t0_01100000));
wire t0_011000000, t0_011000001;
mixer mix_t0_011000000 (.a(t0_0110000000), .b(t0_0110000001), .y(t0_011000000));
wire t0_0110000000, t0_0110000001;
mixer mix_t0_0110000000 (.a(t0_01100000000), .b(t0_01100000001), .y(t0_0110000000));
wire t0_01100000000, t0_01100000001;
mixer mix_t0_01100000000 (.a(t0_011000000000), .b(t0_011000000001), .y(t0_01100000000));
wire t0_011000000000, t0_011000000001;
mixer mix_t0_01100000001 (.a(t0_011000000010), .b(t0_011000000011), .y(t0_01100000001));
wire t0_011000000010, t0_011000000011;
mixer mix_t0_0110000001 (.a(t0_01100000010), .b(t0_01100000011), .y(t0_0110000001));
wire t0_01100000010, t0_01100000011;
mixer mix_t0_01100000010 (.a(t0_011000000100), .b(t0_011000000101), .y(t0_01100000010));
wire t0_011000000100, t0_011000000101;
mixer mix_t0_01100000011 (.a(t0_011000000110), .b(t0_011000000111), .y(t0_01100000011));
wire t0_011000000110, t0_011000000111;
mixer mix_t0_011000001 (.a(t0_0110000010), .b(t0_0110000011), .y(t0_011000001));
wire t0_0110000010, t0_0110000011;
mixer mix_t0_0110000010 (.a(t0_01100000100), .b(t0_01100000101), .y(t0_0110000010));
wire t0_01100000100, t0_01100000101;
mixer mix_t0_01100000100 (.a(t0_011000001000), .b(t0_011000001001), .y(t0_01100000100));
wire t0_011000001000, t0_011000001001;
mixer mix_t0_01100000101 (.a(t0_011000001010), .b(t0_011000001011), .y(t0_01100000101));
wire t0_011000001010, t0_011000001011;
mixer mix_t0_0110000011 (.a(t0_01100000110), .b(t0_01100000111), .y(t0_0110000011));
wire t0_01100000110, t0_01100000111;
mixer mix_t0_01100000110 (.a(t0_011000001100), .b(t0_011000001101), .y(t0_01100000110));
wire t0_011000001100, t0_011000001101;
mixer mix_t0_01100000111 (.a(t0_011000001110), .b(t0_011000001111), .y(t0_01100000111));
wire t0_011000001110, t0_011000001111;
mixer mix_t0_01100001 (.a(t0_011000010), .b(t0_011000011), .y(t0_01100001));
wire t0_011000010, t0_011000011;
mixer mix_t0_011000010 (.a(t0_0110000100), .b(t0_0110000101), .y(t0_011000010));
wire t0_0110000100, t0_0110000101;
mixer mix_t0_0110000100 (.a(t0_01100001000), .b(t0_01100001001), .y(t0_0110000100));
wire t0_01100001000, t0_01100001001;
mixer mix_t0_01100001000 (.a(t0_011000010000), .b(t0_011000010001), .y(t0_01100001000));
wire t0_011000010000, t0_011000010001;
mixer mix_t0_01100001001 (.a(t0_011000010010), .b(t0_011000010011), .y(t0_01100001001));
wire t0_011000010010, t0_011000010011;
mixer mix_t0_0110000101 (.a(t0_01100001010), .b(t0_01100001011), .y(t0_0110000101));
wire t0_01100001010, t0_01100001011;
mixer mix_t0_01100001010 (.a(t0_011000010100), .b(t0_011000010101), .y(t0_01100001010));
wire t0_011000010100, t0_011000010101;
mixer mix_t0_01100001011 (.a(t0_011000010110), .b(t0_011000010111), .y(t0_01100001011));
wire t0_011000010110, t0_011000010111;
mixer mix_t0_011000011 (.a(t0_0110000110), .b(t0_0110000111), .y(t0_011000011));
wire t0_0110000110, t0_0110000111;
mixer mix_t0_0110000110 (.a(t0_01100001100), .b(t0_01100001101), .y(t0_0110000110));
wire t0_01100001100, t0_01100001101;
mixer mix_t0_01100001100 (.a(t0_011000011000), .b(t0_011000011001), .y(t0_01100001100));
wire t0_011000011000, t0_011000011001;
mixer mix_t0_01100001101 (.a(t0_011000011010), .b(t0_011000011011), .y(t0_01100001101));
wire t0_011000011010, t0_011000011011;
mixer mix_t0_0110000111 (.a(t0_01100001110), .b(t0_01100001111), .y(t0_0110000111));
wire t0_01100001110, t0_01100001111;
mixer mix_t0_01100001110 (.a(t0_011000011100), .b(t0_011000011101), .y(t0_01100001110));
wire t0_011000011100, t0_011000011101;
mixer mix_t0_01100001111 (.a(t0_011000011110), .b(t0_011000011111), .y(t0_01100001111));
wire t0_011000011110, t0_011000011111;
mixer mix_t0_0110001 (.a(t0_01100010), .b(t0_01100011), .y(t0_0110001));
wire t0_01100010, t0_01100011;
mixer mix_t0_01100010 (.a(t0_011000100), .b(t0_011000101), .y(t0_01100010));
wire t0_011000100, t0_011000101;
mixer mix_t0_011000100 (.a(t0_0110001000), .b(t0_0110001001), .y(t0_011000100));
wire t0_0110001000, t0_0110001001;
mixer mix_t0_0110001000 (.a(t0_01100010000), .b(t0_01100010001), .y(t0_0110001000));
wire t0_01100010000, t0_01100010001;
mixer mix_t0_01100010000 (.a(t0_011000100000), .b(t0_011000100001), .y(t0_01100010000));
wire t0_011000100000, t0_011000100001;
mixer mix_t0_01100010001 (.a(t0_011000100010), .b(t0_011000100011), .y(t0_01100010001));
wire t0_011000100010, t0_011000100011;
mixer mix_t0_0110001001 (.a(t0_01100010010), .b(t0_01100010011), .y(t0_0110001001));
wire t0_01100010010, t0_01100010011;
mixer mix_t0_01100010010 (.a(t0_011000100100), .b(t0_011000100101), .y(t0_01100010010));
wire t0_011000100100, t0_011000100101;
mixer mix_t0_01100010011 (.a(t0_011000100110), .b(t0_011000100111), .y(t0_01100010011));
wire t0_011000100110, t0_011000100111;
mixer mix_t0_011000101 (.a(t0_0110001010), .b(t0_0110001011), .y(t0_011000101));
wire t0_0110001010, t0_0110001011;
mixer mix_t0_0110001010 (.a(t0_01100010100), .b(t0_01100010101), .y(t0_0110001010));
wire t0_01100010100, t0_01100010101;
mixer mix_t0_01100010100 (.a(t0_011000101000), .b(t0_011000101001), .y(t0_01100010100));
wire t0_011000101000, t0_011000101001;
mixer mix_t0_01100010101 (.a(t0_011000101010), .b(t0_011000101011), .y(t0_01100010101));
wire t0_011000101010, t0_011000101011;
mixer mix_t0_0110001011 (.a(t0_01100010110), .b(t0_01100010111), .y(t0_0110001011));
wire t0_01100010110, t0_01100010111;
mixer mix_t0_01100010110 (.a(t0_011000101100), .b(t0_011000101101), .y(t0_01100010110));
wire t0_011000101100, t0_011000101101;
mixer mix_t0_01100010111 (.a(t0_011000101110), .b(t0_011000101111), .y(t0_01100010111));
wire t0_011000101110, t0_011000101111;
mixer mix_t0_01100011 (.a(t0_011000110), .b(t0_011000111), .y(t0_01100011));
wire t0_011000110, t0_011000111;
mixer mix_t0_011000110 (.a(t0_0110001100), .b(t0_0110001101), .y(t0_011000110));
wire t0_0110001100, t0_0110001101;
mixer mix_t0_0110001100 (.a(t0_01100011000), .b(t0_01100011001), .y(t0_0110001100));
wire t0_01100011000, t0_01100011001;
mixer mix_t0_01100011000 (.a(t0_011000110000), .b(t0_011000110001), .y(t0_01100011000));
wire t0_011000110000, t0_011000110001;
mixer mix_t0_01100011001 (.a(t0_011000110010), .b(t0_011000110011), .y(t0_01100011001));
wire t0_011000110010, t0_011000110011;
mixer mix_t0_0110001101 (.a(t0_01100011010), .b(t0_01100011011), .y(t0_0110001101));
wire t0_01100011010, t0_01100011011;
mixer mix_t0_01100011010 (.a(t0_011000110100), .b(t0_011000110101), .y(t0_01100011010));
wire t0_011000110100, t0_011000110101;
mixer mix_t0_01100011011 (.a(t0_011000110110), .b(t0_011000110111), .y(t0_01100011011));
wire t0_011000110110, t0_011000110111;
mixer mix_t0_011000111 (.a(t0_0110001110), .b(t0_0110001111), .y(t0_011000111));
wire t0_0110001110, t0_0110001111;
mixer mix_t0_0110001110 (.a(t0_01100011100), .b(t0_01100011101), .y(t0_0110001110));
wire t0_01100011100, t0_01100011101;
mixer mix_t0_01100011100 (.a(t0_011000111000), .b(t0_011000111001), .y(t0_01100011100));
wire t0_011000111000, t0_011000111001;
mixer mix_t0_01100011101 (.a(t0_011000111010), .b(t0_011000111011), .y(t0_01100011101));
wire t0_011000111010, t0_011000111011;
mixer mix_t0_0110001111 (.a(t0_01100011110), .b(t0_01100011111), .y(t0_0110001111));
wire t0_01100011110, t0_01100011111;
mixer mix_t0_01100011110 (.a(t0_011000111100), .b(t0_011000111101), .y(t0_01100011110));
wire t0_011000111100, t0_011000111101;
mixer mix_t0_01100011111 (.a(t0_011000111110), .b(t0_011000111111), .y(t0_01100011111));
wire t0_011000111110, t0_011000111111;
mixer mix_t0_011001 (.a(t0_0110010), .b(t0_0110011), .y(t0_011001));
wire t0_0110010, t0_0110011;
mixer mix_t0_0110010 (.a(t0_01100100), .b(t0_01100101), .y(t0_0110010));
wire t0_01100100, t0_01100101;
mixer mix_t0_01100100 (.a(t0_011001000), .b(t0_011001001), .y(t0_01100100));
wire t0_011001000, t0_011001001;
mixer mix_t0_011001000 (.a(t0_0110010000), .b(t0_0110010001), .y(t0_011001000));
wire t0_0110010000, t0_0110010001;
mixer mix_t0_0110010000 (.a(t0_01100100000), .b(t0_01100100001), .y(t0_0110010000));
wire t0_01100100000, t0_01100100001;
mixer mix_t0_01100100000 (.a(t0_011001000000), .b(t0_011001000001), .y(t0_01100100000));
wire t0_011001000000, t0_011001000001;
mixer mix_t0_01100100001 (.a(t0_011001000010), .b(t0_011001000011), .y(t0_01100100001));
wire t0_011001000010, t0_011001000011;
mixer mix_t0_0110010001 (.a(t0_01100100010), .b(t0_01100100011), .y(t0_0110010001));
wire t0_01100100010, t0_01100100011;
mixer mix_t0_01100100010 (.a(t0_011001000100), .b(t0_011001000101), .y(t0_01100100010));
wire t0_011001000100, t0_011001000101;
mixer mix_t0_01100100011 (.a(t0_011001000110), .b(t0_011001000111), .y(t0_01100100011));
wire t0_011001000110, t0_011001000111;
mixer mix_t0_011001001 (.a(t0_0110010010), .b(t0_0110010011), .y(t0_011001001));
wire t0_0110010010, t0_0110010011;
mixer mix_t0_0110010010 (.a(t0_01100100100), .b(t0_01100100101), .y(t0_0110010010));
wire t0_01100100100, t0_01100100101;
mixer mix_t0_01100100100 (.a(t0_011001001000), .b(t0_011001001001), .y(t0_01100100100));
wire t0_011001001000, t0_011001001001;
mixer mix_t0_01100100101 (.a(t0_011001001010), .b(t0_011001001011), .y(t0_01100100101));
wire t0_011001001010, t0_011001001011;
mixer mix_t0_0110010011 (.a(t0_01100100110), .b(t0_01100100111), .y(t0_0110010011));
wire t0_01100100110, t0_01100100111;
mixer mix_t0_01100100110 (.a(t0_011001001100), .b(t0_011001001101), .y(t0_01100100110));
wire t0_011001001100, t0_011001001101;
mixer mix_t0_01100100111 (.a(t0_011001001110), .b(t0_011001001111), .y(t0_01100100111));
wire t0_011001001110, t0_011001001111;
mixer mix_t0_01100101 (.a(t0_011001010), .b(t0_011001011), .y(t0_01100101));
wire t0_011001010, t0_011001011;
mixer mix_t0_011001010 (.a(t0_0110010100), .b(t0_0110010101), .y(t0_011001010));
wire t0_0110010100, t0_0110010101;
mixer mix_t0_0110010100 (.a(t0_01100101000), .b(t0_01100101001), .y(t0_0110010100));
wire t0_01100101000, t0_01100101001;
mixer mix_t0_01100101000 (.a(t0_011001010000), .b(t0_011001010001), .y(t0_01100101000));
wire t0_011001010000, t0_011001010001;
mixer mix_t0_01100101001 (.a(t0_011001010010), .b(t0_011001010011), .y(t0_01100101001));
wire t0_011001010010, t0_011001010011;
mixer mix_t0_0110010101 (.a(t0_01100101010), .b(t0_01100101011), .y(t0_0110010101));
wire t0_01100101010, t0_01100101011;
mixer mix_t0_01100101010 (.a(t0_011001010100), .b(t0_011001010101), .y(t0_01100101010));
wire t0_011001010100, t0_011001010101;
mixer mix_t0_01100101011 (.a(t0_011001010110), .b(t0_011001010111), .y(t0_01100101011));
wire t0_011001010110, t0_011001010111;
mixer mix_t0_011001011 (.a(t0_0110010110), .b(t0_0110010111), .y(t0_011001011));
wire t0_0110010110, t0_0110010111;
mixer mix_t0_0110010110 (.a(t0_01100101100), .b(t0_01100101101), .y(t0_0110010110));
wire t0_01100101100, t0_01100101101;
mixer mix_t0_01100101100 (.a(t0_011001011000), .b(t0_011001011001), .y(t0_01100101100));
wire t0_011001011000, t0_011001011001;
mixer mix_t0_01100101101 (.a(t0_011001011010), .b(t0_011001011011), .y(t0_01100101101));
wire t0_011001011010, t0_011001011011;
mixer mix_t0_0110010111 (.a(t0_01100101110), .b(t0_01100101111), .y(t0_0110010111));
wire t0_01100101110, t0_01100101111;
mixer mix_t0_01100101110 (.a(t0_011001011100), .b(t0_011001011101), .y(t0_01100101110));
wire t0_011001011100, t0_011001011101;
mixer mix_t0_01100101111 (.a(t0_011001011110), .b(t0_011001011111), .y(t0_01100101111));
wire t0_011001011110, t0_011001011111;
mixer mix_t0_0110011 (.a(t0_01100110), .b(t0_01100111), .y(t0_0110011));
wire t0_01100110, t0_01100111;
mixer mix_t0_01100110 (.a(t0_011001100), .b(t0_011001101), .y(t0_01100110));
wire t0_011001100, t0_011001101;
mixer mix_t0_011001100 (.a(t0_0110011000), .b(t0_0110011001), .y(t0_011001100));
wire t0_0110011000, t0_0110011001;
mixer mix_t0_0110011000 (.a(t0_01100110000), .b(t0_01100110001), .y(t0_0110011000));
wire t0_01100110000, t0_01100110001;
mixer mix_t0_01100110000 (.a(t0_011001100000), .b(t0_011001100001), .y(t0_01100110000));
wire t0_011001100000, t0_011001100001;
mixer mix_t0_01100110001 (.a(t0_011001100010), .b(t0_011001100011), .y(t0_01100110001));
wire t0_011001100010, t0_011001100011;
mixer mix_t0_0110011001 (.a(t0_01100110010), .b(t0_01100110011), .y(t0_0110011001));
wire t0_01100110010, t0_01100110011;
mixer mix_t0_01100110010 (.a(t0_011001100100), .b(t0_011001100101), .y(t0_01100110010));
wire t0_011001100100, t0_011001100101;
mixer mix_t0_01100110011 (.a(t0_011001100110), .b(t0_011001100111), .y(t0_01100110011));
wire t0_011001100110, t0_011001100111;
mixer mix_t0_011001101 (.a(t0_0110011010), .b(t0_0110011011), .y(t0_011001101));
wire t0_0110011010, t0_0110011011;
mixer mix_t0_0110011010 (.a(t0_01100110100), .b(t0_01100110101), .y(t0_0110011010));
wire t0_01100110100, t0_01100110101;
mixer mix_t0_01100110100 (.a(t0_011001101000), .b(t0_011001101001), .y(t0_01100110100));
wire t0_011001101000, t0_011001101001;
mixer mix_t0_01100110101 (.a(t0_011001101010), .b(t0_011001101011), .y(t0_01100110101));
wire t0_011001101010, t0_011001101011;
mixer mix_t0_0110011011 (.a(t0_01100110110), .b(t0_01100110111), .y(t0_0110011011));
wire t0_01100110110, t0_01100110111;
mixer mix_t0_01100110110 (.a(t0_011001101100), .b(t0_011001101101), .y(t0_01100110110));
wire t0_011001101100, t0_011001101101;
mixer mix_t0_01100110111 (.a(t0_011001101110), .b(t0_011001101111), .y(t0_01100110111));
wire t0_011001101110, t0_011001101111;
mixer mix_t0_01100111 (.a(t0_011001110), .b(t0_011001111), .y(t0_01100111));
wire t0_011001110, t0_011001111;
mixer mix_t0_011001110 (.a(t0_0110011100), .b(t0_0110011101), .y(t0_011001110));
wire t0_0110011100, t0_0110011101;
mixer mix_t0_0110011100 (.a(t0_01100111000), .b(t0_01100111001), .y(t0_0110011100));
wire t0_01100111000, t0_01100111001;
mixer mix_t0_01100111000 (.a(t0_011001110000), .b(t0_011001110001), .y(t0_01100111000));
wire t0_011001110000, t0_011001110001;
mixer mix_t0_01100111001 (.a(t0_011001110010), .b(t0_011001110011), .y(t0_01100111001));
wire t0_011001110010, t0_011001110011;
mixer mix_t0_0110011101 (.a(t0_01100111010), .b(t0_01100111011), .y(t0_0110011101));
wire t0_01100111010, t0_01100111011;
mixer mix_t0_01100111010 (.a(t0_011001110100), .b(t0_011001110101), .y(t0_01100111010));
wire t0_011001110100, t0_011001110101;
mixer mix_t0_01100111011 (.a(t0_011001110110), .b(t0_011001110111), .y(t0_01100111011));
wire t0_011001110110, t0_011001110111;
mixer mix_t0_011001111 (.a(t0_0110011110), .b(t0_0110011111), .y(t0_011001111));
wire t0_0110011110, t0_0110011111;
mixer mix_t0_0110011110 (.a(t0_01100111100), .b(t0_01100111101), .y(t0_0110011110));
wire t0_01100111100, t0_01100111101;
mixer mix_t0_01100111100 (.a(t0_011001111000), .b(t0_011001111001), .y(t0_01100111100));
wire t0_011001111000, t0_011001111001;
mixer mix_t0_01100111101 (.a(t0_011001111010), .b(t0_011001111011), .y(t0_01100111101));
wire t0_011001111010, t0_011001111011;
mixer mix_t0_0110011111 (.a(t0_01100111110), .b(t0_01100111111), .y(t0_0110011111));
wire t0_01100111110, t0_01100111111;
mixer mix_t0_01100111110 (.a(t0_011001111100), .b(t0_011001111101), .y(t0_01100111110));
wire t0_011001111100, t0_011001111101;
mixer mix_t0_01100111111 (.a(t0_011001111110), .b(t0_011001111111), .y(t0_01100111111));
wire t0_011001111110, t0_011001111111;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_011010 (.a(t0_0110100), .b(t0_0110101), .y(t0_011010));
wire t0_0110100, t0_0110101;
mixer mix_t0_0110100 (.a(t0_01101000), .b(t0_01101001), .y(t0_0110100));
wire t0_01101000, t0_01101001;
mixer mix_t0_01101000 (.a(t0_011010000), .b(t0_011010001), .y(t0_01101000));
wire t0_011010000, t0_011010001;
mixer mix_t0_011010000 (.a(t0_0110100000), .b(t0_0110100001), .y(t0_011010000));
wire t0_0110100000, t0_0110100001;
mixer mix_t0_0110100000 (.a(t0_01101000000), .b(t0_01101000001), .y(t0_0110100000));
wire t0_01101000000, t0_01101000001;
mixer mix_t0_01101000000 (.a(t0_011010000000), .b(t0_011010000001), .y(t0_01101000000));
wire t0_011010000000, t0_011010000001;
mixer mix_t0_01101000001 (.a(t0_011010000010), .b(t0_011010000011), .y(t0_01101000001));
wire t0_011010000010, t0_011010000011;
mixer mix_t0_0110100001 (.a(t0_01101000010), .b(t0_01101000011), .y(t0_0110100001));
wire t0_01101000010, t0_01101000011;
mixer mix_t0_01101000010 (.a(t0_011010000100), .b(t0_011010000101), .y(t0_01101000010));
wire t0_011010000100, t0_011010000101;
mixer mix_t0_01101000011 (.a(t0_011010000110), .b(t0_011010000111), .y(t0_01101000011));
wire t0_011010000110, t0_011010000111;
mixer mix_t0_011010001 (.a(t0_0110100010), .b(t0_0110100011), .y(t0_011010001));
wire t0_0110100010, t0_0110100011;
mixer mix_t0_0110100010 (.a(t0_01101000100), .b(t0_01101000101), .y(t0_0110100010));
wire t0_01101000100, t0_01101000101;
mixer mix_t0_01101000100 (.a(t0_011010001000), .b(t0_011010001001), .y(t0_01101000100));
wire t0_011010001000, t0_011010001001;
mixer mix_t0_01101000101 (.a(t0_011010001010), .b(t0_011010001011), .y(t0_01101000101));
wire t0_011010001010, t0_011010001011;
mixer mix_t0_0110100011 (.a(t0_01101000110), .b(t0_01101000111), .y(t0_0110100011));
wire t0_01101000110, t0_01101000111;
mixer mix_t0_01101000110 (.a(t0_011010001100), .b(t0_011010001101), .y(t0_01101000110));
wire t0_011010001100, t0_011010001101;
mixer mix_t0_01101000111 (.a(t0_011010001110), .b(t0_011010001111), .y(t0_01101000111));
wire t0_011010001110, t0_011010001111;
mixer mix_t0_01101001 (.a(t0_011010010), .b(t0_011010011), .y(t0_01101001));
wire t0_011010010, t0_011010011;
mixer mix_t0_011010010 (.a(t0_0110100100), .b(t0_0110100101), .y(t0_011010010));
wire t0_0110100100, t0_0110100101;
mixer mix_t0_0110100100 (.a(t0_01101001000), .b(t0_01101001001), .y(t0_0110100100));
wire t0_01101001000, t0_01101001001;
mixer mix_t0_01101001000 (.a(t0_011010010000), .b(t0_011010010001), .y(t0_01101001000));
wire t0_011010010000, t0_011010010001;
mixer mix_t0_01101001001 (.a(t0_011010010010), .b(t0_011010010011), .y(t0_01101001001));
wire t0_011010010010, t0_011010010011;
mixer mix_t0_0110100101 (.a(t0_01101001010), .b(t0_01101001011), .y(t0_0110100101));
wire t0_01101001010, t0_01101001011;
mixer mix_t0_01101001010 (.a(t0_011010010100), .b(t0_011010010101), .y(t0_01101001010));
wire t0_011010010100, t0_011010010101;
mixer mix_t0_01101001011 (.a(t0_011010010110), .b(t0_011010010111), .y(t0_01101001011));
wire t0_011010010110, t0_011010010111;
mixer mix_t0_011010011 (.a(t0_0110100110), .b(t0_0110100111), .y(t0_011010011));
wire t0_0110100110, t0_0110100111;
mixer mix_t0_0110100110 (.a(t0_01101001100), .b(t0_01101001101), .y(t0_0110100110));
wire t0_01101001100, t0_01101001101;
mixer mix_t0_01101001100 (.a(t0_011010011000), .b(t0_011010011001), .y(t0_01101001100));
wire t0_011010011000, t0_011010011001;
mixer mix_t0_01101001101 (.a(t0_011010011010), .b(t0_011010011011), .y(t0_01101001101));
wire t0_011010011010, t0_011010011011;
mixer mix_t0_0110100111 (.a(t0_01101001110), .b(t0_01101001111), .y(t0_0110100111));
wire t0_01101001110, t0_01101001111;
mixer mix_t0_01101001110 (.a(t0_011010011100), .b(t0_011010011101), .y(t0_01101001110));
wire t0_011010011100, t0_011010011101;
mixer mix_t0_01101001111 (.a(t0_011010011110), .b(t0_011010011111), .y(t0_01101001111));
wire t0_011010011110, t0_011010011111;
mixer mix_t0_0110101 (.a(t0_01101010), .b(t0_01101011), .y(t0_0110101));
wire t0_01101010, t0_01101011;
mixer mix_t0_01101010 (.a(t0_011010100), .b(t0_011010101), .y(t0_01101010));
wire t0_011010100, t0_011010101;
mixer mix_t0_011010100 (.a(t0_0110101000), .b(t0_0110101001), .y(t0_011010100));
wire t0_0110101000, t0_0110101001;
mixer mix_t0_0110101000 (.a(t0_01101010000), .b(t0_01101010001), .y(t0_0110101000));
wire t0_01101010000, t0_01101010001;
mixer mix_t0_01101010000 (.a(t0_011010100000), .b(t0_011010100001), .y(t0_01101010000));
wire t0_011010100000, t0_011010100001;
mixer mix_t0_01101010001 (.a(t0_011010100010), .b(t0_011010100011), .y(t0_01101010001));
wire t0_011010100010, t0_011010100011;
mixer mix_t0_0110101001 (.a(t0_01101010010), .b(t0_01101010011), .y(t0_0110101001));
wire t0_01101010010, t0_01101010011;
mixer mix_t0_01101010010 (.a(t0_011010100100), .b(t0_011010100101), .y(t0_01101010010));
wire t0_011010100100, t0_011010100101;
mixer mix_t0_01101010011 (.a(t0_011010100110), .b(t0_011010100111), .y(t0_01101010011));
wire t0_011010100110, t0_011010100111;
mixer mix_t0_011010101 (.a(t0_0110101010), .b(t0_0110101011), .y(t0_011010101));
wire t0_0110101010, t0_0110101011;
mixer mix_t0_0110101010 (.a(t0_01101010100), .b(t0_01101010101), .y(t0_0110101010));
wire t0_01101010100, t0_01101010101;
mixer mix_t0_01101010100 (.a(t0_011010101000), .b(t0_011010101001), .y(t0_01101010100));
wire t0_011010101000, t0_011010101001;
mixer mix_t0_01101010101 (.a(t0_011010101010), .b(t0_011010101011), .y(t0_01101010101));
wire t0_011010101010, t0_011010101011;
mixer mix_t0_0110101011 (.a(t0_01101010110), .b(t0_01101010111), .y(t0_0110101011));
wire t0_01101010110, t0_01101010111;
mixer mix_t0_01101010110 (.a(t0_011010101100), .b(t0_011010101101), .y(t0_01101010110));
wire t0_011010101100, t0_011010101101;
mixer mix_t0_01101010111 (.a(t0_011010101110), .b(t0_011010101111), .y(t0_01101010111));
wire t0_011010101110, t0_011010101111;
mixer mix_t0_01101011 (.a(t0_011010110), .b(t0_011010111), .y(t0_01101011));
wire t0_011010110, t0_011010111;
mixer mix_t0_011010110 (.a(t0_0110101100), .b(t0_0110101101), .y(t0_011010110));
wire t0_0110101100, t0_0110101101;
mixer mix_t0_0110101100 (.a(t0_01101011000), .b(t0_01101011001), .y(t0_0110101100));
wire t0_01101011000, t0_01101011001;
mixer mix_t0_01101011000 (.a(t0_011010110000), .b(t0_011010110001), .y(t0_01101011000));
wire t0_011010110000, t0_011010110001;
mixer mix_t0_01101011001 (.a(t0_011010110010), .b(t0_011010110011), .y(t0_01101011001));
wire t0_011010110010, t0_011010110011;
mixer mix_t0_0110101101 (.a(t0_01101011010), .b(t0_01101011011), .y(t0_0110101101));
wire t0_01101011010, t0_01101011011;
mixer mix_t0_01101011010 (.a(t0_011010110100), .b(t0_011010110101), .y(t0_01101011010));
wire t0_011010110100, t0_011010110101;
mixer mix_t0_01101011011 (.a(t0_011010110110), .b(t0_011010110111), .y(t0_01101011011));
wire t0_011010110110, t0_011010110111;
mixer mix_t0_011010111 (.a(t0_0110101110), .b(t0_0110101111), .y(t0_011010111));
wire t0_0110101110, t0_0110101111;
mixer mix_t0_0110101110 (.a(t0_01101011100), .b(t0_01101011101), .y(t0_0110101110));
wire t0_01101011100, t0_01101011101;
mixer mix_t0_01101011100 (.a(t0_011010111000), .b(t0_011010111001), .y(t0_01101011100));
wire t0_011010111000, t0_011010111001;
mixer mix_t0_01101011101 (.a(t0_011010111010), .b(t0_011010111011), .y(t0_01101011101));
wire t0_011010111010, t0_011010111011;
mixer mix_t0_0110101111 (.a(t0_01101011110), .b(t0_01101011111), .y(t0_0110101111));
wire t0_01101011110, t0_01101011111;
mixer mix_t0_01101011110 (.a(t0_011010111100), .b(t0_011010111101), .y(t0_01101011110));
wire t0_011010111100, t0_011010111101;
mixer mix_t0_01101011111 (.a(t0_011010111110), .b(t0_011010111111), .y(t0_01101011111));
wire t0_011010111110, t0_011010111111;
mixer mix_t0_011011 (.a(t0_0110110), .b(t0_0110111), .y(t0_011011));
wire t0_0110110, t0_0110111;
mixer mix_t0_0110110 (.a(t0_01101100), .b(t0_01101101), .y(t0_0110110));
wire t0_01101100, t0_01101101;
mixer mix_t0_01101100 (.a(t0_011011000), .b(t0_011011001), .y(t0_01101100));
wire t0_011011000, t0_011011001;
mixer mix_t0_011011000 (.a(t0_0110110000), .b(t0_0110110001), .y(t0_011011000));
wire t0_0110110000, t0_0110110001;
mixer mix_t0_0110110000 (.a(t0_01101100000), .b(t0_01101100001), .y(t0_0110110000));
wire t0_01101100000, t0_01101100001;
mixer mix_t0_01101100000 (.a(t0_011011000000), .b(t0_011011000001), .y(t0_01101100000));
wire t0_011011000000, t0_011011000001;
mixer mix_t0_01101100001 (.a(t0_011011000010), .b(t0_011011000011), .y(t0_01101100001));
wire t0_011011000010, t0_011011000011;
mixer mix_t0_0110110001 (.a(t0_01101100010), .b(t0_01101100011), .y(t0_0110110001));
wire t0_01101100010, t0_01101100011;
mixer mix_t0_01101100010 (.a(t0_011011000100), .b(t0_011011000101), .y(t0_01101100010));
wire t0_011011000100, t0_011011000101;
mixer mix_t0_01101100011 (.a(t0_011011000110), .b(t0_011011000111), .y(t0_01101100011));
wire t0_011011000110, t0_011011000111;
mixer mix_t0_011011001 (.a(t0_0110110010), .b(t0_0110110011), .y(t0_011011001));
wire t0_0110110010, t0_0110110011;
mixer mix_t0_0110110010 (.a(t0_01101100100), .b(t0_01101100101), .y(t0_0110110010));
wire t0_01101100100, t0_01101100101;
mixer mix_t0_01101100100 (.a(t0_011011001000), .b(t0_011011001001), .y(t0_01101100100));
wire t0_011011001000, t0_011011001001;
mixer mix_t0_01101100101 (.a(t0_011011001010), .b(t0_011011001011), .y(t0_01101100101));
wire t0_011011001010, t0_011011001011;
mixer mix_t0_0110110011 (.a(t0_01101100110), .b(t0_01101100111), .y(t0_0110110011));
wire t0_01101100110, t0_01101100111;
mixer mix_t0_01101100110 (.a(t0_011011001100), .b(t0_011011001101), .y(t0_01101100110));
wire t0_011011001100, t0_011011001101;
mixer mix_t0_01101100111 (.a(t0_011011001110), .b(t0_011011001111), .y(t0_01101100111));
wire t0_011011001110, t0_011011001111;
mixer mix_t0_01101101 (.a(t0_011011010), .b(t0_011011011), .y(t0_01101101));
wire t0_011011010, t0_011011011;
mixer mix_t0_011011010 (.a(t0_0110110100), .b(t0_0110110101), .y(t0_011011010));
wire t0_0110110100, t0_0110110101;
mixer mix_t0_0110110100 (.a(t0_01101101000), .b(t0_01101101001), .y(t0_0110110100));
wire t0_01101101000, t0_01101101001;
mixer mix_t0_01101101000 (.a(t0_011011010000), .b(t0_011011010001), .y(t0_01101101000));
wire t0_011011010000, t0_011011010001;
mixer mix_t0_01101101001 (.a(t0_011011010010), .b(t0_011011010011), .y(t0_01101101001));
wire t0_011011010010, t0_011011010011;
mixer mix_t0_0110110101 (.a(t0_01101101010), .b(t0_01101101011), .y(t0_0110110101));
wire t0_01101101010, t0_01101101011;
mixer mix_t0_01101101010 (.a(t0_011011010100), .b(t0_011011010101), .y(t0_01101101010));
wire t0_011011010100, t0_011011010101;
mixer mix_t0_01101101011 (.a(t0_011011010110), .b(t0_011011010111), .y(t0_01101101011));
wire t0_011011010110, t0_011011010111;
mixer mix_t0_011011011 (.a(t0_0110110110), .b(t0_0110110111), .y(t0_011011011));
wire t0_0110110110, t0_0110110111;
mixer mix_t0_0110110110 (.a(t0_01101101100), .b(t0_01101101101), .y(t0_0110110110));
wire t0_01101101100, t0_01101101101;
mixer mix_t0_01101101100 (.a(t0_011011011000), .b(t0_011011011001), .y(t0_01101101100));
wire t0_011011011000, t0_011011011001;
mixer mix_t0_01101101101 (.a(t0_011011011010), .b(t0_011011011011), .y(t0_01101101101));
wire t0_011011011010, t0_011011011011;
mixer mix_t0_0110110111 (.a(t0_01101101110), .b(t0_01101101111), .y(t0_0110110111));
wire t0_01101101110, t0_01101101111;
mixer mix_t0_01101101110 (.a(t0_011011011100), .b(t0_011011011101), .y(t0_01101101110));
wire t0_011011011100, t0_011011011101;
mixer mix_t0_01101101111 (.a(t0_011011011110), .b(t0_011011011111), .y(t0_01101101111));
wire t0_011011011110, t0_011011011111;
mixer mix_t0_0110111 (.a(t0_01101110), .b(t0_01101111), .y(t0_0110111));
wire t0_01101110, t0_01101111;
mixer mix_t0_01101110 (.a(t0_011011100), .b(t0_011011101), .y(t0_01101110));
wire t0_011011100, t0_011011101;
mixer mix_t0_011011100 (.a(t0_0110111000), .b(t0_0110111001), .y(t0_011011100));
wire t0_0110111000, t0_0110111001;
mixer mix_t0_0110111000 (.a(t0_01101110000), .b(t0_01101110001), .y(t0_0110111000));
wire t0_01101110000, t0_01101110001;
mixer mix_t0_01101110000 (.a(t0_011011100000), .b(t0_011011100001), .y(t0_01101110000));
wire t0_011011100000, t0_011011100001;
mixer mix_t0_01101110001 (.a(t0_011011100010), .b(t0_011011100011), .y(t0_01101110001));
wire t0_011011100010, t0_011011100011;
mixer mix_t0_0110111001 (.a(t0_01101110010), .b(t0_01101110011), .y(t0_0110111001));
wire t0_01101110010, t0_01101110011;
mixer mix_t0_01101110010 (.a(t0_011011100100), .b(t0_011011100101), .y(t0_01101110010));
wire t0_011011100100, t0_011011100101;
mixer mix_t0_01101110011 (.a(t0_011011100110), .b(t0_011011100111), .y(t0_01101110011));
wire t0_011011100110, t0_011011100111;
mixer mix_t0_011011101 (.a(t0_0110111010), .b(t0_0110111011), .y(t0_011011101));
wire t0_0110111010, t0_0110111011;
mixer mix_t0_0110111010 (.a(t0_01101110100), .b(t0_01101110101), .y(t0_0110111010));
wire t0_01101110100, t0_01101110101;
mixer mix_t0_01101110100 (.a(t0_011011101000), .b(t0_011011101001), .y(t0_01101110100));
wire t0_011011101000, t0_011011101001;
mixer mix_t0_01101110101 (.a(t0_011011101010), .b(t0_011011101011), .y(t0_01101110101));
wire t0_011011101010, t0_011011101011;
mixer mix_t0_0110111011 (.a(t0_01101110110), .b(t0_01101110111), .y(t0_0110111011));
wire t0_01101110110, t0_01101110111;
mixer mix_t0_01101110110 (.a(t0_011011101100), .b(t0_011011101101), .y(t0_01101110110));
wire t0_011011101100, t0_011011101101;
mixer mix_t0_01101110111 (.a(t0_011011101110), .b(t0_011011101111), .y(t0_01101110111));
wire t0_011011101110, t0_011011101111;
mixer mix_t0_01101111 (.a(t0_011011110), .b(t0_011011111), .y(t0_01101111));
wire t0_011011110, t0_011011111;
mixer mix_t0_011011110 (.a(t0_0110111100), .b(t0_0110111101), .y(t0_011011110));
wire t0_0110111100, t0_0110111101;
mixer mix_t0_0110111100 (.a(t0_01101111000), .b(t0_01101111001), .y(t0_0110111100));
wire t0_01101111000, t0_01101111001;
mixer mix_t0_01101111000 (.a(t0_011011110000), .b(t0_011011110001), .y(t0_01101111000));
wire t0_011011110000, t0_011011110001;
mixer mix_t0_01101111001 (.a(t0_011011110010), .b(t0_011011110011), .y(t0_01101111001));
wire t0_011011110010, t0_011011110011;
mixer mix_t0_0110111101 (.a(t0_01101111010), .b(t0_01101111011), .y(t0_0110111101));
wire t0_01101111010, t0_01101111011;
mixer mix_t0_01101111010 (.a(t0_011011110100), .b(t0_011011110101), .y(t0_01101111010));
wire t0_011011110100, t0_011011110101;
mixer mix_t0_01101111011 (.a(t0_011011110110), .b(t0_011011110111), .y(t0_01101111011));
wire t0_011011110110, t0_011011110111;
mixer mix_t0_011011111 (.a(t0_0110111110), .b(t0_0110111111), .y(t0_011011111));
wire t0_0110111110, t0_0110111111;
mixer mix_t0_0110111110 (.a(t0_01101111100), .b(t0_01101111101), .y(t0_0110111110));
wire t0_01101111100, t0_01101111101;
mixer mix_t0_01101111100 (.a(t0_011011111000), .b(t0_011011111001), .y(t0_01101111100));
wire t0_011011111000, t0_011011111001;
mixer mix_t0_01101111101 (.a(t0_011011111010), .b(t0_011011111011), .y(t0_01101111101));
wire t0_011011111010, t0_011011111011;
mixer mix_t0_0110111111 (.a(t0_01101111110), .b(t0_01101111111), .y(t0_0110111111));
wire t0_01101111110, t0_01101111111;
mixer mix_t0_01101111110 (.a(t0_011011111100), .b(t0_011011111101), .y(t0_01101111110));
wire t0_011011111100, t0_011011111101;
mixer mix_t0_01101111111 (.a(t0_011011111110), .b(t0_011011111111), .y(t0_01101111111));
wire t0_011011111110, t0_011011111111;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_011100 (.a(t0_0111000), .b(t0_0111001), .y(t0_011100));
wire t0_0111000, t0_0111001;
mixer mix_t0_0111000 (.a(t0_01110000), .b(t0_01110001), .y(t0_0111000));
wire t0_01110000, t0_01110001;
mixer mix_t0_01110000 (.a(t0_011100000), .b(t0_011100001), .y(t0_01110000));
wire t0_011100000, t0_011100001;
mixer mix_t0_011100000 (.a(t0_0111000000), .b(t0_0111000001), .y(t0_011100000));
wire t0_0111000000, t0_0111000001;
mixer mix_t0_0111000000 (.a(t0_01110000000), .b(t0_01110000001), .y(t0_0111000000));
wire t0_01110000000, t0_01110000001;
mixer mix_t0_01110000000 (.a(t0_011100000000), .b(t0_011100000001), .y(t0_01110000000));
wire t0_011100000000, t0_011100000001;
mixer mix_t0_01110000001 (.a(t0_011100000010), .b(t0_011100000011), .y(t0_01110000001));
wire t0_011100000010, t0_011100000011;
mixer mix_t0_0111000001 (.a(t0_01110000010), .b(t0_01110000011), .y(t0_0111000001));
wire t0_01110000010, t0_01110000011;
mixer mix_t0_01110000010 (.a(t0_011100000100), .b(t0_011100000101), .y(t0_01110000010));
wire t0_011100000100, t0_011100000101;
mixer mix_t0_01110000011 (.a(t0_011100000110), .b(t0_011100000111), .y(t0_01110000011));
wire t0_011100000110, t0_011100000111;
mixer mix_t0_011100001 (.a(t0_0111000010), .b(t0_0111000011), .y(t0_011100001));
wire t0_0111000010, t0_0111000011;
mixer mix_t0_0111000010 (.a(t0_01110000100), .b(t0_01110000101), .y(t0_0111000010));
wire t0_01110000100, t0_01110000101;
mixer mix_t0_01110000100 (.a(t0_011100001000), .b(t0_011100001001), .y(t0_01110000100));
wire t0_011100001000, t0_011100001001;
mixer mix_t0_01110000101 (.a(t0_011100001010), .b(t0_011100001011), .y(t0_01110000101));
wire t0_011100001010, t0_011100001011;
mixer mix_t0_0111000011 (.a(t0_01110000110), .b(t0_01110000111), .y(t0_0111000011));
wire t0_01110000110, t0_01110000111;
mixer mix_t0_01110000110 (.a(t0_011100001100), .b(t0_011100001101), .y(t0_01110000110));
wire t0_011100001100, t0_011100001101;
mixer mix_t0_01110000111 (.a(t0_011100001110), .b(t0_011100001111), .y(t0_01110000111));
wire t0_011100001110, t0_011100001111;
mixer mix_t0_01110001 (.a(t0_011100010), .b(t0_011100011), .y(t0_01110001));
wire t0_011100010, t0_011100011;
mixer mix_t0_011100010 (.a(t0_0111000100), .b(t0_0111000101), .y(t0_011100010));
wire t0_0111000100, t0_0111000101;
mixer mix_t0_0111000100 (.a(t0_01110001000), .b(t0_01110001001), .y(t0_0111000100));
wire t0_01110001000, t0_01110001001;
mixer mix_t0_01110001000 (.a(t0_011100010000), .b(t0_011100010001), .y(t0_01110001000));
wire t0_011100010000, t0_011100010001;
mixer mix_t0_01110001001 (.a(t0_011100010010), .b(t0_011100010011), .y(t0_01110001001));
wire t0_011100010010, t0_011100010011;
mixer mix_t0_0111000101 (.a(t0_01110001010), .b(t0_01110001011), .y(t0_0111000101));
wire t0_01110001010, t0_01110001011;
mixer mix_t0_01110001010 (.a(t0_011100010100), .b(t0_011100010101), .y(t0_01110001010));
wire t0_011100010100, t0_011100010101;
mixer mix_t0_01110001011 (.a(t0_011100010110), .b(t0_011100010111), .y(t0_01110001011));
wire t0_011100010110, t0_011100010111;
mixer mix_t0_011100011 (.a(t0_0111000110), .b(t0_0111000111), .y(t0_011100011));
wire t0_0111000110, t0_0111000111;
mixer mix_t0_0111000110 (.a(t0_01110001100), .b(t0_01110001101), .y(t0_0111000110));
wire t0_01110001100, t0_01110001101;
mixer mix_t0_01110001100 (.a(t0_011100011000), .b(t0_011100011001), .y(t0_01110001100));
wire t0_011100011000, t0_011100011001;
mixer mix_t0_01110001101 (.a(t0_011100011010), .b(t0_011100011011), .y(t0_01110001101));
wire t0_011100011010, t0_011100011011;
mixer mix_t0_0111000111 (.a(t0_01110001110), .b(t0_01110001111), .y(t0_0111000111));
wire t0_01110001110, t0_01110001111;
mixer mix_t0_01110001110 (.a(t0_011100011100), .b(t0_011100011101), .y(t0_01110001110));
wire t0_011100011100, t0_011100011101;
mixer mix_t0_01110001111 (.a(t0_011100011110), .b(t0_011100011111), .y(t0_01110001111));
wire t0_011100011110, t0_011100011111;
mixer mix_t0_0111001 (.a(t0_01110010), .b(t0_01110011), .y(t0_0111001));
wire t0_01110010, t0_01110011;
mixer mix_t0_01110010 (.a(t0_011100100), .b(t0_011100101), .y(t0_01110010));
wire t0_011100100, t0_011100101;
mixer mix_t0_011100100 (.a(t0_0111001000), .b(t0_0111001001), .y(t0_011100100));
wire t0_0111001000, t0_0111001001;
mixer mix_t0_0111001000 (.a(t0_01110010000), .b(t0_01110010001), .y(t0_0111001000));
wire t0_01110010000, t0_01110010001;
mixer mix_t0_01110010000 (.a(t0_011100100000), .b(t0_011100100001), .y(t0_01110010000));
wire t0_011100100000, t0_011100100001;
mixer mix_t0_01110010001 (.a(t0_011100100010), .b(t0_011100100011), .y(t0_01110010001));
wire t0_011100100010, t0_011100100011;
mixer mix_t0_0111001001 (.a(t0_01110010010), .b(t0_01110010011), .y(t0_0111001001));
wire t0_01110010010, t0_01110010011;
mixer mix_t0_01110010010 (.a(t0_011100100100), .b(t0_011100100101), .y(t0_01110010010));
wire t0_011100100100, t0_011100100101;
mixer mix_t0_01110010011 (.a(t0_011100100110), .b(t0_011100100111), .y(t0_01110010011));
wire t0_011100100110, t0_011100100111;
mixer mix_t0_011100101 (.a(t0_0111001010), .b(t0_0111001011), .y(t0_011100101));
wire t0_0111001010, t0_0111001011;
mixer mix_t0_0111001010 (.a(t0_01110010100), .b(t0_01110010101), .y(t0_0111001010));
wire t0_01110010100, t0_01110010101;
mixer mix_t0_01110010100 (.a(t0_011100101000), .b(t0_011100101001), .y(t0_01110010100));
wire t0_011100101000, t0_011100101001;
mixer mix_t0_01110010101 (.a(t0_011100101010), .b(t0_011100101011), .y(t0_01110010101));
wire t0_011100101010, t0_011100101011;
mixer mix_t0_0111001011 (.a(t0_01110010110), .b(t0_01110010111), .y(t0_0111001011));
wire t0_01110010110, t0_01110010111;
mixer mix_t0_01110010110 (.a(t0_011100101100), .b(t0_011100101101), .y(t0_01110010110));
wire t0_011100101100, t0_011100101101;
mixer mix_t0_01110010111 (.a(t0_011100101110), .b(t0_011100101111), .y(t0_01110010111));
wire t0_011100101110, t0_011100101111;
mixer mix_t0_01110011 (.a(t0_011100110), .b(t0_011100111), .y(t0_01110011));
wire t0_011100110, t0_011100111;
mixer mix_t0_011100110 (.a(t0_0111001100), .b(t0_0111001101), .y(t0_011100110));
wire t0_0111001100, t0_0111001101;
mixer mix_t0_0111001100 (.a(t0_01110011000), .b(t0_01110011001), .y(t0_0111001100));
wire t0_01110011000, t0_01110011001;
mixer mix_t0_01110011000 (.a(t0_011100110000), .b(t0_011100110001), .y(t0_01110011000));
wire t0_011100110000, t0_011100110001;
mixer mix_t0_01110011001 (.a(t0_011100110010), .b(t0_011100110011), .y(t0_01110011001));
wire t0_011100110010, t0_011100110011;
mixer mix_t0_0111001101 (.a(t0_01110011010), .b(t0_01110011011), .y(t0_0111001101));
wire t0_01110011010, t0_01110011011;
mixer mix_t0_01110011010 (.a(t0_011100110100), .b(t0_011100110101), .y(t0_01110011010));
wire t0_011100110100, t0_011100110101;
mixer mix_t0_01110011011 (.a(t0_011100110110), .b(t0_011100110111), .y(t0_01110011011));
wire t0_011100110110, t0_011100110111;
mixer mix_t0_011100111 (.a(t0_0111001110), .b(t0_0111001111), .y(t0_011100111));
wire t0_0111001110, t0_0111001111;
mixer mix_t0_0111001110 (.a(t0_01110011100), .b(t0_01110011101), .y(t0_0111001110));
wire t0_01110011100, t0_01110011101;
mixer mix_t0_01110011100 (.a(t0_011100111000), .b(t0_011100111001), .y(t0_01110011100));
wire t0_011100111000, t0_011100111001;
mixer mix_t0_01110011101 (.a(t0_011100111010), .b(t0_011100111011), .y(t0_01110011101));
wire t0_011100111010, t0_011100111011;
mixer mix_t0_0111001111 (.a(t0_01110011110), .b(t0_01110011111), .y(t0_0111001111));
wire t0_01110011110, t0_01110011111;
mixer mix_t0_01110011110 (.a(t0_011100111100), .b(t0_011100111101), .y(t0_01110011110));
wire t0_011100111100, t0_011100111101;
mixer mix_t0_01110011111 (.a(t0_011100111110), .b(t0_011100111111), .y(t0_01110011111));
wire t0_011100111110, t0_011100111111;
mixer mix_t0_011101 (.a(t0_0111010), .b(t0_0111011), .y(t0_011101));
wire t0_0111010, t0_0111011;
mixer mix_t0_0111010 (.a(t0_01110100), .b(t0_01110101), .y(t0_0111010));
wire t0_01110100, t0_01110101;
mixer mix_t0_01110100 (.a(t0_011101000), .b(t0_011101001), .y(t0_01110100));
wire t0_011101000, t0_011101001;
mixer mix_t0_011101000 (.a(t0_0111010000), .b(t0_0111010001), .y(t0_011101000));
wire t0_0111010000, t0_0111010001;
mixer mix_t0_0111010000 (.a(t0_01110100000), .b(t0_01110100001), .y(t0_0111010000));
wire t0_01110100000, t0_01110100001;
mixer mix_t0_01110100000 (.a(t0_011101000000), .b(t0_011101000001), .y(t0_01110100000));
wire t0_011101000000, t0_011101000001;
mixer mix_t0_01110100001 (.a(t0_011101000010), .b(t0_011101000011), .y(t0_01110100001));
wire t0_011101000010, t0_011101000011;
mixer mix_t0_0111010001 (.a(t0_01110100010), .b(t0_01110100011), .y(t0_0111010001));
wire t0_01110100010, t0_01110100011;
mixer mix_t0_01110100010 (.a(t0_011101000100), .b(t0_011101000101), .y(t0_01110100010));
wire t0_011101000100, t0_011101000101;
mixer mix_t0_01110100011 (.a(t0_011101000110), .b(t0_011101000111), .y(t0_01110100011));
wire t0_011101000110, t0_011101000111;
mixer mix_t0_011101001 (.a(t0_0111010010), .b(t0_0111010011), .y(t0_011101001));
wire t0_0111010010, t0_0111010011;
mixer mix_t0_0111010010 (.a(t0_01110100100), .b(t0_01110100101), .y(t0_0111010010));
wire t0_01110100100, t0_01110100101;
mixer mix_t0_01110100100 (.a(t0_011101001000), .b(t0_011101001001), .y(t0_01110100100));
wire t0_011101001000, t0_011101001001;
mixer mix_t0_01110100101 (.a(t0_011101001010), .b(t0_011101001011), .y(t0_01110100101));
wire t0_011101001010, t0_011101001011;
mixer mix_t0_0111010011 (.a(t0_01110100110), .b(t0_01110100111), .y(t0_0111010011));
wire t0_01110100110, t0_01110100111;
mixer mix_t0_01110100110 (.a(t0_011101001100), .b(t0_011101001101), .y(t0_01110100110));
wire t0_011101001100, t0_011101001101;
mixer mix_t0_01110100111 (.a(t0_011101001110), .b(t0_011101001111), .y(t0_01110100111));
wire t0_011101001110, t0_011101001111;
mixer mix_t0_01110101 (.a(t0_011101010), .b(t0_011101011), .y(t0_01110101));
wire t0_011101010, t0_011101011;
mixer mix_t0_011101010 (.a(t0_0111010100), .b(t0_0111010101), .y(t0_011101010));
wire t0_0111010100, t0_0111010101;
mixer mix_t0_0111010100 (.a(t0_01110101000), .b(t0_01110101001), .y(t0_0111010100));
wire t0_01110101000, t0_01110101001;
mixer mix_t0_01110101000 (.a(t0_011101010000), .b(t0_011101010001), .y(t0_01110101000));
wire t0_011101010000, t0_011101010001;
mixer mix_t0_01110101001 (.a(t0_011101010010), .b(t0_011101010011), .y(t0_01110101001));
wire t0_011101010010, t0_011101010011;
mixer mix_t0_0111010101 (.a(t0_01110101010), .b(t0_01110101011), .y(t0_0111010101));
wire t0_01110101010, t0_01110101011;
mixer mix_t0_01110101010 (.a(t0_011101010100), .b(t0_011101010101), .y(t0_01110101010));
wire t0_011101010100, t0_011101010101;
mixer mix_t0_01110101011 (.a(t0_011101010110), .b(t0_011101010111), .y(t0_01110101011));
wire t0_011101010110, t0_011101010111;
mixer mix_t0_011101011 (.a(t0_0111010110), .b(t0_0111010111), .y(t0_011101011));
wire t0_0111010110, t0_0111010111;
mixer mix_t0_0111010110 (.a(t0_01110101100), .b(t0_01110101101), .y(t0_0111010110));
wire t0_01110101100, t0_01110101101;
mixer mix_t0_01110101100 (.a(t0_011101011000), .b(t0_011101011001), .y(t0_01110101100));
wire t0_011101011000, t0_011101011001;
mixer mix_t0_01110101101 (.a(t0_011101011010), .b(t0_011101011011), .y(t0_01110101101));
wire t0_011101011010, t0_011101011011;
mixer mix_t0_0111010111 (.a(t0_01110101110), .b(t0_01110101111), .y(t0_0111010111));
wire t0_01110101110, t0_01110101111;
mixer mix_t0_01110101110 (.a(t0_011101011100), .b(t0_011101011101), .y(t0_01110101110));
wire t0_011101011100, t0_011101011101;
mixer mix_t0_01110101111 (.a(t0_011101011110), .b(t0_011101011111), .y(t0_01110101111));
wire t0_011101011110, t0_011101011111;
mixer mix_t0_0111011 (.a(t0_01110110), .b(t0_01110111), .y(t0_0111011));
wire t0_01110110, t0_01110111;
mixer mix_t0_01110110 (.a(t0_011101100), .b(t0_011101101), .y(t0_01110110));
wire t0_011101100, t0_011101101;
mixer mix_t0_011101100 (.a(t0_0111011000), .b(t0_0111011001), .y(t0_011101100));
wire t0_0111011000, t0_0111011001;
mixer mix_t0_0111011000 (.a(t0_01110110000), .b(t0_01110110001), .y(t0_0111011000));
wire t0_01110110000, t0_01110110001;
mixer mix_t0_01110110000 (.a(t0_011101100000), .b(t0_011101100001), .y(t0_01110110000));
wire t0_011101100000, t0_011101100001;
mixer mix_t0_01110110001 (.a(t0_011101100010), .b(t0_011101100011), .y(t0_01110110001));
wire t0_011101100010, t0_011101100011;
mixer mix_t0_0111011001 (.a(t0_01110110010), .b(t0_01110110011), .y(t0_0111011001));
wire t0_01110110010, t0_01110110011;
mixer mix_t0_01110110010 (.a(t0_011101100100), .b(t0_011101100101), .y(t0_01110110010));
wire t0_011101100100, t0_011101100101;
mixer mix_t0_01110110011 (.a(t0_011101100110), .b(t0_011101100111), .y(t0_01110110011));
wire t0_011101100110, t0_011101100111;
mixer mix_t0_011101101 (.a(t0_0111011010), .b(t0_0111011011), .y(t0_011101101));
wire t0_0111011010, t0_0111011011;
mixer mix_t0_0111011010 (.a(t0_01110110100), .b(t0_01110110101), .y(t0_0111011010));
wire t0_01110110100, t0_01110110101;
mixer mix_t0_01110110100 (.a(t0_011101101000), .b(t0_011101101001), .y(t0_01110110100));
wire t0_011101101000, t0_011101101001;
mixer mix_t0_01110110101 (.a(t0_011101101010), .b(t0_011101101011), .y(t0_01110110101));
wire t0_011101101010, t0_011101101011;
mixer mix_t0_0111011011 (.a(t0_01110110110), .b(t0_01110110111), .y(t0_0111011011));
wire t0_01110110110, t0_01110110111;
mixer mix_t0_01110110110 (.a(t0_011101101100), .b(t0_011101101101), .y(t0_01110110110));
wire t0_011101101100, t0_011101101101;
mixer mix_t0_01110110111 (.a(t0_011101101110), .b(t0_011101101111), .y(t0_01110110111));
wire t0_011101101110, t0_011101101111;
mixer mix_t0_01110111 (.a(t0_011101110), .b(t0_011101111), .y(t0_01110111));
wire t0_011101110, t0_011101111;
mixer mix_t0_011101110 (.a(t0_0111011100), .b(t0_0111011101), .y(t0_011101110));
wire t0_0111011100, t0_0111011101;
mixer mix_t0_0111011100 (.a(t0_01110111000), .b(t0_01110111001), .y(t0_0111011100));
wire t0_01110111000, t0_01110111001;
mixer mix_t0_01110111000 (.a(t0_011101110000), .b(t0_011101110001), .y(t0_01110111000));
wire t0_011101110000, t0_011101110001;
mixer mix_t0_01110111001 (.a(t0_011101110010), .b(t0_011101110011), .y(t0_01110111001));
wire t0_011101110010, t0_011101110011;
mixer mix_t0_0111011101 (.a(t0_01110111010), .b(t0_01110111011), .y(t0_0111011101));
wire t0_01110111010, t0_01110111011;
mixer mix_t0_01110111010 (.a(t0_011101110100), .b(t0_011101110101), .y(t0_01110111010));
wire t0_011101110100, t0_011101110101;
mixer mix_t0_01110111011 (.a(t0_011101110110), .b(t0_011101110111), .y(t0_01110111011));
wire t0_011101110110, t0_011101110111;
mixer mix_t0_011101111 (.a(t0_0111011110), .b(t0_0111011111), .y(t0_011101111));
wire t0_0111011110, t0_0111011111;
mixer mix_t0_0111011110 (.a(t0_01110111100), .b(t0_01110111101), .y(t0_0111011110));
wire t0_01110111100, t0_01110111101;
mixer mix_t0_01110111100 (.a(t0_011101111000), .b(t0_011101111001), .y(t0_01110111100));
wire t0_011101111000, t0_011101111001;
mixer mix_t0_01110111101 (.a(t0_011101111010), .b(t0_011101111011), .y(t0_01110111101));
wire t0_011101111010, t0_011101111011;
mixer mix_t0_0111011111 (.a(t0_01110111110), .b(t0_01110111111), .y(t0_0111011111));
wire t0_01110111110, t0_01110111111;
mixer mix_t0_01110111110 (.a(t0_011101111100), .b(t0_011101111101), .y(t0_01110111110));
wire t0_011101111100, t0_011101111101;
mixer mix_t0_01110111111 (.a(t0_011101111110), .b(t0_011101111111), .y(t0_01110111111));
wire t0_011101111110, t0_011101111111;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
mixer mix_t0_011110 (.a(t0_0111100), .b(t0_0111101), .y(t0_011110));
wire t0_0111100, t0_0111101;
mixer mix_t0_0111100 (.a(t0_01111000), .b(t0_01111001), .y(t0_0111100));
wire t0_01111000, t0_01111001;
mixer mix_t0_01111000 (.a(t0_011110000), .b(t0_011110001), .y(t0_01111000));
wire t0_011110000, t0_011110001;
mixer mix_t0_011110000 (.a(t0_0111100000), .b(t0_0111100001), .y(t0_011110000));
wire t0_0111100000, t0_0111100001;
mixer mix_t0_0111100000 (.a(t0_01111000000), .b(t0_01111000001), .y(t0_0111100000));
wire t0_01111000000, t0_01111000001;
mixer mix_t0_01111000000 (.a(t0_011110000000), .b(t0_011110000001), .y(t0_01111000000));
wire t0_011110000000, t0_011110000001;
mixer mix_t0_01111000001 (.a(t0_011110000010), .b(t0_011110000011), .y(t0_01111000001));
wire t0_011110000010, t0_011110000011;
mixer mix_t0_0111100001 (.a(t0_01111000010), .b(t0_01111000011), .y(t0_0111100001));
wire t0_01111000010, t0_01111000011;
mixer mix_t0_01111000010 (.a(t0_011110000100), .b(t0_011110000101), .y(t0_01111000010));
wire t0_011110000100, t0_011110000101;
mixer mix_t0_01111000011 (.a(t0_011110000110), .b(t0_011110000111), .y(t0_01111000011));
wire t0_011110000110, t0_011110000111;
mixer mix_t0_011110001 (.a(t0_0111100010), .b(t0_0111100011), .y(t0_011110001));
wire t0_0111100010, t0_0111100011;
mixer mix_t0_0111100010 (.a(t0_01111000100), .b(t0_01111000101), .y(t0_0111100010));
wire t0_01111000100, t0_01111000101;
mixer mix_t0_01111000100 (.a(t0_011110001000), .b(t0_011110001001), .y(t0_01111000100));
wire t0_011110001000, t0_011110001001;
mixer mix_t0_01111000101 (.a(t0_011110001010), .b(t0_011110001011), .y(t0_01111000101));
wire t0_011110001010, t0_011110001011;
mixer mix_t0_0111100011 (.a(t0_01111000110), .b(t0_01111000111), .y(t0_0111100011));
wire t0_01111000110, t0_01111000111;
mixer mix_t0_01111000110 (.a(t0_011110001100), .b(t0_011110001101), .y(t0_01111000110));
wire t0_011110001100, t0_011110001101;
mixer mix_t0_01111000111 (.a(t0_011110001110), .b(t0_011110001111), .y(t0_01111000111));
wire t0_011110001110, t0_011110001111;
mixer mix_t0_01111001 (.a(t0_011110010), .b(t0_011110011), .y(t0_01111001));
wire t0_011110010, t0_011110011;
mixer mix_t0_011110010 (.a(t0_0111100100), .b(t0_0111100101), .y(t0_011110010));
wire t0_0111100100, t0_0111100101;
mixer mix_t0_0111100100 (.a(t0_01111001000), .b(t0_01111001001), .y(t0_0111100100));
wire t0_01111001000, t0_01111001001;
mixer mix_t0_01111001000 (.a(t0_011110010000), .b(t0_011110010001), .y(t0_01111001000));
wire t0_011110010000, t0_011110010001;
mixer mix_t0_01111001001 (.a(t0_011110010010), .b(t0_011110010011), .y(t0_01111001001));
wire t0_011110010010, t0_011110010011;
mixer mix_t0_0111100101 (.a(t0_01111001010), .b(t0_01111001011), .y(t0_0111100101));
wire t0_01111001010, t0_01111001011;
mixer mix_t0_01111001010 (.a(t0_011110010100), .b(t0_011110010101), .y(t0_01111001010));
wire t0_011110010100, t0_011110010101;
mixer mix_t0_01111001011 (.a(t0_011110010110), .b(t0_011110010111), .y(t0_01111001011));
wire t0_011110010110, t0_011110010111;
mixer mix_t0_011110011 (.a(t0_0111100110), .b(t0_0111100111), .y(t0_011110011));
wire t0_0111100110, t0_0111100111;
mixer mix_t0_0111100110 (.a(t0_01111001100), .b(t0_01111001101), .y(t0_0111100110));
wire t0_01111001100, t0_01111001101;
mixer mix_t0_01111001100 (.a(t0_011110011000), .b(t0_011110011001), .y(t0_01111001100));
wire t0_011110011000, t0_011110011001;
mixer mix_t0_01111001101 (.a(t0_011110011010), .b(t0_011110011011), .y(t0_01111001101));
wire t0_011110011010, t0_011110011011;
mixer mix_t0_0111100111 (.a(t0_01111001110), .b(t0_01111001111), .y(t0_0111100111));
wire t0_01111001110, t0_01111001111;
mixer mix_t0_01111001110 (.a(t0_011110011100), .b(t0_011110011101), .y(t0_01111001110));
wire t0_011110011100, t0_011110011101;
mixer mix_t0_01111001111 (.a(t0_011110011110), .b(t0_011110011111), .y(t0_01111001111));
wire t0_011110011110, t0_011110011111;
mixer mix_t0_0111101 (.a(t0_01111010), .b(t0_01111011), .y(t0_0111101));
wire t0_01111010, t0_01111011;
mixer mix_t0_01111010 (.a(t0_011110100), .b(t0_011110101), .y(t0_01111010));
wire t0_011110100, t0_011110101;
mixer mix_t0_011110100 (.a(t0_0111101000), .b(t0_0111101001), .y(t0_011110100));
wire t0_0111101000, t0_0111101001;
mixer mix_t0_0111101000 (.a(t0_01111010000), .b(t0_01111010001), .y(t0_0111101000));
wire t0_01111010000, t0_01111010001;
mixer mix_t0_01111010000 (.a(t0_011110100000), .b(t0_011110100001), .y(t0_01111010000));
wire t0_011110100000, t0_011110100001;
mixer mix_t0_01111010001 (.a(t0_011110100010), .b(t0_011110100011), .y(t0_01111010001));
wire t0_011110100010, t0_011110100011;
mixer mix_t0_0111101001 (.a(t0_01111010010), .b(t0_01111010011), .y(t0_0111101001));
wire t0_01111010010, t0_01111010011;
mixer mix_t0_01111010010 (.a(t0_011110100100), .b(t0_011110100101), .y(t0_01111010010));
wire t0_011110100100, t0_011110100101;
mixer mix_t0_01111010011 (.a(t0_011110100110), .b(t0_011110100111), .y(t0_01111010011));
wire t0_011110100110, t0_011110100111;
mixer mix_t0_011110101 (.a(t0_0111101010), .b(t0_0111101011), .y(t0_011110101));
wire t0_0111101010, t0_0111101011;
mixer mix_t0_0111101010 (.a(t0_01111010100), .b(t0_01111010101), .y(t0_0111101010));
wire t0_01111010100, t0_01111010101;
mixer mix_t0_01111010100 (.a(t0_011110101000), .b(t0_011110101001), .y(t0_01111010100));
wire t0_011110101000, t0_011110101001;
mixer mix_t0_01111010101 (.a(t0_011110101010), .b(t0_011110101011), .y(t0_01111010101));
wire t0_011110101010, t0_011110101011;
mixer mix_t0_0111101011 (.a(t0_01111010110), .b(t0_01111010111), .y(t0_0111101011));
wire t0_01111010110, t0_01111010111;
mixer mix_t0_01111010110 (.a(t0_011110101100), .b(t0_011110101101), .y(t0_01111010110));
wire t0_011110101100, t0_011110101101;
mixer mix_t0_01111010111 (.a(t0_011110101110), .b(t0_011110101111), .y(t0_01111010111));
wire t0_011110101110, t0_011110101111;
mixer mix_t0_01111011 (.a(t0_011110110), .b(t0_011110111), .y(t0_01111011));
wire t0_011110110, t0_011110111;
mixer mix_t0_011110110 (.a(t0_0111101100), .b(t0_0111101101), .y(t0_011110110));
wire t0_0111101100, t0_0111101101;
mixer mix_t0_0111101100 (.a(t0_01111011000), .b(t0_01111011001), .y(t0_0111101100));
wire t0_01111011000, t0_01111011001;
mixer mix_t0_01111011000 (.a(t0_011110110000), .b(t0_011110110001), .y(t0_01111011000));
wire t0_011110110000, t0_011110110001;
mixer mix_t0_01111011001 (.a(t0_011110110010), .b(t0_011110110011), .y(t0_01111011001));
wire t0_011110110010, t0_011110110011;
mixer mix_t0_0111101101 (.a(t0_01111011010), .b(t0_01111011011), .y(t0_0111101101));
wire t0_01111011010, t0_01111011011;
mixer mix_t0_01111011010 (.a(t0_011110110100), .b(t0_011110110101), .y(t0_01111011010));
wire t0_011110110100, t0_011110110101;
mixer mix_t0_01111011011 (.a(t0_011110110110), .b(t0_011110110111), .y(t0_01111011011));
wire t0_011110110110, t0_011110110111;
mixer mix_t0_011110111 (.a(t0_0111101110), .b(t0_0111101111), .y(t0_011110111));
wire t0_0111101110, t0_0111101111;
mixer mix_t0_0111101110 (.a(t0_01111011100), .b(t0_01111011101), .y(t0_0111101110));
wire t0_01111011100, t0_01111011101;
mixer mix_t0_01111011100 (.a(t0_011110111000), .b(t0_011110111001), .y(t0_01111011100));
wire t0_011110111000, t0_011110111001;
mixer mix_t0_01111011101 (.a(t0_011110111010), .b(t0_011110111011), .y(t0_01111011101));
wire t0_011110111010, t0_011110111011;
mixer mix_t0_0111101111 (.a(t0_01111011110), .b(t0_01111011111), .y(t0_0111101111));
wire t0_01111011110, t0_01111011111;
mixer mix_t0_01111011110 (.a(t0_011110111100), .b(t0_011110111101), .y(t0_01111011110));
wire t0_011110111100, t0_011110111101;
mixer mix_t0_01111011111 (.a(t0_011110111110), .b(t0_011110111111), .y(t0_01111011111));
wire t0_011110111110, t0_011110111111;
mixer mix_t0_011111 (.a(t0_0111110), .b(t0_0111111), .y(t0_011111));
wire t0_0111110, t0_0111111;
mixer mix_t0_0111110 (.a(t0_01111100), .b(t0_01111101), .y(t0_0111110));
wire t0_01111100, t0_01111101;
mixer mix_t0_01111100 (.a(t0_011111000), .b(t0_011111001), .y(t0_01111100));
wire t0_011111000, t0_011111001;
mixer mix_t0_011111000 (.a(t0_0111110000), .b(t0_0111110001), .y(t0_011111000));
wire t0_0111110000, t0_0111110001;
mixer mix_t0_0111110000 (.a(t0_01111100000), .b(t0_01111100001), .y(t0_0111110000));
wire t0_01111100000, t0_01111100001;
mixer mix_t0_01111100000 (.a(t0_011111000000), .b(t0_011111000001), .y(t0_01111100000));
wire t0_011111000000, t0_011111000001;
mixer mix_t0_01111100001 (.a(t0_011111000010), .b(t0_011111000011), .y(t0_01111100001));
wire t0_011111000010, t0_011111000011;
mixer mix_t0_0111110001 (.a(t0_01111100010), .b(t0_01111100011), .y(t0_0111110001));
wire t0_01111100010, t0_01111100011;
mixer mix_t0_01111100010 (.a(t0_011111000100), .b(t0_011111000101), .y(t0_01111100010));
wire t0_011111000100, t0_011111000101;
mixer mix_t0_01111100011 (.a(t0_011111000110), .b(t0_011111000111), .y(t0_01111100011));
wire t0_011111000110, t0_011111000111;
mixer mix_t0_011111001 (.a(t0_0111110010), .b(t0_0111110011), .y(t0_011111001));
wire t0_0111110010, t0_0111110011;
mixer mix_t0_0111110010 (.a(t0_01111100100), .b(t0_01111100101), .y(t0_0111110010));
wire t0_01111100100, t0_01111100101;
mixer mix_t0_01111100100 (.a(t0_011111001000), .b(t0_011111001001), .y(t0_01111100100));
wire t0_011111001000, t0_011111001001;
mixer mix_t0_01111100101 (.a(t0_011111001010), .b(t0_011111001011), .y(t0_01111100101));
wire t0_011111001010, t0_011111001011;
mixer mix_t0_0111110011 (.a(t0_01111100110), .b(t0_01111100111), .y(t0_0111110011));
wire t0_01111100110, t0_01111100111;
mixer mix_t0_01111100110 (.a(t0_011111001100), .b(t0_011111001101), .y(t0_01111100110));
wire t0_011111001100, t0_011111001101;
mixer mix_t0_01111100111 (.a(t0_011111001110), .b(t0_011111001111), .y(t0_01111100111));
wire t0_011111001110, t0_011111001111;
mixer mix_t0_01111101 (.a(t0_011111010), .b(t0_011111011), .y(t0_01111101));
wire t0_011111010, t0_011111011;
mixer mix_t0_011111010 (.a(t0_0111110100), .b(t0_0111110101), .y(t0_011111010));
wire t0_0111110100, t0_0111110101;
mixer mix_t0_0111110100 (.a(t0_01111101000), .b(t0_01111101001), .y(t0_0111110100));
wire t0_01111101000, t0_01111101001;
mixer mix_t0_01111101000 (.a(t0_011111010000), .b(t0_011111010001), .y(t0_01111101000));
wire t0_011111010000, t0_011111010001;
mixer mix_t0_01111101001 (.a(t0_011111010010), .b(t0_011111010011), .y(t0_01111101001));
wire t0_011111010010, t0_011111010011;
mixer mix_t0_0111110101 (.a(t0_01111101010), .b(t0_01111101011), .y(t0_0111110101));
wire t0_01111101010, t0_01111101011;
mixer mix_t0_01111101010 (.a(t0_011111010100), .b(t0_011111010101), .y(t0_01111101010));
wire t0_011111010100, t0_011111010101;
mixer mix_t0_01111101011 (.a(t0_011111010110), .b(t0_011111010111), .y(t0_01111101011));
wire t0_011111010110, t0_011111010111;
mixer mix_t0_011111011 (.a(t0_0111110110), .b(t0_0111110111), .y(t0_011111011));
wire t0_0111110110, t0_0111110111;
mixer mix_t0_0111110110 (.a(t0_01111101100), .b(t0_01111101101), .y(t0_0111110110));
wire t0_01111101100, t0_01111101101;
mixer mix_t0_01111101100 (.a(t0_011111011000), .b(t0_011111011001), .y(t0_01111101100));
wire t0_011111011000, t0_011111011001;
mixer mix_t0_01111101101 (.a(t0_011111011010), .b(t0_011111011011), .y(t0_01111101101));
wire t0_011111011010, t0_011111011011;
mixer mix_t0_0111110111 (.a(t0_01111101110), .b(t0_01111101111), .y(t0_0111110111));
wire t0_01111101110, t0_01111101111;
mixer mix_t0_01111101110 (.a(t0_011111011100), .b(t0_011111011101), .y(t0_01111101110));
wire t0_011111011100, t0_011111011101;
mixer mix_t0_01111101111 (.a(t0_011111011110), .b(t0_011111011111), .y(t0_01111101111));
wire t0_011111011110, t0_011111011111;
mixer mix_t0_0111111 (.a(t0_01111110), .b(t0_01111111), .y(t0_0111111));
wire t0_01111110, t0_01111111;
mixer mix_t0_01111110 (.a(t0_011111100), .b(t0_011111101), .y(t0_01111110));
wire t0_011111100, t0_011111101;
mixer mix_t0_011111100 (.a(t0_0111111000), .b(t0_0111111001), .y(t0_011111100));
wire t0_0111111000, t0_0111111001;
mixer mix_t0_0111111000 (.a(t0_01111110000), .b(t0_01111110001), .y(t0_0111111000));
wire t0_01111110000, t0_01111110001;
mixer mix_t0_01111110000 (.a(t0_011111100000), .b(t0_011111100001), .y(t0_01111110000));
wire t0_011111100000, t0_011111100001;
mixer mix_t0_01111110001 (.a(t0_011111100010), .b(t0_011111100011), .y(t0_01111110001));
wire t0_011111100010, t0_011111100011;
mixer mix_t0_0111111001 (.a(t0_01111110010), .b(t0_01111110011), .y(t0_0111111001));
wire t0_01111110010, t0_01111110011;
mixer mix_t0_01111110010 (.a(t0_011111100100), .b(t0_011111100101), .y(t0_01111110010));
wire t0_011111100100, t0_011111100101;
mixer mix_t0_01111110011 (.a(t0_011111100110), .b(t0_011111100111), .y(t0_01111110011));
wire t0_011111100110, t0_011111100111;
mixer mix_t0_011111101 (.a(t0_0111111010), .b(t0_0111111011), .y(t0_011111101));
wire t0_0111111010, t0_0111111011;
mixer mix_t0_0111111010 (.a(t0_01111110100), .b(t0_01111110101), .y(t0_0111111010));
wire t0_01111110100, t0_01111110101;
mixer mix_t0_01111110100 (.a(t0_011111101000), .b(t0_011111101001), .y(t0_01111110100));
wire t0_011111101000, t0_011111101001;
mixer mix_t0_01111110101 (.a(t0_011111101010), .b(t0_011111101011), .y(t0_01111110101));
wire t0_011111101010, t0_011111101011;
mixer mix_t0_0111111011 (.a(t0_01111110110), .b(t0_01111110111), .y(t0_0111111011));
wire t0_01111110110, t0_01111110111;
mixer mix_t0_01111110110 (.a(t0_011111101100), .b(t0_011111101101), .y(t0_01111110110));
wire t0_011111101100, t0_011111101101;
mixer mix_t0_01111110111 (.a(t0_011111101110), .b(t0_011111101111), .y(t0_01111110111));
wire t0_011111101110, t0_011111101111;
mixer mix_t0_01111111 (.a(t0_011111110), .b(t0_011111111), .y(t0_01111111));
wire t0_011111110, t0_011111111;
mixer mix_t0_011111110 (.a(t0_0111111100), .b(t0_0111111101), .y(t0_011111110));
wire t0_0111111100, t0_0111111101;
mixer mix_t0_0111111100 (.a(t0_01111111000), .b(t0_01111111001), .y(t0_0111111100));
wire t0_01111111000, t0_01111111001;
mixer mix_t0_01111111000 (.a(t0_011111110000), .b(t0_011111110001), .y(t0_01111111000));
wire t0_011111110000, t0_011111110001;
mixer mix_t0_01111111001 (.a(t0_011111110010), .b(t0_011111110011), .y(t0_01111111001));
wire t0_011111110010, t0_011111110011;
mixer mix_t0_0111111101 (.a(t0_01111111010), .b(t0_01111111011), .y(t0_0111111101));
wire t0_01111111010, t0_01111111011;
mixer mix_t0_01111111010 (.a(t0_011111110100), .b(t0_011111110101), .y(t0_01111111010));
wire t0_011111110100, t0_011111110101;
mixer mix_t0_01111111011 (.a(t0_011111110110), .b(t0_011111110111), .y(t0_01111111011));
wire t0_011111110110, t0_011111110111;
mixer mix_t0_011111111 (.a(t0_0111111110), .b(t0_0111111111), .y(t0_011111111));
wire t0_0111111110, t0_0111111111;
mixer mix_t0_0111111110 (.a(t0_01111111100), .b(t0_01111111101), .y(t0_0111111110));
wire t0_01111111100, t0_01111111101;
mixer mix_t0_01111111100 (.a(t0_011111111000), .b(t0_011111111001), .y(t0_01111111100));
wire t0_011111111000, t0_011111111001;
mixer mix_t0_01111111101 (.a(t0_011111111010), .b(t0_011111111011), .y(t0_01111111101));
wire t0_011111111010, t0_011111111011;
mixer mix_t0_0111111111 (.a(t0_01111111110), .b(t0_01111111111), .y(t0_0111111111));
wire t0_01111111110, t0_01111111111;
mixer mix_t0_01111111110 (.a(t0_011111111100), .b(t0_011111111101), .y(t0_01111111110));
wire t0_011111111100, t0_011111111101;
mixer mix_t0_01111111111 (.a(t0_011111111110), .b(t0_011111111111), .y(t0_01111111111));
wire t0_011111111110, t0_011111111111;
wire t0_0;
assign out_0 = t0_0;
assign input_0 = t0_000000000000;
assign input_1 = t0_000000000001;
assign input_2 = t0_000000000010;
assign input_3 = t0_000000000011;
assign input_4 = t0_000000000100;
assign input_5 = t0_000000000101;
assign input_6 = t0_000000000110;
assign input_7 = t0_000000000111;
assign input_8 = t0_000000001000;
assign input_9 = t0_000000001001;
assign input_10 = t0_000000001010;
assign input_11 = t0_000000001011;
assign input_12 = t0_000000001100;
assign input_13 = t0_000000001101;
assign input_14 = t0_000000001110;
assign input_15 = t0_000000001111;
assign input_16 = t0_000000010000;
assign input_17 = t0_000000010001;
assign input_18 = t0_000000010010;
assign input_19 = t0_000000010011;
assign input_20 = t0_000000010100;
assign input_21 = t0_000000010101;
assign input_22 = t0_000000010110;
assign input_23 = t0_000000010111;
assign input_24 = t0_000000011000;
assign input_25 = t0_000000011001;
assign input_26 = t0_000000011010;
assign input_27 = t0_000000011011;
assign input_28 = t0_000000011100;
assign input_29 = t0_000000011101;
assign input_30 = t0_000000011110;
assign input_31 = t0_000000011111;
assign input_32 = t0_000000100000;
assign input_33 = t0_000000100001;
assign input_34 = t0_000000100010;
assign input_35 = t0_000000100011;
assign input_36 = t0_000000100100;
assign input_37 = t0_000000100101;
assign input_38 = t0_000000100110;
assign input_39 = t0_000000100111;
assign input_40 = t0_000000101000;
assign input_41 = t0_000000101001;
assign input_42 = t0_000000101010;
assign input_43 = t0_000000101011;
assign input_44 = t0_000000101100;
assign input_45 = t0_000000101101;
assign input_46 = t0_000000101110;
assign input_47 = t0_000000101111;
assign input_48 = t0_000000110000;
assign input_49 = t0_000000110001;
assign input_50 = t0_000000110010;
assign input_51 = t0_000000110011;
assign input_52 = t0_000000110100;
assign input_53 = t0_000000110101;
assign input_54 = t0_000000110110;
assign input_55 = t0_000000110111;
assign input_56 = t0_000000111000;
assign input_57 = t0_000000111001;
assign input_58 = t0_000000111010;
assign input_59 = t0_000000111011;
assign input_60 = t0_000000111100;
assign input_61 = t0_000000111101;
assign input_62 = t0_000000111110;
assign input_63 = t0_000000111111;
assign input_64 = t0_000001000000;
assign input_65 = t0_000001000001;
assign input_66 = t0_000001000010;
assign input_67 = t0_000001000011;
assign input_68 = t0_000001000100;
assign input_69 = t0_000001000101;
assign input_70 = t0_000001000110;
assign input_71 = t0_000001000111;
assign input_72 = t0_000001001000;
assign input_73 = t0_000001001001;
assign input_74 = t0_000001001010;
assign input_75 = t0_000001001011;
assign input_76 = t0_000001001100;
assign input_77 = t0_000001001101;
assign input_78 = t0_000001001110;
assign input_79 = t0_000001001111;
assign input_80 = t0_000001010000;
assign input_81 = t0_000001010001;
assign input_82 = t0_000001010010;
assign input_83 = t0_000001010011;
assign input_84 = t0_000001010100;
assign input_85 = t0_000001010101;
assign input_86 = t0_000001010110;
assign input_87 = t0_000001010111;
assign input_88 = t0_000001011000;
assign input_89 = t0_000001011001;
assign input_90 = t0_000001011010;
assign input_91 = t0_000001011011;
assign input_92 = t0_000001011100;
assign input_93 = t0_000001011101;
assign input_94 = t0_000001011110;
assign input_95 = t0_000001011111;
assign input_96 = t0_000001100000;
assign input_97 = t0_000001100001;
assign input_98 = t0_000001100010;
assign input_99 = t0_000001100011;
assign input_100 = t0_000001100100;
assign input_101 = t0_000001100101;
assign input_102 = t0_000001100110;
assign input_103 = t0_000001100111;
assign input_104 = t0_000001101000;
assign input_105 = t0_000001101001;
assign input_106 = t0_000001101010;
assign input_107 = t0_000001101011;
assign input_108 = t0_000001101100;
assign input_109 = t0_000001101101;
assign input_110 = t0_000001101110;
assign input_111 = t0_000001101111;
assign input_112 = t0_000001110000;
assign input_113 = t0_000001110001;
assign input_114 = t0_000001110010;
assign input_115 = t0_000001110011;
assign input_116 = t0_000001110100;
assign input_117 = t0_000001110101;
assign input_118 = t0_000001110110;
assign input_119 = t0_000001110111;
assign input_120 = t0_000001111000;
assign input_121 = t0_000001111001;
assign input_122 = t0_000001111010;
assign input_123 = t0_000001111011;
assign input_124 = t0_000001111100;
assign input_125 = t0_000001111101;
assign input_126 = t0_000001111110;
assign input_127 = t0_000001111111;
assign input_128 = t0_000010000000;
assign input_129 = t0_000010000001;
assign input_130 = t0_000010000010;
assign input_131 = t0_000010000011;
assign input_132 = t0_000010000100;
assign input_133 = t0_000010000101;
assign input_134 = t0_000010000110;
assign input_135 = t0_000010000111;
assign input_136 = t0_000010001000;
assign input_137 = t0_000010001001;
assign input_138 = t0_000010001010;
assign input_139 = t0_000010001011;
assign input_140 = t0_000010001100;
assign input_141 = t0_000010001101;
assign input_142 = t0_000010001110;
assign input_143 = t0_000010001111;
assign input_144 = t0_000010010000;
assign input_145 = t0_000010010001;
assign input_146 = t0_000010010010;
assign input_147 = t0_000010010011;
assign input_148 = t0_000010010100;
assign input_149 = t0_000010010101;
assign input_150 = t0_000010010110;
assign input_151 = t0_000010010111;
assign input_152 = t0_000010011000;
assign input_153 = t0_000010011001;
assign input_154 = t0_000010011010;
assign input_155 = t0_000010011011;
assign input_156 = t0_000010011100;
assign input_157 = t0_000010011101;
assign input_158 = t0_000010011110;
assign input_159 = t0_000010011111;
assign input_160 = t0_000010100000;
assign input_161 = t0_000010100001;
assign input_162 = t0_000010100010;
assign input_163 = t0_000010100011;
assign input_164 = t0_000010100100;
assign input_165 = t0_000010100101;
assign input_166 = t0_000010100110;
assign input_167 = t0_000010100111;
assign input_168 = t0_000010101000;
assign input_169 = t0_000010101001;
assign input_170 = t0_000010101010;
assign input_171 = t0_000010101011;
assign input_172 = t0_000010101100;
assign input_173 = t0_000010101101;
assign input_174 = t0_000010101110;
assign input_175 = t0_000010101111;
assign input_176 = t0_000010110000;
assign input_177 = t0_000010110001;
assign input_178 = t0_000010110010;
assign input_179 = t0_000010110011;
assign input_180 = t0_000010110100;
assign input_181 = t0_000010110101;
assign input_182 = t0_000010110110;
assign input_183 = t0_000010110111;
assign input_184 = t0_000010111000;
assign input_185 = t0_000010111001;
assign input_186 = t0_000010111010;
assign input_187 = t0_000010111011;
assign input_188 = t0_000010111100;
assign input_189 = t0_000010111101;
assign input_190 = t0_000010111110;
assign input_191 = t0_000010111111;
assign input_192 = t0_000011000000;
assign input_193 = t0_000011000001;
assign input_194 = t0_000011000010;
assign input_195 = t0_000011000011;
assign input_196 = t0_000011000100;
assign input_197 = t0_000011000101;
assign input_198 = t0_000011000110;
assign input_199 = t0_000011000111;
assign input_200 = t0_000011001000;
assign input_201 = t0_000011001001;
assign input_202 = t0_000011001010;
assign input_203 = t0_000011001011;
assign input_204 = t0_000011001100;
assign input_205 = t0_000011001101;
assign input_206 = t0_000011001110;
assign input_207 = t0_000011001111;
assign input_208 = t0_000011010000;
assign input_209 = t0_000011010001;
assign input_210 = t0_000011010010;
assign input_211 = t0_000011010011;
assign input_212 = t0_000011010100;
assign input_213 = t0_000011010101;
assign input_214 = t0_000011010110;
assign input_215 = t0_000011010111;
assign input_216 = t0_000011011000;
assign input_217 = t0_000011011001;
assign input_218 = t0_000011011010;
assign input_219 = t0_000011011011;
assign input_220 = t0_000011011100;
assign input_221 = t0_000011011101;
assign input_222 = t0_000011011110;
assign input_223 = t0_000011011111;
assign input_224 = t0_000011100000;
assign input_225 = t0_000011100001;
assign input_226 = t0_000011100010;
assign input_227 = t0_000011100011;
assign input_228 = t0_000011100100;
assign input_229 = t0_000011100101;
assign input_230 = t0_000011100110;
assign input_231 = t0_000011100111;
assign input_232 = t0_000011101000;
assign input_233 = t0_000011101001;
assign input_234 = t0_000011101010;
assign input_235 = t0_000011101011;
assign input_236 = t0_000011101100;
assign input_237 = t0_000011101101;
assign input_238 = t0_000011101110;
assign input_239 = t0_000011101111;
assign input_240 = t0_000011110000;
assign input_241 = t0_000011110001;
assign input_242 = t0_000011110010;
assign input_243 = t0_000011110011;
assign input_244 = t0_000011110100;
assign input_245 = t0_000011110101;
assign input_246 = t0_000011110110;
assign input_247 = t0_000011110111;
assign input_248 = t0_000011111000;
assign input_249 = t0_000011111001;
assign input_250 = t0_000011111010;
assign input_251 = t0_000011111011;
assign input_252 = t0_000011111100;
assign input_253 = t0_000011111101;
assign input_254 = t0_000011111110;
assign input_255 = t0_000011111111;
assign input_256 = t0_000100000000;
assign input_257 = t0_000100000001;
assign input_258 = t0_000100000010;
assign input_259 = t0_000100000011;
assign input_260 = t0_000100000100;
assign input_261 = t0_000100000101;
assign input_262 = t0_000100000110;
assign input_263 = t0_000100000111;
assign input_264 = t0_000100001000;
assign input_265 = t0_000100001001;
assign input_266 = t0_000100001010;
assign input_267 = t0_000100001011;
assign input_268 = t0_000100001100;
assign input_269 = t0_000100001101;
assign input_270 = t0_000100001110;
assign input_271 = t0_000100001111;
assign input_272 = t0_000100010000;
assign input_273 = t0_000100010001;
assign input_274 = t0_000100010010;
assign input_275 = t0_000100010011;
assign input_276 = t0_000100010100;
assign input_277 = t0_000100010101;
assign input_278 = t0_000100010110;
assign input_279 = t0_000100010111;
assign input_280 = t0_000100011000;
assign input_281 = t0_000100011001;
assign input_282 = t0_000100011010;
assign input_283 = t0_000100011011;
assign input_284 = t0_000100011100;
assign input_285 = t0_000100011101;
assign input_286 = t0_000100011110;
assign input_287 = t0_000100011111;
assign input_288 = t0_000100100000;
assign input_289 = t0_000100100001;
assign input_290 = t0_000100100010;
assign input_291 = t0_000100100011;
assign input_292 = t0_000100100100;
assign input_293 = t0_000100100101;
assign input_294 = t0_000100100110;
assign input_295 = t0_000100100111;
assign input_296 = t0_000100101000;
assign input_297 = t0_000100101001;
assign input_298 = t0_000100101010;
assign input_299 = t0_000100101011;
assign input_300 = t0_000100101100;
assign input_301 = t0_000100101101;
assign input_302 = t0_000100101110;
assign input_303 = t0_000100101111;
assign input_304 = t0_000100110000;
assign input_305 = t0_000100110001;
assign input_306 = t0_000100110010;
assign input_307 = t0_000100110011;
assign input_308 = t0_000100110100;
assign input_309 = t0_000100110101;
assign input_310 = t0_000100110110;
assign input_311 = t0_000100110111;
assign input_312 = t0_000100111000;
assign input_313 = t0_000100111001;
assign input_314 = t0_000100111010;
assign input_315 = t0_000100111011;
assign input_316 = t0_000100111100;
assign input_317 = t0_000100111101;
assign input_318 = t0_000100111110;
assign input_319 = t0_000100111111;
assign input_320 = t0_000101000000;
assign input_321 = t0_000101000001;
assign input_322 = t0_000101000010;
assign input_323 = t0_000101000011;
assign input_324 = t0_000101000100;
assign input_325 = t0_000101000101;
assign input_326 = t0_000101000110;
assign input_327 = t0_000101000111;
assign input_328 = t0_000101001000;
assign input_329 = t0_000101001001;
assign input_330 = t0_000101001010;
assign input_331 = t0_000101001011;
assign input_332 = t0_000101001100;
assign input_333 = t0_000101001101;
assign input_334 = t0_000101001110;
assign input_335 = t0_000101001111;
assign input_336 = t0_000101010000;
assign input_337 = t0_000101010001;
assign input_338 = t0_000101010010;
assign input_339 = t0_000101010011;
assign input_340 = t0_000101010100;
assign input_341 = t0_000101010101;
assign input_342 = t0_000101010110;
assign input_343 = t0_000101010111;
assign input_344 = t0_000101011000;
assign input_345 = t0_000101011001;
assign input_346 = t0_000101011010;
assign input_347 = t0_000101011011;
assign input_348 = t0_000101011100;
assign input_349 = t0_000101011101;
assign input_350 = t0_000101011110;
assign input_351 = t0_000101011111;
assign input_352 = t0_000101100000;
assign input_353 = t0_000101100001;
assign input_354 = t0_000101100010;
assign input_355 = t0_000101100011;
assign input_356 = t0_000101100100;
assign input_357 = t0_000101100101;
assign input_358 = t0_000101100110;
assign input_359 = t0_000101100111;
assign input_360 = t0_000101101000;
assign input_361 = t0_000101101001;
assign input_362 = t0_000101101010;
assign input_363 = t0_000101101011;
assign input_364 = t0_000101101100;
assign input_365 = t0_000101101101;
assign input_366 = t0_000101101110;
assign input_367 = t0_000101101111;
assign input_368 = t0_000101110000;
assign input_369 = t0_000101110001;
assign input_370 = t0_000101110010;
assign input_371 = t0_000101110011;
assign input_372 = t0_000101110100;
assign input_373 = t0_000101110101;
assign input_374 = t0_000101110110;
assign input_375 = t0_000101110111;
assign input_376 = t0_000101111000;
assign input_377 = t0_000101111001;
assign input_378 = t0_000101111010;
assign input_379 = t0_000101111011;
assign input_380 = t0_000101111100;
assign input_381 = t0_000101111101;
assign input_382 = t0_000101111110;
assign input_383 = t0_000101111111;
assign input_384 = t0_000110000000;
assign input_385 = t0_000110000001;
assign input_386 = t0_000110000010;
assign input_387 = t0_000110000011;
assign input_388 = t0_000110000100;
assign input_389 = t0_000110000101;
assign input_390 = t0_000110000110;
assign input_391 = t0_000110000111;
assign input_392 = t0_000110001000;
assign input_393 = t0_000110001001;
assign input_394 = t0_000110001010;
assign input_395 = t0_000110001011;
assign input_396 = t0_000110001100;
assign input_397 = t0_000110001101;
assign input_398 = t0_000110001110;
assign input_399 = t0_000110001111;
assign input_400 = t0_000110010000;
assign input_401 = t0_000110010001;
assign input_402 = t0_000110010010;
assign input_403 = t0_000110010011;
assign input_404 = t0_000110010100;
assign input_405 = t0_000110010101;
assign input_406 = t0_000110010110;
assign input_407 = t0_000110010111;
assign input_408 = t0_000110011000;
assign input_409 = t0_000110011001;
assign input_410 = t0_000110011010;
assign input_411 = t0_000110011011;
assign input_412 = t0_000110011100;
assign input_413 = t0_000110011101;
assign input_414 = t0_000110011110;
assign input_415 = t0_000110011111;
assign input_416 = t0_000110100000;
assign input_417 = t0_000110100001;
assign input_418 = t0_000110100010;
assign input_419 = t0_000110100011;
assign input_420 = t0_000110100100;
assign input_421 = t0_000110100101;
assign input_422 = t0_000110100110;
assign input_423 = t0_000110100111;
assign input_424 = t0_000110101000;
assign input_425 = t0_000110101001;
assign input_426 = t0_000110101010;
assign input_427 = t0_000110101011;
assign input_428 = t0_000110101100;
assign input_429 = t0_000110101101;
assign input_430 = t0_000110101110;
assign input_431 = t0_000110101111;
assign input_432 = t0_000110110000;
assign input_433 = t0_000110110001;
assign input_434 = t0_000110110010;
assign input_435 = t0_000110110011;
assign input_436 = t0_000110110100;
assign input_437 = t0_000110110101;
assign input_438 = t0_000110110110;
assign input_439 = t0_000110110111;
assign input_440 = t0_000110111000;
assign input_441 = t0_000110111001;
assign input_442 = t0_000110111010;
assign input_443 = t0_000110111011;
assign input_444 = t0_000110111100;
assign input_445 = t0_000110111101;
assign input_446 = t0_000110111110;
assign input_447 = t0_000110111111;
assign input_448 = t0_000111000000;
assign input_449 = t0_000111000001;
assign input_450 = t0_000111000010;
assign input_451 = t0_000111000011;
assign input_452 = t0_000111000100;
assign input_453 = t0_000111000101;
assign input_454 = t0_000111000110;
assign input_455 = t0_000111000111;
assign input_456 = t0_000111001000;
assign input_457 = t0_000111001001;
assign input_458 = t0_000111001010;
assign input_459 = t0_000111001011;
assign input_460 = t0_000111001100;
assign input_461 = t0_000111001101;
assign input_462 = t0_000111001110;
assign input_463 = t0_000111001111;
assign input_464 = t0_000111010000;
assign input_465 = t0_000111010001;
assign input_466 = t0_000111010010;
assign input_467 = t0_000111010011;
assign input_468 = t0_000111010100;
assign input_469 = t0_000111010101;
assign input_470 = t0_000111010110;
assign input_471 = t0_000111010111;
assign input_472 = t0_000111011000;
assign input_473 = t0_000111011001;
assign input_474 = t0_000111011010;
assign input_475 = t0_000111011011;
assign input_476 = t0_000111011100;
assign input_477 = t0_000111011101;
assign input_478 = t0_000111011110;
assign input_479 = t0_000111011111;
assign input_480 = t0_000111100000;
assign input_481 = t0_000111100001;
assign input_482 = t0_000111100010;
assign input_483 = t0_000111100011;
assign input_484 = t0_000111100100;
assign input_485 = t0_000111100101;
assign input_486 = t0_000111100110;
assign input_487 = t0_000111100111;
assign input_488 = t0_000111101000;
assign input_489 = t0_000111101001;
assign input_490 = t0_000111101010;
assign input_491 = t0_000111101011;
assign input_492 = t0_000111101100;
assign input_493 = t0_000111101101;
assign input_494 = t0_000111101110;
assign input_495 = t0_000111101111;
assign input_496 = t0_000111110000;
assign input_497 = t0_000111110001;
assign input_498 = t0_000111110010;
assign input_499 = t0_000111110011;
assign input_500 = t0_000111110100;
assign input_501 = t0_000111110101;
assign input_502 = t0_000111110110;
assign input_503 = t0_000111110111;
assign input_504 = t0_000111111000;
assign input_505 = t0_000111111001;
assign input_506 = t0_000111111010;
assign input_507 = t0_000111111011;
assign input_508 = t0_000111111100;
assign input_509 = t0_000111111101;
assign input_510 = t0_000111111110;
assign input_511 = t0_000111111111;
assign input_512 = t0_001000000000;
assign input_513 = t0_001000000001;
assign input_514 = t0_001000000010;
assign input_515 = t0_001000000011;
assign input_516 = t0_001000000100;
assign input_517 = t0_001000000101;
assign input_518 = t0_001000000110;
assign input_519 = t0_001000000111;
assign input_520 = t0_001000001000;
assign input_521 = t0_001000001001;
assign input_522 = t0_001000001010;
assign input_523 = t0_001000001011;
assign input_524 = t0_001000001100;
assign input_525 = t0_001000001101;
assign input_526 = t0_001000001110;
assign input_527 = t0_001000001111;
assign input_528 = t0_001000010000;
assign input_529 = t0_001000010001;
assign input_530 = t0_001000010010;
assign input_531 = t0_001000010011;
assign input_532 = t0_001000010100;
assign input_533 = t0_001000010101;
assign input_534 = t0_001000010110;
assign input_535 = t0_001000010111;
assign input_536 = t0_001000011000;
assign input_537 = t0_001000011001;
assign input_538 = t0_001000011010;
assign input_539 = t0_001000011011;
assign input_540 = t0_001000011100;
assign input_541 = t0_001000011101;
assign input_542 = t0_001000011110;
assign input_543 = t0_001000011111;
assign input_544 = t0_001000100000;
assign input_545 = t0_001000100001;
assign input_546 = t0_001000100010;
assign input_547 = t0_001000100011;
assign input_548 = t0_001000100100;
assign input_549 = t0_001000100101;
assign input_550 = t0_001000100110;
assign input_551 = t0_001000100111;
assign input_552 = t0_001000101000;
assign input_553 = t0_001000101001;
assign input_554 = t0_001000101010;
assign input_555 = t0_001000101011;
assign input_556 = t0_001000101100;
assign input_557 = t0_001000101101;
assign input_558 = t0_001000101110;
assign input_559 = t0_001000101111;
assign input_560 = t0_001000110000;
assign input_561 = t0_001000110001;
assign input_562 = t0_001000110010;
assign input_563 = t0_001000110011;
assign input_564 = t0_001000110100;
assign input_565 = t0_001000110101;
assign input_566 = t0_001000110110;
assign input_567 = t0_001000110111;
assign input_568 = t0_001000111000;
assign input_569 = t0_001000111001;
assign input_570 = t0_001000111010;
assign input_571 = t0_001000111011;
assign input_572 = t0_001000111100;
assign input_573 = t0_001000111101;
assign input_574 = t0_001000111110;
assign input_575 = t0_001000111111;
assign input_576 = t0_001001000000;
assign input_577 = t0_001001000001;
assign input_578 = t0_001001000010;
assign input_579 = t0_001001000011;
assign input_580 = t0_001001000100;
assign input_581 = t0_001001000101;
assign input_582 = t0_001001000110;
assign input_583 = t0_001001000111;
assign input_584 = t0_001001001000;
assign input_585 = t0_001001001001;
assign input_586 = t0_001001001010;
assign input_587 = t0_001001001011;
assign input_588 = t0_001001001100;
assign input_589 = t0_001001001101;
assign input_590 = t0_001001001110;
assign input_591 = t0_001001001111;
assign input_592 = t0_001001010000;
assign input_593 = t0_001001010001;
assign input_594 = t0_001001010010;
assign input_595 = t0_001001010011;
assign input_596 = t0_001001010100;
assign input_597 = t0_001001010101;
assign input_598 = t0_001001010110;
assign input_599 = t0_001001010111;
assign input_600 = t0_001001011000;
assign input_601 = t0_001001011001;
assign input_602 = t0_001001011010;
assign input_603 = t0_001001011011;
assign input_604 = t0_001001011100;
assign input_605 = t0_001001011101;
assign input_606 = t0_001001011110;
assign input_607 = t0_001001011111;
assign input_608 = t0_001001100000;
assign input_609 = t0_001001100001;
assign input_610 = t0_001001100010;
assign input_611 = t0_001001100011;
assign input_612 = t0_001001100100;
assign input_613 = t0_001001100101;
assign input_614 = t0_001001100110;
assign input_615 = t0_001001100111;
assign input_616 = t0_001001101000;
assign input_617 = t0_001001101001;
assign input_618 = t0_001001101010;
assign input_619 = t0_001001101011;
assign input_620 = t0_001001101100;
assign input_621 = t0_001001101101;
assign input_622 = t0_001001101110;
assign input_623 = t0_001001101111;
assign input_624 = t0_001001110000;
assign input_625 = t0_001001110001;
assign input_626 = t0_001001110010;
assign input_627 = t0_001001110011;
assign input_628 = t0_001001110100;
assign input_629 = t0_001001110101;
assign input_630 = t0_001001110110;
assign input_631 = t0_001001110111;
assign input_632 = t0_001001111000;
assign input_633 = t0_001001111001;
assign input_634 = t0_001001111010;
assign input_635 = t0_001001111011;
assign input_636 = t0_001001111100;
assign input_637 = t0_001001111101;
assign input_638 = t0_001001111110;
assign input_639 = t0_001001111111;
assign input_640 = t0_001010000000;
assign input_641 = t0_001010000001;
assign input_642 = t0_001010000010;
assign input_643 = t0_001010000011;
assign input_644 = t0_001010000100;
assign input_645 = t0_001010000101;
assign input_646 = t0_001010000110;
assign input_647 = t0_001010000111;
assign input_648 = t0_001010001000;
assign input_649 = t0_001010001001;
assign input_650 = t0_001010001010;
assign input_651 = t0_001010001011;
assign input_652 = t0_001010001100;
assign input_653 = t0_001010001101;
assign input_654 = t0_001010001110;
assign input_655 = t0_001010001111;
assign input_656 = t0_001010010000;
assign input_657 = t0_001010010001;
assign input_658 = t0_001010010010;
assign input_659 = t0_001010010011;
assign input_660 = t0_001010010100;
assign input_661 = t0_001010010101;
assign input_662 = t0_001010010110;
assign input_663 = t0_001010010111;
assign input_664 = t0_001010011000;
assign input_665 = t0_001010011001;
assign input_666 = t0_001010011010;
assign input_667 = t0_001010011011;
assign input_668 = t0_001010011100;
assign input_669 = t0_001010011101;
assign input_670 = t0_001010011110;
assign input_671 = t0_001010011111;
assign input_672 = t0_001010100000;
assign input_673 = t0_001010100001;
assign input_674 = t0_001010100010;
assign input_675 = t0_001010100011;
assign input_676 = t0_001010100100;
assign input_677 = t0_001010100101;
assign input_678 = t0_001010100110;
assign input_679 = t0_001010100111;
assign input_680 = t0_001010101000;
assign input_681 = t0_001010101001;
assign input_682 = t0_001010101010;
assign input_683 = t0_001010101011;
assign input_684 = t0_001010101100;
assign input_685 = t0_001010101101;
assign input_686 = t0_001010101110;
assign input_687 = t0_001010101111;
assign input_688 = t0_001010110000;
assign input_689 = t0_001010110001;
assign input_690 = t0_001010110010;
assign input_691 = t0_001010110011;
assign input_692 = t0_001010110100;
assign input_693 = t0_001010110101;
assign input_694 = t0_001010110110;
assign input_695 = t0_001010110111;
assign input_696 = t0_001010111000;
assign input_697 = t0_001010111001;
assign input_698 = t0_001010111010;
assign input_699 = t0_001010111011;
assign input_700 = t0_001010111100;
assign input_701 = t0_001010111101;
assign input_702 = t0_001010111110;
assign input_703 = t0_001010111111;
assign input_704 = t0_001011000000;
assign input_705 = t0_001011000001;
assign input_706 = t0_001011000010;
assign input_707 = t0_001011000011;
assign input_708 = t0_001011000100;
assign input_709 = t0_001011000101;
assign input_710 = t0_001011000110;
assign input_711 = t0_001011000111;
assign input_712 = t0_001011001000;
assign input_713 = t0_001011001001;
assign input_714 = t0_001011001010;
assign input_715 = t0_001011001011;
assign input_716 = t0_001011001100;
assign input_717 = t0_001011001101;
assign input_718 = t0_001011001110;
assign input_719 = t0_001011001111;
assign input_720 = t0_001011010000;
assign input_721 = t0_001011010001;
assign input_722 = t0_001011010010;
assign input_723 = t0_001011010011;
assign input_724 = t0_001011010100;
assign input_725 = t0_001011010101;
assign input_726 = t0_001011010110;
assign input_727 = t0_001011010111;
assign input_728 = t0_001011011000;
assign input_729 = t0_001011011001;
assign input_730 = t0_001011011010;
assign input_731 = t0_001011011011;
assign input_732 = t0_001011011100;
assign input_733 = t0_001011011101;
assign input_734 = t0_001011011110;
assign input_735 = t0_001011011111;
assign input_736 = t0_001011100000;
assign input_737 = t0_001011100001;
assign input_738 = t0_001011100010;
assign input_739 = t0_001011100011;
assign input_740 = t0_001011100100;
assign input_741 = t0_001011100101;
assign input_742 = t0_001011100110;
assign input_743 = t0_001011100111;
assign input_744 = t0_001011101000;
assign input_745 = t0_001011101001;
assign input_746 = t0_001011101010;
assign input_747 = t0_001011101011;
assign input_748 = t0_001011101100;
assign input_749 = t0_001011101101;
assign input_750 = t0_001011101110;
assign input_751 = t0_001011101111;
assign input_752 = t0_001011110000;
assign input_753 = t0_001011110001;
assign input_754 = t0_001011110010;
assign input_755 = t0_001011110011;
assign input_756 = t0_001011110100;
assign input_757 = t0_001011110101;
assign input_758 = t0_001011110110;
assign input_759 = t0_001011110111;
assign input_760 = t0_001011111000;
assign input_761 = t0_001011111001;
assign input_762 = t0_001011111010;
assign input_763 = t0_001011111011;
assign input_764 = t0_001011111100;
assign input_765 = t0_001011111101;
assign input_766 = t0_001011111110;
assign input_767 = t0_001011111111;
assign input_768 = t0_001100000000;
assign input_769 = t0_001100000001;
assign input_770 = t0_001100000010;
assign input_771 = t0_001100000011;
assign input_772 = t0_001100000100;
assign input_773 = t0_001100000101;
assign input_774 = t0_001100000110;
assign input_775 = t0_001100000111;
assign input_776 = t0_001100001000;
assign input_777 = t0_001100001001;
assign input_778 = t0_001100001010;
assign input_779 = t0_001100001011;
assign input_780 = t0_001100001100;
assign input_781 = t0_001100001101;
assign input_782 = t0_001100001110;
assign input_783 = t0_001100001111;
assign input_784 = t0_001100010000;
assign input_785 = t0_001100010001;
assign input_786 = t0_001100010010;
assign input_787 = t0_001100010011;
assign input_788 = t0_001100010100;
assign input_789 = t0_001100010101;
assign input_790 = t0_001100010110;
assign input_791 = t0_001100010111;
assign input_792 = t0_001100011000;
assign input_793 = t0_001100011001;
assign input_794 = t0_001100011010;
assign input_795 = t0_001100011011;
assign input_796 = t0_001100011100;
assign input_797 = t0_001100011101;
assign input_798 = t0_001100011110;
assign input_799 = t0_001100011111;
assign input_800 = t0_001100100000;
assign input_801 = t0_001100100001;
assign input_802 = t0_001100100010;
assign input_803 = t0_001100100011;
assign input_804 = t0_001100100100;
assign input_805 = t0_001100100101;
assign input_806 = t0_001100100110;
assign input_807 = t0_001100100111;
assign input_808 = t0_001100101000;
assign input_809 = t0_001100101001;
assign input_810 = t0_001100101010;
assign input_811 = t0_001100101011;
assign input_812 = t0_001100101100;
assign input_813 = t0_001100101101;
assign input_814 = t0_001100101110;
assign input_815 = t0_001100101111;
assign input_816 = t0_001100110000;
assign input_817 = t0_001100110001;
assign input_818 = t0_001100110010;
assign input_819 = t0_001100110011;
assign input_820 = t0_001100110100;
assign input_821 = t0_001100110101;
assign input_822 = t0_001100110110;
assign input_823 = t0_001100110111;
assign input_824 = t0_001100111000;
assign input_825 = t0_001100111001;
assign input_826 = t0_001100111010;
assign input_827 = t0_001100111011;
assign input_828 = t0_001100111100;
assign input_829 = t0_001100111101;
assign input_830 = t0_001100111110;
assign input_831 = t0_001100111111;
assign input_832 = t0_001101000000;
assign input_833 = t0_001101000001;
assign input_834 = t0_001101000010;
assign input_835 = t0_001101000011;
assign input_836 = t0_001101000100;
assign input_837 = t0_001101000101;
assign input_838 = t0_001101000110;
assign input_839 = t0_001101000111;
assign input_840 = t0_001101001000;
assign input_841 = t0_001101001001;
assign input_842 = t0_001101001010;
assign input_843 = t0_001101001011;
assign input_844 = t0_001101001100;
assign input_845 = t0_001101001101;
assign input_846 = t0_001101001110;
assign input_847 = t0_001101001111;
assign input_848 = t0_001101010000;
assign input_849 = t0_001101010001;
assign input_850 = t0_001101010010;
assign input_851 = t0_001101010011;
assign input_852 = t0_001101010100;
assign input_853 = t0_001101010101;
assign input_854 = t0_001101010110;
assign input_855 = t0_001101010111;
assign input_856 = t0_001101011000;
assign input_857 = t0_001101011001;
assign input_858 = t0_001101011010;
assign input_859 = t0_001101011011;
assign input_860 = t0_001101011100;
assign input_861 = t0_001101011101;
assign input_862 = t0_001101011110;
assign input_863 = t0_001101011111;
assign input_864 = t0_001101100000;
assign input_865 = t0_001101100001;
assign input_866 = t0_001101100010;
assign input_867 = t0_001101100011;
assign input_868 = t0_001101100100;
assign input_869 = t0_001101100101;
assign input_870 = t0_001101100110;
assign input_871 = t0_001101100111;
assign input_872 = t0_001101101000;
assign input_873 = t0_001101101001;
assign input_874 = t0_001101101010;
assign input_875 = t0_001101101011;
assign input_876 = t0_001101101100;
assign input_877 = t0_001101101101;
assign input_878 = t0_001101101110;
assign input_879 = t0_001101101111;
assign input_880 = t0_001101110000;
assign input_881 = t0_001101110001;
assign input_882 = t0_001101110010;
assign input_883 = t0_001101110011;
assign input_884 = t0_001101110100;
assign input_885 = t0_001101110101;
assign input_886 = t0_001101110110;
assign input_887 = t0_001101110111;
assign input_888 = t0_001101111000;
assign input_889 = t0_001101111001;
assign input_890 = t0_001101111010;
assign input_891 = t0_001101111011;
assign input_892 = t0_001101111100;
assign input_893 = t0_001101111101;
assign input_894 = t0_001101111110;
assign input_895 = t0_001101111111;
assign input_896 = t0_001110000000;
assign input_897 = t0_001110000001;
assign input_898 = t0_001110000010;
assign input_899 = t0_001110000011;
assign input_900 = t0_001110000100;
assign input_901 = t0_001110000101;
assign input_902 = t0_001110000110;
assign input_903 = t0_001110000111;
assign input_904 = t0_001110001000;
assign input_905 = t0_001110001001;
assign input_906 = t0_001110001010;
assign input_907 = t0_001110001011;
assign input_908 = t0_001110001100;
assign input_909 = t0_001110001101;
assign input_910 = t0_001110001110;
assign input_911 = t0_001110001111;
assign input_912 = t0_001110010000;
assign input_913 = t0_001110010001;
assign input_914 = t0_001110010010;
assign input_915 = t0_001110010011;
assign input_916 = t0_001110010100;
assign input_917 = t0_001110010101;
assign input_918 = t0_001110010110;
assign input_919 = t0_001110010111;
assign input_920 = t0_001110011000;
assign input_921 = t0_001110011001;
assign input_922 = t0_001110011010;
assign input_923 = t0_001110011011;
assign input_924 = t0_001110011100;
assign input_925 = t0_001110011101;
assign input_926 = t0_001110011110;
assign input_927 = t0_001110011111;
assign input_928 = t0_001110100000;
assign input_929 = t0_001110100001;
assign input_930 = t0_001110100010;
assign input_931 = t0_001110100011;
assign input_932 = t0_001110100100;
assign input_933 = t0_001110100101;
assign input_934 = t0_001110100110;
assign input_935 = t0_001110100111;
assign input_936 = t0_001110101000;
assign input_937 = t0_001110101001;
assign input_938 = t0_001110101010;
assign input_939 = t0_001110101011;
assign input_940 = t0_001110101100;
assign input_941 = t0_001110101101;
assign input_942 = t0_001110101110;
assign input_943 = t0_001110101111;
assign input_944 = t0_001110110000;
assign input_945 = t0_001110110001;
assign input_946 = t0_001110110010;
assign input_947 = t0_001110110011;
assign input_948 = t0_001110110100;
assign input_949 = t0_001110110101;
assign input_950 = t0_001110110110;
assign input_951 = t0_001110110111;
assign input_952 = t0_001110111000;
assign input_953 = t0_001110111001;
assign input_954 = t0_001110111010;
assign input_955 = t0_001110111011;
assign input_956 = t0_001110111100;
assign input_957 = t0_001110111101;
assign input_958 = t0_001110111110;
assign input_959 = t0_001110111111;
assign input_960 = t0_001111000000;
assign input_961 = t0_001111000001;
assign input_962 = t0_001111000010;
assign input_963 = t0_001111000011;
assign input_964 = t0_001111000100;
assign input_965 = t0_001111000101;
assign input_966 = t0_001111000110;
assign input_967 = t0_001111000111;
assign input_968 = t0_001111001000;
assign input_969 = t0_001111001001;
assign input_970 = t0_001111001010;
assign input_971 = t0_001111001011;
assign input_972 = t0_001111001100;
assign input_973 = t0_001111001101;
assign input_974 = t0_001111001110;
assign input_975 = t0_001111001111;
assign input_976 = t0_001111010000;
assign input_977 = t0_001111010001;
assign input_978 = t0_001111010010;
assign input_979 = t0_001111010011;
assign input_980 = t0_001111010100;
assign input_981 = t0_001111010101;
assign input_982 = t0_001111010110;
assign input_983 = t0_001111010111;
assign input_984 = t0_001111011000;
assign input_985 = t0_001111011001;
assign input_986 = t0_001111011010;
assign input_987 = t0_001111011011;
assign input_988 = t0_001111011100;
assign input_989 = t0_001111011101;
assign input_990 = t0_001111011110;
assign input_991 = t0_001111011111;
assign input_992 = t0_001111100000;
assign input_993 = t0_001111100001;
assign input_994 = t0_001111100010;
assign input_995 = t0_001111100011;
assign input_996 = t0_001111100100;
assign input_997 = t0_001111100101;
assign input_998 = t0_001111100110;
assign input_999 = t0_001111100111;
assign input_1000 = t0_001111101000;
assign input_1001 = t0_001111101001;
assign input_1002 = t0_001111101010;
assign input_1003 = t0_001111101011;
assign input_1004 = t0_001111101100;
assign input_1005 = t0_001111101101;
assign input_1006 = t0_001111101110;
assign input_1007 = t0_001111101111;
assign input_1008 = t0_001111110000;
assign input_1009 = t0_001111110001;
assign input_1010 = t0_001111110010;
assign input_1011 = t0_001111110011;
assign input_1012 = t0_001111110100;
assign input_1013 = t0_001111110101;
assign input_1014 = t0_001111110110;
assign input_1015 = t0_001111110111;
assign input_1016 = t0_001111111000;
assign input_1017 = t0_001111111001;
assign input_1018 = t0_001111111010;
assign input_1019 = t0_001111111011;
assign input_1020 = t0_001111111100;
assign input_1021 = t0_001111111101;
assign input_1022 = t0_001111111110;
assign input_1023 = t0_001111111111;
assign input_1024 = t0_010000000000;
assign input_1025 = t0_010000000001;
assign input_1026 = t0_010000000010;
assign input_1027 = t0_010000000011;
assign input_1028 = t0_010000000100;
assign input_1029 = t0_010000000101;
assign input_1030 = t0_010000000110;
assign input_1031 = t0_010000000111;
assign input_1032 = t0_010000001000;
assign input_1033 = t0_010000001001;
assign input_1034 = t0_010000001010;
assign input_1035 = t0_010000001011;
assign input_1036 = t0_010000001100;
assign input_1037 = t0_010000001101;
assign input_1038 = t0_010000001110;
assign input_1039 = t0_010000001111;
assign input_1040 = t0_010000010000;
assign input_1041 = t0_010000010001;
assign input_1042 = t0_010000010010;
assign input_1043 = t0_010000010011;
assign input_1044 = t0_010000010100;
assign input_1045 = t0_010000010101;
assign input_1046 = t0_010000010110;
assign input_1047 = t0_010000010111;
assign input_1048 = t0_010000011000;
assign input_1049 = t0_010000011001;
assign input_1050 = t0_010000011010;
assign input_1051 = t0_010000011011;
assign input_1052 = t0_010000011100;
assign input_1053 = t0_010000011101;
assign input_1054 = t0_010000011110;
assign input_1055 = t0_010000011111;
assign input_1056 = t0_010000100000;
assign input_1057 = t0_010000100001;
assign input_1058 = t0_010000100010;
assign input_1059 = t0_010000100011;
assign input_1060 = t0_010000100100;
assign input_1061 = t0_010000100101;
assign input_1062 = t0_010000100110;
assign input_1063 = t0_010000100111;
assign input_1064 = t0_010000101000;
assign input_1065 = t0_010000101001;
assign input_1066 = t0_010000101010;
assign input_1067 = t0_010000101011;
assign input_1068 = t0_010000101100;
assign input_1069 = t0_010000101101;
assign input_1070 = t0_010000101110;
assign input_1071 = t0_010000101111;
assign input_1072 = t0_010000110000;
assign input_1073 = t0_010000110001;
assign input_1074 = t0_010000110010;
assign input_1075 = t0_010000110011;
assign input_1076 = t0_010000110100;
assign input_1077 = t0_010000110101;
assign input_1078 = t0_010000110110;
assign input_1079 = t0_010000110111;
assign input_1080 = t0_010000111000;
assign input_1081 = t0_010000111001;
assign input_1082 = t0_010000111010;
assign input_1083 = t0_010000111011;
assign input_1084 = t0_010000111100;
assign input_1085 = t0_010000111101;
assign input_1086 = t0_010000111110;
assign input_1087 = t0_010000111111;
assign input_1088 = t0_010001000000;
assign input_1089 = t0_010001000001;
assign input_1090 = t0_010001000010;
assign input_1091 = t0_010001000011;
assign input_1092 = t0_010001000100;
assign input_1093 = t0_010001000101;
assign input_1094 = t0_010001000110;
assign input_1095 = t0_010001000111;
assign input_1096 = t0_010001001000;
assign input_1097 = t0_010001001001;
assign input_1098 = t0_010001001010;
assign input_1099 = t0_010001001011;
assign input_1100 = t0_010001001100;
assign input_1101 = t0_010001001101;
assign input_1102 = t0_010001001110;
assign input_1103 = t0_010001001111;
assign input_1104 = t0_010001010000;
assign input_1105 = t0_010001010001;
assign input_1106 = t0_010001010010;
assign input_1107 = t0_010001010011;
assign input_1108 = t0_010001010100;
assign input_1109 = t0_010001010101;
assign input_1110 = t0_010001010110;
assign input_1111 = t0_010001010111;
assign input_1112 = t0_010001011000;
assign input_1113 = t0_010001011001;
assign input_1114 = t0_010001011010;
assign input_1115 = t0_010001011011;
assign input_1116 = t0_010001011100;
assign input_1117 = t0_010001011101;
assign input_1118 = t0_010001011110;
assign input_1119 = t0_010001011111;
assign input_1120 = t0_010001100000;
assign input_1121 = t0_010001100001;
assign input_1122 = t0_010001100010;
assign input_1123 = t0_010001100011;
assign input_1124 = t0_010001100100;
assign input_1125 = t0_010001100101;
assign input_1126 = t0_010001100110;
assign input_1127 = t0_010001100111;
assign input_1128 = t0_010001101000;
assign input_1129 = t0_010001101001;
assign input_1130 = t0_010001101010;
assign input_1131 = t0_010001101011;
assign input_1132 = t0_010001101100;
assign input_1133 = t0_010001101101;
assign input_1134 = t0_010001101110;
assign input_1135 = t0_010001101111;
assign input_1136 = t0_010001110000;
assign input_1137 = t0_010001110001;
assign input_1138 = t0_010001110010;
assign input_1139 = t0_010001110011;
assign input_1140 = t0_010001110100;
assign input_1141 = t0_010001110101;
assign input_1142 = t0_010001110110;
assign input_1143 = t0_010001110111;
assign input_1144 = t0_010001111000;
assign input_1145 = t0_010001111001;
assign input_1146 = t0_010001111010;
assign input_1147 = t0_010001111011;
assign input_1148 = t0_010001111100;
assign input_1149 = t0_010001111101;
assign input_1150 = t0_010001111110;
assign input_1151 = t0_010001111111;
assign input_1152 = t0_010010000000;
assign input_1153 = t0_010010000001;
assign input_1154 = t0_010010000010;
assign input_1155 = t0_010010000011;
assign input_1156 = t0_010010000100;
assign input_1157 = t0_010010000101;
assign input_1158 = t0_010010000110;
assign input_1159 = t0_010010000111;
assign input_1160 = t0_010010001000;
assign input_1161 = t0_010010001001;
assign input_1162 = t0_010010001010;
assign input_1163 = t0_010010001011;
assign input_1164 = t0_010010001100;
assign input_1165 = t0_010010001101;
assign input_1166 = t0_010010001110;
assign input_1167 = t0_010010001111;
assign input_1168 = t0_010010010000;
assign input_1169 = t0_010010010001;
assign input_1170 = t0_010010010010;
assign input_1171 = t0_010010010011;
assign input_1172 = t0_010010010100;
assign input_1173 = t0_010010010101;
assign input_1174 = t0_010010010110;
assign input_1175 = t0_010010010111;
assign input_1176 = t0_010010011000;
assign input_1177 = t0_010010011001;
assign input_1178 = t0_010010011010;
assign input_1179 = t0_010010011011;
assign input_1180 = t0_010010011100;
assign input_1181 = t0_010010011101;
assign input_1182 = t0_010010011110;
assign input_1183 = t0_010010011111;
assign input_1184 = t0_010010100000;
assign input_1185 = t0_010010100001;
assign input_1186 = t0_010010100010;
assign input_1187 = t0_010010100011;
assign input_1188 = t0_010010100100;
assign input_1189 = t0_010010100101;
assign input_1190 = t0_010010100110;
assign input_1191 = t0_010010100111;
assign input_1192 = t0_010010101000;
assign input_1193 = t0_010010101001;
assign input_1194 = t0_010010101010;
assign input_1195 = t0_010010101011;
assign input_1196 = t0_010010101100;
assign input_1197 = t0_010010101101;
assign input_1198 = t0_010010101110;
assign input_1199 = t0_010010101111;
assign input_1200 = t0_010010110000;
assign input_1201 = t0_010010110001;
assign input_1202 = t0_010010110010;
assign input_1203 = t0_010010110011;
assign input_1204 = t0_010010110100;
assign input_1205 = t0_010010110101;
assign input_1206 = t0_010010110110;
assign input_1207 = t0_010010110111;
assign input_1208 = t0_010010111000;
assign input_1209 = t0_010010111001;
assign input_1210 = t0_010010111010;
assign input_1211 = t0_010010111011;
assign input_1212 = t0_010010111100;
assign input_1213 = t0_010010111101;
assign input_1214 = t0_010010111110;
assign input_1215 = t0_010010111111;
assign input_1216 = t0_010011000000;
assign input_1217 = t0_010011000001;
assign input_1218 = t0_010011000010;
assign input_1219 = t0_010011000011;
assign input_1220 = t0_010011000100;
assign input_1221 = t0_010011000101;
assign input_1222 = t0_010011000110;
assign input_1223 = t0_010011000111;
assign input_1224 = t0_010011001000;
assign input_1225 = t0_010011001001;
assign input_1226 = t0_010011001010;
assign input_1227 = t0_010011001011;
assign input_1228 = t0_010011001100;
assign input_1229 = t0_010011001101;
assign input_1230 = t0_010011001110;
assign input_1231 = t0_010011001111;
assign input_1232 = t0_010011010000;
assign input_1233 = t0_010011010001;
assign input_1234 = t0_010011010010;
assign input_1235 = t0_010011010011;
assign input_1236 = t0_010011010100;
assign input_1237 = t0_010011010101;
assign input_1238 = t0_010011010110;
assign input_1239 = t0_010011010111;
assign input_1240 = t0_010011011000;
assign input_1241 = t0_010011011001;
assign input_1242 = t0_010011011010;
assign input_1243 = t0_010011011011;
assign input_1244 = t0_010011011100;
assign input_1245 = t0_010011011101;
assign input_1246 = t0_010011011110;
assign input_1247 = t0_010011011111;
assign input_1248 = t0_010011100000;
assign input_1249 = t0_010011100001;
assign input_1250 = t0_010011100010;
assign input_1251 = t0_010011100011;
assign input_1252 = t0_010011100100;
assign input_1253 = t0_010011100101;
assign input_1254 = t0_010011100110;
assign input_1255 = t0_010011100111;
assign input_1256 = t0_010011101000;
assign input_1257 = t0_010011101001;
assign input_1258 = t0_010011101010;
assign input_1259 = t0_010011101011;
assign input_1260 = t0_010011101100;
assign input_1261 = t0_010011101101;
assign input_1262 = t0_010011101110;
assign input_1263 = t0_010011101111;
assign input_1264 = t0_010011110000;
assign input_1265 = t0_010011110001;
assign input_1266 = t0_010011110010;
assign input_1267 = t0_010011110011;
assign input_1268 = t0_010011110100;
assign input_1269 = t0_010011110101;
assign input_1270 = t0_010011110110;
assign input_1271 = t0_010011110111;
assign input_1272 = t0_010011111000;
assign input_1273 = t0_010011111001;
assign input_1274 = t0_010011111010;
assign input_1275 = t0_010011111011;
assign input_1276 = t0_010011111100;
assign input_1277 = t0_010011111101;
assign input_1278 = t0_010011111110;
assign input_1279 = t0_010011111111;
assign input_1280 = t0_010100000000;
assign input_1281 = t0_010100000001;
assign input_1282 = t0_010100000010;
assign input_1283 = t0_010100000011;
assign input_1284 = t0_010100000100;
assign input_1285 = t0_010100000101;
assign input_1286 = t0_010100000110;
assign input_1287 = t0_010100000111;
assign input_1288 = t0_010100001000;
assign input_1289 = t0_010100001001;
assign input_1290 = t0_010100001010;
assign input_1291 = t0_010100001011;
assign input_1292 = t0_010100001100;
assign input_1293 = t0_010100001101;
assign input_1294 = t0_010100001110;
assign input_1295 = t0_010100001111;
assign input_1296 = t0_010100010000;
assign input_1297 = t0_010100010001;
assign input_1298 = t0_010100010010;
assign input_1299 = t0_010100010011;
assign input_1300 = t0_010100010100;
assign input_1301 = t0_010100010101;
assign input_1302 = t0_010100010110;
assign input_1303 = t0_010100010111;
assign input_1304 = t0_010100011000;
assign input_1305 = t0_010100011001;
assign input_1306 = t0_010100011010;
assign input_1307 = t0_010100011011;
assign input_1308 = t0_010100011100;
assign input_1309 = t0_010100011101;
assign input_1310 = t0_010100011110;
assign input_1311 = t0_010100011111;
assign input_1312 = t0_010100100000;
assign input_1313 = t0_010100100001;
assign input_1314 = t0_010100100010;
assign input_1315 = t0_010100100011;
assign input_1316 = t0_010100100100;
assign input_1317 = t0_010100100101;
assign input_1318 = t0_010100100110;
assign input_1319 = t0_010100100111;
assign input_1320 = t0_010100101000;
assign input_1321 = t0_010100101001;
assign input_1322 = t0_010100101010;
assign input_1323 = t0_010100101011;
assign input_1324 = t0_010100101100;
assign input_1325 = t0_010100101101;
assign input_1326 = t0_010100101110;
assign input_1327 = t0_010100101111;
assign input_1328 = t0_010100110000;
assign input_1329 = t0_010100110001;
assign input_1330 = t0_010100110010;
assign input_1331 = t0_010100110011;
assign input_1332 = t0_010100110100;
assign input_1333 = t0_010100110101;
assign input_1334 = t0_010100110110;
assign input_1335 = t0_010100110111;
assign input_1336 = t0_010100111000;
assign input_1337 = t0_010100111001;
assign input_1338 = t0_010100111010;
assign input_1339 = t0_010100111011;
assign input_1340 = t0_010100111100;
assign input_1341 = t0_010100111101;
assign input_1342 = t0_010100111110;
assign input_1343 = t0_010100111111;
assign input_1344 = t0_010101000000;
assign input_1345 = t0_010101000001;
assign input_1346 = t0_010101000010;
assign input_1347 = t0_010101000011;
assign input_1348 = t0_010101000100;
assign input_1349 = t0_010101000101;
assign input_1350 = t0_010101000110;
assign input_1351 = t0_010101000111;
assign input_1352 = t0_010101001000;
assign input_1353 = t0_010101001001;
assign input_1354 = t0_010101001010;
assign input_1355 = t0_010101001011;
assign input_1356 = t0_010101001100;
assign input_1357 = t0_010101001101;
assign input_1358 = t0_010101001110;
assign input_1359 = t0_010101001111;
assign input_1360 = t0_010101010000;
assign input_1361 = t0_010101010001;
assign input_1362 = t0_010101010010;
assign input_1363 = t0_010101010011;
assign input_1364 = t0_010101010100;
assign input_1365 = t0_010101010101;
assign input_1366 = t0_010101010110;
assign input_1367 = t0_010101010111;
assign input_1368 = t0_010101011000;
assign input_1369 = t0_010101011001;
assign input_1370 = t0_010101011010;
assign input_1371 = t0_010101011011;
assign input_1372 = t0_010101011100;
assign input_1373 = t0_010101011101;
assign input_1374 = t0_010101011110;
assign input_1375 = t0_010101011111;
assign input_1376 = t0_010101100000;
assign input_1377 = t0_010101100001;
assign input_1378 = t0_010101100010;
assign input_1379 = t0_010101100011;
assign input_1380 = t0_010101100100;
assign input_1381 = t0_010101100101;
assign input_1382 = t0_010101100110;
assign input_1383 = t0_010101100111;
assign input_1384 = t0_010101101000;
assign input_1385 = t0_010101101001;
assign input_1386 = t0_010101101010;
assign input_1387 = t0_010101101011;
assign input_1388 = t0_010101101100;
assign input_1389 = t0_010101101101;
assign input_1390 = t0_010101101110;
assign input_1391 = t0_010101101111;
assign input_1392 = t0_010101110000;
assign input_1393 = t0_010101110001;
assign input_1394 = t0_010101110010;
assign input_1395 = t0_010101110011;
assign input_1396 = t0_010101110100;
assign input_1397 = t0_010101110101;
assign input_1398 = t0_010101110110;
assign input_1399 = t0_010101110111;
assign input_1400 = t0_010101111000;
assign input_1401 = t0_010101111001;
assign input_1402 = t0_010101111010;
assign input_1403 = t0_010101111011;
assign input_1404 = t0_010101111100;
assign input_1405 = t0_010101111101;
assign input_1406 = t0_010101111110;
assign input_1407 = t0_010101111111;
assign input_1408 = t0_010110000000;
assign input_1409 = t0_010110000001;
assign input_1410 = t0_010110000010;
assign input_1411 = t0_010110000011;
assign input_1412 = t0_010110000100;
assign input_1413 = t0_010110000101;
assign input_1414 = t0_010110000110;
assign input_1415 = t0_010110000111;
assign input_1416 = t0_010110001000;
assign input_1417 = t0_010110001001;
assign input_1418 = t0_010110001010;
assign input_1419 = t0_010110001011;
assign input_1420 = t0_010110001100;
assign input_1421 = t0_010110001101;
assign input_1422 = t0_010110001110;
assign input_1423 = t0_010110001111;
assign input_1424 = t0_010110010000;
assign input_1425 = t0_010110010001;
assign input_1426 = t0_010110010010;
assign input_1427 = t0_010110010011;
assign input_1428 = t0_010110010100;
assign input_1429 = t0_010110010101;
assign input_1430 = t0_010110010110;
assign input_1431 = t0_010110010111;
assign input_1432 = t0_010110011000;
assign input_1433 = t0_010110011001;
assign input_1434 = t0_010110011010;
assign input_1435 = t0_010110011011;
assign input_1436 = t0_010110011100;
assign input_1437 = t0_010110011101;
assign input_1438 = t0_010110011110;
assign input_1439 = t0_010110011111;
assign input_1440 = t0_010110100000;
assign input_1441 = t0_010110100001;
assign input_1442 = t0_010110100010;
assign input_1443 = t0_010110100011;
assign input_1444 = t0_010110100100;
assign input_1445 = t0_010110100101;
assign input_1446 = t0_010110100110;
assign input_1447 = t0_010110100111;
assign input_1448 = t0_010110101000;
assign input_1449 = t0_010110101001;
assign input_1450 = t0_010110101010;
assign input_1451 = t0_010110101011;
assign input_1452 = t0_010110101100;
assign input_1453 = t0_010110101101;
assign input_1454 = t0_010110101110;
assign input_1455 = t0_010110101111;
assign input_1456 = t0_010110110000;
assign input_1457 = t0_010110110001;
assign input_1458 = t0_010110110010;
assign input_1459 = t0_010110110011;
assign input_1460 = t0_010110110100;
assign input_1461 = t0_010110110101;
assign input_1462 = t0_010110110110;
assign input_1463 = t0_010110110111;
assign input_1464 = t0_010110111000;
assign input_1465 = t0_010110111001;
assign input_1466 = t0_010110111010;
assign input_1467 = t0_010110111011;
assign input_1468 = t0_010110111100;
assign input_1469 = t0_010110111101;
assign input_1470 = t0_010110111110;
assign input_1471 = t0_010110111111;
assign input_1472 = t0_010111000000;
assign input_1473 = t0_010111000001;
assign input_1474 = t0_010111000010;
assign input_1475 = t0_010111000011;
assign input_1476 = t0_010111000100;
assign input_1477 = t0_010111000101;
assign input_1478 = t0_010111000110;
assign input_1479 = t0_010111000111;
assign input_1480 = t0_010111001000;
assign input_1481 = t0_010111001001;
assign input_1482 = t0_010111001010;
assign input_1483 = t0_010111001011;
assign input_1484 = t0_010111001100;
assign input_1485 = t0_010111001101;
assign input_1486 = t0_010111001110;
assign input_1487 = t0_010111001111;
assign input_1488 = t0_010111010000;
assign input_1489 = t0_010111010001;
assign input_1490 = t0_010111010010;
assign input_1491 = t0_010111010011;
assign input_1492 = t0_010111010100;
assign input_1493 = t0_010111010101;
assign input_1494 = t0_010111010110;
assign input_1495 = t0_010111010111;
assign input_1496 = t0_010111011000;
assign input_1497 = t0_010111011001;
assign input_1498 = t0_010111011010;
assign input_1499 = t0_010111011011;
assign input_1500 = t0_010111011100;
assign input_1501 = t0_010111011101;
assign input_1502 = t0_010111011110;
assign input_1503 = t0_010111011111;
assign input_1504 = t0_010111100000;
assign input_1505 = t0_010111100001;
assign input_1506 = t0_010111100010;
assign input_1507 = t0_010111100011;
assign input_1508 = t0_010111100100;
assign input_1509 = t0_010111100101;
assign input_1510 = t0_010111100110;
assign input_1511 = t0_010111100111;
assign input_1512 = t0_010111101000;
assign input_1513 = t0_010111101001;
assign input_1514 = t0_010111101010;
assign input_1515 = t0_010111101011;
assign input_1516 = t0_010111101100;
assign input_1517 = t0_010111101101;
assign input_1518 = t0_010111101110;
assign input_1519 = t0_010111101111;
assign input_1520 = t0_010111110000;
assign input_1521 = t0_010111110001;
assign input_1522 = t0_010111110010;
assign input_1523 = t0_010111110011;
assign input_1524 = t0_010111110100;
assign input_1525 = t0_010111110101;
assign input_1526 = t0_010111110110;
assign input_1527 = t0_010111110111;
assign input_1528 = t0_010111111000;
assign input_1529 = t0_010111111001;
assign input_1530 = t0_010111111010;
assign input_1531 = t0_010111111011;
assign input_1532 = t0_010111111100;
assign input_1533 = t0_010111111101;
assign input_1534 = t0_010111111110;
assign input_1535 = t0_010111111111;
assign input_1536 = t0_011000000000;
assign input_1537 = t0_011000000001;
assign input_1538 = t0_011000000010;
assign input_1539 = t0_011000000011;
assign input_1540 = t0_011000000100;
assign input_1541 = t0_011000000101;
assign input_1542 = t0_011000000110;
assign input_1543 = t0_011000000111;
assign input_1544 = t0_011000001000;
assign input_1545 = t0_011000001001;
assign input_1546 = t0_011000001010;
assign input_1547 = t0_011000001011;
assign input_1548 = t0_011000001100;
assign input_1549 = t0_011000001101;
assign input_1550 = t0_011000001110;
assign input_1551 = t0_011000001111;
assign input_1552 = t0_011000010000;
assign input_1553 = t0_011000010001;
assign input_1554 = t0_011000010010;
assign input_1555 = t0_011000010011;
assign input_1556 = t0_011000010100;
assign input_1557 = t0_011000010101;
assign input_1558 = t0_011000010110;
assign input_1559 = t0_011000010111;
assign input_1560 = t0_011000011000;
assign input_1561 = t0_011000011001;
assign input_1562 = t0_011000011010;
assign input_1563 = t0_011000011011;
assign input_1564 = t0_011000011100;
assign input_1565 = t0_011000011101;
assign input_1566 = t0_011000011110;
assign input_1567 = t0_011000011111;
assign input_1568 = t0_011000100000;
assign input_1569 = t0_011000100001;
assign input_1570 = t0_011000100010;
assign input_1571 = t0_011000100011;
assign input_1572 = t0_011000100100;
assign input_1573 = t0_011000100101;
assign input_1574 = t0_011000100110;
assign input_1575 = t0_011000100111;
assign input_1576 = t0_011000101000;
assign input_1577 = t0_011000101001;
assign input_1578 = t0_011000101010;
assign input_1579 = t0_011000101011;
assign input_1580 = t0_011000101100;
assign input_1581 = t0_011000101101;
assign input_1582 = t0_011000101110;
assign input_1583 = t0_011000101111;
assign input_1584 = t0_011000110000;
assign input_1585 = t0_011000110001;
assign input_1586 = t0_011000110010;
assign input_1587 = t0_011000110011;
assign input_1588 = t0_011000110100;
assign input_1589 = t0_011000110101;
assign input_1590 = t0_011000110110;
assign input_1591 = t0_011000110111;
assign input_1592 = t0_011000111000;
assign input_1593 = t0_011000111001;
assign input_1594 = t0_011000111010;
assign input_1595 = t0_011000111011;
assign input_1596 = t0_011000111100;
assign input_1597 = t0_011000111101;
assign input_1598 = t0_011000111110;
assign input_1599 = t0_011000111111;
assign input_1600 = t0_011001000000;
assign input_1601 = t0_011001000001;
assign input_1602 = t0_011001000010;
assign input_1603 = t0_011001000011;
assign input_1604 = t0_011001000100;
assign input_1605 = t0_011001000101;
assign input_1606 = t0_011001000110;
assign input_1607 = t0_011001000111;
assign input_1608 = t0_011001001000;
assign input_1609 = t0_011001001001;
assign input_1610 = t0_011001001010;
assign input_1611 = t0_011001001011;
assign input_1612 = t0_011001001100;
assign input_1613 = t0_011001001101;
assign input_1614 = t0_011001001110;
assign input_1615 = t0_011001001111;
assign input_1616 = t0_011001010000;
assign input_1617 = t0_011001010001;
assign input_1618 = t0_011001010010;
assign input_1619 = t0_011001010011;
assign input_1620 = t0_011001010100;
assign input_1621 = t0_011001010101;
assign input_1622 = t0_011001010110;
assign input_1623 = t0_011001010111;
assign input_1624 = t0_011001011000;
assign input_1625 = t0_011001011001;
assign input_1626 = t0_011001011010;
assign input_1627 = t0_011001011011;
assign input_1628 = t0_011001011100;
assign input_1629 = t0_011001011101;
assign input_1630 = t0_011001011110;
assign input_1631 = t0_011001011111;
assign input_1632 = t0_011001100000;
assign input_1633 = t0_011001100001;
assign input_1634 = t0_011001100010;
assign input_1635 = t0_011001100011;
assign input_1636 = t0_011001100100;
assign input_1637 = t0_011001100101;
assign input_1638 = t0_011001100110;
assign input_1639 = t0_011001100111;
assign input_1640 = t0_011001101000;
assign input_1641 = t0_011001101001;
assign input_1642 = t0_011001101010;
assign input_1643 = t0_011001101011;
assign input_1644 = t0_011001101100;
assign input_1645 = t0_011001101101;
assign input_1646 = t0_011001101110;
assign input_1647 = t0_011001101111;
assign input_1648 = t0_011001110000;
assign input_1649 = t0_011001110001;
assign input_1650 = t0_011001110010;
assign input_1651 = t0_011001110011;
assign input_1652 = t0_011001110100;
assign input_1653 = t0_011001110101;
assign input_1654 = t0_011001110110;
assign input_1655 = t0_011001110111;
assign input_1656 = t0_011001111000;
assign input_1657 = t0_011001111001;
assign input_1658 = t0_011001111010;
assign input_1659 = t0_011001111011;
assign input_1660 = t0_011001111100;
assign input_1661 = t0_011001111101;
assign input_1662 = t0_011001111110;
assign input_1663 = t0_011001111111;
assign input_1664 = t0_011010000000;
assign input_1665 = t0_011010000001;
assign input_1666 = t0_011010000010;
assign input_1667 = t0_011010000011;
assign input_1668 = t0_011010000100;
assign input_1669 = t0_011010000101;
assign input_1670 = t0_011010000110;
assign input_1671 = t0_011010000111;
assign input_1672 = t0_011010001000;
assign input_1673 = t0_011010001001;
assign input_1674 = t0_011010001010;
assign input_1675 = t0_011010001011;
assign input_1676 = t0_011010001100;
assign input_1677 = t0_011010001101;
assign input_1678 = t0_011010001110;
assign input_1679 = t0_011010001111;
assign input_1680 = t0_011010010000;
assign input_1681 = t0_011010010001;
assign input_1682 = t0_011010010010;
assign input_1683 = t0_011010010011;
assign input_1684 = t0_011010010100;
assign input_1685 = t0_011010010101;
assign input_1686 = t0_011010010110;
assign input_1687 = t0_011010010111;
assign input_1688 = t0_011010011000;
assign input_1689 = t0_011010011001;
assign input_1690 = t0_011010011010;
assign input_1691 = t0_011010011011;
assign input_1692 = t0_011010011100;
assign input_1693 = t0_011010011101;
assign input_1694 = t0_011010011110;
assign input_1695 = t0_011010011111;
assign input_1696 = t0_011010100000;
assign input_1697 = t0_011010100001;
assign input_1698 = t0_011010100010;
assign input_1699 = t0_011010100011;
assign input_1700 = t0_011010100100;
assign input_1701 = t0_011010100101;
assign input_1702 = t0_011010100110;
assign input_1703 = t0_011010100111;
assign input_1704 = t0_011010101000;
assign input_1705 = t0_011010101001;
assign input_1706 = t0_011010101010;
assign input_1707 = t0_011010101011;
assign input_1708 = t0_011010101100;
assign input_1709 = t0_011010101101;
assign input_1710 = t0_011010101110;
assign input_1711 = t0_011010101111;
assign input_1712 = t0_011010110000;
assign input_1713 = t0_011010110001;
assign input_1714 = t0_011010110010;
assign input_1715 = t0_011010110011;
assign input_1716 = t0_011010110100;
assign input_1717 = t0_011010110101;
assign input_1718 = t0_011010110110;
assign input_1719 = t0_011010110111;
assign input_1720 = t0_011010111000;
assign input_1721 = t0_011010111001;
assign input_1722 = t0_011010111010;
assign input_1723 = t0_011010111011;
assign input_1724 = t0_011010111100;
assign input_1725 = t0_011010111101;
assign input_1726 = t0_011010111110;
assign input_1727 = t0_011010111111;
assign input_1728 = t0_011011000000;
assign input_1729 = t0_011011000001;
assign input_1730 = t0_011011000010;
assign input_1731 = t0_011011000011;
assign input_1732 = t0_011011000100;
assign input_1733 = t0_011011000101;
assign input_1734 = t0_011011000110;
assign input_1735 = t0_011011000111;
assign input_1736 = t0_011011001000;
assign input_1737 = t0_011011001001;
assign input_1738 = t0_011011001010;
assign input_1739 = t0_011011001011;
assign input_1740 = t0_011011001100;
assign input_1741 = t0_011011001101;
assign input_1742 = t0_011011001110;
assign input_1743 = t0_011011001111;
assign input_1744 = t0_011011010000;
assign input_1745 = t0_011011010001;
assign input_1746 = t0_011011010010;
assign input_1747 = t0_011011010011;
assign input_1748 = t0_011011010100;
assign input_1749 = t0_011011010101;
assign input_1750 = t0_011011010110;
assign input_1751 = t0_011011010111;
assign input_1752 = t0_011011011000;
assign input_1753 = t0_011011011001;
assign input_1754 = t0_011011011010;
assign input_1755 = t0_011011011011;
assign input_1756 = t0_011011011100;
assign input_1757 = t0_011011011101;
assign input_1758 = t0_011011011110;
assign input_1759 = t0_011011011111;
assign input_1760 = t0_011011100000;
assign input_1761 = t0_011011100001;
assign input_1762 = t0_011011100010;
assign input_1763 = t0_011011100011;
assign input_1764 = t0_011011100100;
assign input_1765 = t0_011011100101;
assign input_1766 = t0_011011100110;
assign input_1767 = t0_011011100111;
assign input_1768 = t0_011011101000;
assign input_1769 = t0_011011101001;
assign input_1770 = t0_011011101010;
assign input_1771 = t0_011011101011;
assign input_1772 = t0_011011101100;
assign input_1773 = t0_011011101101;
assign input_1774 = t0_011011101110;
assign input_1775 = t0_011011101111;
assign input_1776 = t0_011011110000;
assign input_1777 = t0_011011110001;
assign input_1778 = t0_011011110010;
assign input_1779 = t0_011011110011;
assign input_1780 = t0_011011110100;
assign input_1781 = t0_011011110101;
assign input_1782 = t0_011011110110;
assign input_1783 = t0_011011110111;
assign input_1784 = t0_011011111000;
assign input_1785 = t0_011011111001;
assign input_1786 = t0_011011111010;
assign input_1787 = t0_011011111011;
assign input_1788 = t0_011011111100;
assign input_1789 = t0_011011111101;
assign input_1790 = t0_011011111110;
assign input_1791 = t0_011011111111;
assign input_1792 = t0_011100000000;
assign input_1793 = t0_011100000001;
assign input_1794 = t0_011100000010;
assign input_1795 = t0_011100000011;
assign input_1796 = t0_011100000100;
assign input_1797 = t0_011100000101;
assign input_1798 = t0_011100000110;
assign input_1799 = t0_011100000111;
assign input_1800 = t0_011100001000;
assign input_1801 = t0_011100001001;
assign input_1802 = t0_011100001010;
assign input_1803 = t0_011100001011;
assign input_1804 = t0_011100001100;
assign input_1805 = t0_011100001101;
assign input_1806 = t0_011100001110;
assign input_1807 = t0_011100001111;
assign input_1808 = t0_011100010000;
assign input_1809 = t0_011100010001;
assign input_1810 = t0_011100010010;
assign input_1811 = t0_011100010011;
assign input_1812 = t0_011100010100;
assign input_1813 = t0_011100010101;
assign input_1814 = t0_011100010110;
assign input_1815 = t0_011100010111;
assign input_1816 = t0_011100011000;
assign input_1817 = t0_011100011001;
assign input_1818 = t0_011100011010;
assign input_1819 = t0_011100011011;
assign input_1820 = t0_011100011100;
assign input_1821 = t0_011100011101;
assign input_1822 = t0_011100011110;
assign input_1823 = t0_011100011111;
assign input_1824 = t0_011100100000;
assign input_1825 = t0_011100100001;
assign input_1826 = t0_011100100010;
assign input_1827 = t0_011100100011;
assign input_1828 = t0_011100100100;
assign input_1829 = t0_011100100101;
assign input_1830 = t0_011100100110;
assign input_1831 = t0_011100100111;
assign input_1832 = t0_011100101000;
assign input_1833 = t0_011100101001;
assign input_1834 = t0_011100101010;
assign input_1835 = t0_011100101011;
assign input_1836 = t0_011100101100;
assign input_1837 = t0_011100101101;
assign input_1838 = t0_011100101110;
assign input_1839 = t0_011100101111;
assign input_1840 = t0_011100110000;
assign input_1841 = t0_011100110001;
assign input_1842 = t0_011100110010;
assign input_1843 = t0_011100110011;
assign input_1844 = t0_011100110100;
assign input_1845 = t0_011100110101;
assign input_1846 = t0_011100110110;
assign input_1847 = t0_011100110111;
assign input_1848 = t0_011100111000;
assign input_1849 = t0_011100111001;
assign input_1850 = t0_011100111010;
assign input_1851 = t0_011100111011;
assign input_1852 = t0_011100111100;
assign input_1853 = t0_011100111101;
assign input_1854 = t0_011100111110;
assign input_1855 = t0_011100111111;
assign input_1856 = t0_011101000000;
assign input_1857 = t0_011101000001;
assign input_1858 = t0_011101000010;
assign input_1859 = t0_011101000011;
assign input_1860 = t0_011101000100;
assign input_1861 = t0_011101000101;
assign input_1862 = t0_011101000110;
assign input_1863 = t0_011101000111;
assign input_1864 = t0_011101001000;
assign input_1865 = t0_011101001001;
assign input_1866 = t0_011101001010;
assign input_1867 = t0_011101001011;
assign input_1868 = t0_011101001100;
assign input_1869 = t0_011101001101;
assign input_1870 = t0_011101001110;
assign input_1871 = t0_011101001111;
assign input_1872 = t0_011101010000;
assign input_1873 = t0_011101010001;
assign input_1874 = t0_011101010010;
assign input_1875 = t0_011101010011;
assign input_1876 = t0_011101010100;
assign input_1877 = t0_011101010101;
assign input_1878 = t0_011101010110;
assign input_1879 = t0_011101010111;
assign input_1880 = t0_011101011000;
assign input_1881 = t0_011101011001;
assign input_1882 = t0_011101011010;
assign input_1883 = t0_011101011011;
assign input_1884 = t0_011101011100;
assign input_1885 = t0_011101011101;
assign input_1886 = t0_011101011110;
assign input_1887 = t0_011101011111;
assign input_1888 = t0_011101100000;
assign input_1889 = t0_011101100001;
assign input_1890 = t0_011101100010;
assign input_1891 = t0_011101100011;
assign input_1892 = t0_011101100100;
assign input_1893 = t0_011101100101;
assign input_1894 = t0_011101100110;
assign input_1895 = t0_011101100111;
assign input_1896 = t0_011101101000;
assign input_1897 = t0_011101101001;
assign input_1898 = t0_011101101010;
assign input_1899 = t0_011101101011;
assign input_1900 = t0_011101101100;
assign input_1901 = t0_011101101101;
assign input_1902 = t0_011101101110;
assign input_1903 = t0_011101101111;
assign input_1904 = t0_011101110000;
assign input_1905 = t0_011101110001;
assign input_1906 = t0_011101110010;
assign input_1907 = t0_011101110011;
assign input_1908 = t0_011101110100;
assign input_1909 = t0_011101110101;
assign input_1910 = t0_011101110110;
assign input_1911 = t0_011101110111;
assign input_1912 = t0_011101111000;
assign input_1913 = t0_011101111001;
assign input_1914 = t0_011101111010;
assign input_1915 = t0_011101111011;
assign input_1916 = t0_011101111100;
assign input_1917 = t0_011101111101;
assign input_1918 = t0_011101111110;
assign input_1919 = t0_011101111111;
assign input_1920 = t0_011110000000;
assign input_1921 = t0_011110000001;
assign input_1922 = t0_011110000010;
assign input_1923 = t0_011110000011;
assign input_1924 = t0_011110000100;
assign input_1925 = t0_011110000101;
assign input_1926 = t0_011110000110;
assign input_1927 = t0_011110000111;
assign input_1928 = t0_011110001000;
assign input_1929 = t0_011110001001;
assign input_1930 = t0_011110001010;
assign input_1931 = t0_011110001011;
assign input_1932 = t0_011110001100;
assign input_1933 = t0_011110001101;
assign input_1934 = t0_011110001110;
assign input_1935 = t0_011110001111;
assign input_1936 = t0_011110010000;
assign input_1937 = t0_011110010001;
assign input_1938 = t0_011110010010;
assign input_1939 = t0_011110010011;
assign input_1940 = t0_011110010100;
assign input_1941 = t0_011110010101;
assign input_1942 = t0_011110010110;
assign input_1943 = t0_011110010111;
assign input_1944 = t0_011110011000;
assign input_1945 = t0_011110011001;
assign input_1946 = t0_011110011010;
assign input_1947 = t0_011110011011;
assign input_1948 = t0_011110011100;
assign input_1949 = t0_011110011101;
assign input_1950 = t0_011110011110;
assign input_1951 = t0_011110011111;
assign input_1952 = t0_011110100000;
assign input_1953 = t0_011110100001;
assign input_1954 = t0_011110100010;
assign input_1955 = t0_011110100011;
assign input_1956 = t0_011110100100;
assign input_1957 = t0_011110100101;
assign input_1958 = t0_011110100110;
assign input_1959 = t0_011110100111;
assign input_1960 = t0_011110101000;
assign input_1961 = t0_011110101001;
assign input_1962 = t0_011110101010;
assign input_1963 = t0_011110101011;
assign input_1964 = t0_011110101100;
assign input_1965 = t0_011110101101;
assign input_1966 = t0_011110101110;
assign input_1967 = t0_011110101111;
assign input_1968 = t0_011110110000;
assign input_1969 = t0_011110110001;
assign input_1970 = t0_011110110010;
assign input_1971 = t0_011110110011;
assign input_1972 = t0_011110110100;
assign input_1973 = t0_011110110101;
assign input_1974 = t0_011110110110;
assign input_1975 = t0_011110110111;
assign input_1976 = t0_011110111000;
assign input_1977 = t0_011110111001;
assign input_1978 = t0_011110111010;
assign input_1979 = t0_011110111011;
assign input_1980 = t0_011110111100;
assign input_1981 = t0_011110111101;
assign input_1982 = t0_011110111110;
assign input_1983 = t0_011110111111;
assign input_1984 = t0_011111000000;
assign input_1985 = t0_011111000001;
assign input_1986 = t0_011111000010;
assign input_1987 = t0_011111000011;
assign input_1988 = t0_011111000100;
assign input_1989 = t0_011111000101;
assign input_1990 = t0_011111000110;
assign input_1991 = t0_011111000111;
assign input_1992 = t0_011111001000;
assign input_1993 = t0_011111001001;
assign input_1994 = t0_011111001010;
assign input_1995 = t0_011111001011;
assign input_1996 = t0_011111001100;
assign input_1997 = t0_011111001101;
assign input_1998 = t0_011111001110;
assign input_1999 = t0_011111001111;
assign input_2000 = t0_011111010000;
assign input_2001 = t0_011111010001;
assign input_2002 = t0_011111010010;
assign input_2003 = t0_011111010011;
assign input_2004 = t0_011111010100;
assign input_2005 = t0_011111010101;
assign input_2006 = t0_011111010110;
assign input_2007 = t0_011111010111;
assign input_2008 = t0_011111011000;
assign input_2009 = t0_011111011001;
assign input_2010 = t0_011111011010;
assign input_2011 = t0_011111011011;
assign input_2012 = t0_011111011100;
assign input_2013 = t0_011111011101;
assign input_2014 = t0_011111011110;
assign input_2015 = t0_011111011111;
assign input_2016 = t0_011111100000;
assign input_2017 = t0_011111100001;
assign input_2018 = t0_011111100010;
assign input_2019 = t0_011111100011;
assign input_2020 = t0_011111100100;
assign input_2021 = t0_011111100101;
assign input_2022 = t0_011111100110;
assign input_2023 = t0_011111100111;
assign input_2024 = t0_011111101000;
assign input_2025 = t0_011111101001;
assign input_2026 = t0_011111101010;
assign input_2027 = t0_011111101011;
assign input_2028 = t0_011111101100;
assign input_2029 = t0_011111101101;
assign input_2030 = t0_011111101110;
assign input_2031 = t0_011111101111;
assign input_2032 = t0_011111110000;
assign input_2033 = t0_011111110001;
assign input_2034 = t0_011111110010;
assign input_2035 = t0_011111110011;
assign input_2036 = t0_011111110100;
assign input_2037 = t0_011111110101;
assign input_2038 = t0_011111110110;
assign input_2039 = t0_011111110111;
assign input_2040 = t0_011111111000;
assign input_2041 = t0_011111111001;
assign input_2042 = t0_011111111010;
assign input_2043 = t0_011111111011;
assign input_2044 = t0_011111111100;
assign input_2045 = t0_011111111101;
assign input_2046 = t0_011111111110;
assign input_2047 = t0_011111111111;
endmodule
