module complete_bipartite_96_96 (
inout input_0,inout input_1,inout input_2,inout input_3,inout input_4,inout input_5,inout input_6,inout input_7,inout input_8,inout input_9,inout input_10,inout input_11,inout input_12,inout input_13,inout input_14,inout input_15,inout input_16,inout input_17,inout input_18,inout input_19,inout input_20,inout input_21,inout input_22,inout input_23,inout input_24,inout input_25,inout input_26,inout input_27,inout input_28,inout input_29,inout input_30,inout input_31,inout input_32,inout input_33,inout input_34,inout input_35,inout input_36,inout input_37,inout input_38,inout input_39,inout input_40,inout input_41,inout input_42,inout input_43,inout input_44,inout input_45,inout input_46,inout input_47,inout input_48,inout input_49,inout input_50,inout input_51,inout input_52,inout input_53,inout input_54,inout input_55,inout input_56,inout input_57,inout input_58,inout input_59,inout input_60,inout input_61,inout input_62,inout input_63,inout input_64,inout input_65,inout input_66,inout input_67,inout input_68,inout input_69,inout input_70,inout input_71,inout input_72,inout input_73,inout input_74,inout input_75,inout input_76,inout input_77,inout input_78,inout input_79,inout input_80,inout input_81,inout input_82,inout input_83,inout input_84,inout input_85,inout input_86,inout input_87,inout input_88,inout input_89,inout input_90,inout input_91,inout input_92,inout input_93,inout input_94,inout input_95,inout output_0,inout output_1,inout output_2,inout output_3,inout output_4,inout output_5,inout output_6,inout output_7,inout output_8,inout output_9,inout output_10,inout output_11,inout output_12,inout output_13,inout output_14,inout output_15,inout output_16,inout output_17,inout output_18,inout output_19,inout output_20,inout output_21,inout output_22,inout output_23,inout output_24,inout output_25,inout output_26,inout output_27,inout output_28,inout output_29,inout output_30,inout output_31,inout output_32,inout output_33,inout output_34,inout output_35,inout output_36,inout output_37,inout output_38,inout output_39,inout output_40,inout output_41,inout output_42,inout output_43,inout output_44,inout output_45,inout output_46,inout output_47,inout output_48,inout output_49,inout output_50,inout output_51,inout output_52,inout output_53,inout output_54,inout output_55,inout output_56,inout output_57,inout output_58,inout output_59,inout output_60,inout output_61,inout output_62,inout output_63,inout output_64,inout output_65,inout output_66,inout output_67,inout output_68,inout output_69,inout output_70,inout output_71,inout output_72,inout output_73,inout output_74,inout output_75,inout output_76,inout output_77,inout output_78,inout output_79,inout output_80,inout output_81,inout output_82,inout output_83,inout output_84,inout output_85,inout output_86,inout output_87,inout output_88,inout output_89,inout output_90,inout output_91,inout output_92,inout output_93,inout output_94,inout output_95
);
assign output_0 = input_0;
assign output_1 = input_0;
assign output_2 = input_0;
assign output_3 = input_0;
assign output_4 = input_0;
assign output_5 = input_0;
assign output_6 = input_0;
assign output_7 = input_0;
assign output_8 = input_0;
assign output_9 = input_0;
assign output_10 = input_0;
assign output_11 = input_0;
assign output_12 = input_0;
assign output_13 = input_0;
assign output_14 = input_0;
assign output_15 = input_0;
assign output_16 = input_0;
assign output_17 = input_0;
assign output_18 = input_0;
assign output_19 = input_0;
assign output_20 = input_0;
assign output_21 = input_0;
assign output_22 = input_0;
assign output_23 = input_0;
assign output_24 = input_0;
assign output_25 = input_0;
assign output_26 = input_0;
assign output_27 = input_0;
assign output_28 = input_0;
assign output_29 = input_0;
assign output_30 = input_0;
assign output_31 = input_0;
assign output_32 = input_0;
assign output_33 = input_0;
assign output_34 = input_0;
assign output_35 = input_0;
assign output_36 = input_0;
assign output_37 = input_0;
assign output_38 = input_0;
assign output_39 = input_0;
assign output_40 = input_0;
assign output_41 = input_0;
assign output_42 = input_0;
assign output_43 = input_0;
assign output_44 = input_0;
assign output_45 = input_0;
assign output_46 = input_0;
assign output_47 = input_0;
assign output_48 = input_0;
assign output_49 = input_0;
assign output_50 = input_0;
assign output_51 = input_0;
assign output_52 = input_0;
assign output_53 = input_0;
assign output_54 = input_0;
assign output_55 = input_0;
assign output_56 = input_0;
assign output_57 = input_0;
assign output_58 = input_0;
assign output_59 = input_0;
assign output_60 = input_0;
assign output_61 = input_0;
assign output_62 = input_0;
assign output_63 = input_0;
assign output_64 = input_0;
assign output_65 = input_0;
assign output_66 = input_0;
assign output_67 = input_0;
assign output_68 = input_0;
assign output_69 = input_0;
assign output_70 = input_0;
assign output_71 = input_0;
assign output_72 = input_0;
assign output_73 = input_0;
assign output_74 = input_0;
assign output_75 = input_0;
assign output_76 = input_0;
assign output_77 = input_0;
assign output_78 = input_0;
assign output_79 = input_0;
assign output_80 = input_0;
assign output_81 = input_0;
assign output_82 = input_0;
assign output_83 = input_0;
assign output_84 = input_0;
assign output_85 = input_0;
assign output_86 = input_0;
assign output_87 = input_0;
assign output_88 = input_0;
assign output_89 = input_0;
assign output_90 = input_0;
assign output_91 = input_0;
assign output_92 = input_0;
assign output_93 = input_0;
assign output_94 = input_0;
assign output_95 = input_0;
assign output_0 = input_1;
assign output_1 = input_1;
assign output_2 = input_1;
assign output_3 = input_1;
assign output_4 = input_1;
assign output_5 = input_1;
assign output_6 = input_1;
assign output_7 = input_1;
assign output_8 = input_1;
assign output_9 = input_1;
assign output_10 = input_1;
assign output_11 = input_1;
assign output_12 = input_1;
assign output_13 = input_1;
assign output_14 = input_1;
assign output_15 = input_1;
assign output_16 = input_1;
assign output_17 = input_1;
assign output_18 = input_1;
assign output_19 = input_1;
assign output_20 = input_1;
assign output_21 = input_1;
assign output_22 = input_1;
assign output_23 = input_1;
assign output_24 = input_1;
assign output_25 = input_1;
assign output_26 = input_1;
assign output_27 = input_1;
assign output_28 = input_1;
assign output_29 = input_1;
assign output_30 = input_1;
assign output_31 = input_1;
assign output_32 = input_1;
assign output_33 = input_1;
assign output_34 = input_1;
assign output_35 = input_1;
assign output_36 = input_1;
assign output_37 = input_1;
assign output_38 = input_1;
assign output_39 = input_1;
assign output_40 = input_1;
assign output_41 = input_1;
assign output_42 = input_1;
assign output_43 = input_1;
assign output_44 = input_1;
assign output_45 = input_1;
assign output_46 = input_1;
assign output_47 = input_1;
assign output_48 = input_1;
assign output_49 = input_1;
assign output_50 = input_1;
assign output_51 = input_1;
assign output_52 = input_1;
assign output_53 = input_1;
assign output_54 = input_1;
assign output_55 = input_1;
assign output_56 = input_1;
assign output_57 = input_1;
assign output_58 = input_1;
assign output_59 = input_1;
assign output_60 = input_1;
assign output_61 = input_1;
assign output_62 = input_1;
assign output_63 = input_1;
assign output_64 = input_1;
assign output_65 = input_1;
assign output_66 = input_1;
assign output_67 = input_1;
assign output_68 = input_1;
assign output_69 = input_1;
assign output_70 = input_1;
assign output_71 = input_1;
assign output_72 = input_1;
assign output_73 = input_1;
assign output_74 = input_1;
assign output_75 = input_1;
assign output_76 = input_1;
assign output_77 = input_1;
assign output_78 = input_1;
assign output_79 = input_1;
assign output_80 = input_1;
assign output_81 = input_1;
assign output_82 = input_1;
assign output_83 = input_1;
assign output_84 = input_1;
assign output_85 = input_1;
assign output_86 = input_1;
assign output_87 = input_1;
assign output_88 = input_1;
assign output_89 = input_1;
assign output_90 = input_1;
assign output_91 = input_1;
assign output_92 = input_1;
assign output_93 = input_1;
assign output_94 = input_1;
assign output_95 = input_1;
assign output_0 = input_2;
assign output_1 = input_2;
assign output_2 = input_2;
assign output_3 = input_2;
assign output_4 = input_2;
assign output_5 = input_2;
assign output_6 = input_2;
assign output_7 = input_2;
assign output_8 = input_2;
assign output_9 = input_2;
assign output_10 = input_2;
assign output_11 = input_2;
assign output_12 = input_2;
assign output_13 = input_2;
assign output_14 = input_2;
assign output_15 = input_2;
assign output_16 = input_2;
assign output_17 = input_2;
assign output_18 = input_2;
assign output_19 = input_2;
assign output_20 = input_2;
assign output_21 = input_2;
assign output_22 = input_2;
assign output_23 = input_2;
assign output_24 = input_2;
assign output_25 = input_2;
assign output_26 = input_2;
assign output_27 = input_2;
assign output_28 = input_2;
assign output_29 = input_2;
assign output_30 = input_2;
assign output_31 = input_2;
assign output_32 = input_2;
assign output_33 = input_2;
assign output_34 = input_2;
assign output_35 = input_2;
assign output_36 = input_2;
assign output_37 = input_2;
assign output_38 = input_2;
assign output_39 = input_2;
assign output_40 = input_2;
assign output_41 = input_2;
assign output_42 = input_2;
assign output_43 = input_2;
assign output_44 = input_2;
assign output_45 = input_2;
assign output_46 = input_2;
assign output_47 = input_2;
assign output_48 = input_2;
assign output_49 = input_2;
assign output_50 = input_2;
assign output_51 = input_2;
assign output_52 = input_2;
assign output_53 = input_2;
assign output_54 = input_2;
assign output_55 = input_2;
assign output_56 = input_2;
assign output_57 = input_2;
assign output_58 = input_2;
assign output_59 = input_2;
assign output_60 = input_2;
assign output_61 = input_2;
assign output_62 = input_2;
assign output_63 = input_2;
assign output_64 = input_2;
assign output_65 = input_2;
assign output_66 = input_2;
assign output_67 = input_2;
assign output_68 = input_2;
assign output_69 = input_2;
assign output_70 = input_2;
assign output_71 = input_2;
assign output_72 = input_2;
assign output_73 = input_2;
assign output_74 = input_2;
assign output_75 = input_2;
assign output_76 = input_2;
assign output_77 = input_2;
assign output_78 = input_2;
assign output_79 = input_2;
assign output_80 = input_2;
assign output_81 = input_2;
assign output_82 = input_2;
assign output_83 = input_2;
assign output_84 = input_2;
assign output_85 = input_2;
assign output_86 = input_2;
assign output_87 = input_2;
assign output_88 = input_2;
assign output_89 = input_2;
assign output_90 = input_2;
assign output_91 = input_2;
assign output_92 = input_2;
assign output_93 = input_2;
assign output_94 = input_2;
assign output_95 = input_2;
assign output_0 = input_3;
assign output_1 = input_3;
assign output_2 = input_3;
assign output_3 = input_3;
assign output_4 = input_3;
assign output_5 = input_3;
assign output_6 = input_3;
assign output_7 = input_3;
assign output_8 = input_3;
assign output_9 = input_3;
assign output_10 = input_3;
assign output_11 = input_3;
assign output_12 = input_3;
assign output_13 = input_3;
assign output_14 = input_3;
assign output_15 = input_3;
assign output_16 = input_3;
assign output_17 = input_3;
assign output_18 = input_3;
assign output_19 = input_3;
assign output_20 = input_3;
assign output_21 = input_3;
assign output_22 = input_3;
assign output_23 = input_3;
assign output_24 = input_3;
assign output_25 = input_3;
assign output_26 = input_3;
assign output_27 = input_3;
assign output_28 = input_3;
assign output_29 = input_3;
assign output_30 = input_3;
assign output_31 = input_3;
assign output_32 = input_3;
assign output_33 = input_3;
assign output_34 = input_3;
assign output_35 = input_3;
assign output_36 = input_3;
assign output_37 = input_3;
assign output_38 = input_3;
assign output_39 = input_3;
assign output_40 = input_3;
assign output_41 = input_3;
assign output_42 = input_3;
assign output_43 = input_3;
assign output_44 = input_3;
assign output_45 = input_3;
assign output_46 = input_3;
assign output_47 = input_3;
assign output_48 = input_3;
assign output_49 = input_3;
assign output_50 = input_3;
assign output_51 = input_3;
assign output_52 = input_3;
assign output_53 = input_3;
assign output_54 = input_3;
assign output_55 = input_3;
assign output_56 = input_3;
assign output_57 = input_3;
assign output_58 = input_3;
assign output_59 = input_3;
assign output_60 = input_3;
assign output_61 = input_3;
assign output_62 = input_3;
assign output_63 = input_3;
assign output_64 = input_3;
assign output_65 = input_3;
assign output_66 = input_3;
assign output_67 = input_3;
assign output_68 = input_3;
assign output_69 = input_3;
assign output_70 = input_3;
assign output_71 = input_3;
assign output_72 = input_3;
assign output_73 = input_3;
assign output_74 = input_3;
assign output_75 = input_3;
assign output_76 = input_3;
assign output_77 = input_3;
assign output_78 = input_3;
assign output_79 = input_3;
assign output_80 = input_3;
assign output_81 = input_3;
assign output_82 = input_3;
assign output_83 = input_3;
assign output_84 = input_3;
assign output_85 = input_3;
assign output_86 = input_3;
assign output_87 = input_3;
assign output_88 = input_3;
assign output_89 = input_3;
assign output_90 = input_3;
assign output_91 = input_3;
assign output_92 = input_3;
assign output_93 = input_3;
assign output_94 = input_3;
assign output_95 = input_3;
assign output_0 = input_4;
assign output_1 = input_4;
assign output_2 = input_4;
assign output_3 = input_4;
assign output_4 = input_4;
assign output_5 = input_4;
assign output_6 = input_4;
assign output_7 = input_4;
assign output_8 = input_4;
assign output_9 = input_4;
assign output_10 = input_4;
assign output_11 = input_4;
assign output_12 = input_4;
assign output_13 = input_4;
assign output_14 = input_4;
assign output_15 = input_4;
assign output_16 = input_4;
assign output_17 = input_4;
assign output_18 = input_4;
assign output_19 = input_4;
assign output_20 = input_4;
assign output_21 = input_4;
assign output_22 = input_4;
assign output_23 = input_4;
assign output_24 = input_4;
assign output_25 = input_4;
assign output_26 = input_4;
assign output_27 = input_4;
assign output_28 = input_4;
assign output_29 = input_4;
assign output_30 = input_4;
assign output_31 = input_4;
assign output_32 = input_4;
assign output_33 = input_4;
assign output_34 = input_4;
assign output_35 = input_4;
assign output_36 = input_4;
assign output_37 = input_4;
assign output_38 = input_4;
assign output_39 = input_4;
assign output_40 = input_4;
assign output_41 = input_4;
assign output_42 = input_4;
assign output_43 = input_4;
assign output_44 = input_4;
assign output_45 = input_4;
assign output_46 = input_4;
assign output_47 = input_4;
assign output_48 = input_4;
assign output_49 = input_4;
assign output_50 = input_4;
assign output_51 = input_4;
assign output_52 = input_4;
assign output_53 = input_4;
assign output_54 = input_4;
assign output_55 = input_4;
assign output_56 = input_4;
assign output_57 = input_4;
assign output_58 = input_4;
assign output_59 = input_4;
assign output_60 = input_4;
assign output_61 = input_4;
assign output_62 = input_4;
assign output_63 = input_4;
assign output_64 = input_4;
assign output_65 = input_4;
assign output_66 = input_4;
assign output_67 = input_4;
assign output_68 = input_4;
assign output_69 = input_4;
assign output_70 = input_4;
assign output_71 = input_4;
assign output_72 = input_4;
assign output_73 = input_4;
assign output_74 = input_4;
assign output_75 = input_4;
assign output_76 = input_4;
assign output_77 = input_4;
assign output_78 = input_4;
assign output_79 = input_4;
assign output_80 = input_4;
assign output_81 = input_4;
assign output_82 = input_4;
assign output_83 = input_4;
assign output_84 = input_4;
assign output_85 = input_4;
assign output_86 = input_4;
assign output_87 = input_4;
assign output_88 = input_4;
assign output_89 = input_4;
assign output_90 = input_4;
assign output_91 = input_4;
assign output_92 = input_4;
assign output_93 = input_4;
assign output_94 = input_4;
assign output_95 = input_4;
assign output_0 = input_5;
assign output_1 = input_5;
assign output_2 = input_5;
assign output_3 = input_5;
assign output_4 = input_5;
assign output_5 = input_5;
assign output_6 = input_5;
assign output_7 = input_5;
assign output_8 = input_5;
assign output_9 = input_5;
assign output_10 = input_5;
assign output_11 = input_5;
assign output_12 = input_5;
assign output_13 = input_5;
assign output_14 = input_5;
assign output_15 = input_5;
assign output_16 = input_5;
assign output_17 = input_5;
assign output_18 = input_5;
assign output_19 = input_5;
assign output_20 = input_5;
assign output_21 = input_5;
assign output_22 = input_5;
assign output_23 = input_5;
assign output_24 = input_5;
assign output_25 = input_5;
assign output_26 = input_5;
assign output_27 = input_5;
assign output_28 = input_5;
assign output_29 = input_5;
assign output_30 = input_5;
assign output_31 = input_5;
assign output_32 = input_5;
assign output_33 = input_5;
assign output_34 = input_5;
assign output_35 = input_5;
assign output_36 = input_5;
assign output_37 = input_5;
assign output_38 = input_5;
assign output_39 = input_5;
assign output_40 = input_5;
assign output_41 = input_5;
assign output_42 = input_5;
assign output_43 = input_5;
assign output_44 = input_5;
assign output_45 = input_5;
assign output_46 = input_5;
assign output_47 = input_5;
assign output_48 = input_5;
assign output_49 = input_5;
assign output_50 = input_5;
assign output_51 = input_5;
assign output_52 = input_5;
assign output_53 = input_5;
assign output_54 = input_5;
assign output_55 = input_5;
assign output_56 = input_5;
assign output_57 = input_5;
assign output_58 = input_5;
assign output_59 = input_5;
assign output_60 = input_5;
assign output_61 = input_5;
assign output_62 = input_5;
assign output_63 = input_5;
assign output_64 = input_5;
assign output_65 = input_5;
assign output_66 = input_5;
assign output_67 = input_5;
assign output_68 = input_5;
assign output_69 = input_5;
assign output_70 = input_5;
assign output_71 = input_5;
assign output_72 = input_5;
assign output_73 = input_5;
assign output_74 = input_5;
assign output_75 = input_5;
assign output_76 = input_5;
assign output_77 = input_5;
assign output_78 = input_5;
assign output_79 = input_5;
assign output_80 = input_5;
assign output_81 = input_5;
assign output_82 = input_5;
assign output_83 = input_5;
assign output_84 = input_5;
assign output_85 = input_5;
assign output_86 = input_5;
assign output_87 = input_5;
assign output_88 = input_5;
assign output_89 = input_5;
assign output_90 = input_5;
assign output_91 = input_5;
assign output_92 = input_5;
assign output_93 = input_5;
assign output_94 = input_5;
assign output_95 = input_5;
assign output_0 = input_6;
assign output_1 = input_6;
assign output_2 = input_6;
assign output_3 = input_6;
assign output_4 = input_6;
assign output_5 = input_6;
assign output_6 = input_6;
assign output_7 = input_6;
assign output_8 = input_6;
assign output_9 = input_6;
assign output_10 = input_6;
assign output_11 = input_6;
assign output_12 = input_6;
assign output_13 = input_6;
assign output_14 = input_6;
assign output_15 = input_6;
assign output_16 = input_6;
assign output_17 = input_6;
assign output_18 = input_6;
assign output_19 = input_6;
assign output_20 = input_6;
assign output_21 = input_6;
assign output_22 = input_6;
assign output_23 = input_6;
assign output_24 = input_6;
assign output_25 = input_6;
assign output_26 = input_6;
assign output_27 = input_6;
assign output_28 = input_6;
assign output_29 = input_6;
assign output_30 = input_6;
assign output_31 = input_6;
assign output_32 = input_6;
assign output_33 = input_6;
assign output_34 = input_6;
assign output_35 = input_6;
assign output_36 = input_6;
assign output_37 = input_6;
assign output_38 = input_6;
assign output_39 = input_6;
assign output_40 = input_6;
assign output_41 = input_6;
assign output_42 = input_6;
assign output_43 = input_6;
assign output_44 = input_6;
assign output_45 = input_6;
assign output_46 = input_6;
assign output_47 = input_6;
assign output_48 = input_6;
assign output_49 = input_6;
assign output_50 = input_6;
assign output_51 = input_6;
assign output_52 = input_6;
assign output_53 = input_6;
assign output_54 = input_6;
assign output_55 = input_6;
assign output_56 = input_6;
assign output_57 = input_6;
assign output_58 = input_6;
assign output_59 = input_6;
assign output_60 = input_6;
assign output_61 = input_6;
assign output_62 = input_6;
assign output_63 = input_6;
assign output_64 = input_6;
assign output_65 = input_6;
assign output_66 = input_6;
assign output_67 = input_6;
assign output_68 = input_6;
assign output_69 = input_6;
assign output_70 = input_6;
assign output_71 = input_6;
assign output_72 = input_6;
assign output_73 = input_6;
assign output_74 = input_6;
assign output_75 = input_6;
assign output_76 = input_6;
assign output_77 = input_6;
assign output_78 = input_6;
assign output_79 = input_6;
assign output_80 = input_6;
assign output_81 = input_6;
assign output_82 = input_6;
assign output_83 = input_6;
assign output_84 = input_6;
assign output_85 = input_6;
assign output_86 = input_6;
assign output_87 = input_6;
assign output_88 = input_6;
assign output_89 = input_6;
assign output_90 = input_6;
assign output_91 = input_6;
assign output_92 = input_6;
assign output_93 = input_6;
assign output_94 = input_6;
assign output_95 = input_6;
assign output_0 = input_7;
assign output_1 = input_7;
assign output_2 = input_7;
assign output_3 = input_7;
assign output_4 = input_7;
assign output_5 = input_7;
assign output_6 = input_7;
assign output_7 = input_7;
assign output_8 = input_7;
assign output_9 = input_7;
assign output_10 = input_7;
assign output_11 = input_7;
assign output_12 = input_7;
assign output_13 = input_7;
assign output_14 = input_7;
assign output_15 = input_7;
assign output_16 = input_7;
assign output_17 = input_7;
assign output_18 = input_7;
assign output_19 = input_7;
assign output_20 = input_7;
assign output_21 = input_7;
assign output_22 = input_7;
assign output_23 = input_7;
assign output_24 = input_7;
assign output_25 = input_7;
assign output_26 = input_7;
assign output_27 = input_7;
assign output_28 = input_7;
assign output_29 = input_7;
assign output_30 = input_7;
assign output_31 = input_7;
assign output_32 = input_7;
assign output_33 = input_7;
assign output_34 = input_7;
assign output_35 = input_7;
assign output_36 = input_7;
assign output_37 = input_7;
assign output_38 = input_7;
assign output_39 = input_7;
assign output_40 = input_7;
assign output_41 = input_7;
assign output_42 = input_7;
assign output_43 = input_7;
assign output_44 = input_7;
assign output_45 = input_7;
assign output_46 = input_7;
assign output_47 = input_7;
assign output_48 = input_7;
assign output_49 = input_7;
assign output_50 = input_7;
assign output_51 = input_7;
assign output_52 = input_7;
assign output_53 = input_7;
assign output_54 = input_7;
assign output_55 = input_7;
assign output_56 = input_7;
assign output_57 = input_7;
assign output_58 = input_7;
assign output_59 = input_7;
assign output_60 = input_7;
assign output_61 = input_7;
assign output_62 = input_7;
assign output_63 = input_7;
assign output_64 = input_7;
assign output_65 = input_7;
assign output_66 = input_7;
assign output_67 = input_7;
assign output_68 = input_7;
assign output_69 = input_7;
assign output_70 = input_7;
assign output_71 = input_7;
assign output_72 = input_7;
assign output_73 = input_7;
assign output_74 = input_7;
assign output_75 = input_7;
assign output_76 = input_7;
assign output_77 = input_7;
assign output_78 = input_7;
assign output_79 = input_7;
assign output_80 = input_7;
assign output_81 = input_7;
assign output_82 = input_7;
assign output_83 = input_7;
assign output_84 = input_7;
assign output_85 = input_7;
assign output_86 = input_7;
assign output_87 = input_7;
assign output_88 = input_7;
assign output_89 = input_7;
assign output_90 = input_7;
assign output_91 = input_7;
assign output_92 = input_7;
assign output_93 = input_7;
assign output_94 = input_7;
assign output_95 = input_7;
assign output_0 = input_8;
assign output_1 = input_8;
assign output_2 = input_8;
assign output_3 = input_8;
assign output_4 = input_8;
assign output_5 = input_8;
assign output_6 = input_8;
assign output_7 = input_8;
assign output_8 = input_8;
assign output_9 = input_8;
assign output_10 = input_8;
assign output_11 = input_8;
assign output_12 = input_8;
assign output_13 = input_8;
assign output_14 = input_8;
assign output_15 = input_8;
assign output_16 = input_8;
assign output_17 = input_8;
assign output_18 = input_8;
assign output_19 = input_8;
assign output_20 = input_8;
assign output_21 = input_8;
assign output_22 = input_8;
assign output_23 = input_8;
assign output_24 = input_8;
assign output_25 = input_8;
assign output_26 = input_8;
assign output_27 = input_8;
assign output_28 = input_8;
assign output_29 = input_8;
assign output_30 = input_8;
assign output_31 = input_8;
assign output_32 = input_8;
assign output_33 = input_8;
assign output_34 = input_8;
assign output_35 = input_8;
assign output_36 = input_8;
assign output_37 = input_8;
assign output_38 = input_8;
assign output_39 = input_8;
assign output_40 = input_8;
assign output_41 = input_8;
assign output_42 = input_8;
assign output_43 = input_8;
assign output_44 = input_8;
assign output_45 = input_8;
assign output_46 = input_8;
assign output_47 = input_8;
assign output_48 = input_8;
assign output_49 = input_8;
assign output_50 = input_8;
assign output_51 = input_8;
assign output_52 = input_8;
assign output_53 = input_8;
assign output_54 = input_8;
assign output_55 = input_8;
assign output_56 = input_8;
assign output_57 = input_8;
assign output_58 = input_8;
assign output_59 = input_8;
assign output_60 = input_8;
assign output_61 = input_8;
assign output_62 = input_8;
assign output_63 = input_8;
assign output_64 = input_8;
assign output_65 = input_8;
assign output_66 = input_8;
assign output_67 = input_8;
assign output_68 = input_8;
assign output_69 = input_8;
assign output_70 = input_8;
assign output_71 = input_8;
assign output_72 = input_8;
assign output_73 = input_8;
assign output_74 = input_8;
assign output_75 = input_8;
assign output_76 = input_8;
assign output_77 = input_8;
assign output_78 = input_8;
assign output_79 = input_8;
assign output_80 = input_8;
assign output_81 = input_8;
assign output_82 = input_8;
assign output_83 = input_8;
assign output_84 = input_8;
assign output_85 = input_8;
assign output_86 = input_8;
assign output_87 = input_8;
assign output_88 = input_8;
assign output_89 = input_8;
assign output_90 = input_8;
assign output_91 = input_8;
assign output_92 = input_8;
assign output_93 = input_8;
assign output_94 = input_8;
assign output_95 = input_8;
assign output_0 = input_9;
assign output_1 = input_9;
assign output_2 = input_9;
assign output_3 = input_9;
assign output_4 = input_9;
assign output_5 = input_9;
assign output_6 = input_9;
assign output_7 = input_9;
assign output_8 = input_9;
assign output_9 = input_9;
assign output_10 = input_9;
assign output_11 = input_9;
assign output_12 = input_9;
assign output_13 = input_9;
assign output_14 = input_9;
assign output_15 = input_9;
assign output_16 = input_9;
assign output_17 = input_9;
assign output_18 = input_9;
assign output_19 = input_9;
assign output_20 = input_9;
assign output_21 = input_9;
assign output_22 = input_9;
assign output_23 = input_9;
assign output_24 = input_9;
assign output_25 = input_9;
assign output_26 = input_9;
assign output_27 = input_9;
assign output_28 = input_9;
assign output_29 = input_9;
assign output_30 = input_9;
assign output_31 = input_9;
assign output_32 = input_9;
assign output_33 = input_9;
assign output_34 = input_9;
assign output_35 = input_9;
assign output_36 = input_9;
assign output_37 = input_9;
assign output_38 = input_9;
assign output_39 = input_9;
assign output_40 = input_9;
assign output_41 = input_9;
assign output_42 = input_9;
assign output_43 = input_9;
assign output_44 = input_9;
assign output_45 = input_9;
assign output_46 = input_9;
assign output_47 = input_9;
assign output_48 = input_9;
assign output_49 = input_9;
assign output_50 = input_9;
assign output_51 = input_9;
assign output_52 = input_9;
assign output_53 = input_9;
assign output_54 = input_9;
assign output_55 = input_9;
assign output_56 = input_9;
assign output_57 = input_9;
assign output_58 = input_9;
assign output_59 = input_9;
assign output_60 = input_9;
assign output_61 = input_9;
assign output_62 = input_9;
assign output_63 = input_9;
assign output_64 = input_9;
assign output_65 = input_9;
assign output_66 = input_9;
assign output_67 = input_9;
assign output_68 = input_9;
assign output_69 = input_9;
assign output_70 = input_9;
assign output_71 = input_9;
assign output_72 = input_9;
assign output_73 = input_9;
assign output_74 = input_9;
assign output_75 = input_9;
assign output_76 = input_9;
assign output_77 = input_9;
assign output_78 = input_9;
assign output_79 = input_9;
assign output_80 = input_9;
assign output_81 = input_9;
assign output_82 = input_9;
assign output_83 = input_9;
assign output_84 = input_9;
assign output_85 = input_9;
assign output_86 = input_9;
assign output_87 = input_9;
assign output_88 = input_9;
assign output_89 = input_9;
assign output_90 = input_9;
assign output_91 = input_9;
assign output_92 = input_9;
assign output_93 = input_9;
assign output_94 = input_9;
assign output_95 = input_9;
assign output_0 = input_10;
assign output_1 = input_10;
assign output_2 = input_10;
assign output_3 = input_10;
assign output_4 = input_10;
assign output_5 = input_10;
assign output_6 = input_10;
assign output_7 = input_10;
assign output_8 = input_10;
assign output_9 = input_10;
assign output_10 = input_10;
assign output_11 = input_10;
assign output_12 = input_10;
assign output_13 = input_10;
assign output_14 = input_10;
assign output_15 = input_10;
assign output_16 = input_10;
assign output_17 = input_10;
assign output_18 = input_10;
assign output_19 = input_10;
assign output_20 = input_10;
assign output_21 = input_10;
assign output_22 = input_10;
assign output_23 = input_10;
assign output_24 = input_10;
assign output_25 = input_10;
assign output_26 = input_10;
assign output_27 = input_10;
assign output_28 = input_10;
assign output_29 = input_10;
assign output_30 = input_10;
assign output_31 = input_10;
assign output_32 = input_10;
assign output_33 = input_10;
assign output_34 = input_10;
assign output_35 = input_10;
assign output_36 = input_10;
assign output_37 = input_10;
assign output_38 = input_10;
assign output_39 = input_10;
assign output_40 = input_10;
assign output_41 = input_10;
assign output_42 = input_10;
assign output_43 = input_10;
assign output_44 = input_10;
assign output_45 = input_10;
assign output_46 = input_10;
assign output_47 = input_10;
assign output_48 = input_10;
assign output_49 = input_10;
assign output_50 = input_10;
assign output_51 = input_10;
assign output_52 = input_10;
assign output_53 = input_10;
assign output_54 = input_10;
assign output_55 = input_10;
assign output_56 = input_10;
assign output_57 = input_10;
assign output_58 = input_10;
assign output_59 = input_10;
assign output_60 = input_10;
assign output_61 = input_10;
assign output_62 = input_10;
assign output_63 = input_10;
assign output_64 = input_10;
assign output_65 = input_10;
assign output_66 = input_10;
assign output_67 = input_10;
assign output_68 = input_10;
assign output_69 = input_10;
assign output_70 = input_10;
assign output_71 = input_10;
assign output_72 = input_10;
assign output_73 = input_10;
assign output_74 = input_10;
assign output_75 = input_10;
assign output_76 = input_10;
assign output_77 = input_10;
assign output_78 = input_10;
assign output_79 = input_10;
assign output_80 = input_10;
assign output_81 = input_10;
assign output_82 = input_10;
assign output_83 = input_10;
assign output_84 = input_10;
assign output_85 = input_10;
assign output_86 = input_10;
assign output_87 = input_10;
assign output_88 = input_10;
assign output_89 = input_10;
assign output_90 = input_10;
assign output_91 = input_10;
assign output_92 = input_10;
assign output_93 = input_10;
assign output_94 = input_10;
assign output_95 = input_10;
assign output_0 = input_11;
assign output_1 = input_11;
assign output_2 = input_11;
assign output_3 = input_11;
assign output_4 = input_11;
assign output_5 = input_11;
assign output_6 = input_11;
assign output_7 = input_11;
assign output_8 = input_11;
assign output_9 = input_11;
assign output_10 = input_11;
assign output_11 = input_11;
assign output_12 = input_11;
assign output_13 = input_11;
assign output_14 = input_11;
assign output_15 = input_11;
assign output_16 = input_11;
assign output_17 = input_11;
assign output_18 = input_11;
assign output_19 = input_11;
assign output_20 = input_11;
assign output_21 = input_11;
assign output_22 = input_11;
assign output_23 = input_11;
assign output_24 = input_11;
assign output_25 = input_11;
assign output_26 = input_11;
assign output_27 = input_11;
assign output_28 = input_11;
assign output_29 = input_11;
assign output_30 = input_11;
assign output_31 = input_11;
assign output_32 = input_11;
assign output_33 = input_11;
assign output_34 = input_11;
assign output_35 = input_11;
assign output_36 = input_11;
assign output_37 = input_11;
assign output_38 = input_11;
assign output_39 = input_11;
assign output_40 = input_11;
assign output_41 = input_11;
assign output_42 = input_11;
assign output_43 = input_11;
assign output_44 = input_11;
assign output_45 = input_11;
assign output_46 = input_11;
assign output_47 = input_11;
assign output_48 = input_11;
assign output_49 = input_11;
assign output_50 = input_11;
assign output_51 = input_11;
assign output_52 = input_11;
assign output_53 = input_11;
assign output_54 = input_11;
assign output_55 = input_11;
assign output_56 = input_11;
assign output_57 = input_11;
assign output_58 = input_11;
assign output_59 = input_11;
assign output_60 = input_11;
assign output_61 = input_11;
assign output_62 = input_11;
assign output_63 = input_11;
assign output_64 = input_11;
assign output_65 = input_11;
assign output_66 = input_11;
assign output_67 = input_11;
assign output_68 = input_11;
assign output_69 = input_11;
assign output_70 = input_11;
assign output_71 = input_11;
assign output_72 = input_11;
assign output_73 = input_11;
assign output_74 = input_11;
assign output_75 = input_11;
assign output_76 = input_11;
assign output_77 = input_11;
assign output_78 = input_11;
assign output_79 = input_11;
assign output_80 = input_11;
assign output_81 = input_11;
assign output_82 = input_11;
assign output_83 = input_11;
assign output_84 = input_11;
assign output_85 = input_11;
assign output_86 = input_11;
assign output_87 = input_11;
assign output_88 = input_11;
assign output_89 = input_11;
assign output_90 = input_11;
assign output_91 = input_11;
assign output_92 = input_11;
assign output_93 = input_11;
assign output_94 = input_11;
assign output_95 = input_11;
assign output_0 = input_12;
assign output_1 = input_12;
assign output_2 = input_12;
assign output_3 = input_12;
assign output_4 = input_12;
assign output_5 = input_12;
assign output_6 = input_12;
assign output_7 = input_12;
assign output_8 = input_12;
assign output_9 = input_12;
assign output_10 = input_12;
assign output_11 = input_12;
assign output_12 = input_12;
assign output_13 = input_12;
assign output_14 = input_12;
assign output_15 = input_12;
assign output_16 = input_12;
assign output_17 = input_12;
assign output_18 = input_12;
assign output_19 = input_12;
assign output_20 = input_12;
assign output_21 = input_12;
assign output_22 = input_12;
assign output_23 = input_12;
assign output_24 = input_12;
assign output_25 = input_12;
assign output_26 = input_12;
assign output_27 = input_12;
assign output_28 = input_12;
assign output_29 = input_12;
assign output_30 = input_12;
assign output_31 = input_12;
assign output_32 = input_12;
assign output_33 = input_12;
assign output_34 = input_12;
assign output_35 = input_12;
assign output_36 = input_12;
assign output_37 = input_12;
assign output_38 = input_12;
assign output_39 = input_12;
assign output_40 = input_12;
assign output_41 = input_12;
assign output_42 = input_12;
assign output_43 = input_12;
assign output_44 = input_12;
assign output_45 = input_12;
assign output_46 = input_12;
assign output_47 = input_12;
assign output_48 = input_12;
assign output_49 = input_12;
assign output_50 = input_12;
assign output_51 = input_12;
assign output_52 = input_12;
assign output_53 = input_12;
assign output_54 = input_12;
assign output_55 = input_12;
assign output_56 = input_12;
assign output_57 = input_12;
assign output_58 = input_12;
assign output_59 = input_12;
assign output_60 = input_12;
assign output_61 = input_12;
assign output_62 = input_12;
assign output_63 = input_12;
assign output_64 = input_12;
assign output_65 = input_12;
assign output_66 = input_12;
assign output_67 = input_12;
assign output_68 = input_12;
assign output_69 = input_12;
assign output_70 = input_12;
assign output_71 = input_12;
assign output_72 = input_12;
assign output_73 = input_12;
assign output_74 = input_12;
assign output_75 = input_12;
assign output_76 = input_12;
assign output_77 = input_12;
assign output_78 = input_12;
assign output_79 = input_12;
assign output_80 = input_12;
assign output_81 = input_12;
assign output_82 = input_12;
assign output_83 = input_12;
assign output_84 = input_12;
assign output_85 = input_12;
assign output_86 = input_12;
assign output_87 = input_12;
assign output_88 = input_12;
assign output_89 = input_12;
assign output_90 = input_12;
assign output_91 = input_12;
assign output_92 = input_12;
assign output_93 = input_12;
assign output_94 = input_12;
assign output_95 = input_12;
assign output_0 = input_13;
assign output_1 = input_13;
assign output_2 = input_13;
assign output_3 = input_13;
assign output_4 = input_13;
assign output_5 = input_13;
assign output_6 = input_13;
assign output_7 = input_13;
assign output_8 = input_13;
assign output_9 = input_13;
assign output_10 = input_13;
assign output_11 = input_13;
assign output_12 = input_13;
assign output_13 = input_13;
assign output_14 = input_13;
assign output_15 = input_13;
assign output_16 = input_13;
assign output_17 = input_13;
assign output_18 = input_13;
assign output_19 = input_13;
assign output_20 = input_13;
assign output_21 = input_13;
assign output_22 = input_13;
assign output_23 = input_13;
assign output_24 = input_13;
assign output_25 = input_13;
assign output_26 = input_13;
assign output_27 = input_13;
assign output_28 = input_13;
assign output_29 = input_13;
assign output_30 = input_13;
assign output_31 = input_13;
assign output_32 = input_13;
assign output_33 = input_13;
assign output_34 = input_13;
assign output_35 = input_13;
assign output_36 = input_13;
assign output_37 = input_13;
assign output_38 = input_13;
assign output_39 = input_13;
assign output_40 = input_13;
assign output_41 = input_13;
assign output_42 = input_13;
assign output_43 = input_13;
assign output_44 = input_13;
assign output_45 = input_13;
assign output_46 = input_13;
assign output_47 = input_13;
assign output_48 = input_13;
assign output_49 = input_13;
assign output_50 = input_13;
assign output_51 = input_13;
assign output_52 = input_13;
assign output_53 = input_13;
assign output_54 = input_13;
assign output_55 = input_13;
assign output_56 = input_13;
assign output_57 = input_13;
assign output_58 = input_13;
assign output_59 = input_13;
assign output_60 = input_13;
assign output_61 = input_13;
assign output_62 = input_13;
assign output_63 = input_13;
assign output_64 = input_13;
assign output_65 = input_13;
assign output_66 = input_13;
assign output_67 = input_13;
assign output_68 = input_13;
assign output_69 = input_13;
assign output_70 = input_13;
assign output_71 = input_13;
assign output_72 = input_13;
assign output_73 = input_13;
assign output_74 = input_13;
assign output_75 = input_13;
assign output_76 = input_13;
assign output_77 = input_13;
assign output_78 = input_13;
assign output_79 = input_13;
assign output_80 = input_13;
assign output_81 = input_13;
assign output_82 = input_13;
assign output_83 = input_13;
assign output_84 = input_13;
assign output_85 = input_13;
assign output_86 = input_13;
assign output_87 = input_13;
assign output_88 = input_13;
assign output_89 = input_13;
assign output_90 = input_13;
assign output_91 = input_13;
assign output_92 = input_13;
assign output_93 = input_13;
assign output_94 = input_13;
assign output_95 = input_13;
assign output_0 = input_14;
assign output_1 = input_14;
assign output_2 = input_14;
assign output_3 = input_14;
assign output_4 = input_14;
assign output_5 = input_14;
assign output_6 = input_14;
assign output_7 = input_14;
assign output_8 = input_14;
assign output_9 = input_14;
assign output_10 = input_14;
assign output_11 = input_14;
assign output_12 = input_14;
assign output_13 = input_14;
assign output_14 = input_14;
assign output_15 = input_14;
assign output_16 = input_14;
assign output_17 = input_14;
assign output_18 = input_14;
assign output_19 = input_14;
assign output_20 = input_14;
assign output_21 = input_14;
assign output_22 = input_14;
assign output_23 = input_14;
assign output_24 = input_14;
assign output_25 = input_14;
assign output_26 = input_14;
assign output_27 = input_14;
assign output_28 = input_14;
assign output_29 = input_14;
assign output_30 = input_14;
assign output_31 = input_14;
assign output_32 = input_14;
assign output_33 = input_14;
assign output_34 = input_14;
assign output_35 = input_14;
assign output_36 = input_14;
assign output_37 = input_14;
assign output_38 = input_14;
assign output_39 = input_14;
assign output_40 = input_14;
assign output_41 = input_14;
assign output_42 = input_14;
assign output_43 = input_14;
assign output_44 = input_14;
assign output_45 = input_14;
assign output_46 = input_14;
assign output_47 = input_14;
assign output_48 = input_14;
assign output_49 = input_14;
assign output_50 = input_14;
assign output_51 = input_14;
assign output_52 = input_14;
assign output_53 = input_14;
assign output_54 = input_14;
assign output_55 = input_14;
assign output_56 = input_14;
assign output_57 = input_14;
assign output_58 = input_14;
assign output_59 = input_14;
assign output_60 = input_14;
assign output_61 = input_14;
assign output_62 = input_14;
assign output_63 = input_14;
assign output_64 = input_14;
assign output_65 = input_14;
assign output_66 = input_14;
assign output_67 = input_14;
assign output_68 = input_14;
assign output_69 = input_14;
assign output_70 = input_14;
assign output_71 = input_14;
assign output_72 = input_14;
assign output_73 = input_14;
assign output_74 = input_14;
assign output_75 = input_14;
assign output_76 = input_14;
assign output_77 = input_14;
assign output_78 = input_14;
assign output_79 = input_14;
assign output_80 = input_14;
assign output_81 = input_14;
assign output_82 = input_14;
assign output_83 = input_14;
assign output_84 = input_14;
assign output_85 = input_14;
assign output_86 = input_14;
assign output_87 = input_14;
assign output_88 = input_14;
assign output_89 = input_14;
assign output_90 = input_14;
assign output_91 = input_14;
assign output_92 = input_14;
assign output_93 = input_14;
assign output_94 = input_14;
assign output_95 = input_14;
assign output_0 = input_15;
assign output_1 = input_15;
assign output_2 = input_15;
assign output_3 = input_15;
assign output_4 = input_15;
assign output_5 = input_15;
assign output_6 = input_15;
assign output_7 = input_15;
assign output_8 = input_15;
assign output_9 = input_15;
assign output_10 = input_15;
assign output_11 = input_15;
assign output_12 = input_15;
assign output_13 = input_15;
assign output_14 = input_15;
assign output_15 = input_15;
assign output_16 = input_15;
assign output_17 = input_15;
assign output_18 = input_15;
assign output_19 = input_15;
assign output_20 = input_15;
assign output_21 = input_15;
assign output_22 = input_15;
assign output_23 = input_15;
assign output_24 = input_15;
assign output_25 = input_15;
assign output_26 = input_15;
assign output_27 = input_15;
assign output_28 = input_15;
assign output_29 = input_15;
assign output_30 = input_15;
assign output_31 = input_15;
assign output_32 = input_15;
assign output_33 = input_15;
assign output_34 = input_15;
assign output_35 = input_15;
assign output_36 = input_15;
assign output_37 = input_15;
assign output_38 = input_15;
assign output_39 = input_15;
assign output_40 = input_15;
assign output_41 = input_15;
assign output_42 = input_15;
assign output_43 = input_15;
assign output_44 = input_15;
assign output_45 = input_15;
assign output_46 = input_15;
assign output_47 = input_15;
assign output_48 = input_15;
assign output_49 = input_15;
assign output_50 = input_15;
assign output_51 = input_15;
assign output_52 = input_15;
assign output_53 = input_15;
assign output_54 = input_15;
assign output_55 = input_15;
assign output_56 = input_15;
assign output_57 = input_15;
assign output_58 = input_15;
assign output_59 = input_15;
assign output_60 = input_15;
assign output_61 = input_15;
assign output_62 = input_15;
assign output_63 = input_15;
assign output_64 = input_15;
assign output_65 = input_15;
assign output_66 = input_15;
assign output_67 = input_15;
assign output_68 = input_15;
assign output_69 = input_15;
assign output_70 = input_15;
assign output_71 = input_15;
assign output_72 = input_15;
assign output_73 = input_15;
assign output_74 = input_15;
assign output_75 = input_15;
assign output_76 = input_15;
assign output_77 = input_15;
assign output_78 = input_15;
assign output_79 = input_15;
assign output_80 = input_15;
assign output_81 = input_15;
assign output_82 = input_15;
assign output_83 = input_15;
assign output_84 = input_15;
assign output_85 = input_15;
assign output_86 = input_15;
assign output_87 = input_15;
assign output_88 = input_15;
assign output_89 = input_15;
assign output_90 = input_15;
assign output_91 = input_15;
assign output_92 = input_15;
assign output_93 = input_15;
assign output_94 = input_15;
assign output_95 = input_15;
assign output_0 = input_16;
assign output_1 = input_16;
assign output_2 = input_16;
assign output_3 = input_16;
assign output_4 = input_16;
assign output_5 = input_16;
assign output_6 = input_16;
assign output_7 = input_16;
assign output_8 = input_16;
assign output_9 = input_16;
assign output_10 = input_16;
assign output_11 = input_16;
assign output_12 = input_16;
assign output_13 = input_16;
assign output_14 = input_16;
assign output_15 = input_16;
assign output_16 = input_16;
assign output_17 = input_16;
assign output_18 = input_16;
assign output_19 = input_16;
assign output_20 = input_16;
assign output_21 = input_16;
assign output_22 = input_16;
assign output_23 = input_16;
assign output_24 = input_16;
assign output_25 = input_16;
assign output_26 = input_16;
assign output_27 = input_16;
assign output_28 = input_16;
assign output_29 = input_16;
assign output_30 = input_16;
assign output_31 = input_16;
assign output_32 = input_16;
assign output_33 = input_16;
assign output_34 = input_16;
assign output_35 = input_16;
assign output_36 = input_16;
assign output_37 = input_16;
assign output_38 = input_16;
assign output_39 = input_16;
assign output_40 = input_16;
assign output_41 = input_16;
assign output_42 = input_16;
assign output_43 = input_16;
assign output_44 = input_16;
assign output_45 = input_16;
assign output_46 = input_16;
assign output_47 = input_16;
assign output_48 = input_16;
assign output_49 = input_16;
assign output_50 = input_16;
assign output_51 = input_16;
assign output_52 = input_16;
assign output_53 = input_16;
assign output_54 = input_16;
assign output_55 = input_16;
assign output_56 = input_16;
assign output_57 = input_16;
assign output_58 = input_16;
assign output_59 = input_16;
assign output_60 = input_16;
assign output_61 = input_16;
assign output_62 = input_16;
assign output_63 = input_16;
assign output_64 = input_16;
assign output_65 = input_16;
assign output_66 = input_16;
assign output_67 = input_16;
assign output_68 = input_16;
assign output_69 = input_16;
assign output_70 = input_16;
assign output_71 = input_16;
assign output_72 = input_16;
assign output_73 = input_16;
assign output_74 = input_16;
assign output_75 = input_16;
assign output_76 = input_16;
assign output_77 = input_16;
assign output_78 = input_16;
assign output_79 = input_16;
assign output_80 = input_16;
assign output_81 = input_16;
assign output_82 = input_16;
assign output_83 = input_16;
assign output_84 = input_16;
assign output_85 = input_16;
assign output_86 = input_16;
assign output_87 = input_16;
assign output_88 = input_16;
assign output_89 = input_16;
assign output_90 = input_16;
assign output_91 = input_16;
assign output_92 = input_16;
assign output_93 = input_16;
assign output_94 = input_16;
assign output_95 = input_16;
assign output_0 = input_17;
assign output_1 = input_17;
assign output_2 = input_17;
assign output_3 = input_17;
assign output_4 = input_17;
assign output_5 = input_17;
assign output_6 = input_17;
assign output_7 = input_17;
assign output_8 = input_17;
assign output_9 = input_17;
assign output_10 = input_17;
assign output_11 = input_17;
assign output_12 = input_17;
assign output_13 = input_17;
assign output_14 = input_17;
assign output_15 = input_17;
assign output_16 = input_17;
assign output_17 = input_17;
assign output_18 = input_17;
assign output_19 = input_17;
assign output_20 = input_17;
assign output_21 = input_17;
assign output_22 = input_17;
assign output_23 = input_17;
assign output_24 = input_17;
assign output_25 = input_17;
assign output_26 = input_17;
assign output_27 = input_17;
assign output_28 = input_17;
assign output_29 = input_17;
assign output_30 = input_17;
assign output_31 = input_17;
assign output_32 = input_17;
assign output_33 = input_17;
assign output_34 = input_17;
assign output_35 = input_17;
assign output_36 = input_17;
assign output_37 = input_17;
assign output_38 = input_17;
assign output_39 = input_17;
assign output_40 = input_17;
assign output_41 = input_17;
assign output_42 = input_17;
assign output_43 = input_17;
assign output_44 = input_17;
assign output_45 = input_17;
assign output_46 = input_17;
assign output_47 = input_17;
assign output_48 = input_17;
assign output_49 = input_17;
assign output_50 = input_17;
assign output_51 = input_17;
assign output_52 = input_17;
assign output_53 = input_17;
assign output_54 = input_17;
assign output_55 = input_17;
assign output_56 = input_17;
assign output_57 = input_17;
assign output_58 = input_17;
assign output_59 = input_17;
assign output_60 = input_17;
assign output_61 = input_17;
assign output_62 = input_17;
assign output_63 = input_17;
assign output_64 = input_17;
assign output_65 = input_17;
assign output_66 = input_17;
assign output_67 = input_17;
assign output_68 = input_17;
assign output_69 = input_17;
assign output_70 = input_17;
assign output_71 = input_17;
assign output_72 = input_17;
assign output_73 = input_17;
assign output_74 = input_17;
assign output_75 = input_17;
assign output_76 = input_17;
assign output_77 = input_17;
assign output_78 = input_17;
assign output_79 = input_17;
assign output_80 = input_17;
assign output_81 = input_17;
assign output_82 = input_17;
assign output_83 = input_17;
assign output_84 = input_17;
assign output_85 = input_17;
assign output_86 = input_17;
assign output_87 = input_17;
assign output_88 = input_17;
assign output_89 = input_17;
assign output_90 = input_17;
assign output_91 = input_17;
assign output_92 = input_17;
assign output_93 = input_17;
assign output_94 = input_17;
assign output_95 = input_17;
assign output_0 = input_18;
assign output_1 = input_18;
assign output_2 = input_18;
assign output_3 = input_18;
assign output_4 = input_18;
assign output_5 = input_18;
assign output_6 = input_18;
assign output_7 = input_18;
assign output_8 = input_18;
assign output_9 = input_18;
assign output_10 = input_18;
assign output_11 = input_18;
assign output_12 = input_18;
assign output_13 = input_18;
assign output_14 = input_18;
assign output_15 = input_18;
assign output_16 = input_18;
assign output_17 = input_18;
assign output_18 = input_18;
assign output_19 = input_18;
assign output_20 = input_18;
assign output_21 = input_18;
assign output_22 = input_18;
assign output_23 = input_18;
assign output_24 = input_18;
assign output_25 = input_18;
assign output_26 = input_18;
assign output_27 = input_18;
assign output_28 = input_18;
assign output_29 = input_18;
assign output_30 = input_18;
assign output_31 = input_18;
assign output_32 = input_18;
assign output_33 = input_18;
assign output_34 = input_18;
assign output_35 = input_18;
assign output_36 = input_18;
assign output_37 = input_18;
assign output_38 = input_18;
assign output_39 = input_18;
assign output_40 = input_18;
assign output_41 = input_18;
assign output_42 = input_18;
assign output_43 = input_18;
assign output_44 = input_18;
assign output_45 = input_18;
assign output_46 = input_18;
assign output_47 = input_18;
assign output_48 = input_18;
assign output_49 = input_18;
assign output_50 = input_18;
assign output_51 = input_18;
assign output_52 = input_18;
assign output_53 = input_18;
assign output_54 = input_18;
assign output_55 = input_18;
assign output_56 = input_18;
assign output_57 = input_18;
assign output_58 = input_18;
assign output_59 = input_18;
assign output_60 = input_18;
assign output_61 = input_18;
assign output_62 = input_18;
assign output_63 = input_18;
assign output_64 = input_18;
assign output_65 = input_18;
assign output_66 = input_18;
assign output_67 = input_18;
assign output_68 = input_18;
assign output_69 = input_18;
assign output_70 = input_18;
assign output_71 = input_18;
assign output_72 = input_18;
assign output_73 = input_18;
assign output_74 = input_18;
assign output_75 = input_18;
assign output_76 = input_18;
assign output_77 = input_18;
assign output_78 = input_18;
assign output_79 = input_18;
assign output_80 = input_18;
assign output_81 = input_18;
assign output_82 = input_18;
assign output_83 = input_18;
assign output_84 = input_18;
assign output_85 = input_18;
assign output_86 = input_18;
assign output_87 = input_18;
assign output_88 = input_18;
assign output_89 = input_18;
assign output_90 = input_18;
assign output_91 = input_18;
assign output_92 = input_18;
assign output_93 = input_18;
assign output_94 = input_18;
assign output_95 = input_18;
assign output_0 = input_19;
assign output_1 = input_19;
assign output_2 = input_19;
assign output_3 = input_19;
assign output_4 = input_19;
assign output_5 = input_19;
assign output_6 = input_19;
assign output_7 = input_19;
assign output_8 = input_19;
assign output_9 = input_19;
assign output_10 = input_19;
assign output_11 = input_19;
assign output_12 = input_19;
assign output_13 = input_19;
assign output_14 = input_19;
assign output_15 = input_19;
assign output_16 = input_19;
assign output_17 = input_19;
assign output_18 = input_19;
assign output_19 = input_19;
assign output_20 = input_19;
assign output_21 = input_19;
assign output_22 = input_19;
assign output_23 = input_19;
assign output_24 = input_19;
assign output_25 = input_19;
assign output_26 = input_19;
assign output_27 = input_19;
assign output_28 = input_19;
assign output_29 = input_19;
assign output_30 = input_19;
assign output_31 = input_19;
assign output_32 = input_19;
assign output_33 = input_19;
assign output_34 = input_19;
assign output_35 = input_19;
assign output_36 = input_19;
assign output_37 = input_19;
assign output_38 = input_19;
assign output_39 = input_19;
assign output_40 = input_19;
assign output_41 = input_19;
assign output_42 = input_19;
assign output_43 = input_19;
assign output_44 = input_19;
assign output_45 = input_19;
assign output_46 = input_19;
assign output_47 = input_19;
assign output_48 = input_19;
assign output_49 = input_19;
assign output_50 = input_19;
assign output_51 = input_19;
assign output_52 = input_19;
assign output_53 = input_19;
assign output_54 = input_19;
assign output_55 = input_19;
assign output_56 = input_19;
assign output_57 = input_19;
assign output_58 = input_19;
assign output_59 = input_19;
assign output_60 = input_19;
assign output_61 = input_19;
assign output_62 = input_19;
assign output_63 = input_19;
assign output_64 = input_19;
assign output_65 = input_19;
assign output_66 = input_19;
assign output_67 = input_19;
assign output_68 = input_19;
assign output_69 = input_19;
assign output_70 = input_19;
assign output_71 = input_19;
assign output_72 = input_19;
assign output_73 = input_19;
assign output_74 = input_19;
assign output_75 = input_19;
assign output_76 = input_19;
assign output_77 = input_19;
assign output_78 = input_19;
assign output_79 = input_19;
assign output_80 = input_19;
assign output_81 = input_19;
assign output_82 = input_19;
assign output_83 = input_19;
assign output_84 = input_19;
assign output_85 = input_19;
assign output_86 = input_19;
assign output_87 = input_19;
assign output_88 = input_19;
assign output_89 = input_19;
assign output_90 = input_19;
assign output_91 = input_19;
assign output_92 = input_19;
assign output_93 = input_19;
assign output_94 = input_19;
assign output_95 = input_19;
assign output_0 = input_20;
assign output_1 = input_20;
assign output_2 = input_20;
assign output_3 = input_20;
assign output_4 = input_20;
assign output_5 = input_20;
assign output_6 = input_20;
assign output_7 = input_20;
assign output_8 = input_20;
assign output_9 = input_20;
assign output_10 = input_20;
assign output_11 = input_20;
assign output_12 = input_20;
assign output_13 = input_20;
assign output_14 = input_20;
assign output_15 = input_20;
assign output_16 = input_20;
assign output_17 = input_20;
assign output_18 = input_20;
assign output_19 = input_20;
assign output_20 = input_20;
assign output_21 = input_20;
assign output_22 = input_20;
assign output_23 = input_20;
assign output_24 = input_20;
assign output_25 = input_20;
assign output_26 = input_20;
assign output_27 = input_20;
assign output_28 = input_20;
assign output_29 = input_20;
assign output_30 = input_20;
assign output_31 = input_20;
assign output_32 = input_20;
assign output_33 = input_20;
assign output_34 = input_20;
assign output_35 = input_20;
assign output_36 = input_20;
assign output_37 = input_20;
assign output_38 = input_20;
assign output_39 = input_20;
assign output_40 = input_20;
assign output_41 = input_20;
assign output_42 = input_20;
assign output_43 = input_20;
assign output_44 = input_20;
assign output_45 = input_20;
assign output_46 = input_20;
assign output_47 = input_20;
assign output_48 = input_20;
assign output_49 = input_20;
assign output_50 = input_20;
assign output_51 = input_20;
assign output_52 = input_20;
assign output_53 = input_20;
assign output_54 = input_20;
assign output_55 = input_20;
assign output_56 = input_20;
assign output_57 = input_20;
assign output_58 = input_20;
assign output_59 = input_20;
assign output_60 = input_20;
assign output_61 = input_20;
assign output_62 = input_20;
assign output_63 = input_20;
assign output_64 = input_20;
assign output_65 = input_20;
assign output_66 = input_20;
assign output_67 = input_20;
assign output_68 = input_20;
assign output_69 = input_20;
assign output_70 = input_20;
assign output_71 = input_20;
assign output_72 = input_20;
assign output_73 = input_20;
assign output_74 = input_20;
assign output_75 = input_20;
assign output_76 = input_20;
assign output_77 = input_20;
assign output_78 = input_20;
assign output_79 = input_20;
assign output_80 = input_20;
assign output_81 = input_20;
assign output_82 = input_20;
assign output_83 = input_20;
assign output_84 = input_20;
assign output_85 = input_20;
assign output_86 = input_20;
assign output_87 = input_20;
assign output_88 = input_20;
assign output_89 = input_20;
assign output_90 = input_20;
assign output_91 = input_20;
assign output_92 = input_20;
assign output_93 = input_20;
assign output_94 = input_20;
assign output_95 = input_20;
assign output_0 = input_21;
assign output_1 = input_21;
assign output_2 = input_21;
assign output_3 = input_21;
assign output_4 = input_21;
assign output_5 = input_21;
assign output_6 = input_21;
assign output_7 = input_21;
assign output_8 = input_21;
assign output_9 = input_21;
assign output_10 = input_21;
assign output_11 = input_21;
assign output_12 = input_21;
assign output_13 = input_21;
assign output_14 = input_21;
assign output_15 = input_21;
assign output_16 = input_21;
assign output_17 = input_21;
assign output_18 = input_21;
assign output_19 = input_21;
assign output_20 = input_21;
assign output_21 = input_21;
assign output_22 = input_21;
assign output_23 = input_21;
assign output_24 = input_21;
assign output_25 = input_21;
assign output_26 = input_21;
assign output_27 = input_21;
assign output_28 = input_21;
assign output_29 = input_21;
assign output_30 = input_21;
assign output_31 = input_21;
assign output_32 = input_21;
assign output_33 = input_21;
assign output_34 = input_21;
assign output_35 = input_21;
assign output_36 = input_21;
assign output_37 = input_21;
assign output_38 = input_21;
assign output_39 = input_21;
assign output_40 = input_21;
assign output_41 = input_21;
assign output_42 = input_21;
assign output_43 = input_21;
assign output_44 = input_21;
assign output_45 = input_21;
assign output_46 = input_21;
assign output_47 = input_21;
assign output_48 = input_21;
assign output_49 = input_21;
assign output_50 = input_21;
assign output_51 = input_21;
assign output_52 = input_21;
assign output_53 = input_21;
assign output_54 = input_21;
assign output_55 = input_21;
assign output_56 = input_21;
assign output_57 = input_21;
assign output_58 = input_21;
assign output_59 = input_21;
assign output_60 = input_21;
assign output_61 = input_21;
assign output_62 = input_21;
assign output_63 = input_21;
assign output_64 = input_21;
assign output_65 = input_21;
assign output_66 = input_21;
assign output_67 = input_21;
assign output_68 = input_21;
assign output_69 = input_21;
assign output_70 = input_21;
assign output_71 = input_21;
assign output_72 = input_21;
assign output_73 = input_21;
assign output_74 = input_21;
assign output_75 = input_21;
assign output_76 = input_21;
assign output_77 = input_21;
assign output_78 = input_21;
assign output_79 = input_21;
assign output_80 = input_21;
assign output_81 = input_21;
assign output_82 = input_21;
assign output_83 = input_21;
assign output_84 = input_21;
assign output_85 = input_21;
assign output_86 = input_21;
assign output_87 = input_21;
assign output_88 = input_21;
assign output_89 = input_21;
assign output_90 = input_21;
assign output_91 = input_21;
assign output_92 = input_21;
assign output_93 = input_21;
assign output_94 = input_21;
assign output_95 = input_21;
assign output_0 = input_22;
assign output_1 = input_22;
assign output_2 = input_22;
assign output_3 = input_22;
assign output_4 = input_22;
assign output_5 = input_22;
assign output_6 = input_22;
assign output_7 = input_22;
assign output_8 = input_22;
assign output_9 = input_22;
assign output_10 = input_22;
assign output_11 = input_22;
assign output_12 = input_22;
assign output_13 = input_22;
assign output_14 = input_22;
assign output_15 = input_22;
assign output_16 = input_22;
assign output_17 = input_22;
assign output_18 = input_22;
assign output_19 = input_22;
assign output_20 = input_22;
assign output_21 = input_22;
assign output_22 = input_22;
assign output_23 = input_22;
assign output_24 = input_22;
assign output_25 = input_22;
assign output_26 = input_22;
assign output_27 = input_22;
assign output_28 = input_22;
assign output_29 = input_22;
assign output_30 = input_22;
assign output_31 = input_22;
assign output_32 = input_22;
assign output_33 = input_22;
assign output_34 = input_22;
assign output_35 = input_22;
assign output_36 = input_22;
assign output_37 = input_22;
assign output_38 = input_22;
assign output_39 = input_22;
assign output_40 = input_22;
assign output_41 = input_22;
assign output_42 = input_22;
assign output_43 = input_22;
assign output_44 = input_22;
assign output_45 = input_22;
assign output_46 = input_22;
assign output_47 = input_22;
assign output_48 = input_22;
assign output_49 = input_22;
assign output_50 = input_22;
assign output_51 = input_22;
assign output_52 = input_22;
assign output_53 = input_22;
assign output_54 = input_22;
assign output_55 = input_22;
assign output_56 = input_22;
assign output_57 = input_22;
assign output_58 = input_22;
assign output_59 = input_22;
assign output_60 = input_22;
assign output_61 = input_22;
assign output_62 = input_22;
assign output_63 = input_22;
assign output_64 = input_22;
assign output_65 = input_22;
assign output_66 = input_22;
assign output_67 = input_22;
assign output_68 = input_22;
assign output_69 = input_22;
assign output_70 = input_22;
assign output_71 = input_22;
assign output_72 = input_22;
assign output_73 = input_22;
assign output_74 = input_22;
assign output_75 = input_22;
assign output_76 = input_22;
assign output_77 = input_22;
assign output_78 = input_22;
assign output_79 = input_22;
assign output_80 = input_22;
assign output_81 = input_22;
assign output_82 = input_22;
assign output_83 = input_22;
assign output_84 = input_22;
assign output_85 = input_22;
assign output_86 = input_22;
assign output_87 = input_22;
assign output_88 = input_22;
assign output_89 = input_22;
assign output_90 = input_22;
assign output_91 = input_22;
assign output_92 = input_22;
assign output_93 = input_22;
assign output_94 = input_22;
assign output_95 = input_22;
assign output_0 = input_23;
assign output_1 = input_23;
assign output_2 = input_23;
assign output_3 = input_23;
assign output_4 = input_23;
assign output_5 = input_23;
assign output_6 = input_23;
assign output_7 = input_23;
assign output_8 = input_23;
assign output_9 = input_23;
assign output_10 = input_23;
assign output_11 = input_23;
assign output_12 = input_23;
assign output_13 = input_23;
assign output_14 = input_23;
assign output_15 = input_23;
assign output_16 = input_23;
assign output_17 = input_23;
assign output_18 = input_23;
assign output_19 = input_23;
assign output_20 = input_23;
assign output_21 = input_23;
assign output_22 = input_23;
assign output_23 = input_23;
assign output_24 = input_23;
assign output_25 = input_23;
assign output_26 = input_23;
assign output_27 = input_23;
assign output_28 = input_23;
assign output_29 = input_23;
assign output_30 = input_23;
assign output_31 = input_23;
assign output_32 = input_23;
assign output_33 = input_23;
assign output_34 = input_23;
assign output_35 = input_23;
assign output_36 = input_23;
assign output_37 = input_23;
assign output_38 = input_23;
assign output_39 = input_23;
assign output_40 = input_23;
assign output_41 = input_23;
assign output_42 = input_23;
assign output_43 = input_23;
assign output_44 = input_23;
assign output_45 = input_23;
assign output_46 = input_23;
assign output_47 = input_23;
assign output_48 = input_23;
assign output_49 = input_23;
assign output_50 = input_23;
assign output_51 = input_23;
assign output_52 = input_23;
assign output_53 = input_23;
assign output_54 = input_23;
assign output_55 = input_23;
assign output_56 = input_23;
assign output_57 = input_23;
assign output_58 = input_23;
assign output_59 = input_23;
assign output_60 = input_23;
assign output_61 = input_23;
assign output_62 = input_23;
assign output_63 = input_23;
assign output_64 = input_23;
assign output_65 = input_23;
assign output_66 = input_23;
assign output_67 = input_23;
assign output_68 = input_23;
assign output_69 = input_23;
assign output_70 = input_23;
assign output_71 = input_23;
assign output_72 = input_23;
assign output_73 = input_23;
assign output_74 = input_23;
assign output_75 = input_23;
assign output_76 = input_23;
assign output_77 = input_23;
assign output_78 = input_23;
assign output_79 = input_23;
assign output_80 = input_23;
assign output_81 = input_23;
assign output_82 = input_23;
assign output_83 = input_23;
assign output_84 = input_23;
assign output_85 = input_23;
assign output_86 = input_23;
assign output_87 = input_23;
assign output_88 = input_23;
assign output_89 = input_23;
assign output_90 = input_23;
assign output_91 = input_23;
assign output_92 = input_23;
assign output_93 = input_23;
assign output_94 = input_23;
assign output_95 = input_23;
assign output_0 = input_24;
assign output_1 = input_24;
assign output_2 = input_24;
assign output_3 = input_24;
assign output_4 = input_24;
assign output_5 = input_24;
assign output_6 = input_24;
assign output_7 = input_24;
assign output_8 = input_24;
assign output_9 = input_24;
assign output_10 = input_24;
assign output_11 = input_24;
assign output_12 = input_24;
assign output_13 = input_24;
assign output_14 = input_24;
assign output_15 = input_24;
assign output_16 = input_24;
assign output_17 = input_24;
assign output_18 = input_24;
assign output_19 = input_24;
assign output_20 = input_24;
assign output_21 = input_24;
assign output_22 = input_24;
assign output_23 = input_24;
assign output_24 = input_24;
assign output_25 = input_24;
assign output_26 = input_24;
assign output_27 = input_24;
assign output_28 = input_24;
assign output_29 = input_24;
assign output_30 = input_24;
assign output_31 = input_24;
assign output_32 = input_24;
assign output_33 = input_24;
assign output_34 = input_24;
assign output_35 = input_24;
assign output_36 = input_24;
assign output_37 = input_24;
assign output_38 = input_24;
assign output_39 = input_24;
assign output_40 = input_24;
assign output_41 = input_24;
assign output_42 = input_24;
assign output_43 = input_24;
assign output_44 = input_24;
assign output_45 = input_24;
assign output_46 = input_24;
assign output_47 = input_24;
assign output_48 = input_24;
assign output_49 = input_24;
assign output_50 = input_24;
assign output_51 = input_24;
assign output_52 = input_24;
assign output_53 = input_24;
assign output_54 = input_24;
assign output_55 = input_24;
assign output_56 = input_24;
assign output_57 = input_24;
assign output_58 = input_24;
assign output_59 = input_24;
assign output_60 = input_24;
assign output_61 = input_24;
assign output_62 = input_24;
assign output_63 = input_24;
assign output_64 = input_24;
assign output_65 = input_24;
assign output_66 = input_24;
assign output_67 = input_24;
assign output_68 = input_24;
assign output_69 = input_24;
assign output_70 = input_24;
assign output_71 = input_24;
assign output_72 = input_24;
assign output_73 = input_24;
assign output_74 = input_24;
assign output_75 = input_24;
assign output_76 = input_24;
assign output_77 = input_24;
assign output_78 = input_24;
assign output_79 = input_24;
assign output_80 = input_24;
assign output_81 = input_24;
assign output_82 = input_24;
assign output_83 = input_24;
assign output_84 = input_24;
assign output_85 = input_24;
assign output_86 = input_24;
assign output_87 = input_24;
assign output_88 = input_24;
assign output_89 = input_24;
assign output_90 = input_24;
assign output_91 = input_24;
assign output_92 = input_24;
assign output_93 = input_24;
assign output_94 = input_24;
assign output_95 = input_24;
assign output_0 = input_25;
assign output_1 = input_25;
assign output_2 = input_25;
assign output_3 = input_25;
assign output_4 = input_25;
assign output_5 = input_25;
assign output_6 = input_25;
assign output_7 = input_25;
assign output_8 = input_25;
assign output_9 = input_25;
assign output_10 = input_25;
assign output_11 = input_25;
assign output_12 = input_25;
assign output_13 = input_25;
assign output_14 = input_25;
assign output_15 = input_25;
assign output_16 = input_25;
assign output_17 = input_25;
assign output_18 = input_25;
assign output_19 = input_25;
assign output_20 = input_25;
assign output_21 = input_25;
assign output_22 = input_25;
assign output_23 = input_25;
assign output_24 = input_25;
assign output_25 = input_25;
assign output_26 = input_25;
assign output_27 = input_25;
assign output_28 = input_25;
assign output_29 = input_25;
assign output_30 = input_25;
assign output_31 = input_25;
assign output_32 = input_25;
assign output_33 = input_25;
assign output_34 = input_25;
assign output_35 = input_25;
assign output_36 = input_25;
assign output_37 = input_25;
assign output_38 = input_25;
assign output_39 = input_25;
assign output_40 = input_25;
assign output_41 = input_25;
assign output_42 = input_25;
assign output_43 = input_25;
assign output_44 = input_25;
assign output_45 = input_25;
assign output_46 = input_25;
assign output_47 = input_25;
assign output_48 = input_25;
assign output_49 = input_25;
assign output_50 = input_25;
assign output_51 = input_25;
assign output_52 = input_25;
assign output_53 = input_25;
assign output_54 = input_25;
assign output_55 = input_25;
assign output_56 = input_25;
assign output_57 = input_25;
assign output_58 = input_25;
assign output_59 = input_25;
assign output_60 = input_25;
assign output_61 = input_25;
assign output_62 = input_25;
assign output_63 = input_25;
assign output_64 = input_25;
assign output_65 = input_25;
assign output_66 = input_25;
assign output_67 = input_25;
assign output_68 = input_25;
assign output_69 = input_25;
assign output_70 = input_25;
assign output_71 = input_25;
assign output_72 = input_25;
assign output_73 = input_25;
assign output_74 = input_25;
assign output_75 = input_25;
assign output_76 = input_25;
assign output_77 = input_25;
assign output_78 = input_25;
assign output_79 = input_25;
assign output_80 = input_25;
assign output_81 = input_25;
assign output_82 = input_25;
assign output_83 = input_25;
assign output_84 = input_25;
assign output_85 = input_25;
assign output_86 = input_25;
assign output_87 = input_25;
assign output_88 = input_25;
assign output_89 = input_25;
assign output_90 = input_25;
assign output_91 = input_25;
assign output_92 = input_25;
assign output_93 = input_25;
assign output_94 = input_25;
assign output_95 = input_25;
assign output_0 = input_26;
assign output_1 = input_26;
assign output_2 = input_26;
assign output_3 = input_26;
assign output_4 = input_26;
assign output_5 = input_26;
assign output_6 = input_26;
assign output_7 = input_26;
assign output_8 = input_26;
assign output_9 = input_26;
assign output_10 = input_26;
assign output_11 = input_26;
assign output_12 = input_26;
assign output_13 = input_26;
assign output_14 = input_26;
assign output_15 = input_26;
assign output_16 = input_26;
assign output_17 = input_26;
assign output_18 = input_26;
assign output_19 = input_26;
assign output_20 = input_26;
assign output_21 = input_26;
assign output_22 = input_26;
assign output_23 = input_26;
assign output_24 = input_26;
assign output_25 = input_26;
assign output_26 = input_26;
assign output_27 = input_26;
assign output_28 = input_26;
assign output_29 = input_26;
assign output_30 = input_26;
assign output_31 = input_26;
assign output_32 = input_26;
assign output_33 = input_26;
assign output_34 = input_26;
assign output_35 = input_26;
assign output_36 = input_26;
assign output_37 = input_26;
assign output_38 = input_26;
assign output_39 = input_26;
assign output_40 = input_26;
assign output_41 = input_26;
assign output_42 = input_26;
assign output_43 = input_26;
assign output_44 = input_26;
assign output_45 = input_26;
assign output_46 = input_26;
assign output_47 = input_26;
assign output_48 = input_26;
assign output_49 = input_26;
assign output_50 = input_26;
assign output_51 = input_26;
assign output_52 = input_26;
assign output_53 = input_26;
assign output_54 = input_26;
assign output_55 = input_26;
assign output_56 = input_26;
assign output_57 = input_26;
assign output_58 = input_26;
assign output_59 = input_26;
assign output_60 = input_26;
assign output_61 = input_26;
assign output_62 = input_26;
assign output_63 = input_26;
assign output_64 = input_26;
assign output_65 = input_26;
assign output_66 = input_26;
assign output_67 = input_26;
assign output_68 = input_26;
assign output_69 = input_26;
assign output_70 = input_26;
assign output_71 = input_26;
assign output_72 = input_26;
assign output_73 = input_26;
assign output_74 = input_26;
assign output_75 = input_26;
assign output_76 = input_26;
assign output_77 = input_26;
assign output_78 = input_26;
assign output_79 = input_26;
assign output_80 = input_26;
assign output_81 = input_26;
assign output_82 = input_26;
assign output_83 = input_26;
assign output_84 = input_26;
assign output_85 = input_26;
assign output_86 = input_26;
assign output_87 = input_26;
assign output_88 = input_26;
assign output_89 = input_26;
assign output_90 = input_26;
assign output_91 = input_26;
assign output_92 = input_26;
assign output_93 = input_26;
assign output_94 = input_26;
assign output_95 = input_26;
assign output_0 = input_27;
assign output_1 = input_27;
assign output_2 = input_27;
assign output_3 = input_27;
assign output_4 = input_27;
assign output_5 = input_27;
assign output_6 = input_27;
assign output_7 = input_27;
assign output_8 = input_27;
assign output_9 = input_27;
assign output_10 = input_27;
assign output_11 = input_27;
assign output_12 = input_27;
assign output_13 = input_27;
assign output_14 = input_27;
assign output_15 = input_27;
assign output_16 = input_27;
assign output_17 = input_27;
assign output_18 = input_27;
assign output_19 = input_27;
assign output_20 = input_27;
assign output_21 = input_27;
assign output_22 = input_27;
assign output_23 = input_27;
assign output_24 = input_27;
assign output_25 = input_27;
assign output_26 = input_27;
assign output_27 = input_27;
assign output_28 = input_27;
assign output_29 = input_27;
assign output_30 = input_27;
assign output_31 = input_27;
assign output_32 = input_27;
assign output_33 = input_27;
assign output_34 = input_27;
assign output_35 = input_27;
assign output_36 = input_27;
assign output_37 = input_27;
assign output_38 = input_27;
assign output_39 = input_27;
assign output_40 = input_27;
assign output_41 = input_27;
assign output_42 = input_27;
assign output_43 = input_27;
assign output_44 = input_27;
assign output_45 = input_27;
assign output_46 = input_27;
assign output_47 = input_27;
assign output_48 = input_27;
assign output_49 = input_27;
assign output_50 = input_27;
assign output_51 = input_27;
assign output_52 = input_27;
assign output_53 = input_27;
assign output_54 = input_27;
assign output_55 = input_27;
assign output_56 = input_27;
assign output_57 = input_27;
assign output_58 = input_27;
assign output_59 = input_27;
assign output_60 = input_27;
assign output_61 = input_27;
assign output_62 = input_27;
assign output_63 = input_27;
assign output_64 = input_27;
assign output_65 = input_27;
assign output_66 = input_27;
assign output_67 = input_27;
assign output_68 = input_27;
assign output_69 = input_27;
assign output_70 = input_27;
assign output_71 = input_27;
assign output_72 = input_27;
assign output_73 = input_27;
assign output_74 = input_27;
assign output_75 = input_27;
assign output_76 = input_27;
assign output_77 = input_27;
assign output_78 = input_27;
assign output_79 = input_27;
assign output_80 = input_27;
assign output_81 = input_27;
assign output_82 = input_27;
assign output_83 = input_27;
assign output_84 = input_27;
assign output_85 = input_27;
assign output_86 = input_27;
assign output_87 = input_27;
assign output_88 = input_27;
assign output_89 = input_27;
assign output_90 = input_27;
assign output_91 = input_27;
assign output_92 = input_27;
assign output_93 = input_27;
assign output_94 = input_27;
assign output_95 = input_27;
assign output_0 = input_28;
assign output_1 = input_28;
assign output_2 = input_28;
assign output_3 = input_28;
assign output_4 = input_28;
assign output_5 = input_28;
assign output_6 = input_28;
assign output_7 = input_28;
assign output_8 = input_28;
assign output_9 = input_28;
assign output_10 = input_28;
assign output_11 = input_28;
assign output_12 = input_28;
assign output_13 = input_28;
assign output_14 = input_28;
assign output_15 = input_28;
assign output_16 = input_28;
assign output_17 = input_28;
assign output_18 = input_28;
assign output_19 = input_28;
assign output_20 = input_28;
assign output_21 = input_28;
assign output_22 = input_28;
assign output_23 = input_28;
assign output_24 = input_28;
assign output_25 = input_28;
assign output_26 = input_28;
assign output_27 = input_28;
assign output_28 = input_28;
assign output_29 = input_28;
assign output_30 = input_28;
assign output_31 = input_28;
assign output_32 = input_28;
assign output_33 = input_28;
assign output_34 = input_28;
assign output_35 = input_28;
assign output_36 = input_28;
assign output_37 = input_28;
assign output_38 = input_28;
assign output_39 = input_28;
assign output_40 = input_28;
assign output_41 = input_28;
assign output_42 = input_28;
assign output_43 = input_28;
assign output_44 = input_28;
assign output_45 = input_28;
assign output_46 = input_28;
assign output_47 = input_28;
assign output_48 = input_28;
assign output_49 = input_28;
assign output_50 = input_28;
assign output_51 = input_28;
assign output_52 = input_28;
assign output_53 = input_28;
assign output_54 = input_28;
assign output_55 = input_28;
assign output_56 = input_28;
assign output_57 = input_28;
assign output_58 = input_28;
assign output_59 = input_28;
assign output_60 = input_28;
assign output_61 = input_28;
assign output_62 = input_28;
assign output_63 = input_28;
assign output_64 = input_28;
assign output_65 = input_28;
assign output_66 = input_28;
assign output_67 = input_28;
assign output_68 = input_28;
assign output_69 = input_28;
assign output_70 = input_28;
assign output_71 = input_28;
assign output_72 = input_28;
assign output_73 = input_28;
assign output_74 = input_28;
assign output_75 = input_28;
assign output_76 = input_28;
assign output_77 = input_28;
assign output_78 = input_28;
assign output_79 = input_28;
assign output_80 = input_28;
assign output_81 = input_28;
assign output_82 = input_28;
assign output_83 = input_28;
assign output_84 = input_28;
assign output_85 = input_28;
assign output_86 = input_28;
assign output_87 = input_28;
assign output_88 = input_28;
assign output_89 = input_28;
assign output_90 = input_28;
assign output_91 = input_28;
assign output_92 = input_28;
assign output_93 = input_28;
assign output_94 = input_28;
assign output_95 = input_28;
assign output_0 = input_29;
assign output_1 = input_29;
assign output_2 = input_29;
assign output_3 = input_29;
assign output_4 = input_29;
assign output_5 = input_29;
assign output_6 = input_29;
assign output_7 = input_29;
assign output_8 = input_29;
assign output_9 = input_29;
assign output_10 = input_29;
assign output_11 = input_29;
assign output_12 = input_29;
assign output_13 = input_29;
assign output_14 = input_29;
assign output_15 = input_29;
assign output_16 = input_29;
assign output_17 = input_29;
assign output_18 = input_29;
assign output_19 = input_29;
assign output_20 = input_29;
assign output_21 = input_29;
assign output_22 = input_29;
assign output_23 = input_29;
assign output_24 = input_29;
assign output_25 = input_29;
assign output_26 = input_29;
assign output_27 = input_29;
assign output_28 = input_29;
assign output_29 = input_29;
assign output_30 = input_29;
assign output_31 = input_29;
assign output_32 = input_29;
assign output_33 = input_29;
assign output_34 = input_29;
assign output_35 = input_29;
assign output_36 = input_29;
assign output_37 = input_29;
assign output_38 = input_29;
assign output_39 = input_29;
assign output_40 = input_29;
assign output_41 = input_29;
assign output_42 = input_29;
assign output_43 = input_29;
assign output_44 = input_29;
assign output_45 = input_29;
assign output_46 = input_29;
assign output_47 = input_29;
assign output_48 = input_29;
assign output_49 = input_29;
assign output_50 = input_29;
assign output_51 = input_29;
assign output_52 = input_29;
assign output_53 = input_29;
assign output_54 = input_29;
assign output_55 = input_29;
assign output_56 = input_29;
assign output_57 = input_29;
assign output_58 = input_29;
assign output_59 = input_29;
assign output_60 = input_29;
assign output_61 = input_29;
assign output_62 = input_29;
assign output_63 = input_29;
assign output_64 = input_29;
assign output_65 = input_29;
assign output_66 = input_29;
assign output_67 = input_29;
assign output_68 = input_29;
assign output_69 = input_29;
assign output_70 = input_29;
assign output_71 = input_29;
assign output_72 = input_29;
assign output_73 = input_29;
assign output_74 = input_29;
assign output_75 = input_29;
assign output_76 = input_29;
assign output_77 = input_29;
assign output_78 = input_29;
assign output_79 = input_29;
assign output_80 = input_29;
assign output_81 = input_29;
assign output_82 = input_29;
assign output_83 = input_29;
assign output_84 = input_29;
assign output_85 = input_29;
assign output_86 = input_29;
assign output_87 = input_29;
assign output_88 = input_29;
assign output_89 = input_29;
assign output_90 = input_29;
assign output_91 = input_29;
assign output_92 = input_29;
assign output_93 = input_29;
assign output_94 = input_29;
assign output_95 = input_29;
assign output_0 = input_30;
assign output_1 = input_30;
assign output_2 = input_30;
assign output_3 = input_30;
assign output_4 = input_30;
assign output_5 = input_30;
assign output_6 = input_30;
assign output_7 = input_30;
assign output_8 = input_30;
assign output_9 = input_30;
assign output_10 = input_30;
assign output_11 = input_30;
assign output_12 = input_30;
assign output_13 = input_30;
assign output_14 = input_30;
assign output_15 = input_30;
assign output_16 = input_30;
assign output_17 = input_30;
assign output_18 = input_30;
assign output_19 = input_30;
assign output_20 = input_30;
assign output_21 = input_30;
assign output_22 = input_30;
assign output_23 = input_30;
assign output_24 = input_30;
assign output_25 = input_30;
assign output_26 = input_30;
assign output_27 = input_30;
assign output_28 = input_30;
assign output_29 = input_30;
assign output_30 = input_30;
assign output_31 = input_30;
assign output_32 = input_30;
assign output_33 = input_30;
assign output_34 = input_30;
assign output_35 = input_30;
assign output_36 = input_30;
assign output_37 = input_30;
assign output_38 = input_30;
assign output_39 = input_30;
assign output_40 = input_30;
assign output_41 = input_30;
assign output_42 = input_30;
assign output_43 = input_30;
assign output_44 = input_30;
assign output_45 = input_30;
assign output_46 = input_30;
assign output_47 = input_30;
assign output_48 = input_30;
assign output_49 = input_30;
assign output_50 = input_30;
assign output_51 = input_30;
assign output_52 = input_30;
assign output_53 = input_30;
assign output_54 = input_30;
assign output_55 = input_30;
assign output_56 = input_30;
assign output_57 = input_30;
assign output_58 = input_30;
assign output_59 = input_30;
assign output_60 = input_30;
assign output_61 = input_30;
assign output_62 = input_30;
assign output_63 = input_30;
assign output_64 = input_30;
assign output_65 = input_30;
assign output_66 = input_30;
assign output_67 = input_30;
assign output_68 = input_30;
assign output_69 = input_30;
assign output_70 = input_30;
assign output_71 = input_30;
assign output_72 = input_30;
assign output_73 = input_30;
assign output_74 = input_30;
assign output_75 = input_30;
assign output_76 = input_30;
assign output_77 = input_30;
assign output_78 = input_30;
assign output_79 = input_30;
assign output_80 = input_30;
assign output_81 = input_30;
assign output_82 = input_30;
assign output_83 = input_30;
assign output_84 = input_30;
assign output_85 = input_30;
assign output_86 = input_30;
assign output_87 = input_30;
assign output_88 = input_30;
assign output_89 = input_30;
assign output_90 = input_30;
assign output_91 = input_30;
assign output_92 = input_30;
assign output_93 = input_30;
assign output_94 = input_30;
assign output_95 = input_30;
assign output_0 = input_31;
assign output_1 = input_31;
assign output_2 = input_31;
assign output_3 = input_31;
assign output_4 = input_31;
assign output_5 = input_31;
assign output_6 = input_31;
assign output_7 = input_31;
assign output_8 = input_31;
assign output_9 = input_31;
assign output_10 = input_31;
assign output_11 = input_31;
assign output_12 = input_31;
assign output_13 = input_31;
assign output_14 = input_31;
assign output_15 = input_31;
assign output_16 = input_31;
assign output_17 = input_31;
assign output_18 = input_31;
assign output_19 = input_31;
assign output_20 = input_31;
assign output_21 = input_31;
assign output_22 = input_31;
assign output_23 = input_31;
assign output_24 = input_31;
assign output_25 = input_31;
assign output_26 = input_31;
assign output_27 = input_31;
assign output_28 = input_31;
assign output_29 = input_31;
assign output_30 = input_31;
assign output_31 = input_31;
assign output_32 = input_31;
assign output_33 = input_31;
assign output_34 = input_31;
assign output_35 = input_31;
assign output_36 = input_31;
assign output_37 = input_31;
assign output_38 = input_31;
assign output_39 = input_31;
assign output_40 = input_31;
assign output_41 = input_31;
assign output_42 = input_31;
assign output_43 = input_31;
assign output_44 = input_31;
assign output_45 = input_31;
assign output_46 = input_31;
assign output_47 = input_31;
assign output_48 = input_31;
assign output_49 = input_31;
assign output_50 = input_31;
assign output_51 = input_31;
assign output_52 = input_31;
assign output_53 = input_31;
assign output_54 = input_31;
assign output_55 = input_31;
assign output_56 = input_31;
assign output_57 = input_31;
assign output_58 = input_31;
assign output_59 = input_31;
assign output_60 = input_31;
assign output_61 = input_31;
assign output_62 = input_31;
assign output_63 = input_31;
assign output_64 = input_31;
assign output_65 = input_31;
assign output_66 = input_31;
assign output_67 = input_31;
assign output_68 = input_31;
assign output_69 = input_31;
assign output_70 = input_31;
assign output_71 = input_31;
assign output_72 = input_31;
assign output_73 = input_31;
assign output_74 = input_31;
assign output_75 = input_31;
assign output_76 = input_31;
assign output_77 = input_31;
assign output_78 = input_31;
assign output_79 = input_31;
assign output_80 = input_31;
assign output_81 = input_31;
assign output_82 = input_31;
assign output_83 = input_31;
assign output_84 = input_31;
assign output_85 = input_31;
assign output_86 = input_31;
assign output_87 = input_31;
assign output_88 = input_31;
assign output_89 = input_31;
assign output_90 = input_31;
assign output_91 = input_31;
assign output_92 = input_31;
assign output_93 = input_31;
assign output_94 = input_31;
assign output_95 = input_31;
assign output_0 = input_32;
assign output_1 = input_32;
assign output_2 = input_32;
assign output_3 = input_32;
assign output_4 = input_32;
assign output_5 = input_32;
assign output_6 = input_32;
assign output_7 = input_32;
assign output_8 = input_32;
assign output_9 = input_32;
assign output_10 = input_32;
assign output_11 = input_32;
assign output_12 = input_32;
assign output_13 = input_32;
assign output_14 = input_32;
assign output_15 = input_32;
assign output_16 = input_32;
assign output_17 = input_32;
assign output_18 = input_32;
assign output_19 = input_32;
assign output_20 = input_32;
assign output_21 = input_32;
assign output_22 = input_32;
assign output_23 = input_32;
assign output_24 = input_32;
assign output_25 = input_32;
assign output_26 = input_32;
assign output_27 = input_32;
assign output_28 = input_32;
assign output_29 = input_32;
assign output_30 = input_32;
assign output_31 = input_32;
assign output_32 = input_32;
assign output_33 = input_32;
assign output_34 = input_32;
assign output_35 = input_32;
assign output_36 = input_32;
assign output_37 = input_32;
assign output_38 = input_32;
assign output_39 = input_32;
assign output_40 = input_32;
assign output_41 = input_32;
assign output_42 = input_32;
assign output_43 = input_32;
assign output_44 = input_32;
assign output_45 = input_32;
assign output_46 = input_32;
assign output_47 = input_32;
assign output_48 = input_32;
assign output_49 = input_32;
assign output_50 = input_32;
assign output_51 = input_32;
assign output_52 = input_32;
assign output_53 = input_32;
assign output_54 = input_32;
assign output_55 = input_32;
assign output_56 = input_32;
assign output_57 = input_32;
assign output_58 = input_32;
assign output_59 = input_32;
assign output_60 = input_32;
assign output_61 = input_32;
assign output_62 = input_32;
assign output_63 = input_32;
assign output_64 = input_32;
assign output_65 = input_32;
assign output_66 = input_32;
assign output_67 = input_32;
assign output_68 = input_32;
assign output_69 = input_32;
assign output_70 = input_32;
assign output_71 = input_32;
assign output_72 = input_32;
assign output_73 = input_32;
assign output_74 = input_32;
assign output_75 = input_32;
assign output_76 = input_32;
assign output_77 = input_32;
assign output_78 = input_32;
assign output_79 = input_32;
assign output_80 = input_32;
assign output_81 = input_32;
assign output_82 = input_32;
assign output_83 = input_32;
assign output_84 = input_32;
assign output_85 = input_32;
assign output_86 = input_32;
assign output_87 = input_32;
assign output_88 = input_32;
assign output_89 = input_32;
assign output_90 = input_32;
assign output_91 = input_32;
assign output_92 = input_32;
assign output_93 = input_32;
assign output_94 = input_32;
assign output_95 = input_32;
assign output_0 = input_33;
assign output_1 = input_33;
assign output_2 = input_33;
assign output_3 = input_33;
assign output_4 = input_33;
assign output_5 = input_33;
assign output_6 = input_33;
assign output_7 = input_33;
assign output_8 = input_33;
assign output_9 = input_33;
assign output_10 = input_33;
assign output_11 = input_33;
assign output_12 = input_33;
assign output_13 = input_33;
assign output_14 = input_33;
assign output_15 = input_33;
assign output_16 = input_33;
assign output_17 = input_33;
assign output_18 = input_33;
assign output_19 = input_33;
assign output_20 = input_33;
assign output_21 = input_33;
assign output_22 = input_33;
assign output_23 = input_33;
assign output_24 = input_33;
assign output_25 = input_33;
assign output_26 = input_33;
assign output_27 = input_33;
assign output_28 = input_33;
assign output_29 = input_33;
assign output_30 = input_33;
assign output_31 = input_33;
assign output_32 = input_33;
assign output_33 = input_33;
assign output_34 = input_33;
assign output_35 = input_33;
assign output_36 = input_33;
assign output_37 = input_33;
assign output_38 = input_33;
assign output_39 = input_33;
assign output_40 = input_33;
assign output_41 = input_33;
assign output_42 = input_33;
assign output_43 = input_33;
assign output_44 = input_33;
assign output_45 = input_33;
assign output_46 = input_33;
assign output_47 = input_33;
assign output_48 = input_33;
assign output_49 = input_33;
assign output_50 = input_33;
assign output_51 = input_33;
assign output_52 = input_33;
assign output_53 = input_33;
assign output_54 = input_33;
assign output_55 = input_33;
assign output_56 = input_33;
assign output_57 = input_33;
assign output_58 = input_33;
assign output_59 = input_33;
assign output_60 = input_33;
assign output_61 = input_33;
assign output_62 = input_33;
assign output_63 = input_33;
assign output_64 = input_33;
assign output_65 = input_33;
assign output_66 = input_33;
assign output_67 = input_33;
assign output_68 = input_33;
assign output_69 = input_33;
assign output_70 = input_33;
assign output_71 = input_33;
assign output_72 = input_33;
assign output_73 = input_33;
assign output_74 = input_33;
assign output_75 = input_33;
assign output_76 = input_33;
assign output_77 = input_33;
assign output_78 = input_33;
assign output_79 = input_33;
assign output_80 = input_33;
assign output_81 = input_33;
assign output_82 = input_33;
assign output_83 = input_33;
assign output_84 = input_33;
assign output_85 = input_33;
assign output_86 = input_33;
assign output_87 = input_33;
assign output_88 = input_33;
assign output_89 = input_33;
assign output_90 = input_33;
assign output_91 = input_33;
assign output_92 = input_33;
assign output_93 = input_33;
assign output_94 = input_33;
assign output_95 = input_33;
assign output_0 = input_34;
assign output_1 = input_34;
assign output_2 = input_34;
assign output_3 = input_34;
assign output_4 = input_34;
assign output_5 = input_34;
assign output_6 = input_34;
assign output_7 = input_34;
assign output_8 = input_34;
assign output_9 = input_34;
assign output_10 = input_34;
assign output_11 = input_34;
assign output_12 = input_34;
assign output_13 = input_34;
assign output_14 = input_34;
assign output_15 = input_34;
assign output_16 = input_34;
assign output_17 = input_34;
assign output_18 = input_34;
assign output_19 = input_34;
assign output_20 = input_34;
assign output_21 = input_34;
assign output_22 = input_34;
assign output_23 = input_34;
assign output_24 = input_34;
assign output_25 = input_34;
assign output_26 = input_34;
assign output_27 = input_34;
assign output_28 = input_34;
assign output_29 = input_34;
assign output_30 = input_34;
assign output_31 = input_34;
assign output_32 = input_34;
assign output_33 = input_34;
assign output_34 = input_34;
assign output_35 = input_34;
assign output_36 = input_34;
assign output_37 = input_34;
assign output_38 = input_34;
assign output_39 = input_34;
assign output_40 = input_34;
assign output_41 = input_34;
assign output_42 = input_34;
assign output_43 = input_34;
assign output_44 = input_34;
assign output_45 = input_34;
assign output_46 = input_34;
assign output_47 = input_34;
assign output_48 = input_34;
assign output_49 = input_34;
assign output_50 = input_34;
assign output_51 = input_34;
assign output_52 = input_34;
assign output_53 = input_34;
assign output_54 = input_34;
assign output_55 = input_34;
assign output_56 = input_34;
assign output_57 = input_34;
assign output_58 = input_34;
assign output_59 = input_34;
assign output_60 = input_34;
assign output_61 = input_34;
assign output_62 = input_34;
assign output_63 = input_34;
assign output_64 = input_34;
assign output_65 = input_34;
assign output_66 = input_34;
assign output_67 = input_34;
assign output_68 = input_34;
assign output_69 = input_34;
assign output_70 = input_34;
assign output_71 = input_34;
assign output_72 = input_34;
assign output_73 = input_34;
assign output_74 = input_34;
assign output_75 = input_34;
assign output_76 = input_34;
assign output_77 = input_34;
assign output_78 = input_34;
assign output_79 = input_34;
assign output_80 = input_34;
assign output_81 = input_34;
assign output_82 = input_34;
assign output_83 = input_34;
assign output_84 = input_34;
assign output_85 = input_34;
assign output_86 = input_34;
assign output_87 = input_34;
assign output_88 = input_34;
assign output_89 = input_34;
assign output_90 = input_34;
assign output_91 = input_34;
assign output_92 = input_34;
assign output_93 = input_34;
assign output_94 = input_34;
assign output_95 = input_34;
assign output_0 = input_35;
assign output_1 = input_35;
assign output_2 = input_35;
assign output_3 = input_35;
assign output_4 = input_35;
assign output_5 = input_35;
assign output_6 = input_35;
assign output_7 = input_35;
assign output_8 = input_35;
assign output_9 = input_35;
assign output_10 = input_35;
assign output_11 = input_35;
assign output_12 = input_35;
assign output_13 = input_35;
assign output_14 = input_35;
assign output_15 = input_35;
assign output_16 = input_35;
assign output_17 = input_35;
assign output_18 = input_35;
assign output_19 = input_35;
assign output_20 = input_35;
assign output_21 = input_35;
assign output_22 = input_35;
assign output_23 = input_35;
assign output_24 = input_35;
assign output_25 = input_35;
assign output_26 = input_35;
assign output_27 = input_35;
assign output_28 = input_35;
assign output_29 = input_35;
assign output_30 = input_35;
assign output_31 = input_35;
assign output_32 = input_35;
assign output_33 = input_35;
assign output_34 = input_35;
assign output_35 = input_35;
assign output_36 = input_35;
assign output_37 = input_35;
assign output_38 = input_35;
assign output_39 = input_35;
assign output_40 = input_35;
assign output_41 = input_35;
assign output_42 = input_35;
assign output_43 = input_35;
assign output_44 = input_35;
assign output_45 = input_35;
assign output_46 = input_35;
assign output_47 = input_35;
assign output_48 = input_35;
assign output_49 = input_35;
assign output_50 = input_35;
assign output_51 = input_35;
assign output_52 = input_35;
assign output_53 = input_35;
assign output_54 = input_35;
assign output_55 = input_35;
assign output_56 = input_35;
assign output_57 = input_35;
assign output_58 = input_35;
assign output_59 = input_35;
assign output_60 = input_35;
assign output_61 = input_35;
assign output_62 = input_35;
assign output_63 = input_35;
assign output_64 = input_35;
assign output_65 = input_35;
assign output_66 = input_35;
assign output_67 = input_35;
assign output_68 = input_35;
assign output_69 = input_35;
assign output_70 = input_35;
assign output_71 = input_35;
assign output_72 = input_35;
assign output_73 = input_35;
assign output_74 = input_35;
assign output_75 = input_35;
assign output_76 = input_35;
assign output_77 = input_35;
assign output_78 = input_35;
assign output_79 = input_35;
assign output_80 = input_35;
assign output_81 = input_35;
assign output_82 = input_35;
assign output_83 = input_35;
assign output_84 = input_35;
assign output_85 = input_35;
assign output_86 = input_35;
assign output_87 = input_35;
assign output_88 = input_35;
assign output_89 = input_35;
assign output_90 = input_35;
assign output_91 = input_35;
assign output_92 = input_35;
assign output_93 = input_35;
assign output_94 = input_35;
assign output_95 = input_35;
assign output_0 = input_36;
assign output_1 = input_36;
assign output_2 = input_36;
assign output_3 = input_36;
assign output_4 = input_36;
assign output_5 = input_36;
assign output_6 = input_36;
assign output_7 = input_36;
assign output_8 = input_36;
assign output_9 = input_36;
assign output_10 = input_36;
assign output_11 = input_36;
assign output_12 = input_36;
assign output_13 = input_36;
assign output_14 = input_36;
assign output_15 = input_36;
assign output_16 = input_36;
assign output_17 = input_36;
assign output_18 = input_36;
assign output_19 = input_36;
assign output_20 = input_36;
assign output_21 = input_36;
assign output_22 = input_36;
assign output_23 = input_36;
assign output_24 = input_36;
assign output_25 = input_36;
assign output_26 = input_36;
assign output_27 = input_36;
assign output_28 = input_36;
assign output_29 = input_36;
assign output_30 = input_36;
assign output_31 = input_36;
assign output_32 = input_36;
assign output_33 = input_36;
assign output_34 = input_36;
assign output_35 = input_36;
assign output_36 = input_36;
assign output_37 = input_36;
assign output_38 = input_36;
assign output_39 = input_36;
assign output_40 = input_36;
assign output_41 = input_36;
assign output_42 = input_36;
assign output_43 = input_36;
assign output_44 = input_36;
assign output_45 = input_36;
assign output_46 = input_36;
assign output_47 = input_36;
assign output_48 = input_36;
assign output_49 = input_36;
assign output_50 = input_36;
assign output_51 = input_36;
assign output_52 = input_36;
assign output_53 = input_36;
assign output_54 = input_36;
assign output_55 = input_36;
assign output_56 = input_36;
assign output_57 = input_36;
assign output_58 = input_36;
assign output_59 = input_36;
assign output_60 = input_36;
assign output_61 = input_36;
assign output_62 = input_36;
assign output_63 = input_36;
assign output_64 = input_36;
assign output_65 = input_36;
assign output_66 = input_36;
assign output_67 = input_36;
assign output_68 = input_36;
assign output_69 = input_36;
assign output_70 = input_36;
assign output_71 = input_36;
assign output_72 = input_36;
assign output_73 = input_36;
assign output_74 = input_36;
assign output_75 = input_36;
assign output_76 = input_36;
assign output_77 = input_36;
assign output_78 = input_36;
assign output_79 = input_36;
assign output_80 = input_36;
assign output_81 = input_36;
assign output_82 = input_36;
assign output_83 = input_36;
assign output_84 = input_36;
assign output_85 = input_36;
assign output_86 = input_36;
assign output_87 = input_36;
assign output_88 = input_36;
assign output_89 = input_36;
assign output_90 = input_36;
assign output_91 = input_36;
assign output_92 = input_36;
assign output_93 = input_36;
assign output_94 = input_36;
assign output_95 = input_36;
assign output_0 = input_37;
assign output_1 = input_37;
assign output_2 = input_37;
assign output_3 = input_37;
assign output_4 = input_37;
assign output_5 = input_37;
assign output_6 = input_37;
assign output_7 = input_37;
assign output_8 = input_37;
assign output_9 = input_37;
assign output_10 = input_37;
assign output_11 = input_37;
assign output_12 = input_37;
assign output_13 = input_37;
assign output_14 = input_37;
assign output_15 = input_37;
assign output_16 = input_37;
assign output_17 = input_37;
assign output_18 = input_37;
assign output_19 = input_37;
assign output_20 = input_37;
assign output_21 = input_37;
assign output_22 = input_37;
assign output_23 = input_37;
assign output_24 = input_37;
assign output_25 = input_37;
assign output_26 = input_37;
assign output_27 = input_37;
assign output_28 = input_37;
assign output_29 = input_37;
assign output_30 = input_37;
assign output_31 = input_37;
assign output_32 = input_37;
assign output_33 = input_37;
assign output_34 = input_37;
assign output_35 = input_37;
assign output_36 = input_37;
assign output_37 = input_37;
assign output_38 = input_37;
assign output_39 = input_37;
assign output_40 = input_37;
assign output_41 = input_37;
assign output_42 = input_37;
assign output_43 = input_37;
assign output_44 = input_37;
assign output_45 = input_37;
assign output_46 = input_37;
assign output_47 = input_37;
assign output_48 = input_37;
assign output_49 = input_37;
assign output_50 = input_37;
assign output_51 = input_37;
assign output_52 = input_37;
assign output_53 = input_37;
assign output_54 = input_37;
assign output_55 = input_37;
assign output_56 = input_37;
assign output_57 = input_37;
assign output_58 = input_37;
assign output_59 = input_37;
assign output_60 = input_37;
assign output_61 = input_37;
assign output_62 = input_37;
assign output_63 = input_37;
assign output_64 = input_37;
assign output_65 = input_37;
assign output_66 = input_37;
assign output_67 = input_37;
assign output_68 = input_37;
assign output_69 = input_37;
assign output_70 = input_37;
assign output_71 = input_37;
assign output_72 = input_37;
assign output_73 = input_37;
assign output_74 = input_37;
assign output_75 = input_37;
assign output_76 = input_37;
assign output_77 = input_37;
assign output_78 = input_37;
assign output_79 = input_37;
assign output_80 = input_37;
assign output_81 = input_37;
assign output_82 = input_37;
assign output_83 = input_37;
assign output_84 = input_37;
assign output_85 = input_37;
assign output_86 = input_37;
assign output_87 = input_37;
assign output_88 = input_37;
assign output_89 = input_37;
assign output_90 = input_37;
assign output_91 = input_37;
assign output_92 = input_37;
assign output_93 = input_37;
assign output_94 = input_37;
assign output_95 = input_37;
assign output_0 = input_38;
assign output_1 = input_38;
assign output_2 = input_38;
assign output_3 = input_38;
assign output_4 = input_38;
assign output_5 = input_38;
assign output_6 = input_38;
assign output_7 = input_38;
assign output_8 = input_38;
assign output_9 = input_38;
assign output_10 = input_38;
assign output_11 = input_38;
assign output_12 = input_38;
assign output_13 = input_38;
assign output_14 = input_38;
assign output_15 = input_38;
assign output_16 = input_38;
assign output_17 = input_38;
assign output_18 = input_38;
assign output_19 = input_38;
assign output_20 = input_38;
assign output_21 = input_38;
assign output_22 = input_38;
assign output_23 = input_38;
assign output_24 = input_38;
assign output_25 = input_38;
assign output_26 = input_38;
assign output_27 = input_38;
assign output_28 = input_38;
assign output_29 = input_38;
assign output_30 = input_38;
assign output_31 = input_38;
assign output_32 = input_38;
assign output_33 = input_38;
assign output_34 = input_38;
assign output_35 = input_38;
assign output_36 = input_38;
assign output_37 = input_38;
assign output_38 = input_38;
assign output_39 = input_38;
assign output_40 = input_38;
assign output_41 = input_38;
assign output_42 = input_38;
assign output_43 = input_38;
assign output_44 = input_38;
assign output_45 = input_38;
assign output_46 = input_38;
assign output_47 = input_38;
assign output_48 = input_38;
assign output_49 = input_38;
assign output_50 = input_38;
assign output_51 = input_38;
assign output_52 = input_38;
assign output_53 = input_38;
assign output_54 = input_38;
assign output_55 = input_38;
assign output_56 = input_38;
assign output_57 = input_38;
assign output_58 = input_38;
assign output_59 = input_38;
assign output_60 = input_38;
assign output_61 = input_38;
assign output_62 = input_38;
assign output_63 = input_38;
assign output_64 = input_38;
assign output_65 = input_38;
assign output_66 = input_38;
assign output_67 = input_38;
assign output_68 = input_38;
assign output_69 = input_38;
assign output_70 = input_38;
assign output_71 = input_38;
assign output_72 = input_38;
assign output_73 = input_38;
assign output_74 = input_38;
assign output_75 = input_38;
assign output_76 = input_38;
assign output_77 = input_38;
assign output_78 = input_38;
assign output_79 = input_38;
assign output_80 = input_38;
assign output_81 = input_38;
assign output_82 = input_38;
assign output_83 = input_38;
assign output_84 = input_38;
assign output_85 = input_38;
assign output_86 = input_38;
assign output_87 = input_38;
assign output_88 = input_38;
assign output_89 = input_38;
assign output_90 = input_38;
assign output_91 = input_38;
assign output_92 = input_38;
assign output_93 = input_38;
assign output_94 = input_38;
assign output_95 = input_38;
assign output_0 = input_39;
assign output_1 = input_39;
assign output_2 = input_39;
assign output_3 = input_39;
assign output_4 = input_39;
assign output_5 = input_39;
assign output_6 = input_39;
assign output_7 = input_39;
assign output_8 = input_39;
assign output_9 = input_39;
assign output_10 = input_39;
assign output_11 = input_39;
assign output_12 = input_39;
assign output_13 = input_39;
assign output_14 = input_39;
assign output_15 = input_39;
assign output_16 = input_39;
assign output_17 = input_39;
assign output_18 = input_39;
assign output_19 = input_39;
assign output_20 = input_39;
assign output_21 = input_39;
assign output_22 = input_39;
assign output_23 = input_39;
assign output_24 = input_39;
assign output_25 = input_39;
assign output_26 = input_39;
assign output_27 = input_39;
assign output_28 = input_39;
assign output_29 = input_39;
assign output_30 = input_39;
assign output_31 = input_39;
assign output_32 = input_39;
assign output_33 = input_39;
assign output_34 = input_39;
assign output_35 = input_39;
assign output_36 = input_39;
assign output_37 = input_39;
assign output_38 = input_39;
assign output_39 = input_39;
assign output_40 = input_39;
assign output_41 = input_39;
assign output_42 = input_39;
assign output_43 = input_39;
assign output_44 = input_39;
assign output_45 = input_39;
assign output_46 = input_39;
assign output_47 = input_39;
assign output_48 = input_39;
assign output_49 = input_39;
assign output_50 = input_39;
assign output_51 = input_39;
assign output_52 = input_39;
assign output_53 = input_39;
assign output_54 = input_39;
assign output_55 = input_39;
assign output_56 = input_39;
assign output_57 = input_39;
assign output_58 = input_39;
assign output_59 = input_39;
assign output_60 = input_39;
assign output_61 = input_39;
assign output_62 = input_39;
assign output_63 = input_39;
assign output_64 = input_39;
assign output_65 = input_39;
assign output_66 = input_39;
assign output_67 = input_39;
assign output_68 = input_39;
assign output_69 = input_39;
assign output_70 = input_39;
assign output_71 = input_39;
assign output_72 = input_39;
assign output_73 = input_39;
assign output_74 = input_39;
assign output_75 = input_39;
assign output_76 = input_39;
assign output_77 = input_39;
assign output_78 = input_39;
assign output_79 = input_39;
assign output_80 = input_39;
assign output_81 = input_39;
assign output_82 = input_39;
assign output_83 = input_39;
assign output_84 = input_39;
assign output_85 = input_39;
assign output_86 = input_39;
assign output_87 = input_39;
assign output_88 = input_39;
assign output_89 = input_39;
assign output_90 = input_39;
assign output_91 = input_39;
assign output_92 = input_39;
assign output_93 = input_39;
assign output_94 = input_39;
assign output_95 = input_39;
assign output_0 = input_40;
assign output_1 = input_40;
assign output_2 = input_40;
assign output_3 = input_40;
assign output_4 = input_40;
assign output_5 = input_40;
assign output_6 = input_40;
assign output_7 = input_40;
assign output_8 = input_40;
assign output_9 = input_40;
assign output_10 = input_40;
assign output_11 = input_40;
assign output_12 = input_40;
assign output_13 = input_40;
assign output_14 = input_40;
assign output_15 = input_40;
assign output_16 = input_40;
assign output_17 = input_40;
assign output_18 = input_40;
assign output_19 = input_40;
assign output_20 = input_40;
assign output_21 = input_40;
assign output_22 = input_40;
assign output_23 = input_40;
assign output_24 = input_40;
assign output_25 = input_40;
assign output_26 = input_40;
assign output_27 = input_40;
assign output_28 = input_40;
assign output_29 = input_40;
assign output_30 = input_40;
assign output_31 = input_40;
assign output_32 = input_40;
assign output_33 = input_40;
assign output_34 = input_40;
assign output_35 = input_40;
assign output_36 = input_40;
assign output_37 = input_40;
assign output_38 = input_40;
assign output_39 = input_40;
assign output_40 = input_40;
assign output_41 = input_40;
assign output_42 = input_40;
assign output_43 = input_40;
assign output_44 = input_40;
assign output_45 = input_40;
assign output_46 = input_40;
assign output_47 = input_40;
assign output_48 = input_40;
assign output_49 = input_40;
assign output_50 = input_40;
assign output_51 = input_40;
assign output_52 = input_40;
assign output_53 = input_40;
assign output_54 = input_40;
assign output_55 = input_40;
assign output_56 = input_40;
assign output_57 = input_40;
assign output_58 = input_40;
assign output_59 = input_40;
assign output_60 = input_40;
assign output_61 = input_40;
assign output_62 = input_40;
assign output_63 = input_40;
assign output_64 = input_40;
assign output_65 = input_40;
assign output_66 = input_40;
assign output_67 = input_40;
assign output_68 = input_40;
assign output_69 = input_40;
assign output_70 = input_40;
assign output_71 = input_40;
assign output_72 = input_40;
assign output_73 = input_40;
assign output_74 = input_40;
assign output_75 = input_40;
assign output_76 = input_40;
assign output_77 = input_40;
assign output_78 = input_40;
assign output_79 = input_40;
assign output_80 = input_40;
assign output_81 = input_40;
assign output_82 = input_40;
assign output_83 = input_40;
assign output_84 = input_40;
assign output_85 = input_40;
assign output_86 = input_40;
assign output_87 = input_40;
assign output_88 = input_40;
assign output_89 = input_40;
assign output_90 = input_40;
assign output_91 = input_40;
assign output_92 = input_40;
assign output_93 = input_40;
assign output_94 = input_40;
assign output_95 = input_40;
assign output_0 = input_41;
assign output_1 = input_41;
assign output_2 = input_41;
assign output_3 = input_41;
assign output_4 = input_41;
assign output_5 = input_41;
assign output_6 = input_41;
assign output_7 = input_41;
assign output_8 = input_41;
assign output_9 = input_41;
assign output_10 = input_41;
assign output_11 = input_41;
assign output_12 = input_41;
assign output_13 = input_41;
assign output_14 = input_41;
assign output_15 = input_41;
assign output_16 = input_41;
assign output_17 = input_41;
assign output_18 = input_41;
assign output_19 = input_41;
assign output_20 = input_41;
assign output_21 = input_41;
assign output_22 = input_41;
assign output_23 = input_41;
assign output_24 = input_41;
assign output_25 = input_41;
assign output_26 = input_41;
assign output_27 = input_41;
assign output_28 = input_41;
assign output_29 = input_41;
assign output_30 = input_41;
assign output_31 = input_41;
assign output_32 = input_41;
assign output_33 = input_41;
assign output_34 = input_41;
assign output_35 = input_41;
assign output_36 = input_41;
assign output_37 = input_41;
assign output_38 = input_41;
assign output_39 = input_41;
assign output_40 = input_41;
assign output_41 = input_41;
assign output_42 = input_41;
assign output_43 = input_41;
assign output_44 = input_41;
assign output_45 = input_41;
assign output_46 = input_41;
assign output_47 = input_41;
assign output_48 = input_41;
assign output_49 = input_41;
assign output_50 = input_41;
assign output_51 = input_41;
assign output_52 = input_41;
assign output_53 = input_41;
assign output_54 = input_41;
assign output_55 = input_41;
assign output_56 = input_41;
assign output_57 = input_41;
assign output_58 = input_41;
assign output_59 = input_41;
assign output_60 = input_41;
assign output_61 = input_41;
assign output_62 = input_41;
assign output_63 = input_41;
assign output_64 = input_41;
assign output_65 = input_41;
assign output_66 = input_41;
assign output_67 = input_41;
assign output_68 = input_41;
assign output_69 = input_41;
assign output_70 = input_41;
assign output_71 = input_41;
assign output_72 = input_41;
assign output_73 = input_41;
assign output_74 = input_41;
assign output_75 = input_41;
assign output_76 = input_41;
assign output_77 = input_41;
assign output_78 = input_41;
assign output_79 = input_41;
assign output_80 = input_41;
assign output_81 = input_41;
assign output_82 = input_41;
assign output_83 = input_41;
assign output_84 = input_41;
assign output_85 = input_41;
assign output_86 = input_41;
assign output_87 = input_41;
assign output_88 = input_41;
assign output_89 = input_41;
assign output_90 = input_41;
assign output_91 = input_41;
assign output_92 = input_41;
assign output_93 = input_41;
assign output_94 = input_41;
assign output_95 = input_41;
assign output_0 = input_42;
assign output_1 = input_42;
assign output_2 = input_42;
assign output_3 = input_42;
assign output_4 = input_42;
assign output_5 = input_42;
assign output_6 = input_42;
assign output_7 = input_42;
assign output_8 = input_42;
assign output_9 = input_42;
assign output_10 = input_42;
assign output_11 = input_42;
assign output_12 = input_42;
assign output_13 = input_42;
assign output_14 = input_42;
assign output_15 = input_42;
assign output_16 = input_42;
assign output_17 = input_42;
assign output_18 = input_42;
assign output_19 = input_42;
assign output_20 = input_42;
assign output_21 = input_42;
assign output_22 = input_42;
assign output_23 = input_42;
assign output_24 = input_42;
assign output_25 = input_42;
assign output_26 = input_42;
assign output_27 = input_42;
assign output_28 = input_42;
assign output_29 = input_42;
assign output_30 = input_42;
assign output_31 = input_42;
assign output_32 = input_42;
assign output_33 = input_42;
assign output_34 = input_42;
assign output_35 = input_42;
assign output_36 = input_42;
assign output_37 = input_42;
assign output_38 = input_42;
assign output_39 = input_42;
assign output_40 = input_42;
assign output_41 = input_42;
assign output_42 = input_42;
assign output_43 = input_42;
assign output_44 = input_42;
assign output_45 = input_42;
assign output_46 = input_42;
assign output_47 = input_42;
assign output_48 = input_42;
assign output_49 = input_42;
assign output_50 = input_42;
assign output_51 = input_42;
assign output_52 = input_42;
assign output_53 = input_42;
assign output_54 = input_42;
assign output_55 = input_42;
assign output_56 = input_42;
assign output_57 = input_42;
assign output_58 = input_42;
assign output_59 = input_42;
assign output_60 = input_42;
assign output_61 = input_42;
assign output_62 = input_42;
assign output_63 = input_42;
assign output_64 = input_42;
assign output_65 = input_42;
assign output_66 = input_42;
assign output_67 = input_42;
assign output_68 = input_42;
assign output_69 = input_42;
assign output_70 = input_42;
assign output_71 = input_42;
assign output_72 = input_42;
assign output_73 = input_42;
assign output_74 = input_42;
assign output_75 = input_42;
assign output_76 = input_42;
assign output_77 = input_42;
assign output_78 = input_42;
assign output_79 = input_42;
assign output_80 = input_42;
assign output_81 = input_42;
assign output_82 = input_42;
assign output_83 = input_42;
assign output_84 = input_42;
assign output_85 = input_42;
assign output_86 = input_42;
assign output_87 = input_42;
assign output_88 = input_42;
assign output_89 = input_42;
assign output_90 = input_42;
assign output_91 = input_42;
assign output_92 = input_42;
assign output_93 = input_42;
assign output_94 = input_42;
assign output_95 = input_42;
assign output_0 = input_43;
assign output_1 = input_43;
assign output_2 = input_43;
assign output_3 = input_43;
assign output_4 = input_43;
assign output_5 = input_43;
assign output_6 = input_43;
assign output_7 = input_43;
assign output_8 = input_43;
assign output_9 = input_43;
assign output_10 = input_43;
assign output_11 = input_43;
assign output_12 = input_43;
assign output_13 = input_43;
assign output_14 = input_43;
assign output_15 = input_43;
assign output_16 = input_43;
assign output_17 = input_43;
assign output_18 = input_43;
assign output_19 = input_43;
assign output_20 = input_43;
assign output_21 = input_43;
assign output_22 = input_43;
assign output_23 = input_43;
assign output_24 = input_43;
assign output_25 = input_43;
assign output_26 = input_43;
assign output_27 = input_43;
assign output_28 = input_43;
assign output_29 = input_43;
assign output_30 = input_43;
assign output_31 = input_43;
assign output_32 = input_43;
assign output_33 = input_43;
assign output_34 = input_43;
assign output_35 = input_43;
assign output_36 = input_43;
assign output_37 = input_43;
assign output_38 = input_43;
assign output_39 = input_43;
assign output_40 = input_43;
assign output_41 = input_43;
assign output_42 = input_43;
assign output_43 = input_43;
assign output_44 = input_43;
assign output_45 = input_43;
assign output_46 = input_43;
assign output_47 = input_43;
assign output_48 = input_43;
assign output_49 = input_43;
assign output_50 = input_43;
assign output_51 = input_43;
assign output_52 = input_43;
assign output_53 = input_43;
assign output_54 = input_43;
assign output_55 = input_43;
assign output_56 = input_43;
assign output_57 = input_43;
assign output_58 = input_43;
assign output_59 = input_43;
assign output_60 = input_43;
assign output_61 = input_43;
assign output_62 = input_43;
assign output_63 = input_43;
assign output_64 = input_43;
assign output_65 = input_43;
assign output_66 = input_43;
assign output_67 = input_43;
assign output_68 = input_43;
assign output_69 = input_43;
assign output_70 = input_43;
assign output_71 = input_43;
assign output_72 = input_43;
assign output_73 = input_43;
assign output_74 = input_43;
assign output_75 = input_43;
assign output_76 = input_43;
assign output_77 = input_43;
assign output_78 = input_43;
assign output_79 = input_43;
assign output_80 = input_43;
assign output_81 = input_43;
assign output_82 = input_43;
assign output_83 = input_43;
assign output_84 = input_43;
assign output_85 = input_43;
assign output_86 = input_43;
assign output_87 = input_43;
assign output_88 = input_43;
assign output_89 = input_43;
assign output_90 = input_43;
assign output_91 = input_43;
assign output_92 = input_43;
assign output_93 = input_43;
assign output_94 = input_43;
assign output_95 = input_43;
assign output_0 = input_44;
assign output_1 = input_44;
assign output_2 = input_44;
assign output_3 = input_44;
assign output_4 = input_44;
assign output_5 = input_44;
assign output_6 = input_44;
assign output_7 = input_44;
assign output_8 = input_44;
assign output_9 = input_44;
assign output_10 = input_44;
assign output_11 = input_44;
assign output_12 = input_44;
assign output_13 = input_44;
assign output_14 = input_44;
assign output_15 = input_44;
assign output_16 = input_44;
assign output_17 = input_44;
assign output_18 = input_44;
assign output_19 = input_44;
assign output_20 = input_44;
assign output_21 = input_44;
assign output_22 = input_44;
assign output_23 = input_44;
assign output_24 = input_44;
assign output_25 = input_44;
assign output_26 = input_44;
assign output_27 = input_44;
assign output_28 = input_44;
assign output_29 = input_44;
assign output_30 = input_44;
assign output_31 = input_44;
assign output_32 = input_44;
assign output_33 = input_44;
assign output_34 = input_44;
assign output_35 = input_44;
assign output_36 = input_44;
assign output_37 = input_44;
assign output_38 = input_44;
assign output_39 = input_44;
assign output_40 = input_44;
assign output_41 = input_44;
assign output_42 = input_44;
assign output_43 = input_44;
assign output_44 = input_44;
assign output_45 = input_44;
assign output_46 = input_44;
assign output_47 = input_44;
assign output_48 = input_44;
assign output_49 = input_44;
assign output_50 = input_44;
assign output_51 = input_44;
assign output_52 = input_44;
assign output_53 = input_44;
assign output_54 = input_44;
assign output_55 = input_44;
assign output_56 = input_44;
assign output_57 = input_44;
assign output_58 = input_44;
assign output_59 = input_44;
assign output_60 = input_44;
assign output_61 = input_44;
assign output_62 = input_44;
assign output_63 = input_44;
assign output_64 = input_44;
assign output_65 = input_44;
assign output_66 = input_44;
assign output_67 = input_44;
assign output_68 = input_44;
assign output_69 = input_44;
assign output_70 = input_44;
assign output_71 = input_44;
assign output_72 = input_44;
assign output_73 = input_44;
assign output_74 = input_44;
assign output_75 = input_44;
assign output_76 = input_44;
assign output_77 = input_44;
assign output_78 = input_44;
assign output_79 = input_44;
assign output_80 = input_44;
assign output_81 = input_44;
assign output_82 = input_44;
assign output_83 = input_44;
assign output_84 = input_44;
assign output_85 = input_44;
assign output_86 = input_44;
assign output_87 = input_44;
assign output_88 = input_44;
assign output_89 = input_44;
assign output_90 = input_44;
assign output_91 = input_44;
assign output_92 = input_44;
assign output_93 = input_44;
assign output_94 = input_44;
assign output_95 = input_44;
assign output_0 = input_45;
assign output_1 = input_45;
assign output_2 = input_45;
assign output_3 = input_45;
assign output_4 = input_45;
assign output_5 = input_45;
assign output_6 = input_45;
assign output_7 = input_45;
assign output_8 = input_45;
assign output_9 = input_45;
assign output_10 = input_45;
assign output_11 = input_45;
assign output_12 = input_45;
assign output_13 = input_45;
assign output_14 = input_45;
assign output_15 = input_45;
assign output_16 = input_45;
assign output_17 = input_45;
assign output_18 = input_45;
assign output_19 = input_45;
assign output_20 = input_45;
assign output_21 = input_45;
assign output_22 = input_45;
assign output_23 = input_45;
assign output_24 = input_45;
assign output_25 = input_45;
assign output_26 = input_45;
assign output_27 = input_45;
assign output_28 = input_45;
assign output_29 = input_45;
assign output_30 = input_45;
assign output_31 = input_45;
assign output_32 = input_45;
assign output_33 = input_45;
assign output_34 = input_45;
assign output_35 = input_45;
assign output_36 = input_45;
assign output_37 = input_45;
assign output_38 = input_45;
assign output_39 = input_45;
assign output_40 = input_45;
assign output_41 = input_45;
assign output_42 = input_45;
assign output_43 = input_45;
assign output_44 = input_45;
assign output_45 = input_45;
assign output_46 = input_45;
assign output_47 = input_45;
assign output_48 = input_45;
assign output_49 = input_45;
assign output_50 = input_45;
assign output_51 = input_45;
assign output_52 = input_45;
assign output_53 = input_45;
assign output_54 = input_45;
assign output_55 = input_45;
assign output_56 = input_45;
assign output_57 = input_45;
assign output_58 = input_45;
assign output_59 = input_45;
assign output_60 = input_45;
assign output_61 = input_45;
assign output_62 = input_45;
assign output_63 = input_45;
assign output_64 = input_45;
assign output_65 = input_45;
assign output_66 = input_45;
assign output_67 = input_45;
assign output_68 = input_45;
assign output_69 = input_45;
assign output_70 = input_45;
assign output_71 = input_45;
assign output_72 = input_45;
assign output_73 = input_45;
assign output_74 = input_45;
assign output_75 = input_45;
assign output_76 = input_45;
assign output_77 = input_45;
assign output_78 = input_45;
assign output_79 = input_45;
assign output_80 = input_45;
assign output_81 = input_45;
assign output_82 = input_45;
assign output_83 = input_45;
assign output_84 = input_45;
assign output_85 = input_45;
assign output_86 = input_45;
assign output_87 = input_45;
assign output_88 = input_45;
assign output_89 = input_45;
assign output_90 = input_45;
assign output_91 = input_45;
assign output_92 = input_45;
assign output_93 = input_45;
assign output_94 = input_45;
assign output_95 = input_45;
assign output_0 = input_46;
assign output_1 = input_46;
assign output_2 = input_46;
assign output_3 = input_46;
assign output_4 = input_46;
assign output_5 = input_46;
assign output_6 = input_46;
assign output_7 = input_46;
assign output_8 = input_46;
assign output_9 = input_46;
assign output_10 = input_46;
assign output_11 = input_46;
assign output_12 = input_46;
assign output_13 = input_46;
assign output_14 = input_46;
assign output_15 = input_46;
assign output_16 = input_46;
assign output_17 = input_46;
assign output_18 = input_46;
assign output_19 = input_46;
assign output_20 = input_46;
assign output_21 = input_46;
assign output_22 = input_46;
assign output_23 = input_46;
assign output_24 = input_46;
assign output_25 = input_46;
assign output_26 = input_46;
assign output_27 = input_46;
assign output_28 = input_46;
assign output_29 = input_46;
assign output_30 = input_46;
assign output_31 = input_46;
assign output_32 = input_46;
assign output_33 = input_46;
assign output_34 = input_46;
assign output_35 = input_46;
assign output_36 = input_46;
assign output_37 = input_46;
assign output_38 = input_46;
assign output_39 = input_46;
assign output_40 = input_46;
assign output_41 = input_46;
assign output_42 = input_46;
assign output_43 = input_46;
assign output_44 = input_46;
assign output_45 = input_46;
assign output_46 = input_46;
assign output_47 = input_46;
assign output_48 = input_46;
assign output_49 = input_46;
assign output_50 = input_46;
assign output_51 = input_46;
assign output_52 = input_46;
assign output_53 = input_46;
assign output_54 = input_46;
assign output_55 = input_46;
assign output_56 = input_46;
assign output_57 = input_46;
assign output_58 = input_46;
assign output_59 = input_46;
assign output_60 = input_46;
assign output_61 = input_46;
assign output_62 = input_46;
assign output_63 = input_46;
assign output_64 = input_46;
assign output_65 = input_46;
assign output_66 = input_46;
assign output_67 = input_46;
assign output_68 = input_46;
assign output_69 = input_46;
assign output_70 = input_46;
assign output_71 = input_46;
assign output_72 = input_46;
assign output_73 = input_46;
assign output_74 = input_46;
assign output_75 = input_46;
assign output_76 = input_46;
assign output_77 = input_46;
assign output_78 = input_46;
assign output_79 = input_46;
assign output_80 = input_46;
assign output_81 = input_46;
assign output_82 = input_46;
assign output_83 = input_46;
assign output_84 = input_46;
assign output_85 = input_46;
assign output_86 = input_46;
assign output_87 = input_46;
assign output_88 = input_46;
assign output_89 = input_46;
assign output_90 = input_46;
assign output_91 = input_46;
assign output_92 = input_46;
assign output_93 = input_46;
assign output_94 = input_46;
assign output_95 = input_46;
assign output_0 = input_47;
assign output_1 = input_47;
assign output_2 = input_47;
assign output_3 = input_47;
assign output_4 = input_47;
assign output_5 = input_47;
assign output_6 = input_47;
assign output_7 = input_47;
assign output_8 = input_47;
assign output_9 = input_47;
assign output_10 = input_47;
assign output_11 = input_47;
assign output_12 = input_47;
assign output_13 = input_47;
assign output_14 = input_47;
assign output_15 = input_47;
assign output_16 = input_47;
assign output_17 = input_47;
assign output_18 = input_47;
assign output_19 = input_47;
assign output_20 = input_47;
assign output_21 = input_47;
assign output_22 = input_47;
assign output_23 = input_47;
assign output_24 = input_47;
assign output_25 = input_47;
assign output_26 = input_47;
assign output_27 = input_47;
assign output_28 = input_47;
assign output_29 = input_47;
assign output_30 = input_47;
assign output_31 = input_47;
assign output_32 = input_47;
assign output_33 = input_47;
assign output_34 = input_47;
assign output_35 = input_47;
assign output_36 = input_47;
assign output_37 = input_47;
assign output_38 = input_47;
assign output_39 = input_47;
assign output_40 = input_47;
assign output_41 = input_47;
assign output_42 = input_47;
assign output_43 = input_47;
assign output_44 = input_47;
assign output_45 = input_47;
assign output_46 = input_47;
assign output_47 = input_47;
assign output_48 = input_47;
assign output_49 = input_47;
assign output_50 = input_47;
assign output_51 = input_47;
assign output_52 = input_47;
assign output_53 = input_47;
assign output_54 = input_47;
assign output_55 = input_47;
assign output_56 = input_47;
assign output_57 = input_47;
assign output_58 = input_47;
assign output_59 = input_47;
assign output_60 = input_47;
assign output_61 = input_47;
assign output_62 = input_47;
assign output_63 = input_47;
assign output_64 = input_47;
assign output_65 = input_47;
assign output_66 = input_47;
assign output_67 = input_47;
assign output_68 = input_47;
assign output_69 = input_47;
assign output_70 = input_47;
assign output_71 = input_47;
assign output_72 = input_47;
assign output_73 = input_47;
assign output_74 = input_47;
assign output_75 = input_47;
assign output_76 = input_47;
assign output_77 = input_47;
assign output_78 = input_47;
assign output_79 = input_47;
assign output_80 = input_47;
assign output_81 = input_47;
assign output_82 = input_47;
assign output_83 = input_47;
assign output_84 = input_47;
assign output_85 = input_47;
assign output_86 = input_47;
assign output_87 = input_47;
assign output_88 = input_47;
assign output_89 = input_47;
assign output_90 = input_47;
assign output_91 = input_47;
assign output_92 = input_47;
assign output_93 = input_47;
assign output_94 = input_47;
assign output_95 = input_47;
assign output_0 = input_48;
assign output_1 = input_48;
assign output_2 = input_48;
assign output_3 = input_48;
assign output_4 = input_48;
assign output_5 = input_48;
assign output_6 = input_48;
assign output_7 = input_48;
assign output_8 = input_48;
assign output_9 = input_48;
assign output_10 = input_48;
assign output_11 = input_48;
assign output_12 = input_48;
assign output_13 = input_48;
assign output_14 = input_48;
assign output_15 = input_48;
assign output_16 = input_48;
assign output_17 = input_48;
assign output_18 = input_48;
assign output_19 = input_48;
assign output_20 = input_48;
assign output_21 = input_48;
assign output_22 = input_48;
assign output_23 = input_48;
assign output_24 = input_48;
assign output_25 = input_48;
assign output_26 = input_48;
assign output_27 = input_48;
assign output_28 = input_48;
assign output_29 = input_48;
assign output_30 = input_48;
assign output_31 = input_48;
assign output_32 = input_48;
assign output_33 = input_48;
assign output_34 = input_48;
assign output_35 = input_48;
assign output_36 = input_48;
assign output_37 = input_48;
assign output_38 = input_48;
assign output_39 = input_48;
assign output_40 = input_48;
assign output_41 = input_48;
assign output_42 = input_48;
assign output_43 = input_48;
assign output_44 = input_48;
assign output_45 = input_48;
assign output_46 = input_48;
assign output_47 = input_48;
assign output_48 = input_48;
assign output_49 = input_48;
assign output_50 = input_48;
assign output_51 = input_48;
assign output_52 = input_48;
assign output_53 = input_48;
assign output_54 = input_48;
assign output_55 = input_48;
assign output_56 = input_48;
assign output_57 = input_48;
assign output_58 = input_48;
assign output_59 = input_48;
assign output_60 = input_48;
assign output_61 = input_48;
assign output_62 = input_48;
assign output_63 = input_48;
assign output_64 = input_48;
assign output_65 = input_48;
assign output_66 = input_48;
assign output_67 = input_48;
assign output_68 = input_48;
assign output_69 = input_48;
assign output_70 = input_48;
assign output_71 = input_48;
assign output_72 = input_48;
assign output_73 = input_48;
assign output_74 = input_48;
assign output_75 = input_48;
assign output_76 = input_48;
assign output_77 = input_48;
assign output_78 = input_48;
assign output_79 = input_48;
assign output_80 = input_48;
assign output_81 = input_48;
assign output_82 = input_48;
assign output_83 = input_48;
assign output_84 = input_48;
assign output_85 = input_48;
assign output_86 = input_48;
assign output_87 = input_48;
assign output_88 = input_48;
assign output_89 = input_48;
assign output_90 = input_48;
assign output_91 = input_48;
assign output_92 = input_48;
assign output_93 = input_48;
assign output_94 = input_48;
assign output_95 = input_48;
assign output_0 = input_49;
assign output_1 = input_49;
assign output_2 = input_49;
assign output_3 = input_49;
assign output_4 = input_49;
assign output_5 = input_49;
assign output_6 = input_49;
assign output_7 = input_49;
assign output_8 = input_49;
assign output_9 = input_49;
assign output_10 = input_49;
assign output_11 = input_49;
assign output_12 = input_49;
assign output_13 = input_49;
assign output_14 = input_49;
assign output_15 = input_49;
assign output_16 = input_49;
assign output_17 = input_49;
assign output_18 = input_49;
assign output_19 = input_49;
assign output_20 = input_49;
assign output_21 = input_49;
assign output_22 = input_49;
assign output_23 = input_49;
assign output_24 = input_49;
assign output_25 = input_49;
assign output_26 = input_49;
assign output_27 = input_49;
assign output_28 = input_49;
assign output_29 = input_49;
assign output_30 = input_49;
assign output_31 = input_49;
assign output_32 = input_49;
assign output_33 = input_49;
assign output_34 = input_49;
assign output_35 = input_49;
assign output_36 = input_49;
assign output_37 = input_49;
assign output_38 = input_49;
assign output_39 = input_49;
assign output_40 = input_49;
assign output_41 = input_49;
assign output_42 = input_49;
assign output_43 = input_49;
assign output_44 = input_49;
assign output_45 = input_49;
assign output_46 = input_49;
assign output_47 = input_49;
assign output_48 = input_49;
assign output_49 = input_49;
assign output_50 = input_49;
assign output_51 = input_49;
assign output_52 = input_49;
assign output_53 = input_49;
assign output_54 = input_49;
assign output_55 = input_49;
assign output_56 = input_49;
assign output_57 = input_49;
assign output_58 = input_49;
assign output_59 = input_49;
assign output_60 = input_49;
assign output_61 = input_49;
assign output_62 = input_49;
assign output_63 = input_49;
assign output_64 = input_49;
assign output_65 = input_49;
assign output_66 = input_49;
assign output_67 = input_49;
assign output_68 = input_49;
assign output_69 = input_49;
assign output_70 = input_49;
assign output_71 = input_49;
assign output_72 = input_49;
assign output_73 = input_49;
assign output_74 = input_49;
assign output_75 = input_49;
assign output_76 = input_49;
assign output_77 = input_49;
assign output_78 = input_49;
assign output_79 = input_49;
assign output_80 = input_49;
assign output_81 = input_49;
assign output_82 = input_49;
assign output_83 = input_49;
assign output_84 = input_49;
assign output_85 = input_49;
assign output_86 = input_49;
assign output_87 = input_49;
assign output_88 = input_49;
assign output_89 = input_49;
assign output_90 = input_49;
assign output_91 = input_49;
assign output_92 = input_49;
assign output_93 = input_49;
assign output_94 = input_49;
assign output_95 = input_49;
assign output_0 = input_50;
assign output_1 = input_50;
assign output_2 = input_50;
assign output_3 = input_50;
assign output_4 = input_50;
assign output_5 = input_50;
assign output_6 = input_50;
assign output_7 = input_50;
assign output_8 = input_50;
assign output_9 = input_50;
assign output_10 = input_50;
assign output_11 = input_50;
assign output_12 = input_50;
assign output_13 = input_50;
assign output_14 = input_50;
assign output_15 = input_50;
assign output_16 = input_50;
assign output_17 = input_50;
assign output_18 = input_50;
assign output_19 = input_50;
assign output_20 = input_50;
assign output_21 = input_50;
assign output_22 = input_50;
assign output_23 = input_50;
assign output_24 = input_50;
assign output_25 = input_50;
assign output_26 = input_50;
assign output_27 = input_50;
assign output_28 = input_50;
assign output_29 = input_50;
assign output_30 = input_50;
assign output_31 = input_50;
assign output_32 = input_50;
assign output_33 = input_50;
assign output_34 = input_50;
assign output_35 = input_50;
assign output_36 = input_50;
assign output_37 = input_50;
assign output_38 = input_50;
assign output_39 = input_50;
assign output_40 = input_50;
assign output_41 = input_50;
assign output_42 = input_50;
assign output_43 = input_50;
assign output_44 = input_50;
assign output_45 = input_50;
assign output_46 = input_50;
assign output_47 = input_50;
assign output_48 = input_50;
assign output_49 = input_50;
assign output_50 = input_50;
assign output_51 = input_50;
assign output_52 = input_50;
assign output_53 = input_50;
assign output_54 = input_50;
assign output_55 = input_50;
assign output_56 = input_50;
assign output_57 = input_50;
assign output_58 = input_50;
assign output_59 = input_50;
assign output_60 = input_50;
assign output_61 = input_50;
assign output_62 = input_50;
assign output_63 = input_50;
assign output_64 = input_50;
assign output_65 = input_50;
assign output_66 = input_50;
assign output_67 = input_50;
assign output_68 = input_50;
assign output_69 = input_50;
assign output_70 = input_50;
assign output_71 = input_50;
assign output_72 = input_50;
assign output_73 = input_50;
assign output_74 = input_50;
assign output_75 = input_50;
assign output_76 = input_50;
assign output_77 = input_50;
assign output_78 = input_50;
assign output_79 = input_50;
assign output_80 = input_50;
assign output_81 = input_50;
assign output_82 = input_50;
assign output_83 = input_50;
assign output_84 = input_50;
assign output_85 = input_50;
assign output_86 = input_50;
assign output_87 = input_50;
assign output_88 = input_50;
assign output_89 = input_50;
assign output_90 = input_50;
assign output_91 = input_50;
assign output_92 = input_50;
assign output_93 = input_50;
assign output_94 = input_50;
assign output_95 = input_50;
assign output_0 = input_51;
assign output_1 = input_51;
assign output_2 = input_51;
assign output_3 = input_51;
assign output_4 = input_51;
assign output_5 = input_51;
assign output_6 = input_51;
assign output_7 = input_51;
assign output_8 = input_51;
assign output_9 = input_51;
assign output_10 = input_51;
assign output_11 = input_51;
assign output_12 = input_51;
assign output_13 = input_51;
assign output_14 = input_51;
assign output_15 = input_51;
assign output_16 = input_51;
assign output_17 = input_51;
assign output_18 = input_51;
assign output_19 = input_51;
assign output_20 = input_51;
assign output_21 = input_51;
assign output_22 = input_51;
assign output_23 = input_51;
assign output_24 = input_51;
assign output_25 = input_51;
assign output_26 = input_51;
assign output_27 = input_51;
assign output_28 = input_51;
assign output_29 = input_51;
assign output_30 = input_51;
assign output_31 = input_51;
assign output_32 = input_51;
assign output_33 = input_51;
assign output_34 = input_51;
assign output_35 = input_51;
assign output_36 = input_51;
assign output_37 = input_51;
assign output_38 = input_51;
assign output_39 = input_51;
assign output_40 = input_51;
assign output_41 = input_51;
assign output_42 = input_51;
assign output_43 = input_51;
assign output_44 = input_51;
assign output_45 = input_51;
assign output_46 = input_51;
assign output_47 = input_51;
assign output_48 = input_51;
assign output_49 = input_51;
assign output_50 = input_51;
assign output_51 = input_51;
assign output_52 = input_51;
assign output_53 = input_51;
assign output_54 = input_51;
assign output_55 = input_51;
assign output_56 = input_51;
assign output_57 = input_51;
assign output_58 = input_51;
assign output_59 = input_51;
assign output_60 = input_51;
assign output_61 = input_51;
assign output_62 = input_51;
assign output_63 = input_51;
assign output_64 = input_51;
assign output_65 = input_51;
assign output_66 = input_51;
assign output_67 = input_51;
assign output_68 = input_51;
assign output_69 = input_51;
assign output_70 = input_51;
assign output_71 = input_51;
assign output_72 = input_51;
assign output_73 = input_51;
assign output_74 = input_51;
assign output_75 = input_51;
assign output_76 = input_51;
assign output_77 = input_51;
assign output_78 = input_51;
assign output_79 = input_51;
assign output_80 = input_51;
assign output_81 = input_51;
assign output_82 = input_51;
assign output_83 = input_51;
assign output_84 = input_51;
assign output_85 = input_51;
assign output_86 = input_51;
assign output_87 = input_51;
assign output_88 = input_51;
assign output_89 = input_51;
assign output_90 = input_51;
assign output_91 = input_51;
assign output_92 = input_51;
assign output_93 = input_51;
assign output_94 = input_51;
assign output_95 = input_51;
assign output_0 = input_52;
assign output_1 = input_52;
assign output_2 = input_52;
assign output_3 = input_52;
assign output_4 = input_52;
assign output_5 = input_52;
assign output_6 = input_52;
assign output_7 = input_52;
assign output_8 = input_52;
assign output_9 = input_52;
assign output_10 = input_52;
assign output_11 = input_52;
assign output_12 = input_52;
assign output_13 = input_52;
assign output_14 = input_52;
assign output_15 = input_52;
assign output_16 = input_52;
assign output_17 = input_52;
assign output_18 = input_52;
assign output_19 = input_52;
assign output_20 = input_52;
assign output_21 = input_52;
assign output_22 = input_52;
assign output_23 = input_52;
assign output_24 = input_52;
assign output_25 = input_52;
assign output_26 = input_52;
assign output_27 = input_52;
assign output_28 = input_52;
assign output_29 = input_52;
assign output_30 = input_52;
assign output_31 = input_52;
assign output_32 = input_52;
assign output_33 = input_52;
assign output_34 = input_52;
assign output_35 = input_52;
assign output_36 = input_52;
assign output_37 = input_52;
assign output_38 = input_52;
assign output_39 = input_52;
assign output_40 = input_52;
assign output_41 = input_52;
assign output_42 = input_52;
assign output_43 = input_52;
assign output_44 = input_52;
assign output_45 = input_52;
assign output_46 = input_52;
assign output_47 = input_52;
assign output_48 = input_52;
assign output_49 = input_52;
assign output_50 = input_52;
assign output_51 = input_52;
assign output_52 = input_52;
assign output_53 = input_52;
assign output_54 = input_52;
assign output_55 = input_52;
assign output_56 = input_52;
assign output_57 = input_52;
assign output_58 = input_52;
assign output_59 = input_52;
assign output_60 = input_52;
assign output_61 = input_52;
assign output_62 = input_52;
assign output_63 = input_52;
assign output_64 = input_52;
assign output_65 = input_52;
assign output_66 = input_52;
assign output_67 = input_52;
assign output_68 = input_52;
assign output_69 = input_52;
assign output_70 = input_52;
assign output_71 = input_52;
assign output_72 = input_52;
assign output_73 = input_52;
assign output_74 = input_52;
assign output_75 = input_52;
assign output_76 = input_52;
assign output_77 = input_52;
assign output_78 = input_52;
assign output_79 = input_52;
assign output_80 = input_52;
assign output_81 = input_52;
assign output_82 = input_52;
assign output_83 = input_52;
assign output_84 = input_52;
assign output_85 = input_52;
assign output_86 = input_52;
assign output_87 = input_52;
assign output_88 = input_52;
assign output_89 = input_52;
assign output_90 = input_52;
assign output_91 = input_52;
assign output_92 = input_52;
assign output_93 = input_52;
assign output_94 = input_52;
assign output_95 = input_52;
assign output_0 = input_53;
assign output_1 = input_53;
assign output_2 = input_53;
assign output_3 = input_53;
assign output_4 = input_53;
assign output_5 = input_53;
assign output_6 = input_53;
assign output_7 = input_53;
assign output_8 = input_53;
assign output_9 = input_53;
assign output_10 = input_53;
assign output_11 = input_53;
assign output_12 = input_53;
assign output_13 = input_53;
assign output_14 = input_53;
assign output_15 = input_53;
assign output_16 = input_53;
assign output_17 = input_53;
assign output_18 = input_53;
assign output_19 = input_53;
assign output_20 = input_53;
assign output_21 = input_53;
assign output_22 = input_53;
assign output_23 = input_53;
assign output_24 = input_53;
assign output_25 = input_53;
assign output_26 = input_53;
assign output_27 = input_53;
assign output_28 = input_53;
assign output_29 = input_53;
assign output_30 = input_53;
assign output_31 = input_53;
assign output_32 = input_53;
assign output_33 = input_53;
assign output_34 = input_53;
assign output_35 = input_53;
assign output_36 = input_53;
assign output_37 = input_53;
assign output_38 = input_53;
assign output_39 = input_53;
assign output_40 = input_53;
assign output_41 = input_53;
assign output_42 = input_53;
assign output_43 = input_53;
assign output_44 = input_53;
assign output_45 = input_53;
assign output_46 = input_53;
assign output_47 = input_53;
assign output_48 = input_53;
assign output_49 = input_53;
assign output_50 = input_53;
assign output_51 = input_53;
assign output_52 = input_53;
assign output_53 = input_53;
assign output_54 = input_53;
assign output_55 = input_53;
assign output_56 = input_53;
assign output_57 = input_53;
assign output_58 = input_53;
assign output_59 = input_53;
assign output_60 = input_53;
assign output_61 = input_53;
assign output_62 = input_53;
assign output_63 = input_53;
assign output_64 = input_53;
assign output_65 = input_53;
assign output_66 = input_53;
assign output_67 = input_53;
assign output_68 = input_53;
assign output_69 = input_53;
assign output_70 = input_53;
assign output_71 = input_53;
assign output_72 = input_53;
assign output_73 = input_53;
assign output_74 = input_53;
assign output_75 = input_53;
assign output_76 = input_53;
assign output_77 = input_53;
assign output_78 = input_53;
assign output_79 = input_53;
assign output_80 = input_53;
assign output_81 = input_53;
assign output_82 = input_53;
assign output_83 = input_53;
assign output_84 = input_53;
assign output_85 = input_53;
assign output_86 = input_53;
assign output_87 = input_53;
assign output_88 = input_53;
assign output_89 = input_53;
assign output_90 = input_53;
assign output_91 = input_53;
assign output_92 = input_53;
assign output_93 = input_53;
assign output_94 = input_53;
assign output_95 = input_53;
assign output_0 = input_54;
assign output_1 = input_54;
assign output_2 = input_54;
assign output_3 = input_54;
assign output_4 = input_54;
assign output_5 = input_54;
assign output_6 = input_54;
assign output_7 = input_54;
assign output_8 = input_54;
assign output_9 = input_54;
assign output_10 = input_54;
assign output_11 = input_54;
assign output_12 = input_54;
assign output_13 = input_54;
assign output_14 = input_54;
assign output_15 = input_54;
assign output_16 = input_54;
assign output_17 = input_54;
assign output_18 = input_54;
assign output_19 = input_54;
assign output_20 = input_54;
assign output_21 = input_54;
assign output_22 = input_54;
assign output_23 = input_54;
assign output_24 = input_54;
assign output_25 = input_54;
assign output_26 = input_54;
assign output_27 = input_54;
assign output_28 = input_54;
assign output_29 = input_54;
assign output_30 = input_54;
assign output_31 = input_54;
assign output_32 = input_54;
assign output_33 = input_54;
assign output_34 = input_54;
assign output_35 = input_54;
assign output_36 = input_54;
assign output_37 = input_54;
assign output_38 = input_54;
assign output_39 = input_54;
assign output_40 = input_54;
assign output_41 = input_54;
assign output_42 = input_54;
assign output_43 = input_54;
assign output_44 = input_54;
assign output_45 = input_54;
assign output_46 = input_54;
assign output_47 = input_54;
assign output_48 = input_54;
assign output_49 = input_54;
assign output_50 = input_54;
assign output_51 = input_54;
assign output_52 = input_54;
assign output_53 = input_54;
assign output_54 = input_54;
assign output_55 = input_54;
assign output_56 = input_54;
assign output_57 = input_54;
assign output_58 = input_54;
assign output_59 = input_54;
assign output_60 = input_54;
assign output_61 = input_54;
assign output_62 = input_54;
assign output_63 = input_54;
assign output_64 = input_54;
assign output_65 = input_54;
assign output_66 = input_54;
assign output_67 = input_54;
assign output_68 = input_54;
assign output_69 = input_54;
assign output_70 = input_54;
assign output_71 = input_54;
assign output_72 = input_54;
assign output_73 = input_54;
assign output_74 = input_54;
assign output_75 = input_54;
assign output_76 = input_54;
assign output_77 = input_54;
assign output_78 = input_54;
assign output_79 = input_54;
assign output_80 = input_54;
assign output_81 = input_54;
assign output_82 = input_54;
assign output_83 = input_54;
assign output_84 = input_54;
assign output_85 = input_54;
assign output_86 = input_54;
assign output_87 = input_54;
assign output_88 = input_54;
assign output_89 = input_54;
assign output_90 = input_54;
assign output_91 = input_54;
assign output_92 = input_54;
assign output_93 = input_54;
assign output_94 = input_54;
assign output_95 = input_54;
assign output_0 = input_55;
assign output_1 = input_55;
assign output_2 = input_55;
assign output_3 = input_55;
assign output_4 = input_55;
assign output_5 = input_55;
assign output_6 = input_55;
assign output_7 = input_55;
assign output_8 = input_55;
assign output_9 = input_55;
assign output_10 = input_55;
assign output_11 = input_55;
assign output_12 = input_55;
assign output_13 = input_55;
assign output_14 = input_55;
assign output_15 = input_55;
assign output_16 = input_55;
assign output_17 = input_55;
assign output_18 = input_55;
assign output_19 = input_55;
assign output_20 = input_55;
assign output_21 = input_55;
assign output_22 = input_55;
assign output_23 = input_55;
assign output_24 = input_55;
assign output_25 = input_55;
assign output_26 = input_55;
assign output_27 = input_55;
assign output_28 = input_55;
assign output_29 = input_55;
assign output_30 = input_55;
assign output_31 = input_55;
assign output_32 = input_55;
assign output_33 = input_55;
assign output_34 = input_55;
assign output_35 = input_55;
assign output_36 = input_55;
assign output_37 = input_55;
assign output_38 = input_55;
assign output_39 = input_55;
assign output_40 = input_55;
assign output_41 = input_55;
assign output_42 = input_55;
assign output_43 = input_55;
assign output_44 = input_55;
assign output_45 = input_55;
assign output_46 = input_55;
assign output_47 = input_55;
assign output_48 = input_55;
assign output_49 = input_55;
assign output_50 = input_55;
assign output_51 = input_55;
assign output_52 = input_55;
assign output_53 = input_55;
assign output_54 = input_55;
assign output_55 = input_55;
assign output_56 = input_55;
assign output_57 = input_55;
assign output_58 = input_55;
assign output_59 = input_55;
assign output_60 = input_55;
assign output_61 = input_55;
assign output_62 = input_55;
assign output_63 = input_55;
assign output_64 = input_55;
assign output_65 = input_55;
assign output_66 = input_55;
assign output_67 = input_55;
assign output_68 = input_55;
assign output_69 = input_55;
assign output_70 = input_55;
assign output_71 = input_55;
assign output_72 = input_55;
assign output_73 = input_55;
assign output_74 = input_55;
assign output_75 = input_55;
assign output_76 = input_55;
assign output_77 = input_55;
assign output_78 = input_55;
assign output_79 = input_55;
assign output_80 = input_55;
assign output_81 = input_55;
assign output_82 = input_55;
assign output_83 = input_55;
assign output_84 = input_55;
assign output_85 = input_55;
assign output_86 = input_55;
assign output_87 = input_55;
assign output_88 = input_55;
assign output_89 = input_55;
assign output_90 = input_55;
assign output_91 = input_55;
assign output_92 = input_55;
assign output_93 = input_55;
assign output_94 = input_55;
assign output_95 = input_55;
assign output_0 = input_56;
assign output_1 = input_56;
assign output_2 = input_56;
assign output_3 = input_56;
assign output_4 = input_56;
assign output_5 = input_56;
assign output_6 = input_56;
assign output_7 = input_56;
assign output_8 = input_56;
assign output_9 = input_56;
assign output_10 = input_56;
assign output_11 = input_56;
assign output_12 = input_56;
assign output_13 = input_56;
assign output_14 = input_56;
assign output_15 = input_56;
assign output_16 = input_56;
assign output_17 = input_56;
assign output_18 = input_56;
assign output_19 = input_56;
assign output_20 = input_56;
assign output_21 = input_56;
assign output_22 = input_56;
assign output_23 = input_56;
assign output_24 = input_56;
assign output_25 = input_56;
assign output_26 = input_56;
assign output_27 = input_56;
assign output_28 = input_56;
assign output_29 = input_56;
assign output_30 = input_56;
assign output_31 = input_56;
assign output_32 = input_56;
assign output_33 = input_56;
assign output_34 = input_56;
assign output_35 = input_56;
assign output_36 = input_56;
assign output_37 = input_56;
assign output_38 = input_56;
assign output_39 = input_56;
assign output_40 = input_56;
assign output_41 = input_56;
assign output_42 = input_56;
assign output_43 = input_56;
assign output_44 = input_56;
assign output_45 = input_56;
assign output_46 = input_56;
assign output_47 = input_56;
assign output_48 = input_56;
assign output_49 = input_56;
assign output_50 = input_56;
assign output_51 = input_56;
assign output_52 = input_56;
assign output_53 = input_56;
assign output_54 = input_56;
assign output_55 = input_56;
assign output_56 = input_56;
assign output_57 = input_56;
assign output_58 = input_56;
assign output_59 = input_56;
assign output_60 = input_56;
assign output_61 = input_56;
assign output_62 = input_56;
assign output_63 = input_56;
assign output_64 = input_56;
assign output_65 = input_56;
assign output_66 = input_56;
assign output_67 = input_56;
assign output_68 = input_56;
assign output_69 = input_56;
assign output_70 = input_56;
assign output_71 = input_56;
assign output_72 = input_56;
assign output_73 = input_56;
assign output_74 = input_56;
assign output_75 = input_56;
assign output_76 = input_56;
assign output_77 = input_56;
assign output_78 = input_56;
assign output_79 = input_56;
assign output_80 = input_56;
assign output_81 = input_56;
assign output_82 = input_56;
assign output_83 = input_56;
assign output_84 = input_56;
assign output_85 = input_56;
assign output_86 = input_56;
assign output_87 = input_56;
assign output_88 = input_56;
assign output_89 = input_56;
assign output_90 = input_56;
assign output_91 = input_56;
assign output_92 = input_56;
assign output_93 = input_56;
assign output_94 = input_56;
assign output_95 = input_56;
assign output_0 = input_57;
assign output_1 = input_57;
assign output_2 = input_57;
assign output_3 = input_57;
assign output_4 = input_57;
assign output_5 = input_57;
assign output_6 = input_57;
assign output_7 = input_57;
assign output_8 = input_57;
assign output_9 = input_57;
assign output_10 = input_57;
assign output_11 = input_57;
assign output_12 = input_57;
assign output_13 = input_57;
assign output_14 = input_57;
assign output_15 = input_57;
assign output_16 = input_57;
assign output_17 = input_57;
assign output_18 = input_57;
assign output_19 = input_57;
assign output_20 = input_57;
assign output_21 = input_57;
assign output_22 = input_57;
assign output_23 = input_57;
assign output_24 = input_57;
assign output_25 = input_57;
assign output_26 = input_57;
assign output_27 = input_57;
assign output_28 = input_57;
assign output_29 = input_57;
assign output_30 = input_57;
assign output_31 = input_57;
assign output_32 = input_57;
assign output_33 = input_57;
assign output_34 = input_57;
assign output_35 = input_57;
assign output_36 = input_57;
assign output_37 = input_57;
assign output_38 = input_57;
assign output_39 = input_57;
assign output_40 = input_57;
assign output_41 = input_57;
assign output_42 = input_57;
assign output_43 = input_57;
assign output_44 = input_57;
assign output_45 = input_57;
assign output_46 = input_57;
assign output_47 = input_57;
assign output_48 = input_57;
assign output_49 = input_57;
assign output_50 = input_57;
assign output_51 = input_57;
assign output_52 = input_57;
assign output_53 = input_57;
assign output_54 = input_57;
assign output_55 = input_57;
assign output_56 = input_57;
assign output_57 = input_57;
assign output_58 = input_57;
assign output_59 = input_57;
assign output_60 = input_57;
assign output_61 = input_57;
assign output_62 = input_57;
assign output_63 = input_57;
assign output_64 = input_57;
assign output_65 = input_57;
assign output_66 = input_57;
assign output_67 = input_57;
assign output_68 = input_57;
assign output_69 = input_57;
assign output_70 = input_57;
assign output_71 = input_57;
assign output_72 = input_57;
assign output_73 = input_57;
assign output_74 = input_57;
assign output_75 = input_57;
assign output_76 = input_57;
assign output_77 = input_57;
assign output_78 = input_57;
assign output_79 = input_57;
assign output_80 = input_57;
assign output_81 = input_57;
assign output_82 = input_57;
assign output_83 = input_57;
assign output_84 = input_57;
assign output_85 = input_57;
assign output_86 = input_57;
assign output_87 = input_57;
assign output_88 = input_57;
assign output_89 = input_57;
assign output_90 = input_57;
assign output_91 = input_57;
assign output_92 = input_57;
assign output_93 = input_57;
assign output_94 = input_57;
assign output_95 = input_57;
assign output_0 = input_58;
assign output_1 = input_58;
assign output_2 = input_58;
assign output_3 = input_58;
assign output_4 = input_58;
assign output_5 = input_58;
assign output_6 = input_58;
assign output_7 = input_58;
assign output_8 = input_58;
assign output_9 = input_58;
assign output_10 = input_58;
assign output_11 = input_58;
assign output_12 = input_58;
assign output_13 = input_58;
assign output_14 = input_58;
assign output_15 = input_58;
assign output_16 = input_58;
assign output_17 = input_58;
assign output_18 = input_58;
assign output_19 = input_58;
assign output_20 = input_58;
assign output_21 = input_58;
assign output_22 = input_58;
assign output_23 = input_58;
assign output_24 = input_58;
assign output_25 = input_58;
assign output_26 = input_58;
assign output_27 = input_58;
assign output_28 = input_58;
assign output_29 = input_58;
assign output_30 = input_58;
assign output_31 = input_58;
assign output_32 = input_58;
assign output_33 = input_58;
assign output_34 = input_58;
assign output_35 = input_58;
assign output_36 = input_58;
assign output_37 = input_58;
assign output_38 = input_58;
assign output_39 = input_58;
assign output_40 = input_58;
assign output_41 = input_58;
assign output_42 = input_58;
assign output_43 = input_58;
assign output_44 = input_58;
assign output_45 = input_58;
assign output_46 = input_58;
assign output_47 = input_58;
assign output_48 = input_58;
assign output_49 = input_58;
assign output_50 = input_58;
assign output_51 = input_58;
assign output_52 = input_58;
assign output_53 = input_58;
assign output_54 = input_58;
assign output_55 = input_58;
assign output_56 = input_58;
assign output_57 = input_58;
assign output_58 = input_58;
assign output_59 = input_58;
assign output_60 = input_58;
assign output_61 = input_58;
assign output_62 = input_58;
assign output_63 = input_58;
assign output_64 = input_58;
assign output_65 = input_58;
assign output_66 = input_58;
assign output_67 = input_58;
assign output_68 = input_58;
assign output_69 = input_58;
assign output_70 = input_58;
assign output_71 = input_58;
assign output_72 = input_58;
assign output_73 = input_58;
assign output_74 = input_58;
assign output_75 = input_58;
assign output_76 = input_58;
assign output_77 = input_58;
assign output_78 = input_58;
assign output_79 = input_58;
assign output_80 = input_58;
assign output_81 = input_58;
assign output_82 = input_58;
assign output_83 = input_58;
assign output_84 = input_58;
assign output_85 = input_58;
assign output_86 = input_58;
assign output_87 = input_58;
assign output_88 = input_58;
assign output_89 = input_58;
assign output_90 = input_58;
assign output_91 = input_58;
assign output_92 = input_58;
assign output_93 = input_58;
assign output_94 = input_58;
assign output_95 = input_58;
assign output_0 = input_59;
assign output_1 = input_59;
assign output_2 = input_59;
assign output_3 = input_59;
assign output_4 = input_59;
assign output_5 = input_59;
assign output_6 = input_59;
assign output_7 = input_59;
assign output_8 = input_59;
assign output_9 = input_59;
assign output_10 = input_59;
assign output_11 = input_59;
assign output_12 = input_59;
assign output_13 = input_59;
assign output_14 = input_59;
assign output_15 = input_59;
assign output_16 = input_59;
assign output_17 = input_59;
assign output_18 = input_59;
assign output_19 = input_59;
assign output_20 = input_59;
assign output_21 = input_59;
assign output_22 = input_59;
assign output_23 = input_59;
assign output_24 = input_59;
assign output_25 = input_59;
assign output_26 = input_59;
assign output_27 = input_59;
assign output_28 = input_59;
assign output_29 = input_59;
assign output_30 = input_59;
assign output_31 = input_59;
assign output_32 = input_59;
assign output_33 = input_59;
assign output_34 = input_59;
assign output_35 = input_59;
assign output_36 = input_59;
assign output_37 = input_59;
assign output_38 = input_59;
assign output_39 = input_59;
assign output_40 = input_59;
assign output_41 = input_59;
assign output_42 = input_59;
assign output_43 = input_59;
assign output_44 = input_59;
assign output_45 = input_59;
assign output_46 = input_59;
assign output_47 = input_59;
assign output_48 = input_59;
assign output_49 = input_59;
assign output_50 = input_59;
assign output_51 = input_59;
assign output_52 = input_59;
assign output_53 = input_59;
assign output_54 = input_59;
assign output_55 = input_59;
assign output_56 = input_59;
assign output_57 = input_59;
assign output_58 = input_59;
assign output_59 = input_59;
assign output_60 = input_59;
assign output_61 = input_59;
assign output_62 = input_59;
assign output_63 = input_59;
assign output_64 = input_59;
assign output_65 = input_59;
assign output_66 = input_59;
assign output_67 = input_59;
assign output_68 = input_59;
assign output_69 = input_59;
assign output_70 = input_59;
assign output_71 = input_59;
assign output_72 = input_59;
assign output_73 = input_59;
assign output_74 = input_59;
assign output_75 = input_59;
assign output_76 = input_59;
assign output_77 = input_59;
assign output_78 = input_59;
assign output_79 = input_59;
assign output_80 = input_59;
assign output_81 = input_59;
assign output_82 = input_59;
assign output_83 = input_59;
assign output_84 = input_59;
assign output_85 = input_59;
assign output_86 = input_59;
assign output_87 = input_59;
assign output_88 = input_59;
assign output_89 = input_59;
assign output_90 = input_59;
assign output_91 = input_59;
assign output_92 = input_59;
assign output_93 = input_59;
assign output_94 = input_59;
assign output_95 = input_59;
assign output_0 = input_60;
assign output_1 = input_60;
assign output_2 = input_60;
assign output_3 = input_60;
assign output_4 = input_60;
assign output_5 = input_60;
assign output_6 = input_60;
assign output_7 = input_60;
assign output_8 = input_60;
assign output_9 = input_60;
assign output_10 = input_60;
assign output_11 = input_60;
assign output_12 = input_60;
assign output_13 = input_60;
assign output_14 = input_60;
assign output_15 = input_60;
assign output_16 = input_60;
assign output_17 = input_60;
assign output_18 = input_60;
assign output_19 = input_60;
assign output_20 = input_60;
assign output_21 = input_60;
assign output_22 = input_60;
assign output_23 = input_60;
assign output_24 = input_60;
assign output_25 = input_60;
assign output_26 = input_60;
assign output_27 = input_60;
assign output_28 = input_60;
assign output_29 = input_60;
assign output_30 = input_60;
assign output_31 = input_60;
assign output_32 = input_60;
assign output_33 = input_60;
assign output_34 = input_60;
assign output_35 = input_60;
assign output_36 = input_60;
assign output_37 = input_60;
assign output_38 = input_60;
assign output_39 = input_60;
assign output_40 = input_60;
assign output_41 = input_60;
assign output_42 = input_60;
assign output_43 = input_60;
assign output_44 = input_60;
assign output_45 = input_60;
assign output_46 = input_60;
assign output_47 = input_60;
assign output_48 = input_60;
assign output_49 = input_60;
assign output_50 = input_60;
assign output_51 = input_60;
assign output_52 = input_60;
assign output_53 = input_60;
assign output_54 = input_60;
assign output_55 = input_60;
assign output_56 = input_60;
assign output_57 = input_60;
assign output_58 = input_60;
assign output_59 = input_60;
assign output_60 = input_60;
assign output_61 = input_60;
assign output_62 = input_60;
assign output_63 = input_60;
assign output_64 = input_60;
assign output_65 = input_60;
assign output_66 = input_60;
assign output_67 = input_60;
assign output_68 = input_60;
assign output_69 = input_60;
assign output_70 = input_60;
assign output_71 = input_60;
assign output_72 = input_60;
assign output_73 = input_60;
assign output_74 = input_60;
assign output_75 = input_60;
assign output_76 = input_60;
assign output_77 = input_60;
assign output_78 = input_60;
assign output_79 = input_60;
assign output_80 = input_60;
assign output_81 = input_60;
assign output_82 = input_60;
assign output_83 = input_60;
assign output_84 = input_60;
assign output_85 = input_60;
assign output_86 = input_60;
assign output_87 = input_60;
assign output_88 = input_60;
assign output_89 = input_60;
assign output_90 = input_60;
assign output_91 = input_60;
assign output_92 = input_60;
assign output_93 = input_60;
assign output_94 = input_60;
assign output_95 = input_60;
assign output_0 = input_61;
assign output_1 = input_61;
assign output_2 = input_61;
assign output_3 = input_61;
assign output_4 = input_61;
assign output_5 = input_61;
assign output_6 = input_61;
assign output_7 = input_61;
assign output_8 = input_61;
assign output_9 = input_61;
assign output_10 = input_61;
assign output_11 = input_61;
assign output_12 = input_61;
assign output_13 = input_61;
assign output_14 = input_61;
assign output_15 = input_61;
assign output_16 = input_61;
assign output_17 = input_61;
assign output_18 = input_61;
assign output_19 = input_61;
assign output_20 = input_61;
assign output_21 = input_61;
assign output_22 = input_61;
assign output_23 = input_61;
assign output_24 = input_61;
assign output_25 = input_61;
assign output_26 = input_61;
assign output_27 = input_61;
assign output_28 = input_61;
assign output_29 = input_61;
assign output_30 = input_61;
assign output_31 = input_61;
assign output_32 = input_61;
assign output_33 = input_61;
assign output_34 = input_61;
assign output_35 = input_61;
assign output_36 = input_61;
assign output_37 = input_61;
assign output_38 = input_61;
assign output_39 = input_61;
assign output_40 = input_61;
assign output_41 = input_61;
assign output_42 = input_61;
assign output_43 = input_61;
assign output_44 = input_61;
assign output_45 = input_61;
assign output_46 = input_61;
assign output_47 = input_61;
assign output_48 = input_61;
assign output_49 = input_61;
assign output_50 = input_61;
assign output_51 = input_61;
assign output_52 = input_61;
assign output_53 = input_61;
assign output_54 = input_61;
assign output_55 = input_61;
assign output_56 = input_61;
assign output_57 = input_61;
assign output_58 = input_61;
assign output_59 = input_61;
assign output_60 = input_61;
assign output_61 = input_61;
assign output_62 = input_61;
assign output_63 = input_61;
assign output_64 = input_61;
assign output_65 = input_61;
assign output_66 = input_61;
assign output_67 = input_61;
assign output_68 = input_61;
assign output_69 = input_61;
assign output_70 = input_61;
assign output_71 = input_61;
assign output_72 = input_61;
assign output_73 = input_61;
assign output_74 = input_61;
assign output_75 = input_61;
assign output_76 = input_61;
assign output_77 = input_61;
assign output_78 = input_61;
assign output_79 = input_61;
assign output_80 = input_61;
assign output_81 = input_61;
assign output_82 = input_61;
assign output_83 = input_61;
assign output_84 = input_61;
assign output_85 = input_61;
assign output_86 = input_61;
assign output_87 = input_61;
assign output_88 = input_61;
assign output_89 = input_61;
assign output_90 = input_61;
assign output_91 = input_61;
assign output_92 = input_61;
assign output_93 = input_61;
assign output_94 = input_61;
assign output_95 = input_61;
assign output_0 = input_62;
assign output_1 = input_62;
assign output_2 = input_62;
assign output_3 = input_62;
assign output_4 = input_62;
assign output_5 = input_62;
assign output_6 = input_62;
assign output_7 = input_62;
assign output_8 = input_62;
assign output_9 = input_62;
assign output_10 = input_62;
assign output_11 = input_62;
assign output_12 = input_62;
assign output_13 = input_62;
assign output_14 = input_62;
assign output_15 = input_62;
assign output_16 = input_62;
assign output_17 = input_62;
assign output_18 = input_62;
assign output_19 = input_62;
assign output_20 = input_62;
assign output_21 = input_62;
assign output_22 = input_62;
assign output_23 = input_62;
assign output_24 = input_62;
assign output_25 = input_62;
assign output_26 = input_62;
assign output_27 = input_62;
assign output_28 = input_62;
assign output_29 = input_62;
assign output_30 = input_62;
assign output_31 = input_62;
assign output_32 = input_62;
assign output_33 = input_62;
assign output_34 = input_62;
assign output_35 = input_62;
assign output_36 = input_62;
assign output_37 = input_62;
assign output_38 = input_62;
assign output_39 = input_62;
assign output_40 = input_62;
assign output_41 = input_62;
assign output_42 = input_62;
assign output_43 = input_62;
assign output_44 = input_62;
assign output_45 = input_62;
assign output_46 = input_62;
assign output_47 = input_62;
assign output_48 = input_62;
assign output_49 = input_62;
assign output_50 = input_62;
assign output_51 = input_62;
assign output_52 = input_62;
assign output_53 = input_62;
assign output_54 = input_62;
assign output_55 = input_62;
assign output_56 = input_62;
assign output_57 = input_62;
assign output_58 = input_62;
assign output_59 = input_62;
assign output_60 = input_62;
assign output_61 = input_62;
assign output_62 = input_62;
assign output_63 = input_62;
assign output_64 = input_62;
assign output_65 = input_62;
assign output_66 = input_62;
assign output_67 = input_62;
assign output_68 = input_62;
assign output_69 = input_62;
assign output_70 = input_62;
assign output_71 = input_62;
assign output_72 = input_62;
assign output_73 = input_62;
assign output_74 = input_62;
assign output_75 = input_62;
assign output_76 = input_62;
assign output_77 = input_62;
assign output_78 = input_62;
assign output_79 = input_62;
assign output_80 = input_62;
assign output_81 = input_62;
assign output_82 = input_62;
assign output_83 = input_62;
assign output_84 = input_62;
assign output_85 = input_62;
assign output_86 = input_62;
assign output_87 = input_62;
assign output_88 = input_62;
assign output_89 = input_62;
assign output_90 = input_62;
assign output_91 = input_62;
assign output_92 = input_62;
assign output_93 = input_62;
assign output_94 = input_62;
assign output_95 = input_62;
assign output_0 = input_63;
assign output_1 = input_63;
assign output_2 = input_63;
assign output_3 = input_63;
assign output_4 = input_63;
assign output_5 = input_63;
assign output_6 = input_63;
assign output_7 = input_63;
assign output_8 = input_63;
assign output_9 = input_63;
assign output_10 = input_63;
assign output_11 = input_63;
assign output_12 = input_63;
assign output_13 = input_63;
assign output_14 = input_63;
assign output_15 = input_63;
assign output_16 = input_63;
assign output_17 = input_63;
assign output_18 = input_63;
assign output_19 = input_63;
assign output_20 = input_63;
assign output_21 = input_63;
assign output_22 = input_63;
assign output_23 = input_63;
assign output_24 = input_63;
assign output_25 = input_63;
assign output_26 = input_63;
assign output_27 = input_63;
assign output_28 = input_63;
assign output_29 = input_63;
assign output_30 = input_63;
assign output_31 = input_63;
assign output_32 = input_63;
assign output_33 = input_63;
assign output_34 = input_63;
assign output_35 = input_63;
assign output_36 = input_63;
assign output_37 = input_63;
assign output_38 = input_63;
assign output_39 = input_63;
assign output_40 = input_63;
assign output_41 = input_63;
assign output_42 = input_63;
assign output_43 = input_63;
assign output_44 = input_63;
assign output_45 = input_63;
assign output_46 = input_63;
assign output_47 = input_63;
assign output_48 = input_63;
assign output_49 = input_63;
assign output_50 = input_63;
assign output_51 = input_63;
assign output_52 = input_63;
assign output_53 = input_63;
assign output_54 = input_63;
assign output_55 = input_63;
assign output_56 = input_63;
assign output_57 = input_63;
assign output_58 = input_63;
assign output_59 = input_63;
assign output_60 = input_63;
assign output_61 = input_63;
assign output_62 = input_63;
assign output_63 = input_63;
assign output_64 = input_63;
assign output_65 = input_63;
assign output_66 = input_63;
assign output_67 = input_63;
assign output_68 = input_63;
assign output_69 = input_63;
assign output_70 = input_63;
assign output_71 = input_63;
assign output_72 = input_63;
assign output_73 = input_63;
assign output_74 = input_63;
assign output_75 = input_63;
assign output_76 = input_63;
assign output_77 = input_63;
assign output_78 = input_63;
assign output_79 = input_63;
assign output_80 = input_63;
assign output_81 = input_63;
assign output_82 = input_63;
assign output_83 = input_63;
assign output_84 = input_63;
assign output_85 = input_63;
assign output_86 = input_63;
assign output_87 = input_63;
assign output_88 = input_63;
assign output_89 = input_63;
assign output_90 = input_63;
assign output_91 = input_63;
assign output_92 = input_63;
assign output_93 = input_63;
assign output_94 = input_63;
assign output_95 = input_63;
assign output_0 = input_64;
assign output_1 = input_64;
assign output_2 = input_64;
assign output_3 = input_64;
assign output_4 = input_64;
assign output_5 = input_64;
assign output_6 = input_64;
assign output_7 = input_64;
assign output_8 = input_64;
assign output_9 = input_64;
assign output_10 = input_64;
assign output_11 = input_64;
assign output_12 = input_64;
assign output_13 = input_64;
assign output_14 = input_64;
assign output_15 = input_64;
assign output_16 = input_64;
assign output_17 = input_64;
assign output_18 = input_64;
assign output_19 = input_64;
assign output_20 = input_64;
assign output_21 = input_64;
assign output_22 = input_64;
assign output_23 = input_64;
assign output_24 = input_64;
assign output_25 = input_64;
assign output_26 = input_64;
assign output_27 = input_64;
assign output_28 = input_64;
assign output_29 = input_64;
assign output_30 = input_64;
assign output_31 = input_64;
assign output_32 = input_64;
assign output_33 = input_64;
assign output_34 = input_64;
assign output_35 = input_64;
assign output_36 = input_64;
assign output_37 = input_64;
assign output_38 = input_64;
assign output_39 = input_64;
assign output_40 = input_64;
assign output_41 = input_64;
assign output_42 = input_64;
assign output_43 = input_64;
assign output_44 = input_64;
assign output_45 = input_64;
assign output_46 = input_64;
assign output_47 = input_64;
assign output_48 = input_64;
assign output_49 = input_64;
assign output_50 = input_64;
assign output_51 = input_64;
assign output_52 = input_64;
assign output_53 = input_64;
assign output_54 = input_64;
assign output_55 = input_64;
assign output_56 = input_64;
assign output_57 = input_64;
assign output_58 = input_64;
assign output_59 = input_64;
assign output_60 = input_64;
assign output_61 = input_64;
assign output_62 = input_64;
assign output_63 = input_64;
assign output_64 = input_64;
assign output_65 = input_64;
assign output_66 = input_64;
assign output_67 = input_64;
assign output_68 = input_64;
assign output_69 = input_64;
assign output_70 = input_64;
assign output_71 = input_64;
assign output_72 = input_64;
assign output_73 = input_64;
assign output_74 = input_64;
assign output_75 = input_64;
assign output_76 = input_64;
assign output_77 = input_64;
assign output_78 = input_64;
assign output_79 = input_64;
assign output_80 = input_64;
assign output_81 = input_64;
assign output_82 = input_64;
assign output_83 = input_64;
assign output_84 = input_64;
assign output_85 = input_64;
assign output_86 = input_64;
assign output_87 = input_64;
assign output_88 = input_64;
assign output_89 = input_64;
assign output_90 = input_64;
assign output_91 = input_64;
assign output_92 = input_64;
assign output_93 = input_64;
assign output_94 = input_64;
assign output_95 = input_64;
assign output_0 = input_65;
assign output_1 = input_65;
assign output_2 = input_65;
assign output_3 = input_65;
assign output_4 = input_65;
assign output_5 = input_65;
assign output_6 = input_65;
assign output_7 = input_65;
assign output_8 = input_65;
assign output_9 = input_65;
assign output_10 = input_65;
assign output_11 = input_65;
assign output_12 = input_65;
assign output_13 = input_65;
assign output_14 = input_65;
assign output_15 = input_65;
assign output_16 = input_65;
assign output_17 = input_65;
assign output_18 = input_65;
assign output_19 = input_65;
assign output_20 = input_65;
assign output_21 = input_65;
assign output_22 = input_65;
assign output_23 = input_65;
assign output_24 = input_65;
assign output_25 = input_65;
assign output_26 = input_65;
assign output_27 = input_65;
assign output_28 = input_65;
assign output_29 = input_65;
assign output_30 = input_65;
assign output_31 = input_65;
assign output_32 = input_65;
assign output_33 = input_65;
assign output_34 = input_65;
assign output_35 = input_65;
assign output_36 = input_65;
assign output_37 = input_65;
assign output_38 = input_65;
assign output_39 = input_65;
assign output_40 = input_65;
assign output_41 = input_65;
assign output_42 = input_65;
assign output_43 = input_65;
assign output_44 = input_65;
assign output_45 = input_65;
assign output_46 = input_65;
assign output_47 = input_65;
assign output_48 = input_65;
assign output_49 = input_65;
assign output_50 = input_65;
assign output_51 = input_65;
assign output_52 = input_65;
assign output_53 = input_65;
assign output_54 = input_65;
assign output_55 = input_65;
assign output_56 = input_65;
assign output_57 = input_65;
assign output_58 = input_65;
assign output_59 = input_65;
assign output_60 = input_65;
assign output_61 = input_65;
assign output_62 = input_65;
assign output_63 = input_65;
assign output_64 = input_65;
assign output_65 = input_65;
assign output_66 = input_65;
assign output_67 = input_65;
assign output_68 = input_65;
assign output_69 = input_65;
assign output_70 = input_65;
assign output_71 = input_65;
assign output_72 = input_65;
assign output_73 = input_65;
assign output_74 = input_65;
assign output_75 = input_65;
assign output_76 = input_65;
assign output_77 = input_65;
assign output_78 = input_65;
assign output_79 = input_65;
assign output_80 = input_65;
assign output_81 = input_65;
assign output_82 = input_65;
assign output_83 = input_65;
assign output_84 = input_65;
assign output_85 = input_65;
assign output_86 = input_65;
assign output_87 = input_65;
assign output_88 = input_65;
assign output_89 = input_65;
assign output_90 = input_65;
assign output_91 = input_65;
assign output_92 = input_65;
assign output_93 = input_65;
assign output_94 = input_65;
assign output_95 = input_65;
assign output_0 = input_66;
assign output_1 = input_66;
assign output_2 = input_66;
assign output_3 = input_66;
assign output_4 = input_66;
assign output_5 = input_66;
assign output_6 = input_66;
assign output_7 = input_66;
assign output_8 = input_66;
assign output_9 = input_66;
assign output_10 = input_66;
assign output_11 = input_66;
assign output_12 = input_66;
assign output_13 = input_66;
assign output_14 = input_66;
assign output_15 = input_66;
assign output_16 = input_66;
assign output_17 = input_66;
assign output_18 = input_66;
assign output_19 = input_66;
assign output_20 = input_66;
assign output_21 = input_66;
assign output_22 = input_66;
assign output_23 = input_66;
assign output_24 = input_66;
assign output_25 = input_66;
assign output_26 = input_66;
assign output_27 = input_66;
assign output_28 = input_66;
assign output_29 = input_66;
assign output_30 = input_66;
assign output_31 = input_66;
assign output_32 = input_66;
assign output_33 = input_66;
assign output_34 = input_66;
assign output_35 = input_66;
assign output_36 = input_66;
assign output_37 = input_66;
assign output_38 = input_66;
assign output_39 = input_66;
assign output_40 = input_66;
assign output_41 = input_66;
assign output_42 = input_66;
assign output_43 = input_66;
assign output_44 = input_66;
assign output_45 = input_66;
assign output_46 = input_66;
assign output_47 = input_66;
assign output_48 = input_66;
assign output_49 = input_66;
assign output_50 = input_66;
assign output_51 = input_66;
assign output_52 = input_66;
assign output_53 = input_66;
assign output_54 = input_66;
assign output_55 = input_66;
assign output_56 = input_66;
assign output_57 = input_66;
assign output_58 = input_66;
assign output_59 = input_66;
assign output_60 = input_66;
assign output_61 = input_66;
assign output_62 = input_66;
assign output_63 = input_66;
assign output_64 = input_66;
assign output_65 = input_66;
assign output_66 = input_66;
assign output_67 = input_66;
assign output_68 = input_66;
assign output_69 = input_66;
assign output_70 = input_66;
assign output_71 = input_66;
assign output_72 = input_66;
assign output_73 = input_66;
assign output_74 = input_66;
assign output_75 = input_66;
assign output_76 = input_66;
assign output_77 = input_66;
assign output_78 = input_66;
assign output_79 = input_66;
assign output_80 = input_66;
assign output_81 = input_66;
assign output_82 = input_66;
assign output_83 = input_66;
assign output_84 = input_66;
assign output_85 = input_66;
assign output_86 = input_66;
assign output_87 = input_66;
assign output_88 = input_66;
assign output_89 = input_66;
assign output_90 = input_66;
assign output_91 = input_66;
assign output_92 = input_66;
assign output_93 = input_66;
assign output_94 = input_66;
assign output_95 = input_66;
assign output_0 = input_67;
assign output_1 = input_67;
assign output_2 = input_67;
assign output_3 = input_67;
assign output_4 = input_67;
assign output_5 = input_67;
assign output_6 = input_67;
assign output_7 = input_67;
assign output_8 = input_67;
assign output_9 = input_67;
assign output_10 = input_67;
assign output_11 = input_67;
assign output_12 = input_67;
assign output_13 = input_67;
assign output_14 = input_67;
assign output_15 = input_67;
assign output_16 = input_67;
assign output_17 = input_67;
assign output_18 = input_67;
assign output_19 = input_67;
assign output_20 = input_67;
assign output_21 = input_67;
assign output_22 = input_67;
assign output_23 = input_67;
assign output_24 = input_67;
assign output_25 = input_67;
assign output_26 = input_67;
assign output_27 = input_67;
assign output_28 = input_67;
assign output_29 = input_67;
assign output_30 = input_67;
assign output_31 = input_67;
assign output_32 = input_67;
assign output_33 = input_67;
assign output_34 = input_67;
assign output_35 = input_67;
assign output_36 = input_67;
assign output_37 = input_67;
assign output_38 = input_67;
assign output_39 = input_67;
assign output_40 = input_67;
assign output_41 = input_67;
assign output_42 = input_67;
assign output_43 = input_67;
assign output_44 = input_67;
assign output_45 = input_67;
assign output_46 = input_67;
assign output_47 = input_67;
assign output_48 = input_67;
assign output_49 = input_67;
assign output_50 = input_67;
assign output_51 = input_67;
assign output_52 = input_67;
assign output_53 = input_67;
assign output_54 = input_67;
assign output_55 = input_67;
assign output_56 = input_67;
assign output_57 = input_67;
assign output_58 = input_67;
assign output_59 = input_67;
assign output_60 = input_67;
assign output_61 = input_67;
assign output_62 = input_67;
assign output_63 = input_67;
assign output_64 = input_67;
assign output_65 = input_67;
assign output_66 = input_67;
assign output_67 = input_67;
assign output_68 = input_67;
assign output_69 = input_67;
assign output_70 = input_67;
assign output_71 = input_67;
assign output_72 = input_67;
assign output_73 = input_67;
assign output_74 = input_67;
assign output_75 = input_67;
assign output_76 = input_67;
assign output_77 = input_67;
assign output_78 = input_67;
assign output_79 = input_67;
assign output_80 = input_67;
assign output_81 = input_67;
assign output_82 = input_67;
assign output_83 = input_67;
assign output_84 = input_67;
assign output_85 = input_67;
assign output_86 = input_67;
assign output_87 = input_67;
assign output_88 = input_67;
assign output_89 = input_67;
assign output_90 = input_67;
assign output_91 = input_67;
assign output_92 = input_67;
assign output_93 = input_67;
assign output_94 = input_67;
assign output_95 = input_67;
assign output_0 = input_68;
assign output_1 = input_68;
assign output_2 = input_68;
assign output_3 = input_68;
assign output_4 = input_68;
assign output_5 = input_68;
assign output_6 = input_68;
assign output_7 = input_68;
assign output_8 = input_68;
assign output_9 = input_68;
assign output_10 = input_68;
assign output_11 = input_68;
assign output_12 = input_68;
assign output_13 = input_68;
assign output_14 = input_68;
assign output_15 = input_68;
assign output_16 = input_68;
assign output_17 = input_68;
assign output_18 = input_68;
assign output_19 = input_68;
assign output_20 = input_68;
assign output_21 = input_68;
assign output_22 = input_68;
assign output_23 = input_68;
assign output_24 = input_68;
assign output_25 = input_68;
assign output_26 = input_68;
assign output_27 = input_68;
assign output_28 = input_68;
assign output_29 = input_68;
assign output_30 = input_68;
assign output_31 = input_68;
assign output_32 = input_68;
assign output_33 = input_68;
assign output_34 = input_68;
assign output_35 = input_68;
assign output_36 = input_68;
assign output_37 = input_68;
assign output_38 = input_68;
assign output_39 = input_68;
assign output_40 = input_68;
assign output_41 = input_68;
assign output_42 = input_68;
assign output_43 = input_68;
assign output_44 = input_68;
assign output_45 = input_68;
assign output_46 = input_68;
assign output_47 = input_68;
assign output_48 = input_68;
assign output_49 = input_68;
assign output_50 = input_68;
assign output_51 = input_68;
assign output_52 = input_68;
assign output_53 = input_68;
assign output_54 = input_68;
assign output_55 = input_68;
assign output_56 = input_68;
assign output_57 = input_68;
assign output_58 = input_68;
assign output_59 = input_68;
assign output_60 = input_68;
assign output_61 = input_68;
assign output_62 = input_68;
assign output_63 = input_68;
assign output_64 = input_68;
assign output_65 = input_68;
assign output_66 = input_68;
assign output_67 = input_68;
assign output_68 = input_68;
assign output_69 = input_68;
assign output_70 = input_68;
assign output_71 = input_68;
assign output_72 = input_68;
assign output_73 = input_68;
assign output_74 = input_68;
assign output_75 = input_68;
assign output_76 = input_68;
assign output_77 = input_68;
assign output_78 = input_68;
assign output_79 = input_68;
assign output_80 = input_68;
assign output_81 = input_68;
assign output_82 = input_68;
assign output_83 = input_68;
assign output_84 = input_68;
assign output_85 = input_68;
assign output_86 = input_68;
assign output_87 = input_68;
assign output_88 = input_68;
assign output_89 = input_68;
assign output_90 = input_68;
assign output_91 = input_68;
assign output_92 = input_68;
assign output_93 = input_68;
assign output_94 = input_68;
assign output_95 = input_68;
assign output_0 = input_69;
assign output_1 = input_69;
assign output_2 = input_69;
assign output_3 = input_69;
assign output_4 = input_69;
assign output_5 = input_69;
assign output_6 = input_69;
assign output_7 = input_69;
assign output_8 = input_69;
assign output_9 = input_69;
assign output_10 = input_69;
assign output_11 = input_69;
assign output_12 = input_69;
assign output_13 = input_69;
assign output_14 = input_69;
assign output_15 = input_69;
assign output_16 = input_69;
assign output_17 = input_69;
assign output_18 = input_69;
assign output_19 = input_69;
assign output_20 = input_69;
assign output_21 = input_69;
assign output_22 = input_69;
assign output_23 = input_69;
assign output_24 = input_69;
assign output_25 = input_69;
assign output_26 = input_69;
assign output_27 = input_69;
assign output_28 = input_69;
assign output_29 = input_69;
assign output_30 = input_69;
assign output_31 = input_69;
assign output_32 = input_69;
assign output_33 = input_69;
assign output_34 = input_69;
assign output_35 = input_69;
assign output_36 = input_69;
assign output_37 = input_69;
assign output_38 = input_69;
assign output_39 = input_69;
assign output_40 = input_69;
assign output_41 = input_69;
assign output_42 = input_69;
assign output_43 = input_69;
assign output_44 = input_69;
assign output_45 = input_69;
assign output_46 = input_69;
assign output_47 = input_69;
assign output_48 = input_69;
assign output_49 = input_69;
assign output_50 = input_69;
assign output_51 = input_69;
assign output_52 = input_69;
assign output_53 = input_69;
assign output_54 = input_69;
assign output_55 = input_69;
assign output_56 = input_69;
assign output_57 = input_69;
assign output_58 = input_69;
assign output_59 = input_69;
assign output_60 = input_69;
assign output_61 = input_69;
assign output_62 = input_69;
assign output_63 = input_69;
assign output_64 = input_69;
assign output_65 = input_69;
assign output_66 = input_69;
assign output_67 = input_69;
assign output_68 = input_69;
assign output_69 = input_69;
assign output_70 = input_69;
assign output_71 = input_69;
assign output_72 = input_69;
assign output_73 = input_69;
assign output_74 = input_69;
assign output_75 = input_69;
assign output_76 = input_69;
assign output_77 = input_69;
assign output_78 = input_69;
assign output_79 = input_69;
assign output_80 = input_69;
assign output_81 = input_69;
assign output_82 = input_69;
assign output_83 = input_69;
assign output_84 = input_69;
assign output_85 = input_69;
assign output_86 = input_69;
assign output_87 = input_69;
assign output_88 = input_69;
assign output_89 = input_69;
assign output_90 = input_69;
assign output_91 = input_69;
assign output_92 = input_69;
assign output_93 = input_69;
assign output_94 = input_69;
assign output_95 = input_69;
assign output_0 = input_70;
assign output_1 = input_70;
assign output_2 = input_70;
assign output_3 = input_70;
assign output_4 = input_70;
assign output_5 = input_70;
assign output_6 = input_70;
assign output_7 = input_70;
assign output_8 = input_70;
assign output_9 = input_70;
assign output_10 = input_70;
assign output_11 = input_70;
assign output_12 = input_70;
assign output_13 = input_70;
assign output_14 = input_70;
assign output_15 = input_70;
assign output_16 = input_70;
assign output_17 = input_70;
assign output_18 = input_70;
assign output_19 = input_70;
assign output_20 = input_70;
assign output_21 = input_70;
assign output_22 = input_70;
assign output_23 = input_70;
assign output_24 = input_70;
assign output_25 = input_70;
assign output_26 = input_70;
assign output_27 = input_70;
assign output_28 = input_70;
assign output_29 = input_70;
assign output_30 = input_70;
assign output_31 = input_70;
assign output_32 = input_70;
assign output_33 = input_70;
assign output_34 = input_70;
assign output_35 = input_70;
assign output_36 = input_70;
assign output_37 = input_70;
assign output_38 = input_70;
assign output_39 = input_70;
assign output_40 = input_70;
assign output_41 = input_70;
assign output_42 = input_70;
assign output_43 = input_70;
assign output_44 = input_70;
assign output_45 = input_70;
assign output_46 = input_70;
assign output_47 = input_70;
assign output_48 = input_70;
assign output_49 = input_70;
assign output_50 = input_70;
assign output_51 = input_70;
assign output_52 = input_70;
assign output_53 = input_70;
assign output_54 = input_70;
assign output_55 = input_70;
assign output_56 = input_70;
assign output_57 = input_70;
assign output_58 = input_70;
assign output_59 = input_70;
assign output_60 = input_70;
assign output_61 = input_70;
assign output_62 = input_70;
assign output_63 = input_70;
assign output_64 = input_70;
assign output_65 = input_70;
assign output_66 = input_70;
assign output_67 = input_70;
assign output_68 = input_70;
assign output_69 = input_70;
assign output_70 = input_70;
assign output_71 = input_70;
assign output_72 = input_70;
assign output_73 = input_70;
assign output_74 = input_70;
assign output_75 = input_70;
assign output_76 = input_70;
assign output_77 = input_70;
assign output_78 = input_70;
assign output_79 = input_70;
assign output_80 = input_70;
assign output_81 = input_70;
assign output_82 = input_70;
assign output_83 = input_70;
assign output_84 = input_70;
assign output_85 = input_70;
assign output_86 = input_70;
assign output_87 = input_70;
assign output_88 = input_70;
assign output_89 = input_70;
assign output_90 = input_70;
assign output_91 = input_70;
assign output_92 = input_70;
assign output_93 = input_70;
assign output_94 = input_70;
assign output_95 = input_70;
assign output_0 = input_71;
assign output_1 = input_71;
assign output_2 = input_71;
assign output_3 = input_71;
assign output_4 = input_71;
assign output_5 = input_71;
assign output_6 = input_71;
assign output_7 = input_71;
assign output_8 = input_71;
assign output_9 = input_71;
assign output_10 = input_71;
assign output_11 = input_71;
assign output_12 = input_71;
assign output_13 = input_71;
assign output_14 = input_71;
assign output_15 = input_71;
assign output_16 = input_71;
assign output_17 = input_71;
assign output_18 = input_71;
assign output_19 = input_71;
assign output_20 = input_71;
assign output_21 = input_71;
assign output_22 = input_71;
assign output_23 = input_71;
assign output_24 = input_71;
assign output_25 = input_71;
assign output_26 = input_71;
assign output_27 = input_71;
assign output_28 = input_71;
assign output_29 = input_71;
assign output_30 = input_71;
assign output_31 = input_71;
assign output_32 = input_71;
assign output_33 = input_71;
assign output_34 = input_71;
assign output_35 = input_71;
assign output_36 = input_71;
assign output_37 = input_71;
assign output_38 = input_71;
assign output_39 = input_71;
assign output_40 = input_71;
assign output_41 = input_71;
assign output_42 = input_71;
assign output_43 = input_71;
assign output_44 = input_71;
assign output_45 = input_71;
assign output_46 = input_71;
assign output_47 = input_71;
assign output_48 = input_71;
assign output_49 = input_71;
assign output_50 = input_71;
assign output_51 = input_71;
assign output_52 = input_71;
assign output_53 = input_71;
assign output_54 = input_71;
assign output_55 = input_71;
assign output_56 = input_71;
assign output_57 = input_71;
assign output_58 = input_71;
assign output_59 = input_71;
assign output_60 = input_71;
assign output_61 = input_71;
assign output_62 = input_71;
assign output_63 = input_71;
assign output_64 = input_71;
assign output_65 = input_71;
assign output_66 = input_71;
assign output_67 = input_71;
assign output_68 = input_71;
assign output_69 = input_71;
assign output_70 = input_71;
assign output_71 = input_71;
assign output_72 = input_71;
assign output_73 = input_71;
assign output_74 = input_71;
assign output_75 = input_71;
assign output_76 = input_71;
assign output_77 = input_71;
assign output_78 = input_71;
assign output_79 = input_71;
assign output_80 = input_71;
assign output_81 = input_71;
assign output_82 = input_71;
assign output_83 = input_71;
assign output_84 = input_71;
assign output_85 = input_71;
assign output_86 = input_71;
assign output_87 = input_71;
assign output_88 = input_71;
assign output_89 = input_71;
assign output_90 = input_71;
assign output_91 = input_71;
assign output_92 = input_71;
assign output_93 = input_71;
assign output_94 = input_71;
assign output_95 = input_71;
assign output_0 = input_72;
assign output_1 = input_72;
assign output_2 = input_72;
assign output_3 = input_72;
assign output_4 = input_72;
assign output_5 = input_72;
assign output_6 = input_72;
assign output_7 = input_72;
assign output_8 = input_72;
assign output_9 = input_72;
assign output_10 = input_72;
assign output_11 = input_72;
assign output_12 = input_72;
assign output_13 = input_72;
assign output_14 = input_72;
assign output_15 = input_72;
assign output_16 = input_72;
assign output_17 = input_72;
assign output_18 = input_72;
assign output_19 = input_72;
assign output_20 = input_72;
assign output_21 = input_72;
assign output_22 = input_72;
assign output_23 = input_72;
assign output_24 = input_72;
assign output_25 = input_72;
assign output_26 = input_72;
assign output_27 = input_72;
assign output_28 = input_72;
assign output_29 = input_72;
assign output_30 = input_72;
assign output_31 = input_72;
assign output_32 = input_72;
assign output_33 = input_72;
assign output_34 = input_72;
assign output_35 = input_72;
assign output_36 = input_72;
assign output_37 = input_72;
assign output_38 = input_72;
assign output_39 = input_72;
assign output_40 = input_72;
assign output_41 = input_72;
assign output_42 = input_72;
assign output_43 = input_72;
assign output_44 = input_72;
assign output_45 = input_72;
assign output_46 = input_72;
assign output_47 = input_72;
assign output_48 = input_72;
assign output_49 = input_72;
assign output_50 = input_72;
assign output_51 = input_72;
assign output_52 = input_72;
assign output_53 = input_72;
assign output_54 = input_72;
assign output_55 = input_72;
assign output_56 = input_72;
assign output_57 = input_72;
assign output_58 = input_72;
assign output_59 = input_72;
assign output_60 = input_72;
assign output_61 = input_72;
assign output_62 = input_72;
assign output_63 = input_72;
assign output_64 = input_72;
assign output_65 = input_72;
assign output_66 = input_72;
assign output_67 = input_72;
assign output_68 = input_72;
assign output_69 = input_72;
assign output_70 = input_72;
assign output_71 = input_72;
assign output_72 = input_72;
assign output_73 = input_72;
assign output_74 = input_72;
assign output_75 = input_72;
assign output_76 = input_72;
assign output_77 = input_72;
assign output_78 = input_72;
assign output_79 = input_72;
assign output_80 = input_72;
assign output_81 = input_72;
assign output_82 = input_72;
assign output_83 = input_72;
assign output_84 = input_72;
assign output_85 = input_72;
assign output_86 = input_72;
assign output_87 = input_72;
assign output_88 = input_72;
assign output_89 = input_72;
assign output_90 = input_72;
assign output_91 = input_72;
assign output_92 = input_72;
assign output_93 = input_72;
assign output_94 = input_72;
assign output_95 = input_72;
assign output_0 = input_73;
assign output_1 = input_73;
assign output_2 = input_73;
assign output_3 = input_73;
assign output_4 = input_73;
assign output_5 = input_73;
assign output_6 = input_73;
assign output_7 = input_73;
assign output_8 = input_73;
assign output_9 = input_73;
assign output_10 = input_73;
assign output_11 = input_73;
assign output_12 = input_73;
assign output_13 = input_73;
assign output_14 = input_73;
assign output_15 = input_73;
assign output_16 = input_73;
assign output_17 = input_73;
assign output_18 = input_73;
assign output_19 = input_73;
assign output_20 = input_73;
assign output_21 = input_73;
assign output_22 = input_73;
assign output_23 = input_73;
assign output_24 = input_73;
assign output_25 = input_73;
assign output_26 = input_73;
assign output_27 = input_73;
assign output_28 = input_73;
assign output_29 = input_73;
assign output_30 = input_73;
assign output_31 = input_73;
assign output_32 = input_73;
assign output_33 = input_73;
assign output_34 = input_73;
assign output_35 = input_73;
assign output_36 = input_73;
assign output_37 = input_73;
assign output_38 = input_73;
assign output_39 = input_73;
assign output_40 = input_73;
assign output_41 = input_73;
assign output_42 = input_73;
assign output_43 = input_73;
assign output_44 = input_73;
assign output_45 = input_73;
assign output_46 = input_73;
assign output_47 = input_73;
assign output_48 = input_73;
assign output_49 = input_73;
assign output_50 = input_73;
assign output_51 = input_73;
assign output_52 = input_73;
assign output_53 = input_73;
assign output_54 = input_73;
assign output_55 = input_73;
assign output_56 = input_73;
assign output_57 = input_73;
assign output_58 = input_73;
assign output_59 = input_73;
assign output_60 = input_73;
assign output_61 = input_73;
assign output_62 = input_73;
assign output_63 = input_73;
assign output_64 = input_73;
assign output_65 = input_73;
assign output_66 = input_73;
assign output_67 = input_73;
assign output_68 = input_73;
assign output_69 = input_73;
assign output_70 = input_73;
assign output_71 = input_73;
assign output_72 = input_73;
assign output_73 = input_73;
assign output_74 = input_73;
assign output_75 = input_73;
assign output_76 = input_73;
assign output_77 = input_73;
assign output_78 = input_73;
assign output_79 = input_73;
assign output_80 = input_73;
assign output_81 = input_73;
assign output_82 = input_73;
assign output_83 = input_73;
assign output_84 = input_73;
assign output_85 = input_73;
assign output_86 = input_73;
assign output_87 = input_73;
assign output_88 = input_73;
assign output_89 = input_73;
assign output_90 = input_73;
assign output_91 = input_73;
assign output_92 = input_73;
assign output_93 = input_73;
assign output_94 = input_73;
assign output_95 = input_73;
assign output_0 = input_74;
assign output_1 = input_74;
assign output_2 = input_74;
assign output_3 = input_74;
assign output_4 = input_74;
assign output_5 = input_74;
assign output_6 = input_74;
assign output_7 = input_74;
assign output_8 = input_74;
assign output_9 = input_74;
assign output_10 = input_74;
assign output_11 = input_74;
assign output_12 = input_74;
assign output_13 = input_74;
assign output_14 = input_74;
assign output_15 = input_74;
assign output_16 = input_74;
assign output_17 = input_74;
assign output_18 = input_74;
assign output_19 = input_74;
assign output_20 = input_74;
assign output_21 = input_74;
assign output_22 = input_74;
assign output_23 = input_74;
assign output_24 = input_74;
assign output_25 = input_74;
assign output_26 = input_74;
assign output_27 = input_74;
assign output_28 = input_74;
assign output_29 = input_74;
assign output_30 = input_74;
assign output_31 = input_74;
assign output_32 = input_74;
assign output_33 = input_74;
assign output_34 = input_74;
assign output_35 = input_74;
assign output_36 = input_74;
assign output_37 = input_74;
assign output_38 = input_74;
assign output_39 = input_74;
assign output_40 = input_74;
assign output_41 = input_74;
assign output_42 = input_74;
assign output_43 = input_74;
assign output_44 = input_74;
assign output_45 = input_74;
assign output_46 = input_74;
assign output_47 = input_74;
assign output_48 = input_74;
assign output_49 = input_74;
assign output_50 = input_74;
assign output_51 = input_74;
assign output_52 = input_74;
assign output_53 = input_74;
assign output_54 = input_74;
assign output_55 = input_74;
assign output_56 = input_74;
assign output_57 = input_74;
assign output_58 = input_74;
assign output_59 = input_74;
assign output_60 = input_74;
assign output_61 = input_74;
assign output_62 = input_74;
assign output_63 = input_74;
assign output_64 = input_74;
assign output_65 = input_74;
assign output_66 = input_74;
assign output_67 = input_74;
assign output_68 = input_74;
assign output_69 = input_74;
assign output_70 = input_74;
assign output_71 = input_74;
assign output_72 = input_74;
assign output_73 = input_74;
assign output_74 = input_74;
assign output_75 = input_74;
assign output_76 = input_74;
assign output_77 = input_74;
assign output_78 = input_74;
assign output_79 = input_74;
assign output_80 = input_74;
assign output_81 = input_74;
assign output_82 = input_74;
assign output_83 = input_74;
assign output_84 = input_74;
assign output_85 = input_74;
assign output_86 = input_74;
assign output_87 = input_74;
assign output_88 = input_74;
assign output_89 = input_74;
assign output_90 = input_74;
assign output_91 = input_74;
assign output_92 = input_74;
assign output_93 = input_74;
assign output_94 = input_74;
assign output_95 = input_74;
assign output_0 = input_75;
assign output_1 = input_75;
assign output_2 = input_75;
assign output_3 = input_75;
assign output_4 = input_75;
assign output_5 = input_75;
assign output_6 = input_75;
assign output_7 = input_75;
assign output_8 = input_75;
assign output_9 = input_75;
assign output_10 = input_75;
assign output_11 = input_75;
assign output_12 = input_75;
assign output_13 = input_75;
assign output_14 = input_75;
assign output_15 = input_75;
assign output_16 = input_75;
assign output_17 = input_75;
assign output_18 = input_75;
assign output_19 = input_75;
assign output_20 = input_75;
assign output_21 = input_75;
assign output_22 = input_75;
assign output_23 = input_75;
assign output_24 = input_75;
assign output_25 = input_75;
assign output_26 = input_75;
assign output_27 = input_75;
assign output_28 = input_75;
assign output_29 = input_75;
assign output_30 = input_75;
assign output_31 = input_75;
assign output_32 = input_75;
assign output_33 = input_75;
assign output_34 = input_75;
assign output_35 = input_75;
assign output_36 = input_75;
assign output_37 = input_75;
assign output_38 = input_75;
assign output_39 = input_75;
assign output_40 = input_75;
assign output_41 = input_75;
assign output_42 = input_75;
assign output_43 = input_75;
assign output_44 = input_75;
assign output_45 = input_75;
assign output_46 = input_75;
assign output_47 = input_75;
assign output_48 = input_75;
assign output_49 = input_75;
assign output_50 = input_75;
assign output_51 = input_75;
assign output_52 = input_75;
assign output_53 = input_75;
assign output_54 = input_75;
assign output_55 = input_75;
assign output_56 = input_75;
assign output_57 = input_75;
assign output_58 = input_75;
assign output_59 = input_75;
assign output_60 = input_75;
assign output_61 = input_75;
assign output_62 = input_75;
assign output_63 = input_75;
assign output_64 = input_75;
assign output_65 = input_75;
assign output_66 = input_75;
assign output_67 = input_75;
assign output_68 = input_75;
assign output_69 = input_75;
assign output_70 = input_75;
assign output_71 = input_75;
assign output_72 = input_75;
assign output_73 = input_75;
assign output_74 = input_75;
assign output_75 = input_75;
assign output_76 = input_75;
assign output_77 = input_75;
assign output_78 = input_75;
assign output_79 = input_75;
assign output_80 = input_75;
assign output_81 = input_75;
assign output_82 = input_75;
assign output_83 = input_75;
assign output_84 = input_75;
assign output_85 = input_75;
assign output_86 = input_75;
assign output_87 = input_75;
assign output_88 = input_75;
assign output_89 = input_75;
assign output_90 = input_75;
assign output_91 = input_75;
assign output_92 = input_75;
assign output_93 = input_75;
assign output_94 = input_75;
assign output_95 = input_75;
assign output_0 = input_76;
assign output_1 = input_76;
assign output_2 = input_76;
assign output_3 = input_76;
assign output_4 = input_76;
assign output_5 = input_76;
assign output_6 = input_76;
assign output_7 = input_76;
assign output_8 = input_76;
assign output_9 = input_76;
assign output_10 = input_76;
assign output_11 = input_76;
assign output_12 = input_76;
assign output_13 = input_76;
assign output_14 = input_76;
assign output_15 = input_76;
assign output_16 = input_76;
assign output_17 = input_76;
assign output_18 = input_76;
assign output_19 = input_76;
assign output_20 = input_76;
assign output_21 = input_76;
assign output_22 = input_76;
assign output_23 = input_76;
assign output_24 = input_76;
assign output_25 = input_76;
assign output_26 = input_76;
assign output_27 = input_76;
assign output_28 = input_76;
assign output_29 = input_76;
assign output_30 = input_76;
assign output_31 = input_76;
assign output_32 = input_76;
assign output_33 = input_76;
assign output_34 = input_76;
assign output_35 = input_76;
assign output_36 = input_76;
assign output_37 = input_76;
assign output_38 = input_76;
assign output_39 = input_76;
assign output_40 = input_76;
assign output_41 = input_76;
assign output_42 = input_76;
assign output_43 = input_76;
assign output_44 = input_76;
assign output_45 = input_76;
assign output_46 = input_76;
assign output_47 = input_76;
assign output_48 = input_76;
assign output_49 = input_76;
assign output_50 = input_76;
assign output_51 = input_76;
assign output_52 = input_76;
assign output_53 = input_76;
assign output_54 = input_76;
assign output_55 = input_76;
assign output_56 = input_76;
assign output_57 = input_76;
assign output_58 = input_76;
assign output_59 = input_76;
assign output_60 = input_76;
assign output_61 = input_76;
assign output_62 = input_76;
assign output_63 = input_76;
assign output_64 = input_76;
assign output_65 = input_76;
assign output_66 = input_76;
assign output_67 = input_76;
assign output_68 = input_76;
assign output_69 = input_76;
assign output_70 = input_76;
assign output_71 = input_76;
assign output_72 = input_76;
assign output_73 = input_76;
assign output_74 = input_76;
assign output_75 = input_76;
assign output_76 = input_76;
assign output_77 = input_76;
assign output_78 = input_76;
assign output_79 = input_76;
assign output_80 = input_76;
assign output_81 = input_76;
assign output_82 = input_76;
assign output_83 = input_76;
assign output_84 = input_76;
assign output_85 = input_76;
assign output_86 = input_76;
assign output_87 = input_76;
assign output_88 = input_76;
assign output_89 = input_76;
assign output_90 = input_76;
assign output_91 = input_76;
assign output_92 = input_76;
assign output_93 = input_76;
assign output_94 = input_76;
assign output_95 = input_76;
assign output_0 = input_77;
assign output_1 = input_77;
assign output_2 = input_77;
assign output_3 = input_77;
assign output_4 = input_77;
assign output_5 = input_77;
assign output_6 = input_77;
assign output_7 = input_77;
assign output_8 = input_77;
assign output_9 = input_77;
assign output_10 = input_77;
assign output_11 = input_77;
assign output_12 = input_77;
assign output_13 = input_77;
assign output_14 = input_77;
assign output_15 = input_77;
assign output_16 = input_77;
assign output_17 = input_77;
assign output_18 = input_77;
assign output_19 = input_77;
assign output_20 = input_77;
assign output_21 = input_77;
assign output_22 = input_77;
assign output_23 = input_77;
assign output_24 = input_77;
assign output_25 = input_77;
assign output_26 = input_77;
assign output_27 = input_77;
assign output_28 = input_77;
assign output_29 = input_77;
assign output_30 = input_77;
assign output_31 = input_77;
assign output_32 = input_77;
assign output_33 = input_77;
assign output_34 = input_77;
assign output_35 = input_77;
assign output_36 = input_77;
assign output_37 = input_77;
assign output_38 = input_77;
assign output_39 = input_77;
assign output_40 = input_77;
assign output_41 = input_77;
assign output_42 = input_77;
assign output_43 = input_77;
assign output_44 = input_77;
assign output_45 = input_77;
assign output_46 = input_77;
assign output_47 = input_77;
assign output_48 = input_77;
assign output_49 = input_77;
assign output_50 = input_77;
assign output_51 = input_77;
assign output_52 = input_77;
assign output_53 = input_77;
assign output_54 = input_77;
assign output_55 = input_77;
assign output_56 = input_77;
assign output_57 = input_77;
assign output_58 = input_77;
assign output_59 = input_77;
assign output_60 = input_77;
assign output_61 = input_77;
assign output_62 = input_77;
assign output_63 = input_77;
assign output_64 = input_77;
assign output_65 = input_77;
assign output_66 = input_77;
assign output_67 = input_77;
assign output_68 = input_77;
assign output_69 = input_77;
assign output_70 = input_77;
assign output_71 = input_77;
assign output_72 = input_77;
assign output_73 = input_77;
assign output_74 = input_77;
assign output_75 = input_77;
assign output_76 = input_77;
assign output_77 = input_77;
assign output_78 = input_77;
assign output_79 = input_77;
assign output_80 = input_77;
assign output_81 = input_77;
assign output_82 = input_77;
assign output_83 = input_77;
assign output_84 = input_77;
assign output_85 = input_77;
assign output_86 = input_77;
assign output_87 = input_77;
assign output_88 = input_77;
assign output_89 = input_77;
assign output_90 = input_77;
assign output_91 = input_77;
assign output_92 = input_77;
assign output_93 = input_77;
assign output_94 = input_77;
assign output_95 = input_77;
assign output_0 = input_78;
assign output_1 = input_78;
assign output_2 = input_78;
assign output_3 = input_78;
assign output_4 = input_78;
assign output_5 = input_78;
assign output_6 = input_78;
assign output_7 = input_78;
assign output_8 = input_78;
assign output_9 = input_78;
assign output_10 = input_78;
assign output_11 = input_78;
assign output_12 = input_78;
assign output_13 = input_78;
assign output_14 = input_78;
assign output_15 = input_78;
assign output_16 = input_78;
assign output_17 = input_78;
assign output_18 = input_78;
assign output_19 = input_78;
assign output_20 = input_78;
assign output_21 = input_78;
assign output_22 = input_78;
assign output_23 = input_78;
assign output_24 = input_78;
assign output_25 = input_78;
assign output_26 = input_78;
assign output_27 = input_78;
assign output_28 = input_78;
assign output_29 = input_78;
assign output_30 = input_78;
assign output_31 = input_78;
assign output_32 = input_78;
assign output_33 = input_78;
assign output_34 = input_78;
assign output_35 = input_78;
assign output_36 = input_78;
assign output_37 = input_78;
assign output_38 = input_78;
assign output_39 = input_78;
assign output_40 = input_78;
assign output_41 = input_78;
assign output_42 = input_78;
assign output_43 = input_78;
assign output_44 = input_78;
assign output_45 = input_78;
assign output_46 = input_78;
assign output_47 = input_78;
assign output_48 = input_78;
assign output_49 = input_78;
assign output_50 = input_78;
assign output_51 = input_78;
assign output_52 = input_78;
assign output_53 = input_78;
assign output_54 = input_78;
assign output_55 = input_78;
assign output_56 = input_78;
assign output_57 = input_78;
assign output_58 = input_78;
assign output_59 = input_78;
assign output_60 = input_78;
assign output_61 = input_78;
assign output_62 = input_78;
assign output_63 = input_78;
assign output_64 = input_78;
assign output_65 = input_78;
assign output_66 = input_78;
assign output_67 = input_78;
assign output_68 = input_78;
assign output_69 = input_78;
assign output_70 = input_78;
assign output_71 = input_78;
assign output_72 = input_78;
assign output_73 = input_78;
assign output_74 = input_78;
assign output_75 = input_78;
assign output_76 = input_78;
assign output_77 = input_78;
assign output_78 = input_78;
assign output_79 = input_78;
assign output_80 = input_78;
assign output_81 = input_78;
assign output_82 = input_78;
assign output_83 = input_78;
assign output_84 = input_78;
assign output_85 = input_78;
assign output_86 = input_78;
assign output_87 = input_78;
assign output_88 = input_78;
assign output_89 = input_78;
assign output_90 = input_78;
assign output_91 = input_78;
assign output_92 = input_78;
assign output_93 = input_78;
assign output_94 = input_78;
assign output_95 = input_78;
assign output_0 = input_79;
assign output_1 = input_79;
assign output_2 = input_79;
assign output_3 = input_79;
assign output_4 = input_79;
assign output_5 = input_79;
assign output_6 = input_79;
assign output_7 = input_79;
assign output_8 = input_79;
assign output_9 = input_79;
assign output_10 = input_79;
assign output_11 = input_79;
assign output_12 = input_79;
assign output_13 = input_79;
assign output_14 = input_79;
assign output_15 = input_79;
assign output_16 = input_79;
assign output_17 = input_79;
assign output_18 = input_79;
assign output_19 = input_79;
assign output_20 = input_79;
assign output_21 = input_79;
assign output_22 = input_79;
assign output_23 = input_79;
assign output_24 = input_79;
assign output_25 = input_79;
assign output_26 = input_79;
assign output_27 = input_79;
assign output_28 = input_79;
assign output_29 = input_79;
assign output_30 = input_79;
assign output_31 = input_79;
assign output_32 = input_79;
assign output_33 = input_79;
assign output_34 = input_79;
assign output_35 = input_79;
assign output_36 = input_79;
assign output_37 = input_79;
assign output_38 = input_79;
assign output_39 = input_79;
assign output_40 = input_79;
assign output_41 = input_79;
assign output_42 = input_79;
assign output_43 = input_79;
assign output_44 = input_79;
assign output_45 = input_79;
assign output_46 = input_79;
assign output_47 = input_79;
assign output_48 = input_79;
assign output_49 = input_79;
assign output_50 = input_79;
assign output_51 = input_79;
assign output_52 = input_79;
assign output_53 = input_79;
assign output_54 = input_79;
assign output_55 = input_79;
assign output_56 = input_79;
assign output_57 = input_79;
assign output_58 = input_79;
assign output_59 = input_79;
assign output_60 = input_79;
assign output_61 = input_79;
assign output_62 = input_79;
assign output_63 = input_79;
assign output_64 = input_79;
assign output_65 = input_79;
assign output_66 = input_79;
assign output_67 = input_79;
assign output_68 = input_79;
assign output_69 = input_79;
assign output_70 = input_79;
assign output_71 = input_79;
assign output_72 = input_79;
assign output_73 = input_79;
assign output_74 = input_79;
assign output_75 = input_79;
assign output_76 = input_79;
assign output_77 = input_79;
assign output_78 = input_79;
assign output_79 = input_79;
assign output_80 = input_79;
assign output_81 = input_79;
assign output_82 = input_79;
assign output_83 = input_79;
assign output_84 = input_79;
assign output_85 = input_79;
assign output_86 = input_79;
assign output_87 = input_79;
assign output_88 = input_79;
assign output_89 = input_79;
assign output_90 = input_79;
assign output_91 = input_79;
assign output_92 = input_79;
assign output_93 = input_79;
assign output_94 = input_79;
assign output_95 = input_79;
assign output_0 = input_80;
assign output_1 = input_80;
assign output_2 = input_80;
assign output_3 = input_80;
assign output_4 = input_80;
assign output_5 = input_80;
assign output_6 = input_80;
assign output_7 = input_80;
assign output_8 = input_80;
assign output_9 = input_80;
assign output_10 = input_80;
assign output_11 = input_80;
assign output_12 = input_80;
assign output_13 = input_80;
assign output_14 = input_80;
assign output_15 = input_80;
assign output_16 = input_80;
assign output_17 = input_80;
assign output_18 = input_80;
assign output_19 = input_80;
assign output_20 = input_80;
assign output_21 = input_80;
assign output_22 = input_80;
assign output_23 = input_80;
assign output_24 = input_80;
assign output_25 = input_80;
assign output_26 = input_80;
assign output_27 = input_80;
assign output_28 = input_80;
assign output_29 = input_80;
assign output_30 = input_80;
assign output_31 = input_80;
assign output_32 = input_80;
assign output_33 = input_80;
assign output_34 = input_80;
assign output_35 = input_80;
assign output_36 = input_80;
assign output_37 = input_80;
assign output_38 = input_80;
assign output_39 = input_80;
assign output_40 = input_80;
assign output_41 = input_80;
assign output_42 = input_80;
assign output_43 = input_80;
assign output_44 = input_80;
assign output_45 = input_80;
assign output_46 = input_80;
assign output_47 = input_80;
assign output_48 = input_80;
assign output_49 = input_80;
assign output_50 = input_80;
assign output_51 = input_80;
assign output_52 = input_80;
assign output_53 = input_80;
assign output_54 = input_80;
assign output_55 = input_80;
assign output_56 = input_80;
assign output_57 = input_80;
assign output_58 = input_80;
assign output_59 = input_80;
assign output_60 = input_80;
assign output_61 = input_80;
assign output_62 = input_80;
assign output_63 = input_80;
assign output_64 = input_80;
assign output_65 = input_80;
assign output_66 = input_80;
assign output_67 = input_80;
assign output_68 = input_80;
assign output_69 = input_80;
assign output_70 = input_80;
assign output_71 = input_80;
assign output_72 = input_80;
assign output_73 = input_80;
assign output_74 = input_80;
assign output_75 = input_80;
assign output_76 = input_80;
assign output_77 = input_80;
assign output_78 = input_80;
assign output_79 = input_80;
assign output_80 = input_80;
assign output_81 = input_80;
assign output_82 = input_80;
assign output_83 = input_80;
assign output_84 = input_80;
assign output_85 = input_80;
assign output_86 = input_80;
assign output_87 = input_80;
assign output_88 = input_80;
assign output_89 = input_80;
assign output_90 = input_80;
assign output_91 = input_80;
assign output_92 = input_80;
assign output_93 = input_80;
assign output_94 = input_80;
assign output_95 = input_80;
assign output_0 = input_81;
assign output_1 = input_81;
assign output_2 = input_81;
assign output_3 = input_81;
assign output_4 = input_81;
assign output_5 = input_81;
assign output_6 = input_81;
assign output_7 = input_81;
assign output_8 = input_81;
assign output_9 = input_81;
assign output_10 = input_81;
assign output_11 = input_81;
assign output_12 = input_81;
assign output_13 = input_81;
assign output_14 = input_81;
assign output_15 = input_81;
assign output_16 = input_81;
assign output_17 = input_81;
assign output_18 = input_81;
assign output_19 = input_81;
assign output_20 = input_81;
assign output_21 = input_81;
assign output_22 = input_81;
assign output_23 = input_81;
assign output_24 = input_81;
assign output_25 = input_81;
assign output_26 = input_81;
assign output_27 = input_81;
assign output_28 = input_81;
assign output_29 = input_81;
assign output_30 = input_81;
assign output_31 = input_81;
assign output_32 = input_81;
assign output_33 = input_81;
assign output_34 = input_81;
assign output_35 = input_81;
assign output_36 = input_81;
assign output_37 = input_81;
assign output_38 = input_81;
assign output_39 = input_81;
assign output_40 = input_81;
assign output_41 = input_81;
assign output_42 = input_81;
assign output_43 = input_81;
assign output_44 = input_81;
assign output_45 = input_81;
assign output_46 = input_81;
assign output_47 = input_81;
assign output_48 = input_81;
assign output_49 = input_81;
assign output_50 = input_81;
assign output_51 = input_81;
assign output_52 = input_81;
assign output_53 = input_81;
assign output_54 = input_81;
assign output_55 = input_81;
assign output_56 = input_81;
assign output_57 = input_81;
assign output_58 = input_81;
assign output_59 = input_81;
assign output_60 = input_81;
assign output_61 = input_81;
assign output_62 = input_81;
assign output_63 = input_81;
assign output_64 = input_81;
assign output_65 = input_81;
assign output_66 = input_81;
assign output_67 = input_81;
assign output_68 = input_81;
assign output_69 = input_81;
assign output_70 = input_81;
assign output_71 = input_81;
assign output_72 = input_81;
assign output_73 = input_81;
assign output_74 = input_81;
assign output_75 = input_81;
assign output_76 = input_81;
assign output_77 = input_81;
assign output_78 = input_81;
assign output_79 = input_81;
assign output_80 = input_81;
assign output_81 = input_81;
assign output_82 = input_81;
assign output_83 = input_81;
assign output_84 = input_81;
assign output_85 = input_81;
assign output_86 = input_81;
assign output_87 = input_81;
assign output_88 = input_81;
assign output_89 = input_81;
assign output_90 = input_81;
assign output_91 = input_81;
assign output_92 = input_81;
assign output_93 = input_81;
assign output_94 = input_81;
assign output_95 = input_81;
assign output_0 = input_82;
assign output_1 = input_82;
assign output_2 = input_82;
assign output_3 = input_82;
assign output_4 = input_82;
assign output_5 = input_82;
assign output_6 = input_82;
assign output_7 = input_82;
assign output_8 = input_82;
assign output_9 = input_82;
assign output_10 = input_82;
assign output_11 = input_82;
assign output_12 = input_82;
assign output_13 = input_82;
assign output_14 = input_82;
assign output_15 = input_82;
assign output_16 = input_82;
assign output_17 = input_82;
assign output_18 = input_82;
assign output_19 = input_82;
assign output_20 = input_82;
assign output_21 = input_82;
assign output_22 = input_82;
assign output_23 = input_82;
assign output_24 = input_82;
assign output_25 = input_82;
assign output_26 = input_82;
assign output_27 = input_82;
assign output_28 = input_82;
assign output_29 = input_82;
assign output_30 = input_82;
assign output_31 = input_82;
assign output_32 = input_82;
assign output_33 = input_82;
assign output_34 = input_82;
assign output_35 = input_82;
assign output_36 = input_82;
assign output_37 = input_82;
assign output_38 = input_82;
assign output_39 = input_82;
assign output_40 = input_82;
assign output_41 = input_82;
assign output_42 = input_82;
assign output_43 = input_82;
assign output_44 = input_82;
assign output_45 = input_82;
assign output_46 = input_82;
assign output_47 = input_82;
assign output_48 = input_82;
assign output_49 = input_82;
assign output_50 = input_82;
assign output_51 = input_82;
assign output_52 = input_82;
assign output_53 = input_82;
assign output_54 = input_82;
assign output_55 = input_82;
assign output_56 = input_82;
assign output_57 = input_82;
assign output_58 = input_82;
assign output_59 = input_82;
assign output_60 = input_82;
assign output_61 = input_82;
assign output_62 = input_82;
assign output_63 = input_82;
assign output_64 = input_82;
assign output_65 = input_82;
assign output_66 = input_82;
assign output_67 = input_82;
assign output_68 = input_82;
assign output_69 = input_82;
assign output_70 = input_82;
assign output_71 = input_82;
assign output_72 = input_82;
assign output_73 = input_82;
assign output_74 = input_82;
assign output_75 = input_82;
assign output_76 = input_82;
assign output_77 = input_82;
assign output_78 = input_82;
assign output_79 = input_82;
assign output_80 = input_82;
assign output_81 = input_82;
assign output_82 = input_82;
assign output_83 = input_82;
assign output_84 = input_82;
assign output_85 = input_82;
assign output_86 = input_82;
assign output_87 = input_82;
assign output_88 = input_82;
assign output_89 = input_82;
assign output_90 = input_82;
assign output_91 = input_82;
assign output_92 = input_82;
assign output_93 = input_82;
assign output_94 = input_82;
assign output_95 = input_82;
assign output_0 = input_83;
assign output_1 = input_83;
assign output_2 = input_83;
assign output_3 = input_83;
assign output_4 = input_83;
assign output_5 = input_83;
assign output_6 = input_83;
assign output_7 = input_83;
assign output_8 = input_83;
assign output_9 = input_83;
assign output_10 = input_83;
assign output_11 = input_83;
assign output_12 = input_83;
assign output_13 = input_83;
assign output_14 = input_83;
assign output_15 = input_83;
assign output_16 = input_83;
assign output_17 = input_83;
assign output_18 = input_83;
assign output_19 = input_83;
assign output_20 = input_83;
assign output_21 = input_83;
assign output_22 = input_83;
assign output_23 = input_83;
assign output_24 = input_83;
assign output_25 = input_83;
assign output_26 = input_83;
assign output_27 = input_83;
assign output_28 = input_83;
assign output_29 = input_83;
assign output_30 = input_83;
assign output_31 = input_83;
assign output_32 = input_83;
assign output_33 = input_83;
assign output_34 = input_83;
assign output_35 = input_83;
assign output_36 = input_83;
assign output_37 = input_83;
assign output_38 = input_83;
assign output_39 = input_83;
assign output_40 = input_83;
assign output_41 = input_83;
assign output_42 = input_83;
assign output_43 = input_83;
assign output_44 = input_83;
assign output_45 = input_83;
assign output_46 = input_83;
assign output_47 = input_83;
assign output_48 = input_83;
assign output_49 = input_83;
assign output_50 = input_83;
assign output_51 = input_83;
assign output_52 = input_83;
assign output_53 = input_83;
assign output_54 = input_83;
assign output_55 = input_83;
assign output_56 = input_83;
assign output_57 = input_83;
assign output_58 = input_83;
assign output_59 = input_83;
assign output_60 = input_83;
assign output_61 = input_83;
assign output_62 = input_83;
assign output_63 = input_83;
assign output_64 = input_83;
assign output_65 = input_83;
assign output_66 = input_83;
assign output_67 = input_83;
assign output_68 = input_83;
assign output_69 = input_83;
assign output_70 = input_83;
assign output_71 = input_83;
assign output_72 = input_83;
assign output_73 = input_83;
assign output_74 = input_83;
assign output_75 = input_83;
assign output_76 = input_83;
assign output_77 = input_83;
assign output_78 = input_83;
assign output_79 = input_83;
assign output_80 = input_83;
assign output_81 = input_83;
assign output_82 = input_83;
assign output_83 = input_83;
assign output_84 = input_83;
assign output_85 = input_83;
assign output_86 = input_83;
assign output_87 = input_83;
assign output_88 = input_83;
assign output_89 = input_83;
assign output_90 = input_83;
assign output_91 = input_83;
assign output_92 = input_83;
assign output_93 = input_83;
assign output_94 = input_83;
assign output_95 = input_83;
assign output_0 = input_84;
assign output_1 = input_84;
assign output_2 = input_84;
assign output_3 = input_84;
assign output_4 = input_84;
assign output_5 = input_84;
assign output_6 = input_84;
assign output_7 = input_84;
assign output_8 = input_84;
assign output_9 = input_84;
assign output_10 = input_84;
assign output_11 = input_84;
assign output_12 = input_84;
assign output_13 = input_84;
assign output_14 = input_84;
assign output_15 = input_84;
assign output_16 = input_84;
assign output_17 = input_84;
assign output_18 = input_84;
assign output_19 = input_84;
assign output_20 = input_84;
assign output_21 = input_84;
assign output_22 = input_84;
assign output_23 = input_84;
assign output_24 = input_84;
assign output_25 = input_84;
assign output_26 = input_84;
assign output_27 = input_84;
assign output_28 = input_84;
assign output_29 = input_84;
assign output_30 = input_84;
assign output_31 = input_84;
assign output_32 = input_84;
assign output_33 = input_84;
assign output_34 = input_84;
assign output_35 = input_84;
assign output_36 = input_84;
assign output_37 = input_84;
assign output_38 = input_84;
assign output_39 = input_84;
assign output_40 = input_84;
assign output_41 = input_84;
assign output_42 = input_84;
assign output_43 = input_84;
assign output_44 = input_84;
assign output_45 = input_84;
assign output_46 = input_84;
assign output_47 = input_84;
assign output_48 = input_84;
assign output_49 = input_84;
assign output_50 = input_84;
assign output_51 = input_84;
assign output_52 = input_84;
assign output_53 = input_84;
assign output_54 = input_84;
assign output_55 = input_84;
assign output_56 = input_84;
assign output_57 = input_84;
assign output_58 = input_84;
assign output_59 = input_84;
assign output_60 = input_84;
assign output_61 = input_84;
assign output_62 = input_84;
assign output_63 = input_84;
assign output_64 = input_84;
assign output_65 = input_84;
assign output_66 = input_84;
assign output_67 = input_84;
assign output_68 = input_84;
assign output_69 = input_84;
assign output_70 = input_84;
assign output_71 = input_84;
assign output_72 = input_84;
assign output_73 = input_84;
assign output_74 = input_84;
assign output_75 = input_84;
assign output_76 = input_84;
assign output_77 = input_84;
assign output_78 = input_84;
assign output_79 = input_84;
assign output_80 = input_84;
assign output_81 = input_84;
assign output_82 = input_84;
assign output_83 = input_84;
assign output_84 = input_84;
assign output_85 = input_84;
assign output_86 = input_84;
assign output_87 = input_84;
assign output_88 = input_84;
assign output_89 = input_84;
assign output_90 = input_84;
assign output_91 = input_84;
assign output_92 = input_84;
assign output_93 = input_84;
assign output_94 = input_84;
assign output_95 = input_84;
assign output_0 = input_85;
assign output_1 = input_85;
assign output_2 = input_85;
assign output_3 = input_85;
assign output_4 = input_85;
assign output_5 = input_85;
assign output_6 = input_85;
assign output_7 = input_85;
assign output_8 = input_85;
assign output_9 = input_85;
assign output_10 = input_85;
assign output_11 = input_85;
assign output_12 = input_85;
assign output_13 = input_85;
assign output_14 = input_85;
assign output_15 = input_85;
assign output_16 = input_85;
assign output_17 = input_85;
assign output_18 = input_85;
assign output_19 = input_85;
assign output_20 = input_85;
assign output_21 = input_85;
assign output_22 = input_85;
assign output_23 = input_85;
assign output_24 = input_85;
assign output_25 = input_85;
assign output_26 = input_85;
assign output_27 = input_85;
assign output_28 = input_85;
assign output_29 = input_85;
assign output_30 = input_85;
assign output_31 = input_85;
assign output_32 = input_85;
assign output_33 = input_85;
assign output_34 = input_85;
assign output_35 = input_85;
assign output_36 = input_85;
assign output_37 = input_85;
assign output_38 = input_85;
assign output_39 = input_85;
assign output_40 = input_85;
assign output_41 = input_85;
assign output_42 = input_85;
assign output_43 = input_85;
assign output_44 = input_85;
assign output_45 = input_85;
assign output_46 = input_85;
assign output_47 = input_85;
assign output_48 = input_85;
assign output_49 = input_85;
assign output_50 = input_85;
assign output_51 = input_85;
assign output_52 = input_85;
assign output_53 = input_85;
assign output_54 = input_85;
assign output_55 = input_85;
assign output_56 = input_85;
assign output_57 = input_85;
assign output_58 = input_85;
assign output_59 = input_85;
assign output_60 = input_85;
assign output_61 = input_85;
assign output_62 = input_85;
assign output_63 = input_85;
assign output_64 = input_85;
assign output_65 = input_85;
assign output_66 = input_85;
assign output_67 = input_85;
assign output_68 = input_85;
assign output_69 = input_85;
assign output_70 = input_85;
assign output_71 = input_85;
assign output_72 = input_85;
assign output_73 = input_85;
assign output_74 = input_85;
assign output_75 = input_85;
assign output_76 = input_85;
assign output_77 = input_85;
assign output_78 = input_85;
assign output_79 = input_85;
assign output_80 = input_85;
assign output_81 = input_85;
assign output_82 = input_85;
assign output_83 = input_85;
assign output_84 = input_85;
assign output_85 = input_85;
assign output_86 = input_85;
assign output_87 = input_85;
assign output_88 = input_85;
assign output_89 = input_85;
assign output_90 = input_85;
assign output_91 = input_85;
assign output_92 = input_85;
assign output_93 = input_85;
assign output_94 = input_85;
assign output_95 = input_85;
assign output_0 = input_86;
assign output_1 = input_86;
assign output_2 = input_86;
assign output_3 = input_86;
assign output_4 = input_86;
assign output_5 = input_86;
assign output_6 = input_86;
assign output_7 = input_86;
assign output_8 = input_86;
assign output_9 = input_86;
assign output_10 = input_86;
assign output_11 = input_86;
assign output_12 = input_86;
assign output_13 = input_86;
assign output_14 = input_86;
assign output_15 = input_86;
assign output_16 = input_86;
assign output_17 = input_86;
assign output_18 = input_86;
assign output_19 = input_86;
assign output_20 = input_86;
assign output_21 = input_86;
assign output_22 = input_86;
assign output_23 = input_86;
assign output_24 = input_86;
assign output_25 = input_86;
assign output_26 = input_86;
assign output_27 = input_86;
assign output_28 = input_86;
assign output_29 = input_86;
assign output_30 = input_86;
assign output_31 = input_86;
assign output_32 = input_86;
assign output_33 = input_86;
assign output_34 = input_86;
assign output_35 = input_86;
assign output_36 = input_86;
assign output_37 = input_86;
assign output_38 = input_86;
assign output_39 = input_86;
assign output_40 = input_86;
assign output_41 = input_86;
assign output_42 = input_86;
assign output_43 = input_86;
assign output_44 = input_86;
assign output_45 = input_86;
assign output_46 = input_86;
assign output_47 = input_86;
assign output_48 = input_86;
assign output_49 = input_86;
assign output_50 = input_86;
assign output_51 = input_86;
assign output_52 = input_86;
assign output_53 = input_86;
assign output_54 = input_86;
assign output_55 = input_86;
assign output_56 = input_86;
assign output_57 = input_86;
assign output_58 = input_86;
assign output_59 = input_86;
assign output_60 = input_86;
assign output_61 = input_86;
assign output_62 = input_86;
assign output_63 = input_86;
assign output_64 = input_86;
assign output_65 = input_86;
assign output_66 = input_86;
assign output_67 = input_86;
assign output_68 = input_86;
assign output_69 = input_86;
assign output_70 = input_86;
assign output_71 = input_86;
assign output_72 = input_86;
assign output_73 = input_86;
assign output_74 = input_86;
assign output_75 = input_86;
assign output_76 = input_86;
assign output_77 = input_86;
assign output_78 = input_86;
assign output_79 = input_86;
assign output_80 = input_86;
assign output_81 = input_86;
assign output_82 = input_86;
assign output_83 = input_86;
assign output_84 = input_86;
assign output_85 = input_86;
assign output_86 = input_86;
assign output_87 = input_86;
assign output_88 = input_86;
assign output_89 = input_86;
assign output_90 = input_86;
assign output_91 = input_86;
assign output_92 = input_86;
assign output_93 = input_86;
assign output_94 = input_86;
assign output_95 = input_86;
assign output_0 = input_87;
assign output_1 = input_87;
assign output_2 = input_87;
assign output_3 = input_87;
assign output_4 = input_87;
assign output_5 = input_87;
assign output_6 = input_87;
assign output_7 = input_87;
assign output_8 = input_87;
assign output_9 = input_87;
assign output_10 = input_87;
assign output_11 = input_87;
assign output_12 = input_87;
assign output_13 = input_87;
assign output_14 = input_87;
assign output_15 = input_87;
assign output_16 = input_87;
assign output_17 = input_87;
assign output_18 = input_87;
assign output_19 = input_87;
assign output_20 = input_87;
assign output_21 = input_87;
assign output_22 = input_87;
assign output_23 = input_87;
assign output_24 = input_87;
assign output_25 = input_87;
assign output_26 = input_87;
assign output_27 = input_87;
assign output_28 = input_87;
assign output_29 = input_87;
assign output_30 = input_87;
assign output_31 = input_87;
assign output_32 = input_87;
assign output_33 = input_87;
assign output_34 = input_87;
assign output_35 = input_87;
assign output_36 = input_87;
assign output_37 = input_87;
assign output_38 = input_87;
assign output_39 = input_87;
assign output_40 = input_87;
assign output_41 = input_87;
assign output_42 = input_87;
assign output_43 = input_87;
assign output_44 = input_87;
assign output_45 = input_87;
assign output_46 = input_87;
assign output_47 = input_87;
assign output_48 = input_87;
assign output_49 = input_87;
assign output_50 = input_87;
assign output_51 = input_87;
assign output_52 = input_87;
assign output_53 = input_87;
assign output_54 = input_87;
assign output_55 = input_87;
assign output_56 = input_87;
assign output_57 = input_87;
assign output_58 = input_87;
assign output_59 = input_87;
assign output_60 = input_87;
assign output_61 = input_87;
assign output_62 = input_87;
assign output_63 = input_87;
assign output_64 = input_87;
assign output_65 = input_87;
assign output_66 = input_87;
assign output_67 = input_87;
assign output_68 = input_87;
assign output_69 = input_87;
assign output_70 = input_87;
assign output_71 = input_87;
assign output_72 = input_87;
assign output_73 = input_87;
assign output_74 = input_87;
assign output_75 = input_87;
assign output_76 = input_87;
assign output_77 = input_87;
assign output_78 = input_87;
assign output_79 = input_87;
assign output_80 = input_87;
assign output_81 = input_87;
assign output_82 = input_87;
assign output_83 = input_87;
assign output_84 = input_87;
assign output_85 = input_87;
assign output_86 = input_87;
assign output_87 = input_87;
assign output_88 = input_87;
assign output_89 = input_87;
assign output_90 = input_87;
assign output_91 = input_87;
assign output_92 = input_87;
assign output_93 = input_87;
assign output_94 = input_87;
assign output_95 = input_87;
assign output_0 = input_88;
assign output_1 = input_88;
assign output_2 = input_88;
assign output_3 = input_88;
assign output_4 = input_88;
assign output_5 = input_88;
assign output_6 = input_88;
assign output_7 = input_88;
assign output_8 = input_88;
assign output_9 = input_88;
assign output_10 = input_88;
assign output_11 = input_88;
assign output_12 = input_88;
assign output_13 = input_88;
assign output_14 = input_88;
assign output_15 = input_88;
assign output_16 = input_88;
assign output_17 = input_88;
assign output_18 = input_88;
assign output_19 = input_88;
assign output_20 = input_88;
assign output_21 = input_88;
assign output_22 = input_88;
assign output_23 = input_88;
assign output_24 = input_88;
assign output_25 = input_88;
assign output_26 = input_88;
assign output_27 = input_88;
assign output_28 = input_88;
assign output_29 = input_88;
assign output_30 = input_88;
assign output_31 = input_88;
assign output_32 = input_88;
assign output_33 = input_88;
assign output_34 = input_88;
assign output_35 = input_88;
assign output_36 = input_88;
assign output_37 = input_88;
assign output_38 = input_88;
assign output_39 = input_88;
assign output_40 = input_88;
assign output_41 = input_88;
assign output_42 = input_88;
assign output_43 = input_88;
assign output_44 = input_88;
assign output_45 = input_88;
assign output_46 = input_88;
assign output_47 = input_88;
assign output_48 = input_88;
assign output_49 = input_88;
assign output_50 = input_88;
assign output_51 = input_88;
assign output_52 = input_88;
assign output_53 = input_88;
assign output_54 = input_88;
assign output_55 = input_88;
assign output_56 = input_88;
assign output_57 = input_88;
assign output_58 = input_88;
assign output_59 = input_88;
assign output_60 = input_88;
assign output_61 = input_88;
assign output_62 = input_88;
assign output_63 = input_88;
assign output_64 = input_88;
assign output_65 = input_88;
assign output_66 = input_88;
assign output_67 = input_88;
assign output_68 = input_88;
assign output_69 = input_88;
assign output_70 = input_88;
assign output_71 = input_88;
assign output_72 = input_88;
assign output_73 = input_88;
assign output_74 = input_88;
assign output_75 = input_88;
assign output_76 = input_88;
assign output_77 = input_88;
assign output_78 = input_88;
assign output_79 = input_88;
assign output_80 = input_88;
assign output_81 = input_88;
assign output_82 = input_88;
assign output_83 = input_88;
assign output_84 = input_88;
assign output_85 = input_88;
assign output_86 = input_88;
assign output_87 = input_88;
assign output_88 = input_88;
assign output_89 = input_88;
assign output_90 = input_88;
assign output_91 = input_88;
assign output_92 = input_88;
assign output_93 = input_88;
assign output_94 = input_88;
assign output_95 = input_88;
assign output_0 = input_89;
assign output_1 = input_89;
assign output_2 = input_89;
assign output_3 = input_89;
assign output_4 = input_89;
assign output_5 = input_89;
assign output_6 = input_89;
assign output_7 = input_89;
assign output_8 = input_89;
assign output_9 = input_89;
assign output_10 = input_89;
assign output_11 = input_89;
assign output_12 = input_89;
assign output_13 = input_89;
assign output_14 = input_89;
assign output_15 = input_89;
assign output_16 = input_89;
assign output_17 = input_89;
assign output_18 = input_89;
assign output_19 = input_89;
assign output_20 = input_89;
assign output_21 = input_89;
assign output_22 = input_89;
assign output_23 = input_89;
assign output_24 = input_89;
assign output_25 = input_89;
assign output_26 = input_89;
assign output_27 = input_89;
assign output_28 = input_89;
assign output_29 = input_89;
assign output_30 = input_89;
assign output_31 = input_89;
assign output_32 = input_89;
assign output_33 = input_89;
assign output_34 = input_89;
assign output_35 = input_89;
assign output_36 = input_89;
assign output_37 = input_89;
assign output_38 = input_89;
assign output_39 = input_89;
assign output_40 = input_89;
assign output_41 = input_89;
assign output_42 = input_89;
assign output_43 = input_89;
assign output_44 = input_89;
assign output_45 = input_89;
assign output_46 = input_89;
assign output_47 = input_89;
assign output_48 = input_89;
assign output_49 = input_89;
assign output_50 = input_89;
assign output_51 = input_89;
assign output_52 = input_89;
assign output_53 = input_89;
assign output_54 = input_89;
assign output_55 = input_89;
assign output_56 = input_89;
assign output_57 = input_89;
assign output_58 = input_89;
assign output_59 = input_89;
assign output_60 = input_89;
assign output_61 = input_89;
assign output_62 = input_89;
assign output_63 = input_89;
assign output_64 = input_89;
assign output_65 = input_89;
assign output_66 = input_89;
assign output_67 = input_89;
assign output_68 = input_89;
assign output_69 = input_89;
assign output_70 = input_89;
assign output_71 = input_89;
assign output_72 = input_89;
assign output_73 = input_89;
assign output_74 = input_89;
assign output_75 = input_89;
assign output_76 = input_89;
assign output_77 = input_89;
assign output_78 = input_89;
assign output_79 = input_89;
assign output_80 = input_89;
assign output_81 = input_89;
assign output_82 = input_89;
assign output_83 = input_89;
assign output_84 = input_89;
assign output_85 = input_89;
assign output_86 = input_89;
assign output_87 = input_89;
assign output_88 = input_89;
assign output_89 = input_89;
assign output_90 = input_89;
assign output_91 = input_89;
assign output_92 = input_89;
assign output_93 = input_89;
assign output_94 = input_89;
assign output_95 = input_89;
assign output_0 = input_90;
assign output_1 = input_90;
assign output_2 = input_90;
assign output_3 = input_90;
assign output_4 = input_90;
assign output_5 = input_90;
assign output_6 = input_90;
assign output_7 = input_90;
assign output_8 = input_90;
assign output_9 = input_90;
assign output_10 = input_90;
assign output_11 = input_90;
assign output_12 = input_90;
assign output_13 = input_90;
assign output_14 = input_90;
assign output_15 = input_90;
assign output_16 = input_90;
assign output_17 = input_90;
assign output_18 = input_90;
assign output_19 = input_90;
assign output_20 = input_90;
assign output_21 = input_90;
assign output_22 = input_90;
assign output_23 = input_90;
assign output_24 = input_90;
assign output_25 = input_90;
assign output_26 = input_90;
assign output_27 = input_90;
assign output_28 = input_90;
assign output_29 = input_90;
assign output_30 = input_90;
assign output_31 = input_90;
assign output_32 = input_90;
assign output_33 = input_90;
assign output_34 = input_90;
assign output_35 = input_90;
assign output_36 = input_90;
assign output_37 = input_90;
assign output_38 = input_90;
assign output_39 = input_90;
assign output_40 = input_90;
assign output_41 = input_90;
assign output_42 = input_90;
assign output_43 = input_90;
assign output_44 = input_90;
assign output_45 = input_90;
assign output_46 = input_90;
assign output_47 = input_90;
assign output_48 = input_90;
assign output_49 = input_90;
assign output_50 = input_90;
assign output_51 = input_90;
assign output_52 = input_90;
assign output_53 = input_90;
assign output_54 = input_90;
assign output_55 = input_90;
assign output_56 = input_90;
assign output_57 = input_90;
assign output_58 = input_90;
assign output_59 = input_90;
assign output_60 = input_90;
assign output_61 = input_90;
assign output_62 = input_90;
assign output_63 = input_90;
assign output_64 = input_90;
assign output_65 = input_90;
assign output_66 = input_90;
assign output_67 = input_90;
assign output_68 = input_90;
assign output_69 = input_90;
assign output_70 = input_90;
assign output_71 = input_90;
assign output_72 = input_90;
assign output_73 = input_90;
assign output_74 = input_90;
assign output_75 = input_90;
assign output_76 = input_90;
assign output_77 = input_90;
assign output_78 = input_90;
assign output_79 = input_90;
assign output_80 = input_90;
assign output_81 = input_90;
assign output_82 = input_90;
assign output_83 = input_90;
assign output_84 = input_90;
assign output_85 = input_90;
assign output_86 = input_90;
assign output_87 = input_90;
assign output_88 = input_90;
assign output_89 = input_90;
assign output_90 = input_90;
assign output_91 = input_90;
assign output_92 = input_90;
assign output_93 = input_90;
assign output_94 = input_90;
assign output_95 = input_90;
assign output_0 = input_91;
assign output_1 = input_91;
assign output_2 = input_91;
assign output_3 = input_91;
assign output_4 = input_91;
assign output_5 = input_91;
assign output_6 = input_91;
assign output_7 = input_91;
assign output_8 = input_91;
assign output_9 = input_91;
assign output_10 = input_91;
assign output_11 = input_91;
assign output_12 = input_91;
assign output_13 = input_91;
assign output_14 = input_91;
assign output_15 = input_91;
assign output_16 = input_91;
assign output_17 = input_91;
assign output_18 = input_91;
assign output_19 = input_91;
assign output_20 = input_91;
assign output_21 = input_91;
assign output_22 = input_91;
assign output_23 = input_91;
assign output_24 = input_91;
assign output_25 = input_91;
assign output_26 = input_91;
assign output_27 = input_91;
assign output_28 = input_91;
assign output_29 = input_91;
assign output_30 = input_91;
assign output_31 = input_91;
assign output_32 = input_91;
assign output_33 = input_91;
assign output_34 = input_91;
assign output_35 = input_91;
assign output_36 = input_91;
assign output_37 = input_91;
assign output_38 = input_91;
assign output_39 = input_91;
assign output_40 = input_91;
assign output_41 = input_91;
assign output_42 = input_91;
assign output_43 = input_91;
assign output_44 = input_91;
assign output_45 = input_91;
assign output_46 = input_91;
assign output_47 = input_91;
assign output_48 = input_91;
assign output_49 = input_91;
assign output_50 = input_91;
assign output_51 = input_91;
assign output_52 = input_91;
assign output_53 = input_91;
assign output_54 = input_91;
assign output_55 = input_91;
assign output_56 = input_91;
assign output_57 = input_91;
assign output_58 = input_91;
assign output_59 = input_91;
assign output_60 = input_91;
assign output_61 = input_91;
assign output_62 = input_91;
assign output_63 = input_91;
assign output_64 = input_91;
assign output_65 = input_91;
assign output_66 = input_91;
assign output_67 = input_91;
assign output_68 = input_91;
assign output_69 = input_91;
assign output_70 = input_91;
assign output_71 = input_91;
assign output_72 = input_91;
assign output_73 = input_91;
assign output_74 = input_91;
assign output_75 = input_91;
assign output_76 = input_91;
assign output_77 = input_91;
assign output_78 = input_91;
assign output_79 = input_91;
assign output_80 = input_91;
assign output_81 = input_91;
assign output_82 = input_91;
assign output_83 = input_91;
assign output_84 = input_91;
assign output_85 = input_91;
assign output_86 = input_91;
assign output_87 = input_91;
assign output_88 = input_91;
assign output_89 = input_91;
assign output_90 = input_91;
assign output_91 = input_91;
assign output_92 = input_91;
assign output_93 = input_91;
assign output_94 = input_91;
assign output_95 = input_91;
assign output_0 = input_92;
assign output_1 = input_92;
assign output_2 = input_92;
assign output_3 = input_92;
assign output_4 = input_92;
assign output_5 = input_92;
assign output_6 = input_92;
assign output_7 = input_92;
assign output_8 = input_92;
assign output_9 = input_92;
assign output_10 = input_92;
assign output_11 = input_92;
assign output_12 = input_92;
assign output_13 = input_92;
assign output_14 = input_92;
assign output_15 = input_92;
assign output_16 = input_92;
assign output_17 = input_92;
assign output_18 = input_92;
assign output_19 = input_92;
assign output_20 = input_92;
assign output_21 = input_92;
assign output_22 = input_92;
assign output_23 = input_92;
assign output_24 = input_92;
assign output_25 = input_92;
assign output_26 = input_92;
assign output_27 = input_92;
assign output_28 = input_92;
assign output_29 = input_92;
assign output_30 = input_92;
assign output_31 = input_92;
assign output_32 = input_92;
assign output_33 = input_92;
assign output_34 = input_92;
assign output_35 = input_92;
assign output_36 = input_92;
assign output_37 = input_92;
assign output_38 = input_92;
assign output_39 = input_92;
assign output_40 = input_92;
assign output_41 = input_92;
assign output_42 = input_92;
assign output_43 = input_92;
assign output_44 = input_92;
assign output_45 = input_92;
assign output_46 = input_92;
assign output_47 = input_92;
assign output_48 = input_92;
assign output_49 = input_92;
assign output_50 = input_92;
assign output_51 = input_92;
assign output_52 = input_92;
assign output_53 = input_92;
assign output_54 = input_92;
assign output_55 = input_92;
assign output_56 = input_92;
assign output_57 = input_92;
assign output_58 = input_92;
assign output_59 = input_92;
assign output_60 = input_92;
assign output_61 = input_92;
assign output_62 = input_92;
assign output_63 = input_92;
assign output_64 = input_92;
assign output_65 = input_92;
assign output_66 = input_92;
assign output_67 = input_92;
assign output_68 = input_92;
assign output_69 = input_92;
assign output_70 = input_92;
assign output_71 = input_92;
assign output_72 = input_92;
assign output_73 = input_92;
assign output_74 = input_92;
assign output_75 = input_92;
assign output_76 = input_92;
assign output_77 = input_92;
assign output_78 = input_92;
assign output_79 = input_92;
assign output_80 = input_92;
assign output_81 = input_92;
assign output_82 = input_92;
assign output_83 = input_92;
assign output_84 = input_92;
assign output_85 = input_92;
assign output_86 = input_92;
assign output_87 = input_92;
assign output_88 = input_92;
assign output_89 = input_92;
assign output_90 = input_92;
assign output_91 = input_92;
assign output_92 = input_92;
assign output_93 = input_92;
assign output_94 = input_92;
assign output_95 = input_92;
assign output_0 = input_93;
assign output_1 = input_93;
assign output_2 = input_93;
assign output_3 = input_93;
assign output_4 = input_93;
assign output_5 = input_93;
assign output_6 = input_93;
assign output_7 = input_93;
assign output_8 = input_93;
assign output_9 = input_93;
assign output_10 = input_93;
assign output_11 = input_93;
assign output_12 = input_93;
assign output_13 = input_93;
assign output_14 = input_93;
assign output_15 = input_93;
assign output_16 = input_93;
assign output_17 = input_93;
assign output_18 = input_93;
assign output_19 = input_93;
assign output_20 = input_93;
assign output_21 = input_93;
assign output_22 = input_93;
assign output_23 = input_93;
assign output_24 = input_93;
assign output_25 = input_93;
assign output_26 = input_93;
assign output_27 = input_93;
assign output_28 = input_93;
assign output_29 = input_93;
assign output_30 = input_93;
assign output_31 = input_93;
assign output_32 = input_93;
assign output_33 = input_93;
assign output_34 = input_93;
assign output_35 = input_93;
assign output_36 = input_93;
assign output_37 = input_93;
assign output_38 = input_93;
assign output_39 = input_93;
assign output_40 = input_93;
assign output_41 = input_93;
assign output_42 = input_93;
assign output_43 = input_93;
assign output_44 = input_93;
assign output_45 = input_93;
assign output_46 = input_93;
assign output_47 = input_93;
assign output_48 = input_93;
assign output_49 = input_93;
assign output_50 = input_93;
assign output_51 = input_93;
assign output_52 = input_93;
assign output_53 = input_93;
assign output_54 = input_93;
assign output_55 = input_93;
assign output_56 = input_93;
assign output_57 = input_93;
assign output_58 = input_93;
assign output_59 = input_93;
assign output_60 = input_93;
assign output_61 = input_93;
assign output_62 = input_93;
assign output_63 = input_93;
assign output_64 = input_93;
assign output_65 = input_93;
assign output_66 = input_93;
assign output_67 = input_93;
assign output_68 = input_93;
assign output_69 = input_93;
assign output_70 = input_93;
assign output_71 = input_93;
assign output_72 = input_93;
assign output_73 = input_93;
assign output_74 = input_93;
assign output_75 = input_93;
assign output_76 = input_93;
assign output_77 = input_93;
assign output_78 = input_93;
assign output_79 = input_93;
assign output_80 = input_93;
assign output_81 = input_93;
assign output_82 = input_93;
assign output_83 = input_93;
assign output_84 = input_93;
assign output_85 = input_93;
assign output_86 = input_93;
assign output_87 = input_93;
assign output_88 = input_93;
assign output_89 = input_93;
assign output_90 = input_93;
assign output_91 = input_93;
assign output_92 = input_93;
assign output_93 = input_93;
assign output_94 = input_93;
assign output_95 = input_93;
assign output_0 = input_94;
assign output_1 = input_94;
assign output_2 = input_94;
assign output_3 = input_94;
assign output_4 = input_94;
assign output_5 = input_94;
assign output_6 = input_94;
assign output_7 = input_94;
assign output_8 = input_94;
assign output_9 = input_94;
assign output_10 = input_94;
assign output_11 = input_94;
assign output_12 = input_94;
assign output_13 = input_94;
assign output_14 = input_94;
assign output_15 = input_94;
assign output_16 = input_94;
assign output_17 = input_94;
assign output_18 = input_94;
assign output_19 = input_94;
assign output_20 = input_94;
assign output_21 = input_94;
assign output_22 = input_94;
assign output_23 = input_94;
assign output_24 = input_94;
assign output_25 = input_94;
assign output_26 = input_94;
assign output_27 = input_94;
assign output_28 = input_94;
assign output_29 = input_94;
assign output_30 = input_94;
assign output_31 = input_94;
assign output_32 = input_94;
assign output_33 = input_94;
assign output_34 = input_94;
assign output_35 = input_94;
assign output_36 = input_94;
assign output_37 = input_94;
assign output_38 = input_94;
assign output_39 = input_94;
assign output_40 = input_94;
assign output_41 = input_94;
assign output_42 = input_94;
assign output_43 = input_94;
assign output_44 = input_94;
assign output_45 = input_94;
assign output_46 = input_94;
assign output_47 = input_94;
assign output_48 = input_94;
assign output_49 = input_94;
assign output_50 = input_94;
assign output_51 = input_94;
assign output_52 = input_94;
assign output_53 = input_94;
assign output_54 = input_94;
assign output_55 = input_94;
assign output_56 = input_94;
assign output_57 = input_94;
assign output_58 = input_94;
assign output_59 = input_94;
assign output_60 = input_94;
assign output_61 = input_94;
assign output_62 = input_94;
assign output_63 = input_94;
assign output_64 = input_94;
assign output_65 = input_94;
assign output_66 = input_94;
assign output_67 = input_94;
assign output_68 = input_94;
assign output_69 = input_94;
assign output_70 = input_94;
assign output_71 = input_94;
assign output_72 = input_94;
assign output_73 = input_94;
assign output_74 = input_94;
assign output_75 = input_94;
assign output_76 = input_94;
assign output_77 = input_94;
assign output_78 = input_94;
assign output_79 = input_94;
assign output_80 = input_94;
assign output_81 = input_94;
assign output_82 = input_94;
assign output_83 = input_94;
assign output_84 = input_94;
assign output_85 = input_94;
assign output_86 = input_94;
assign output_87 = input_94;
assign output_88 = input_94;
assign output_89 = input_94;
assign output_90 = input_94;
assign output_91 = input_94;
assign output_92 = input_94;
assign output_93 = input_94;
assign output_94 = input_94;
assign output_95 = input_94;
assign output_0 = input_95;
assign output_1 = input_95;
assign output_2 = input_95;
assign output_3 = input_95;
assign output_4 = input_95;
assign output_5 = input_95;
assign output_6 = input_95;
assign output_7 = input_95;
assign output_8 = input_95;
assign output_9 = input_95;
assign output_10 = input_95;
assign output_11 = input_95;
assign output_12 = input_95;
assign output_13 = input_95;
assign output_14 = input_95;
assign output_15 = input_95;
assign output_16 = input_95;
assign output_17 = input_95;
assign output_18 = input_95;
assign output_19 = input_95;
assign output_20 = input_95;
assign output_21 = input_95;
assign output_22 = input_95;
assign output_23 = input_95;
assign output_24 = input_95;
assign output_25 = input_95;
assign output_26 = input_95;
assign output_27 = input_95;
assign output_28 = input_95;
assign output_29 = input_95;
assign output_30 = input_95;
assign output_31 = input_95;
assign output_32 = input_95;
assign output_33 = input_95;
assign output_34 = input_95;
assign output_35 = input_95;
assign output_36 = input_95;
assign output_37 = input_95;
assign output_38 = input_95;
assign output_39 = input_95;
assign output_40 = input_95;
assign output_41 = input_95;
assign output_42 = input_95;
assign output_43 = input_95;
assign output_44 = input_95;
assign output_45 = input_95;
assign output_46 = input_95;
assign output_47 = input_95;
assign output_48 = input_95;
assign output_49 = input_95;
assign output_50 = input_95;
assign output_51 = input_95;
assign output_52 = input_95;
assign output_53 = input_95;
assign output_54 = input_95;
assign output_55 = input_95;
assign output_56 = input_95;
assign output_57 = input_95;
assign output_58 = input_95;
assign output_59 = input_95;
assign output_60 = input_95;
assign output_61 = input_95;
assign output_62 = input_95;
assign output_63 = input_95;
assign output_64 = input_95;
assign output_65 = input_95;
assign output_66 = input_95;
assign output_67 = input_95;
assign output_68 = input_95;
assign output_69 = input_95;
assign output_70 = input_95;
assign output_71 = input_95;
assign output_72 = input_95;
assign output_73 = input_95;
assign output_74 = input_95;
assign output_75 = input_95;
assign output_76 = input_95;
assign output_77 = input_95;
assign output_78 = input_95;
assign output_79 = input_95;
assign output_80 = input_95;
assign output_81 = input_95;
assign output_82 = input_95;
assign output_83 = input_95;
assign output_84 = input_95;
assign output_85 = input_95;
assign output_86 = input_95;
assign output_87 = input_95;
assign output_88 = input_95;
assign output_89 = input_95;
assign output_90 = input_95;
assign output_91 = input_95;
assign output_92 = input_95;
assign output_93 = input_95;
assign output_94 = input_95;
assign output_95 = input_95;
endmodule
