module fanout2_braid_16_8 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,output output_8,output output_9,output output_10,output output_11,output output_12,output output_13,output output_14,output output_15,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_9_0, output_9_1, output_8_0;
mixer gate_output_8_0(.a(output_9_0), .b(output_9_1), .y(output_8_0));
wire output_10_0, output_10_1, output_9_0;
mixer gate_output_9_0(.a(output_10_0), .b(output_10_1), .y(output_9_0));
wire output_11_0, output_11_1, output_10_0;
mixer gate_output_10_0(.a(output_11_0), .b(output_11_1), .y(output_10_0));
wire output_12_0, output_12_1, output_11_0;
mixer gate_output_11_0(.a(output_12_0), .b(output_12_1), .y(output_11_0));
wire output_13_0, output_13_1, output_12_0;
mixer gate_output_12_0(.a(output_13_0), .b(output_13_1), .y(output_12_0));
wire output_14_0, output_14_1, output_13_0;
mixer gate_output_13_0(.a(output_14_0), .b(output_14_1), .y(output_13_0));
wire output_15_0, output_15_1, output_14_0;
mixer gate_output_14_0(.a(output_15_0), .b(output_15_1), .y(output_14_0));
wire output_16_0, output_16_1, output_15_0;
mixer gate_output_15_0(.a(output_16_0), .b(output_16_1), .y(output_15_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_9_1, output_9_2, output_8_1;
mixer gate_output_8_1(.a(output_9_1), .b(output_9_2), .y(output_8_1));
wire output_10_1, output_10_2, output_9_1;
mixer gate_output_9_1(.a(output_10_1), .b(output_10_2), .y(output_9_1));
wire output_11_1, output_11_2, output_10_1;
mixer gate_output_10_1(.a(output_11_1), .b(output_11_2), .y(output_10_1));
wire output_12_1, output_12_2, output_11_1;
mixer gate_output_11_1(.a(output_12_1), .b(output_12_2), .y(output_11_1));
wire output_13_1, output_13_2, output_12_1;
mixer gate_output_12_1(.a(output_13_1), .b(output_13_2), .y(output_12_1));
wire output_14_1, output_14_2, output_13_1;
mixer gate_output_13_1(.a(output_14_1), .b(output_14_2), .y(output_13_1));
wire output_15_1, output_15_2, output_14_1;
mixer gate_output_14_1(.a(output_15_1), .b(output_15_2), .y(output_14_1));
wire output_16_1, output_16_2, output_15_1;
mixer gate_output_15_1(.a(output_16_1), .b(output_16_2), .y(output_15_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_9_2, output_9_3, output_8_2;
mixer gate_output_8_2(.a(output_9_2), .b(output_9_3), .y(output_8_2));
wire output_10_2, output_10_3, output_9_2;
mixer gate_output_9_2(.a(output_10_2), .b(output_10_3), .y(output_9_2));
wire output_11_2, output_11_3, output_10_2;
mixer gate_output_10_2(.a(output_11_2), .b(output_11_3), .y(output_10_2));
wire output_12_2, output_12_3, output_11_2;
mixer gate_output_11_2(.a(output_12_2), .b(output_12_3), .y(output_11_2));
wire output_13_2, output_13_3, output_12_2;
mixer gate_output_12_2(.a(output_13_2), .b(output_13_3), .y(output_12_2));
wire output_14_2, output_14_3, output_13_2;
mixer gate_output_13_2(.a(output_14_2), .b(output_14_3), .y(output_13_2));
wire output_15_2, output_15_3, output_14_2;
mixer gate_output_14_2(.a(output_15_2), .b(output_15_3), .y(output_14_2));
wire output_16_2, output_16_3, output_15_2;
mixer gate_output_15_2(.a(output_16_2), .b(output_16_3), .y(output_15_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_9_3, output_9_4, output_8_3;
mixer gate_output_8_3(.a(output_9_3), .b(output_9_4), .y(output_8_3));
wire output_10_3, output_10_4, output_9_3;
mixer gate_output_9_3(.a(output_10_3), .b(output_10_4), .y(output_9_3));
wire output_11_3, output_11_4, output_10_3;
mixer gate_output_10_3(.a(output_11_3), .b(output_11_4), .y(output_10_3));
wire output_12_3, output_12_4, output_11_3;
mixer gate_output_11_3(.a(output_12_3), .b(output_12_4), .y(output_11_3));
wire output_13_3, output_13_4, output_12_3;
mixer gate_output_12_3(.a(output_13_3), .b(output_13_4), .y(output_12_3));
wire output_14_3, output_14_4, output_13_3;
mixer gate_output_13_3(.a(output_14_3), .b(output_14_4), .y(output_13_3));
wire output_15_3, output_15_4, output_14_3;
mixer gate_output_14_3(.a(output_15_3), .b(output_15_4), .y(output_14_3));
wire output_16_3, output_16_4, output_15_3;
mixer gate_output_15_3(.a(output_16_3), .b(output_16_4), .y(output_15_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_9_4, output_9_5, output_8_4;
mixer gate_output_8_4(.a(output_9_4), .b(output_9_5), .y(output_8_4));
wire output_10_4, output_10_5, output_9_4;
mixer gate_output_9_4(.a(output_10_4), .b(output_10_5), .y(output_9_4));
wire output_11_4, output_11_5, output_10_4;
mixer gate_output_10_4(.a(output_11_4), .b(output_11_5), .y(output_10_4));
wire output_12_4, output_12_5, output_11_4;
mixer gate_output_11_4(.a(output_12_4), .b(output_12_5), .y(output_11_4));
wire output_13_4, output_13_5, output_12_4;
mixer gate_output_12_4(.a(output_13_4), .b(output_13_5), .y(output_12_4));
wire output_14_4, output_14_5, output_13_4;
mixer gate_output_13_4(.a(output_14_4), .b(output_14_5), .y(output_13_4));
wire output_15_4, output_15_5, output_14_4;
mixer gate_output_14_4(.a(output_15_4), .b(output_15_5), .y(output_14_4));
wire output_16_4, output_16_5, output_15_4;
mixer gate_output_15_4(.a(output_16_4), .b(output_16_5), .y(output_15_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_9_5, output_9_6, output_8_5;
mixer gate_output_8_5(.a(output_9_5), .b(output_9_6), .y(output_8_5));
wire output_10_5, output_10_6, output_9_5;
mixer gate_output_9_5(.a(output_10_5), .b(output_10_6), .y(output_9_5));
wire output_11_5, output_11_6, output_10_5;
mixer gate_output_10_5(.a(output_11_5), .b(output_11_6), .y(output_10_5));
wire output_12_5, output_12_6, output_11_5;
mixer gate_output_11_5(.a(output_12_5), .b(output_12_6), .y(output_11_5));
wire output_13_5, output_13_6, output_12_5;
mixer gate_output_12_5(.a(output_13_5), .b(output_13_6), .y(output_12_5));
wire output_14_5, output_14_6, output_13_5;
mixer gate_output_13_5(.a(output_14_5), .b(output_14_6), .y(output_13_5));
wire output_15_5, output_15_6, output_14_5;
mixer gate_output_14_5(.a(output_15_5), .b(output_15_6), .y(output_14_5));
wire output_16_5, output_16_6, output_15_5;
mixer gate_output_15_5(.a(output_16_5), .b(output_16_6), .y(output_15_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_9_6, output_9_7, output_8_6;
mixer gate_output_8_6(.a(output_9_6), .b(output_9_7), .y(output_8_6));
wire output_10_6, output_10_7, output_9_6;
mixer gate_output_9_6(.a(output_10_6), .b(output_10_7), .y(output_9_6));
wire output_11_6, output_11_7, output_10_6;
mixer gate_output_10_6(.a(output_11_6), .b(output_11_7), .y(output_10_6));
wire output_12_6, output_12_7, output_11_6;
mixer gate_output_11_6(.a(output_12_6), .b(output_12_7), .y(output_11_6));
wire output_13_6, output_13_7, output_12_6;
mixer gate_output_12_6(.a(output_13_6), .b(output_13_7), .y(output_12_6));
wire output_14_6, output_14_7, output_13_6;
mixer gate_output_13_6(.a(output_14_6), .b(output_14_7), .y(output_13_6));
wire output_15_6, output_15_7, output_14_6;
mixer gate_output_14_6(.a(output_15_6), .b(output_15_7), .y(output_14_6));
wire output_16_6, output_16_7, output_15_6;
mixer gate_output_15_6(.a(output_16_6), .b(output_16_7), .y(output_15_6));
wire output_1_7, output_1_8, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_8), .y(output_0_7));
wire output_2_7, output_2_8, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_8), .y(output_1_7));
wire output_3_7, output_3_8, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_8), .y(output_2_7));
wire output_4_7, output_4_8, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_8), .y(output_3_7));
wire output_5_7, output_5_8, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_8), .y(output_4_7));
wire output_6_7, output_6_8, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_8), .y(output_5_7));
wire output_7_7, output_7_8, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_8), .y(output_6_7));
wire output_8_7, output_8_8, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_8), .y(output_7_7));
wire output_9_7, output_9_8, output_8_7;
mixer gate_output_8_7(.a(output_9_7), .b(output_9_8), .y(output_8_7));
wire output_10_7, output_10_8, output_9_7;
mixer gate_output_9_7(.a(output_10_7), .b(output_10_8), .y(output_9_7));
wire output_11_7, output_11_8, output_10_7;
mixer gate_output_10_7(.a(output_11_7), .b(output_11_8), .y(output_10_7));
wire output_12_7, output_12_8, output_11_7;
mixer gate_output_11_7(.a(output_12_7), .b(output_12_8), .y(output_11_7));
wire output_13_7, output_13_8, output_12_7;
mixer gate_output_12_7(.a(output_13_7), .b(output_13_8), .y(output_12_7));
wire output_14_7, output_14_8, output_13_7;
mixer gate_output_13_7(.a(output_14_7), .b(output_14_8), .y(output_13_7));
wire output_15_7, output_15_8, output_14_7;
mixer gate_output_14_7(.a(output_15_7), .b(output_15_8), .y(output_14_7));
wire output_16_7, output_16_8, output_15_7;
mixer gate_output_15_7(.a(output_16_7), .b(output_16_8), .y(output_15_7));
assign output_0 = output_0_0;
wire output_0_8;
assign output_0_8 = input_0;
assign output_1 = output_1_0;
wire output_1_8;
assign output_1_8 = input_1;
assign output_2 = output_2_0;
wire output_2_8;
assign output_2_8 = input_2;
assign output_3 = output_3_0;
wire output_3_8;
assign output_3_8 = input_3;
assign output_4 = output_4_0;
wire output_4_8;
assign output_4_8 = input_4;
assign output_5 = output_5_0;
wire output_5_8;
assign output_5_8 = input_5;
assign output_6 = output_6_0;
wire output_6_8;
assign output_6_8 = input_6;
assign output_7 = output_7_0;
wire output_7_8;
assign output_7_8 = input_7;
assign output_8 = output_8_0;
wire output_8_8;
assign output_8_8 = input_8;
assign output_9 = output_9_0;
wire output_9_8;
assign output_9_8 = input_9;
assign output_10 = output_10_0;
wire output_10_8;
assign output_10_8 = input_10;
assign output_11 = output_11_0;
wire output_11_8;
assign output_11_8 = input_11;
assign output_12 = output_12_0;
wire output_12_8;
assign output_12_8 = input_12;
assign output_13 = output_13_0;
wire output_13_8;
assign output_13_8 = input_13;
assign output_14 = output_14_0;
wire output_14_8;
assign output_14_8 = input_14;
assign output_15 = output_15_0;
wire output_15_8;
assign output_15_8 = input_15;
endmodule
