module binary_tree_1_5 (
output out_0,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
wire t0_0;
assign out_0 = t0_0;
assign input_0 = t0_000000;
assign input_1 = t0_000001;
assign input_2 = t0_000010;
assign input_3 = t0_000011;
assign input_4 = t0_000100;
assign input_5 = t0_000101;
assign input_6 = t0_000110;
assign input_7 = t0_000111;
assign input_8 = t0_001000;
assign input_9 = t0_001001;
assign input_10 = t0_001010;
assign input_11 = t0_001011;
assign input_12 = t0_001100;
assign input_13 = t0_001101;
assign input_14 = t0_001110;
assign input_15 = t0_001111;
assign input_16 = t0_010000;
assign input_17 = t0_010001;
assign input_18 = t0_010010;
assign input_19 = t0_010011;
assign input_20 = t0_010100;
assign input_21 = t0_010101;
assign input_22 = t0_010110;
assign input_23 = t0_010111;
assign input_24 = t0_011000;
assign input_25 = t0_011001;
assign input_26 = t0_011010;
assign input_27 = t0_011011;
assign input_28 = t0_011100;
assign input_29 = t0_011101;
assign input_30 = t0_011110;
assign input_31 = t0_011111;
endmodule
