module binary_tree_8_8 (
output out_0,output out_1,output out_2,output out_3,output out_4,output out_5,output out_6,output out_7,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15,input input_16,input input_17,input input_18,input input_19,input input_20,input input_21,input input_22,input input_23,input input_24,input input_25,input input_26,input input_27,input input_28,input input_29,input input_30,input input_31,input input_32,input input_33,input input_34,input input_35,input input_36,input input_37,input input_38,input input_39,input input_40,input input_41,input input_42,input input_43,input input_44,input input_45,input input_46,input input_47,input input_48,input input_49,input input_50,input input_51,input input_52,input input_53,input input_54,input input_55,input input_56,input input_57,input input_58,input input_59,input input_60,input input_61,input input_62,input input_63,input input_64,input input_65,input input_66,input input_67,input input_68,input input_69,input input_70,input input_71,input input_72,input input_73,input input_74,input input_75,input input_76,input input_77,input input_78,input input_79,input input_80,input input_81,input input_82,input input_83,input input_84,input input_85,input input_86,input input_87,input input_88,input input_89,input input_90,input input_91,input input_92,input input_93,input input_94,input input_95,input input_96,input input_97,input input_98,input input_99,input input_100,input input_101,input input_102,input input_103,input input_104,input input_105,input input_106,input input_107,input input_108,input input_109,input input_110,input input_111,input input_112,input input_113,input input_114,input input_115,input input_116,input input_117,input input_118,input input_119,input input_120,input input_121,input input_122,input input_123,input input_124,input input_125,input input_126,input input_127,input input_128,input input_129,input input_130,input input_131,input input_132,input input_133,input input_134,input input_135,input input_136,input input_137,input input_138,input input_139,input input_140,input input_141,input input_142,input input_143,input input_144,input input_145,input input_146,input input_147,input input_148,input input_149,input input_150,input input_151,input input_152,input input_153,input input_154,input input_155,input input_156,input input_157,input input_158,input input_159,input input_160,input input_161,input input_162,input input_163,input input_164,input input_165,input input_166,input input_167,input input_168,input input_169,input input_170,input input_171,input input_172,input input_173,input input_174,input input_175,input input_176,input input_177,input input_178,input input_179,input input_180,input input_181,input input_182,input input_183,input input_184,input input_185,input input_186,input input_187,input input_188,input input_189,input input_190,input input_191,input input_192,input input_193,input input_194,input input_195,input input_196,input input_197,input input_198,input input_199,input input_200,input input_201,input input_202,input input_203,input input_204,input input_205,input input_206,input input_207,input input_208,input input_209,input input_210,input input_211,input input_212,input input_213,input input_214,input input_215,input input_216,input input_217,input input_218,input input_219,input input_220,input input_221,input input_222,input input_223,input input_224,input input_225,input input_226,input input_227,input input_228,input input_229,input input_230,input input_231,input input_232,input input_233,input input_234,input input_235,input input_236,input input_237,input input_238,input input_239,input input_240,input input_241,input input_242,input input_243,input input_244,input input_245,input input_246,input input_247,input input_248,input input_249,input input_250,input input_251,input input_252,input input_253,input input_254,input input_255,input input_256,input input_257,input input_258,input input_259,input input_260,input input_261,input input_262,input input_263,input input_264,input input_265,input input_266,input input_267,input input_268,input input_269,input input_270,input input_271,input input_272,input input_273,input input_274,input input_275,input input_276,input input_277,input input_278,input input_279,input input_280,input input_281,input input_282,input input_283,input input_284,input input_285,input input_286,input input_287,input input_288,input input_289,input input_290,input input_291,input input_292,input input_293,input input_294,input input_295,input input_296,input input_297,input input_298,input input_299,input input_300,input input_301,input input_302,input input_303,input input_304,input input_305,input input_306,input input_307,input input_308,input input_309,input input_310,input input_311,input input_312,input input_313,input input_314,input input_315,input input_316,input input_317,input input_318,input input_319,input input_320,input input_321,input input_322,input input_323,input input_324,input input_325,input input_326,input input_327,input input_328,input input_329,input input_330,input input_331,input input_332,input input_333,input input_334,input input_335,input input_336,input input_337,input input_338,input input_339,input input_340,input input_341,input input_342,input input_343,input input_344,input input_345,input input_346,input input_347,input input_348,input input_349,input input_350,input input_351,input input_352,input input_353,input input_354,input input_355,input input_356,input input_357,input input_358,input input_359,input input_360,input input_361,input input_362,input input_363,input input_364,input input_365,input input_366,input input_367,input input_368,input input_369,input input_370,input input_371,input input_372,input input_373,input input_374,input input_375,input input_376,input input_377,input input_378,input input_379,input input_380,input input_381,input input_382,input input_383,input input_384,input input_385,input input_386,input input_387,input input_388,input input_389,input input_390,input input_391,input input_392,input input_393,input input_394,input input_395,input input_396,input input_397,input input_398,input input_399,input input_400,input input_401,input input_402,input input_403,input input_404,input input_405,input input_406,input input_407,input input_408,input input_409,input input_410,input input_411,input input_412,input input_413,input input_414,input input_415,input input_416,input input_417,input input_418,input input_419,input input_420,input input_421,input input_422,input input_423,input input_424,input input_425,input input_426,input input_427,input input_428,input input_429,input input_430,input input_431,input input_432,input input_433,input input_434,input input_435,input input_436,input input_437,input input_438,input input_439,input input_440,input input_441,input input_442,input input_443,input input_444,input input_445,input input_446,input input_447,input input_448,input input_449,input input_450,input input_451,input input_452,input input_453,input input_454,input input_455,input input_456,input input_457,input input_458,input input_459,input input_460,input input_461,input input_462,input input_463,input input_464,input input_465,input input_466,input input_467,input input_468,input input_469,input input_470,input input_471,input input_472,input input_473,input input_474,input input_475,input input_476,input input_477,input input_478,input input_479,input input_480,input input_481,input input_482,input input_483,input input_484,input input_485,input input_486,input input_487,input input_488,input input_489,input input_490,input input_491,input input_492,input input_493,input input_494,input input_495,input input_496,input input_497,input input_498,input input_499,input input_500,input input_501,input input_502,input input_503,input input_504,input input_505,input input_506,input input_507,input input_508,input input_509,input input_510,input input_511,input input_512,input input_513,input input_514,input input_515,input input_516,input input_517,input input_518,input input_519,input input_520,input input_521,input input_522,input input_523,input input_524,input input_525,input input_526,input input_527,input input_528,input input_529,input input_530,input input_531,input input_532,input input_533,input input_534,input input_535,input input_536,input input_537,input input_538,input input_539,input input_540,input input_541,input input_542,input input_543,input input_544,input input_545,input input_546,input input_547,input input_548,input input_549,input input_550,input input_551,input input_552,input input_553,input input_554,input input_555,input input_556,input input_557,input input_558,input input_559,input input_560,input input_561,input input_562,input input_563,input input_564,input input_565,input input_566,input input_567,input input_568,input input_569,input input_570,input input_571,input input_572,input input_573,input input_574,input input_575,input input_576,input input_577,input input_578,input input_579,input input_580,input input_581,input input_582,input input_583,input input_584,input input_585,input input_586,input input_587,input input_588,input input_589,input input_590,input input_591,input input_592,input input_593,input input_594,input input_595,input input_596,input input_597,input input_598,input input_599,input input_600,input input_601,input input_602,input input_603,input input_604,input input_605,input input_606,input input_607,input input_608,input input_609,input input_610,input input_611,input input_612,input input_613,input input_614,input input_615,input input_616,input input_617,input input_618,input input_619,input input_620,input input_621,input input_622,input input_623,input input_624,input input_625,input input_626,input input_627,input input_628,input input_629,input input_630,input input_631,input input_632,input input_633,input input_634,input input_635,input input_636,input input_637,input input_638,input input_639,input input_640,input input_641,input input_642,input input_643,input input_644,input input_645,input input_646,input input_647,input input_648,input input_649,input input_650,input input_651,input input_652,input input_653,input input_654,input input_655,input input_656,input input_657,input input_658,input input_659,input input_660,input input_661,input input_662,input input_663,input input_664,input input_665,input input_666,input input_667,input input_668,input input_669,input input_670,input input_671,input input_672,input input_673,input input_674,input input_675,input input_676,input input_677,input input_678,input input_679,input input_680,input input_681,input input_682,input input_683,input input_684,input input_685,input input_686,input input_687,input input_688,input input_689,input input_690,input input_691,input input_692,input input_693,input input_694,input input_695,input input_696,input input_697,input input_698,input input_699,input input_700,input input_701,input input_702,input input_703,input input_704,input input_705,input input_706,input input_707,input input_708,input input_709,input input_710,input input_711,input input_712,input input_713,input input_714,input input_715,input input_716,input input_717,input input_718,input input_719,input input_720,input input_721,input input_722,input input_723,input input_724,input input_725,input input_726,input input_727,input input_728,input input_729,input input_730,input input_731,input input_732,input input_733,input input_734,input input_735,input input_736,input input_737,input input_738,input input_739,input input_740,input input_741,input input_742,input input_743,input input_744,input input_745,input input_746,input input_747,input input_748,input input_749,input input_750,input input_751,input input_752,input input_753,input input_754,input input_755,input input_756,input input_757,input input_758,input input_759,input input_760,input input_761,input input_762,input input_763,input input_764,input input_765,input input_766,input input_767,input input_768,input input_769,input input_770,input input_771,input input_772,input input_773,input input_774,input input_775,input input_776,input input_777,input input_778,input input_779,input input_780,input input_781,input input_782,input input_783,input input_784,input input_785,input input_786,input input_787,input input_788,input input_789,input input_790,input input_791,input input_792,input input_793,input input_794,input input_795,input input_796,input input_797,input input_798,input input_799,input input_800,input input_801,input input_802,input input_803,input input_804,input input_805,input input_806,input input_807,input input_808,input input_809,input input_810,input input_811,input input_812,input input_813,input input_814,input input_815,input input_816,input input_817,input input_818,input input_819,input input_820,input input_821,input input_822,input input_823,input input_824,input input_825,input input_826,input input_827,input input_828,input input_829,input input_830,input input_831,input input_832,input input_833,input input_834,input input_835,input input_836,input input_837,input input_838,input input_839,input input_840,input input_841,input input_842,input input_843,input input_844,input input_845,input input_846,input input_847,input input_848,input input_849,input input_850,input input_851,input input_852,input input_853,input input_854,input input_855,input input_856,input input_857,input input_858,input input_859,input input_860,input input_861,input input_862,input input_863,input input_864,input input_865,input input_866,input input_867,input input_868,input input_869,input input_870,input input_871,input input_872,input input_873,input input_874,input input_875,input input_876,input input_877,input input_878,input input_879,input input_880,input input_881,input input_882,input input_883,input input_884,input input_885,input input_886,input input_887,input input_888,input input_889,input input_890,input input_891,input input_892,input input_893,input input_894,input input_895,input input_896,input input_897,input input_898,input input_899,input input_900,input input_901,input input_902,input input_903,input input_904,input input_905,input input_906,input input_907,input input_908,input input_909,input input_910,input input_911,input input_912,input input_913,input input_914,input input_915,input input_916,input input_917,input input_918,input input_919,input input_920,input input_921,input input_922,input input_923,input input_924,input input_925,input input_926,input input_927,input input_928,input input_929,input input_930,input input_931,input input_932,input input_933,input input_934,input input_935,input input_936,input input_937,input input_938,input input_939,input input_940,input input_941,input input_942,input input_943,input input_944,input input_945,input input_946,input input_947,input input_948,input input_949,input input_950,input input_951,input input_952,input input_953,input input_954,input input_955,input input_956,input input_957,input input_958,input input_959,input input_960,input input_961,input input_962,input input_963,input input_964,input input_965,input input_966,input input_967,input input_968,input input_969,input input_970,input input_971,input input_972,input input_973,input input_974,input input_975,input input_976,input input_977,input input_978,input input_979,input input_980,input input_981,input input_982,input input_983,input input_984,input input_985,input input_986,input input_987,input input_988,input input_989,input input_990,input input_991,input input_992,input input_993,input input_994,input input_995,input input_996,input input_997,input input_998,input input_999,input input_1000,input input_1001,input input_1002,input input_1003,input input_1004,input input_1005,input input_1006,input input_1007,input input_1008,input input_1009,input input_1010,input input_1011,input input_1012,input input_1013,input input_1014,input input_1015,input input_1016,input input_1017,input input_1018,input input_1019,input input_1020,input input_1021,input input_1022,input input_1023,input input_1024,input input_1025,input input_1026,input input_1027,input input_1028,input input_1029,input input_1030,input input_1031,input input_1032,input input_1033,input input_1034,input input_1035,input input_1036,input input_1037,input input_1038,input input_1039,input input_1040,input input_1041,input input_1042,input input_1043,input input_1044,input input_1045,input input_1046,input input_1047,input input_1048,input input_1049,input input_1050,input input_1051,input input_1052,input input_1053,input input_1054,input input_1055,input input_1056,input input_1057,input input_1058,input input_1059,input input_1060,input input_1061,input input_1062,input input_1063,input input_1064,input input_1065,input input_1066,input input_1067,input input_1068,input input_1069,input input_1070,input input_1071,input input_1072,input input_1073,input input_1074,input input_1075,input input_1076,input input_1077,input input_1078,input input_1079,input input_1080,input input_1081,input input_1082,input input_1083,input input_1084,input input_1085,input input_1086,input input_1087,input input_1088,input input_1089,input input_1090,input input_1091,input input_1092,input input_1093,input input_1094,input input_1095,input input_1096,input input_1097,input input_1098,input input_1099,input input_1100,input input_1101,input input_1102,input input_1103,input input_1104,input input_1105,input input_1106,input input_1107,input input_1108,input input_1109,input input_1110,input input_1111,input input_1112,input input_1113,input input_1114,input input_1115,input input_1116,input input_1117,input input_1118,input input_1119,input input_1120,input input_1121,input input_1122,input input_1123,input input_1124,input input_1125,input input_1126,input input_1127,input input_1128,input input_1129,input input_1130,input input_1131,input input_1132,input input_1133,input input_1134,input input_1135,input input_1136,input input_1137,input input_1138,input input_1139,input input_1140,input input_1141,input input_1142,input input_1143,input input_1144,input input_1145,input input_1146,input input_1147,input input_1148,input input_1149,input input_1150,input input_1151,input input_1152,input input_1153,input input_1154,input input_1155,input input_1156,input input_1157,input input_1158,input input_1159,input input_1160,input input_1161,input input_1162,input input_1163,input input_1164,input input_1165,input input_1166,input input_1167,input input_1168,input input_1169,input input_1170,input input_1171,input input_1172,input input_1173,input input_1174,input input_1175,input input_1176,input input_1177,input input_1178,input input_1179,input input_1180,input input_1181,input input_1182,input input_1183,input input_1184,input input_1185,input input_1186,input input_1187,input input_1188,input input_1189,input input_1190,input input_1191,input input_1192,input input_1193,input input_1194,input input_1195,input input_1196,input input_1197,input input_1198,input input_1199,input input_1200,input input_1201,input input_1202,input input_1203,input input_1204,input input_1205,input input_1206,input input_1207,input input_1208,input input_1209,input input_1210,input input_1211,input input_1212,input input_1213,input input_1214,input input_1215,input input_1216,input input_1217,input input_1218,input input_1219,input input_1220,input input_1221,input input_1222,input input_1223,input input_1224,input input_1225,input input_1226,input input_1227,input input_1228,input input_1229,input input_1230,input input_1231,input input_1232,input input_1233,input input_1234,input input_1235,input input_1236,input input_1237,input input_1238,input input_1239,input input_1240,input input_1241,input input_1242,input input_1243,input input_1244,input input_1245,input input_1246,input input_1247,input input_1248,input input_1249,input input_1250,input input_1251,input input_1252,input input_1253,input input_1254,input input_1255,input input_1256,input input_1257,input input_1258,input input_1259,input input_1260,input input_1261,input input_1262,input input_1263,input input_1264,input input_1265,input input_1266,input input_1267,input input_1268,input input_1269,input input_1270,input input_1271,input input_1272,input input_1273,input input_1274,input input_1275,input input_1276,input input_1277,input input_1278,input input_1279,input input_1280,input input_1281,input input_1282,input input_1283,input input_1284,input input_1285,input input_1286,input input_1287,input input_1288,input input_1289,input input_1290,input input_1291,input input_1292,input input_1293,input input_1294,input input_1295,input input_1296,input input_1297,input input_1298,input input_1299,input input_1300,input input_1301,input input_1302,input input_1303,input input_1304,input input_1305,input input_1306,input input_1307,input input_1308,input input_1309,input input_1310,input input_1311,input input_1312,input input_1313,input input_1314,input input_1315,input input_1316,input input_1317,input input_1318,input input_1319,input input_1320,input input_1321,input input_1322,input input_1323,input input_1324,input input_1325,input input_1326,input input_1327,input input_1328,input input_1329,input input_1330,input input_1331,input input_1332,input input_1333,input input_1334,input input_1335,input input_1336,input input_1337,input input_1338,input input_1339,input input_1340,input input_1341,input input_1342,input input_1343,input input_1344,input input_1345,input input_1346,input input_1347,input input_1348,input input_1349,input input_1350,input input_1351,input input_1352,input input_1353,input input_1354,input input_1355,input input_1356,input input_1357,input input_1358,input input_1359,input input_1360,input input_1361,input input_1362,input input_1363,input input_1364,input input_1365,input input_1366,input input_1367,input input_1368,input input_1369,input input_1370,input input_1371,input input_1372,input input_1373,input input_1374,input input_1375,input input_1376,input input_1377,input input_1378,input input_1379,input input_1380,input input_1381,input input_1382,input input_1383,input input_1384,input input_1385,input input_1386,input input_1387,input input_1388,input input_1389,input input_1390,input input_1391,input input_1392,input input_1393,input input_1394,input input_1395,input input_1396,input input_1397,input input_1398,input input_1399,input input_1400,input input_1401,input input_1402,input input_1403,input input_1404,input input_1405,input input_1406,input input_1407,input input_1408,input input_1409,input input_1410,input input_1411,input input_1412,input input_1413,input input_1414,input input_1415,input input_1416,input input_1417,input input_1418,input input_1419,input input_1420,input input_1421,input input_1422,input input_1423,input input_1424,input input_1425,input input_1426,input input_1427,input input_1428,input input_1429,input input_1430,input input_1431,input input_1432,input input_1433,input input_1434,input input_1435,input input_1436,input input_1437,input input_1438,input input_1439,input input_1440,input input_1441,input input_1442,input input_1443,input input_1444,input input_1445,input input_1446,input input_1447,input input_1448,input input_1449,input input_1450,input input_1451,input input_1452,input input_1453,input input_1454,input input_1455,input input_1456,input input_1457,input input_1458,input input_1459,input input_1460,input input_1461,input input_1462,input input_1463,input input_1464,input input_1465,input input_1466,input input_1467,input input_1468,input input_1469,input input_1470,input input_1471,input input_1472,input input_1473,input input_1474,input input_1475,input input_1476,input input_1477,input input_1478,input input_1479,input input_1480,input input_1481,input input_1482,input input_1483,input input_1484,input input_1485,input input_1486,input input_1487,input input_1488,input input_1489,input input_1490,input input_1491,input input_1492,input input_1493,input input_1494,input input_1495,input input_1496,input input_1497,input input_1498,input input_1499,input input_1500,input input_1501,input input_1502,input input_1503,input input_1504,input input_1505,input input_1506,input input_1507,input input_1508,input input_1509,input input_1510,input input_1511,input input_1512,input input_1513,input input_1514,input input_1515,input input_1516,input input_1517,input input_1518,input input_1519,input input_1520,input input_1521,input input_1522,input input_1523,input input_1524,input input_1525,input input_1526,input input_1527,input input_1528,input input_1529,input input_1530,input input_1531,input input_1532,input input_1533,input input_1534,input input_1535,input input_1536,input input_1537,input input_1538,input input_1539,input input_1540,input input_1541,input input_1542,input input_1543,input input_1544,input input_1545,input input_1546,input input_1547,input input_1548,input input_1549,input input_1550,input input_1551,input input_1552,input input_1553,input input_1554,input input_1555,input input_1556,input input_1557,input input_1558,input input_1559,input input_1560,input input_1561,input input_1562,input input_1563,input input_1564,input input_1565,input input_1566,input input_1567,input input_1568,input input_1569,input input_1570,input input_1571,input input_1572,input input_1573,input input_1574,input input_1575,input input_1576,input input_1577,input input_1578,input input_1579,input input_1580,input input_1581,input input_1582,input input_1583,input input_1584,input input_1585,input input_1586,input input_1587,input input_1588,input input_1589,input input_1590,input input_1591,input input_1592,input input_1593,input input_1594,input input_1595,input input_1596,input input_1597,input input_1598,input input_1599,input input_1600,input input_1601,input input_1602,input input_1603,input input_1604,input input_1605,input input_1606,input input_1607,input input_1608,input input_1609,input input_1610,input input_1611,input input_1612,input input_1613,input input_1614,input input_1615,input input_1616,input input_1617,input input_1618,input input_1619,input input_1620,input input_1621,input input_1622,input input_1623,input input_1624,input input_1625,input input_1626,input input_1627,input input_1628,input input_1629,input input_1630,input input_1631,input input_1632,input input_1633,input input_1634,input input_1635,input input_1636,input input_1637,input input_1638,input input_1639,input input_1640,input input_1641,input input_1642,input input_1643,input input_1644,input input_1645,input input_1646,input input_1647,input input_1648,input input_1649,input input_1650,input input_1651,input input_1652,input input_1653,input input_1654,input input_1655,input input_1656,input input_1657,input input_1658,input input_1659,input input_1660,input input_1661,input input_1662,input input_1663,input input_1664,input input_1665,input input_1666,input input_1667,input input_1668,input input_1669,input input_1670,input input_1671,input input_1672,input input_1673,input input_1674,input input_1675,input input_1676,input input_1677,input input_1678,input input_1679,input input_1680,input input_1681,input input_1682,input input_1683,input input_1684,input input_1685,input input_1686,input input_1687,input input_1688,input input_1689,input input_1690,input input_1691,input input_1692,input input_1693,input input_1694,input input_1695,input input_1696,input input_1697,input input_1698,input input_1699,input input_1700,input input_1701,input input_1702,input input_1703,input input_1704,input input_1705,input input_1706,input input_1707,input input_1708,input input_1709,input input_1710,input input_1711,input input_1712,input input_1713,input input_1714,input input_1715,input input_1716,input input_1717,input input_1718,input input_1719,input input_1720,input input_1721,input input_1722,input input_1723,input input_1724,input input_1725,input input_1726,input input_1727,input input_1728,input input_1729,input input_1730,input input_1731,input input_1732,input input_1733,input input_1734,input input_1735,input input_1736,input input_1737,input input_1738,input input_1739,input input_1740,input input_1741,input input_1742,input input_1743,input input_1744,input input_1745,input input_1746,input input_1747,input input_1748,input input_1749,input input_1750,input input_1751,input input_1752,input input_1753,input input_1754,input input_1755,input input_1756,input input_1757,input input_1758,input input_1759,input input_1760,input input_1761,input input_1762,input input_1763,input input_1764,input input_1765,input input_1766,input input_1767,input input_1768,input input_1769,input input_1770,input input_1771,input input_1772,input input_1773,input input_1774,input input_1775,input input_1776,input input_1777,input input_1778,input input_1779,input input_1780,input input_1781,input input_1782,input input_1783,input input_1784,input input_1785,input input_1786,input input_1787,input input_1788,input input_1789,input input_1790,input input_1791,input input_1792,input input_1793,input input_1794,input input_1795,input input_1796,input input_1797,input input_1798,input input_1799,input input_1800,input input_1801,input input_1802,input input_1803,input input_1804,input input_1805,input input_1806,input input_1807,input input_1808,input input_1809,input input_1810,input input_1811,input input_1812,input input_1813,input input_1814,input input_1815,input input_1816,input input_1817,input input_1818,input input_1819,input input_1820,input input_1821,input input_1822,input input_1823,input input_1824,input input_1825,input input_1826,input input_1827,input input_1828,input input_1829,input input_1830,input input_1831,input input_1832,input input_1833,input input_1834,input input_1835,input input_1836,input input_1837,input input_1838,input input_1839,input input_1840,input input_1841,input input_1842,input input_1843,input input_1844,input input_1845,input input_1846,input input_1847,input input_1848,input input_1849,input input_1850,input input_1851,input input_1852,input input_1853,input input_1854,input input_1855,input input_1856,input input_1857,input input_1858,input input_1859,input input_1860,input input_1861,input input_1862,input input_1863,input input_1864,input input_1865,input input_1866,input input_1867,input input_1868,input input_1869,input input_1870,input input_1871,input input_1872,input input_1873,input input_1874,input input_1875,input input_1876,input input_1877,input input_1878,input input_1879,input input_1880,input input_1881,input input_1882,input input_1883,input input_1884,input input_1885,input input_1886,input input_1887,input input_1888,input input_1889,input input_1890,input input_1891,input input_1892,input input_1893,input input_1894,input input_1895,input input_1896,input input_1897,input input_1898,input input_1899,input input_1900,input input_1901,input input_1902,input input_1903,input input_1904,input input_1905,input input_1906,input input_1907,input input_1908,input input_1909,input input_1910,input input_1911,input input_1912,input input_1913,input input_1914,input input_1915,input input_1916,input input_1917,input input_1918,input input_1919,input input_1920,input input_1921,input input_1922,input input_1923,input input_1924,input input_1925,input input_1926,input input_1927,input input_1928,input input_1929,input input_1930,input input_1931,input input_1932,input input_1933,input input_1934,input input_1935,input input_1936,input input_1937,input input_1938,input input_1939,input input_1940,input input_1941,input input_1942,input input_1943,input input_1944,input input_1945,input input_1946,input input_1947,input input_1948,input input_1949,input input_1950,input input_1951,input input_1952,input input_1953,input input_1954,input input_1955,input input_1956,input input_1957,input input_1958,input input_1959,input input_1960,input input_1961,input input_1962,input input_1963,input input_1964,input input_1965,input input_1966,input input_1967,input input_1968,input input_1969,input input_1970,input input_1971,input input_1972,input input_1973,input input_1974,input input_1975,input input_1976,input input_1977,input input_1978,input input_1979,input input_1980,input input_1981,input input_1982,input input_1983,input input_1984,input input_1985,input input_1986,input input_1987,input input_1988,input input_1989,input input_1990,input input_1991,input input_1992,input input_1993,input input_1994,input input_1995,input input_1996,input input_1997,input input_1998,input input_1999,input input_2000,input input_2001,input input_2002,input input_2003,input input_2004,input input_2005,input input_2006,input input_2007,input input_2008,input input_2009,input input_2010,input input_2011,input input_2012,input input_2013,input input_2014,input input_2015,input input_2016,input input_2017,input input_2018,input input_2019,input input_2020,input input_2021,input input_2022,input input_2023,input input_2024,input input_2025,input input_2026,input input_2027,input input_2028,input input_2029,input input_2030,input input_2031,input input_2032,input input_2033,input input_2034,input input_2035,input input_2036,input input_2037,input input_2038,input input_2039,input input_2040,input input_2041,input input_2042,input input_2043,input input_2044,input input_2045,input input_2046,input input_2047
);
mixer mix_t0_0 (.a(t0_00), .b(t0_01), .y(t0_0));
wire t0_00, t0_01;
mixer mix_t0_00 (.a(t0_000), .b(t0_001), .y(t0_00));
wire t0_000, t0_001;
mixer mix_t0_000 (.a(t0_0000), .b(t0_0001), .y(t0_000));
wire t0_0000, t0_0001;
mixer mix_t0_0000 (.a(t0_00000), .b(t0_00001), .y(t0_0000));
wire t0_00000, t0_00001;
mixer mix_t0_00000 (.a(t0_000000), .b(t0_000001), .y(t0_00000));
wire t0_000000, t0_000001;
mixer mix_t0_000000 (.a(t0_0000000), .b(t0_0000001), .y(t0_000000));
wire t0_0000000, t0_0000001;
mixer mix_t0_0000000 (.a(t0_00000000), .b(t0_00000001), .y(t0_0000000));
wire t0_00000000, t0_00000001;
mixer mix_t0_00000000 (.a(t0_000000000), .b(t0_000000001), .y(t0_00000000));
wire t0_000000000, t0_000000001;
mixer mix_t0_00000001 (.a(t0_000000010), .b(t0_000000011), .y(t0_00000001));
wire t0_000000010, t0_000000011;
mixer mix_t0_0000001 (.a(t0_00000010), .b(t0_00000011), .y(t0_0000001));
wire t0_00000010, t0_00000011;
mixer mix_t0_00000010 (.a(t0_000000100), .b(t0_000000101), .y(t0_00000010));
wire t0_000000100, t0_000000101;
mixer mix_t0_00000011 (.a(t0_000000110), .b(t0_000000111), .y(t0_00000011));
wire t0_000000110, t0_000000111;
mixer mix_t0_000001 (.a(t0_0000010), .b(t0_0000011), .y(t0_000001));
wire t0_0000010, t0_0000011;
mixer mix_t0_0000010 (.a(t0_00000100), .b(t0_00000101), .y(t0_0000010));
wire t0_00000100, t0_00000101;
mixer mix_t0_00000100 (.a(t0_000001000), .b(t0_000001001), .y(t0_00000100));
wire t0_000001000, t0_000001001;
mixer mix_t0_00000101 (.a(t0_000001010), .b(t0_000001011), .y(t0_00000101));
wire t0_000001010, t0_000001011;
mixer mix_t0_0000011 (.a(t0_00000110), .b(t0_00000111), .y(t0_0000011));
wire t0_00000110, t0_00000111;
mixer mix_t0_00000110 (.a(t0_000001100), .b(t0_000001101), .y(t0_00000110));
wire t0_000001100, t0_000001101;
mixer mix_t0_00000111 (.a(t0_000001110), .b(t0_000001111), .y(t0_00000111));
wire t0_000001110, t0_000001111;
mixer mix_t0_00001 (.a(t0_000010), .b(t0_000011), .y(t0_00001));
wire t0_000010, t0_000011;
mixer mix_t0_000010 (.a(t0_0000100), .b(t0_0000101), .y(t0_000010));
wire t0_0000100, t0_0000101;
mixer mix_t0_0000100 (.a(t0_00001000), .b(t0_00001001), .y(t0_0000100));
wire t0_00001000, t0_00001001;
mixer mix_t0_00001000 (.a(t0_000010000), .b(t0_000010001), .y(t0_00001000));
wire t0_000010000, t0_000010001;
mixer mix_t0_00001001 (.a(t0_000010010), .b(t0_000010011), .y(t0_00001001));
wire t0_000010010, t0_000010011;
mixer mix_t0_0000101 (.a(t0_00001010), .b(t0_00001011), .y(t0_0000101));
wire t0_00001010, t0_00001011;
mixer mix_t0_00001010 (.a(t0_000010100), .b(t0_000010101), .y(t0_00001010));
wire t0_000010100, t0_000010101;
mixer mix_t0_00001011 (.a(t0_000010110), .b(t0_000010111), .y(t0_00001011));
wire t0_000010110, t0_000010111;
mixer mix_t0_000011 (.a(t0_0000110), .b(t0_0000111), .y(t0_000011));
wire t0_0000110, t0_0000111;
mixer mix_t0_0000110 (.a(t0_00001100), .b(t0_00001101), .y(t0_0000110));
wire t0_00001100, t0_00001101;
mixer mix_t0_00001100 (.a(t0_000011000), .b(t0_000011001), .y(t0_00001100));
wire t0_000011000, t0_000011001;
mixer mix_t0_00001101 (.a(t0_000011010), .b(t0_000011011), .y(t0_00001101));
wire t0_000011010, t0_000011011;
mixer mix_t0_0000111 (.a(t0_00001110), .b(t0_00001111), .y(t0_0000111));
wire t0_00001110, t0_00001111;
mixer mix_t0_00001110 (.a(t0_000011100), .b(t0_000011101), .y(t0_00001110));
wire t0_000011100, t0_000011101;
mixer mix_t0_00001111 (.a(t0_000011110), .b(t0_000011111), .y(t0_00001111));
wire t0_000011110, t0_000011111;
mixer mix_t0_0001 (.a(t0_00010), .b(t0_00011), .y(t0_0001));
wire t0_00010, t0_00011;
mixer mix_t0_00010 (.a(t0_000100), .b(t0_000101), .y(t0_00010));
wire t0_000100, t0_000101;
mixer mix_t0_000100 (.a(t0_0001000), .b(t0_0001001), .y(t0_000100));
wire t0_0001000, t0_0001001;
mixer mix_t0_0001000 (.a(t0_00010000), .b(t0_00010001), .y(t0_0001000));
wire t0_00010000, t0_00010001;
mixer mix_t0_00010000 (.a(t0_000100000), .b(t0_000100001), .y(t0_00010000));
wire t0_000100000, t0_000100001;
mixer mix_t0_00010001 (.a(t0_000100010), .b(t0_000100011), .y(t0_00010001));
wire t0_000100010, t0_000100011;
mixer mix_t0_0001001 (.a(t0_00010010), .b(t0_00010011), .y(t0_0001001));
wire t0_00010010, t0_00010011;
mixer mix_t0_00010010 (.a(t0_000100100), .b(t0_000100101), .y(t0_00010010));
wire t0_000100100, t0_000100101;
mixer mix_t0_00010011 (.a(t0_000100110), .b(t0_000100111), .y(t0_00010011));
wire t0_000100110, t0_000100111;
mixer mix_t0_000101 (.a(t0_0001010), .b(t0_0001011), .y(t0_000101));
wire t0_0001010, t0_0001011;
mixer mix_t0_0001010 (.a(t0_00010100), .b(t0_00010101), .y(t0_0001010));
wire t0_00010100, t0_00010101;
mixer mix_t0_00010100 (.a(t0_000101000), .b(t0_000101001), .y(t0_00010100));
wire t0_000101000, t0_000101001;
mixer mix_t0_00010101 (.a(t0_000101010), .b(t0_000101011), .y(t0_00010101));
wire t0_000101010, t0_000101011;
mixer mix_t0_0001011 (.a(t0_00010110), .b(t0_00010111), .y(t0_0001011));
wire t0_00010110, t0_00010111;
mixer mix_t0_00010110 (.a(t0_000101100), .b(t0_000101101), .y(t0_00010110));
wire t0_000101100, t0_000101101;
mixer mix_t0_00010111 (.a(t0_000101110), .b(t0_000101111), .y(t0_00010111));
wire t0_000101110, t0_000101111;
mixer mix_t0_00011 (.a(t0_000110), .b(t0_000111), .y(t0_00011));
wire t0_000110, t0_000111;
mixer mix_t0_000110 (.a(t0_0001100), .b(t0_0001101), .y(t0_000110));
wire t0_0001100, t0_0001101;
mixer mix_t0_0001100 (.a(t0_00011000), .b(t0_00011001), .y(t0_0001100));
wire t0_00011000, t0_00011001;
mixer mix_t0_00011000 (.a(t0_000110000), .b(t0_000110001), .y(t0_00011000));
wire t0_000110000, t0_000110001;
mixer mix_t0_00011001 (.a(t0_000110010), .b(t0_000110011), .y(t0_00011001));
wire t0_000110010, t0_000110011;
mixer mix_t0_0001101 (.a(t0_00011010), .b(t0_00011011), .y(t0_0001101));
wire t0_00011010, t0_00011011;
mixer mix_t0_00011010 (.a(t0_000110100), .b(t0_000110101), .y(t0_00011010));
wire t0_000110100, t0_000110101;
mixer mix_t0_00011011 (.a(t0_000110110), .b(t0_000110111), .y(t0_00011011));
wire t0_000110110, t0_000110111;
mixer mix_t0_000111 (.a(t0_0001110), .b(t0_0001111), .y(t0_000111));
wire t0_0001110, t0_0001111;
mixer mix_t0_0001110 (.a(t0_00011100), .b(t0_00011101), .y(t0_0001110));
wire t0_00011100, t0_00011101;
mixer mix_t0_00011100 (.a(t0_000111000), .b(t0_000111001), .y(t0_00011100));
wire t0_000111000, t0_000111001;
mixer mix_t0_00011101 (.a(t0_000111010), .b(t0_000111011), .y(t0_00011101));
wire t0_000111010, t0_000111011;
mixer mix_t0_0001111 (.a(t0_00011110), .b(t0_00011111), .y(t0_0001111));
wire t0_00011110, t0_00011111;
mixer mix_t0_00011110 (.a(t0_000111100), .b(t0_000111101), .y(t0_00011110));
wire t0_000111100, t0_000111101;
mixer mix_t0_00011111 (.a(t0_000111110), .b(t0_000111111), .y(t0_00011111));
wire t0_000111110, t0_000111111;
mixer mix_t0_001 (.a(t0_0010), .b(t0_0011), .y(t0_001));
wire t0_0010, t0_0011;
mixer mix_t0_0010 (.a(t0_00100), .b(t0_00101), .y(t0_0010));
wire t0_00100, t0_00101;
mixer mix_t0_00100 (.a(t0_001000), .b(t0_001001), .y(t0_00100));
wire t0_001000, t0_001001;
mixer mix_t0_001000 (.a(t0_0010000), .b(t0_0010001), .y(t0_001000));
wire t0_0010000, t0_0010001;
mixer mix_t0_0010000 (.a(t0_00100000), .b(t0_00100001), .y(t0_0010000));
wire t0_00100000, t0_00100001;
mixer mix_t0_00100000 (.a(t0_001000000), .b(t0_001000001), .y(t0_00100000));
wire t0_001000000, t0_001000001;
mixer mix_t0_00100001 (.a(t0_001000010), .b(t0_001000011), .y(t0_00100001));
wire t0_001000010, t0_001000011;
mixer mix_t0_0010001 (.a(t0_00100010), .b(t0_00100011), .y(t0_0010001));
wire t0_00100010, t0_00100011;
mixer mix_t0_00100010 (.a(t0_001000100), .b(t0_001000101), .y(t0_00100010));
wire t0_001000100, t0_001000101;
mixer mix_t0_00100011 (.a(t0_001000110), .b(t0_001000111), .y(t0_00100011));
wire t0_001000110, t0_001000111;
mixer mix_t0_001001 (.a(t0_0010010), .b(t0_0010011), .y(t0_001001));
wire t0_0010010, t0_0010011;
mixer mix_t0_0010010 (.a(t0_00100100), .b(t0_00100101), .y(t0_0010010));
wire t0_00100100, t0_00100101;
mixer mix_t0_00100100 (.a(t0_001001000), .b(t0_001001001), .y(t0_00100100));
wire t0_001001000, t0_001001001;
mixer mix_t0_00100101 (.a(t0_001001010), .b(t0_001001011), .y(t0_00100101));
wire t0_001001010, t0_001001011;
mixer mix_t0_0010011 (.a(t0_00100110), .b(t0_00100111), .y(t0_0010011));
wire t0_00100110, t0_00100111;
mixer mix_t0_00100110 (.a(t0_001001100), .b(t0_001001101), .y(t0_00100110));
wire t0_001001100, t0_001001101;
mixer mix_t0_00100111 (.a(t0_001001110), .b(t0_001001111), .y(t0_00100111));
wire t0_001001110, t0_001001111;
mixer mix_t0_00101 (.a(t0_001010), .b(t0_001011), .y(t0_00101));
wire t0_001010, t0_001011;
mixer mix_t0_001010 (.a(t0_0010100), .b(t0_0010101), .y(t0_001010));
wire t0_0010100, t0_0010101;
mixer mix_t0_0010100 (.a(t0_00101000), .b(t0_00101001), .y(t0_0010100));
wire t0_00101000, t0_00101001;
mixer mix_t0_00101000 (.a(t0_001010000), .b(t0_001010001), .y(t0_00101000));
wire t0_001010000, t0_001010001;
mixer mix_t0_00101001 (.a(t0_001010010), .b(t0_001010011), .y(t0_00101001));
wire t0_001010010, t0_001010011;
mixer mix_t0_0010101 (.a(t0_00101010), .b(t0_00101011), .y(t0_0010101));
wire t0_00101010, t0_00101011;
mixer mix_t0_00101010 (.a(t0_001010100), .b(t0_001010101), .y(t0_00101010));
wire t0_001010100, t0_001010101;
mixer mix_t0_00101011 (.a(t0_001010110), .b(t0_001010111), .y(t0_00101011));
wire t0_001010110, t0_001010111;
mixer mix_t0_001011 (.a(t0_0010110), .b(t0_0010111), .y(t0_001011));
wire t0_0010110, t0_0010111;
mixer mix_t0_0010110 (.a(t0_00101100), .b(t0_00101101), .y(t0_0010110));
wire t0_00101100, t0_00101101;
mixer mix_t0_00101100 (.a(t0_001011000), .b(t0_001011001), .y(t0_00101100));
wire t0_001011000, t0_001011001;
mixer mix_t0_00101101 (.a(t0_001011010), .b(t0_001011011), .y(t0_00101101));
wire t0_001011010, t0_001011011;
mixer mix_t0_0010111 (.a(t0_00101110), .b(t0_00101111), .y(t0_0010111));
wire t0_00101110, t0_00101111;
mixer mix_t0_00101110 (.a(t0_001011100), .b(t0_001011101), .y(t0_00101110));
wire t0_001011100, t0_001011101;
mixer mix_t0_00101111 (.a(t0_001011110), .b(t0_001011111), .y(t0_00101111));
wire t0_001011110, t0_001011111;
mixer mix_t0_0011 (.a(t0_00110), .b(t0_00111), .y(t0_0011));
wire t0_00110, t0_00111;
mixer mix_t0_00110 (.a(t0_001100), .b(t0_001101), .y(t0_00110));
wire t0_001100, t0_001101;
mixer mix_t0_001100 (.a(t0_0011000), .b(t0_0011001), .y(t0_001100));
wire t0_0011000, t0_0011001;
mixer mix_t0_0011000 (.a(t0_00110000), .b(t0_00110001), .y(t0_0011000));
wire t0_00110000, t0_00110001;
mixer mix_t0_00110000 (.a(t0_001100000), .b(t0_001100001), .y(t0_00110000));
wire t0_001100000, t0_001100001;
mixer mix_t0_00110001 (.a(t0_001100010), .b(t0_001100011), .y(t0_00110001));
wire t0_001100010, t0_001100011;
mixer mix_t0_0011001 (.a(t0_00110010), .b(t0_00110011), .y(t0_0011001));
wire t0_00110010, t0_00110011;
mixer mix_t0_00110010 (.a(t0_001100100), .b(t0_001100101), .y(t0_00110010));
wire t0_001100100, t0_001100101;
mixer mix_t0_00110011 (.a(t0_001100110), .b(t0_001100111), .y(t0_00110011));
wire t0_001100110, t0_001100111;
mixer mix_t0_001101 (.a(t0_0011010), .b(t0_0011011), .y(t0_001101));
wire t0_0011010, t0_0011011;
mixer mix_t0_0011010 (.a(t0_00110100), .b(t0_00110101), .y(t0_0011010));
wire t0_00110100, t0_00110101;
mixer mix_t0_00110100 (.a(t0_001101000), .b(t0_001101001), .y(t0_00110100));
wire t0_001101000, t0_001101001;
mixer mix_t0_00110101 (.a(t0_001101010), .b(t0_001101011), .y(t0_00110101));
wire t0_001101010, t0_001101011;
mixer mix_t0_0011011 (.a(t0_00110110), .b(t0_00110111), .y(t0_0011011));
wire t0_00110110, t0_00110111;
mixer mix_t0_00110110 (.a(t0_001101100), .b(t0_001101101), .y(t0_00110110));
wire t0_001101100, t0_001101101;
mixer mix_t0_00110111 (.a(t0_001101110), .b(t0_001101111), .y(t0_00110111));
wire t0_001101110, t0_001101111;
mixer mix_t0_00111 (.a(t0_001110), .b(t0_001111), .y(t0_00111));
wire t0_001110, t0_001111;
mixer mix_t0_001110 (.a(t0_0011100), .b(t0_0011101), .y(t0_001110));
wire t0_0011100, t0_0011101;
mixer mix_t0_0011100 (.a(t0_00111000), .b(t0_00111001), .y(t0_0011100));
wire t0_00111000, t0_00111001;
mixer mix_t0_00111000 (.a(t0_001110000), .b(t0_001110001), .y(t0_00111000));
wire t0_001110000, t0_001110001;
mixer mix_t0_00111001 (.a(t0_001110010), .b(t0_001110011), .y(t0_00111001));
wire t0_001110010, t0_001110011;
mixer mix_t0_0011101 (.a(t0_00111010), .b(t0_00111011), .y(t0_0011101));
wire t0_00111010, t0_00111011;
mixer mix_t0_00111010 (.a(t0_001110100), .b(t0_001110101), .y(t0_00111010));
wire t0_001110100, t0_001110101;
mixer mix_t0_00111011 (.a(t0_001110110), .b(t0_001110111), .y(t0_00111011));
wire t0_001110110, t0_001110111;
mixer mix_t0_001111 (.a(t0_0011110), .b(t0_0011111), .y(t0_001111));
wire t0_0011110, t0_0011111;
mixer mix_t0_0011110 (.a(t0_00111100), .b(t0_00111101), .y(t0_0011110));
wire t0_00111100, t0_00111101;
mixer mix_t0_00111100 (.a(t0_001111000), .b(t0_001111001), .y(t0_00111100));
wire t0_001111000, t0_001111001;
mixer mix_t0_00111101 (.a(t0_001111010), .b(t0_001111011), .y(t0_00111101));
wire t0_001111010, t0_001111011;
mixer mix_t0_0011111 (.a(t0_00111110), .b(t0_00111111), .y(t0_0011111));
wire t0_00111110, t0_00111111;
mixer mix_t0_00111110 (.a(t0_001111100), .b(t0_001111101), .y(t0_00111110));
wire t0_001111100, t0_001111101;
mixer mix_t0_00111111 (.a(t0_001111110), .b(t0_001111111), .y(t0_00111111));
wire t0_001111110, t0_001111111;
mixer mix_t0_01 (.a(t0_010), .b(t0_011), .y(t0_01));
wire t0_010, t0_011;
mixer mix_t0_010 (.a(t0_0100), .b(t0_0101), .y(t0_010));
wire t0_0100, t0_0101;
mixer mix_t0_0100 (.a(t0_01000), .b(t0_01001), .y(t0_0100));
wire t0_01000, t0_01001;
mixer mix_t0_01000 (.a(t0_010000), .b(t0_010001), .y(t0_01000));
wire t0_010000, t0_010001;
mixer mix_t0_010000 (.a(t0_0100000), .b(t0_0100001), .y(t0_010000));
wire t0_0100000, t0_0100001;
mixer mix_t0_0100000 (.a(t0_01000000), .b(t0_01000001), .y(t0_0100000));
wire t0_01000000, t0_01000001;
mixer mix_t0_01000000 (.a(t0_010000000), .b(t0_010000001), .y(t0_01000000));
wire t0_010000000, t0_010000001;
mixer mix_t0_01000001 (.a(t0_010000010), .b(t0_010000011), .y(t0_01000001));
wire t0_010000010, t0_010000011;
mixer mix_t0_0100001 (.a(t0_01000010), .b(t0_01000011), .y(t0_0100001));
wire t0_01000010, t0_01000011;
mixer mix_t0_01000010 (.a(t0_010000100), .b(t0_010000101), .y(t0_01000010));
wire t0_010000100, t0_010000101;
mixer mix_t0_01000011 (.a(t0_010000110), .b(t0_010000111), .y(t0_01000011));
wire t0_010000110, t0_010000111;
mixer mix_t0_010001 (.a(t0_0100010), .b(t0_0100011), .y(t0_010001));
wire t0_0100010, t0_0100011;
mixer mix_t0_0100010 (.a(t0_01000100), .b(t0_01000101), .y(t0_0100010));
wire t0_01000100, t0_01000101;
mixer mix_t0_01000100 (.a(t0_010001000), .b(t0_010001001), .y(t0_01000100));
wire t0_010001000, t0_010001001;
mixer mix_t0_01000101 (.a(t0_010001010), .b(t0_010001011), .y(t0_01000101));
wire t0_010001010, t0_010001011;
mixer mix_t0_0100011 (.a(t0_01000110), .b(t0_01000111), .y(t0_0100011));
wire t0_01000110, t0_01000111;
mixer mix_t0_01000110 (.a(t0_010001100), .b(t0_010001101), .y(t0_01000110));
wire t0_010001100, t0_010001101;
mixer mix_t0_01000111 (.a(t0_010001110), .b(t0_010001111), .y(t0_01000111));
wire t0_010001110, t0_010001111;
mixer mix_t0_01001 (.a(t0_010010), .b(t0_010011), .y(t0_01001));
wire t0_010010, t0_010011;
mixer mix_t0_010010 (.a(t0_0100100), .b(t0_0100101), .y(t0_010010));
wire t0_0100100, t0_0100101;
mixer mix_t0_0100100 (.a(t0_01001000), .b(t0_01001001), .y(t0_0100100));
wire t0_01001000, t0_01001001;
mixer mix_t0_01001000 (.a(t0_010010000), .b(t0_010010001), .y(t0_01001000));
wire t0_010010000, t0_010010001;
mixer mix_t0_01001001 (.a(t0_010010010), .b(t0_010010011), .y(t0_01001001));
wire t0_010010010, t0_010010011;
mixer mix_t0_0100101 (.a(t0_01001010), .b(t0_01001011), .y(t0_0100101));
wire t0_01001010, t0_01001011;
mixer mix_t0_01001010 (.a(t0_010010100), .b(t0_010010101), .y(t0_01001010));
wire t0_010010100, t0_010010101;
mixer mix_t0_01001011 (.a(t0_010010110), .b(t0_010010111), .y(t0_01001011));
wire t0_010010110, t0_010010111;
mixer mix_t0_010011 (.a(t0_0100110), .b(t0_0100111), .y(t0_010011));
wire t0_0100110, t0_0100111;
mixer mix_t0_0100110 (.a(t0_01001100), .b(t0_01001101), .y(t0_0100110));
wire t0_01001100, t0_01001101;
mixer mix_t0_01001100 (.a(t0_010011000), .b(t0_010011001), .y(t0_01001100));
wire t0_010011000, t0_010011001;
mixer mix_t0_01001101 (.a(t0_010011010), .b(t0_010011011), .y(t0_01001101));
wire t0_010011010, t0_010011011;
mixer mix_t0_0100111 (.a(t0_01001110), .b(t0_01001111), .y(t0_0100111));
wire t0_01001110, t0_01001111;
mixer mix_t0_01001110 (.a(t0_010011100), .b(t0_010011101), .y(t0_01001110));
wire t0_010011100, t0_010011101;
mixer mix_t0_01001111 (.a(t0_010011110), .b(t0_010011111), .y(t0_01001111));
wire t0_010011110, t0_010011111;
mixer mix_t0_0101 (.a(t0_01010), .b(t0_01011), .y(t0_0101));
wire t0_01010, t0_01011;
mixer mix_t0_01010 (.a(t0_010100), .b(t0_010101), .y(t0_01010));
wire t0_010100, t0_010101;
mixer mix_t0_010100 (.a(t0_0101000), .b(t0_0101001), .y(t0_010100));
wire t0_0101000, t0_0101001;
mixer mix_t0_0101000 (.a(t0_01010000), .b(t0_01010001), .y(t0_0101000));
wire t0_01010000, t0_01010001;
mixer mix_t0_01010000 (.a(t0_010100000), .b(t0_010100001), .y(t0_01010000));
wire t0_010100000, t0_010100001;
mixer mix_t0_01010001 (.a(t0_010100010), .b(t0_010100011), .y(t0_01010001));
wire t0_010100010, t0_010100011;
mixer mix_t0_0101001 (.a(t0_01010010), .b(t0_01010011), .y(t0_0101001));
wire t0_01010010, t0_01010011;
mixer mix_t0_01010010 (.a(t0_010100100), .b(t0_010100101), .y(t0_01010010));
wire t0_010100100, t0_010100101;
mixer mix_t0_01010011 (.a(t0_010100110), .b(t0_010100111), .y(t0_01010011));
wire t0_010100110, t0_010100111;
mixer mix_t0_010101 (.a(t0_0101010), .b(t0_0101011), .y(t0_010101));
wire t0_0101010, t0_0101011;
mixer mix_t0_0101010 (.a(t0_01010100), .b(t0_01010101), .y(t0_0101010));
wire t0_01010100, t0_01010101;
mixer mix_t0_01010100 (.a(t0_010101000), .b(t0_010101001), .y(t0_01010100));
wire t0_010101000, t0_010101001;
mixer mix_t0_01010101 (.a(t0_010101010), .b(t0_010101011), .y(t0_01010101));
wire t0_010101010, t0_010101011;
mixer mix_t0_0101011 (.a(t0_01010110), .b(t0_01010111), .y(t0_0101011));
wire t0_01010110, t0_01010111;
mixer mix_t0_01010110 (.a(t0_010101100), .b(t0_010101101), .y(t0_01010110));
wire t0_010101100, t0_010101101;
mixer mix_t0_01010111 (.a(t0_010101110), .b(t0_010101111), .y(t0_01010111));
wire t0_010101110, t0_010101111;
mixer mix_t0_01011 (.a(t0_010110), .b(t0_010111), .y(t0_01011));
wire t0_010110, t0_010111;
mixer mix_t0_010110 (.a(t0_0101100), .b(t0_0101101), .y(t0_010110));
wire t0_0101100, t0_0101101;
mixer mix_t0_0101100 (.a(t0_01011000), .b(t0_01011001), .y(t0_0101100));
wire t0_01011000, t0_01011001;
mixer mix_t0_01011000 (.a(t0_010110000), .b(t0_010110001), .y(t0_01011000));
wire t0_010110000, t0_010110001;
mixer mix_t0_01011001 (.a(t0_010110010), .b(t0_010110011), .y(t0_01011001));
wire t0_010110010, t0_010110011;
mixer mix_t0_0101101 (.a(t0_01011010), .b(t0_01011011), .y(t0_0101101));
wire t0_01011010, t0_01011011;
mixer mix_t0_01011010 (.a(t0_010110100), .b(t0_010110101), .y(t0_01011010));
wire t0_010110100, t0_010110101;
mixer mix_t0_01011011 (.a(t0_010110110), .b(t0_010110111), .y(t0_01011011));
wire t0_010110110, t0_010110111;
mixer mix_t0_010111 (.a(t0_0101110), .b(t0_0101111), .y(t0_010111));
wire t0_0101110, t0_0101111;
mixer mix_t0_0101110 (.a(t0_01011100), .b(t0_01011101), .y(t0_0101110));
wire t0_01011100, t0_01011101;
mixer mix_t0_01011100 (.a(t0_010111000), .b(t0_010111001), .y(t0_01011100));
wire t0_010111000, t0_010111001;
mixer mix_t0_01011101 (.a(t0_010111010), .b(t0_010111011), .y(t0_01011101));
wire t0_010111010, t0_010111011;
mixer mix_t0_0101111 (.a(t0_01011110), .b(t0_01011111), .y(t0_0101111));
wire t0_01011110, t0_01011111;
mixer mix_t0_01011110 (.a(t0_010111100), .b(t0_010111101), .y(t0_01011110));
wire t0_010111100, t0_010111101;
mixer mix_t0_01011111 (.a(t0_010111110), .b(t0_010111111), .y(t0_01011111));
wire t0_010111110, t0_010111111;
mixer mix_t0_011 (.a(t0_0110), .b(t0_0111), .y(t0_011));
wire t0_0110, t0_0111;
mixer mix_t0_0110 (.a(t0_01100), .b(t0_01101), .y(t0_0110));
wire t0_01100, t0_01101;
mixer mix_t0_01100 (.a(t0_011000), .b(t0_011001), .y(t0_01100));
wire t0_011000, t0_011001;
mixer mix_t0_011000 (.a(t0_0110000), .b(t0_0110001), .y(t0_011000));
wire t0_0110000, t0_0110001;
mixer mix_t0_0110000 (.a(t0_01100000), .b(t0_01100001), .y(t0_0110000));
wire t0_01100000, t0_01100001;
mixer mix_t0_01100000 (.a(t0_011000000), .b(t0_011000001), .y(t0_01100000));
wire t0_011000000, t0_011000001;
mixer mix_t0_01100001 (.a(t0_011000010), .b(t0_011000011), .y(t0_01100001));
wire t0_011000010, t0_011000011;
mixer mix_t0_0110001 (.a(t0_01100010), .b(t0_01100011), .y(t0_0110001));
wire t0_01100010, t0_01100011;
mixer mix_t0_01100010 (.a(t0_011000100), .b(t0_011000101), .y(t0_01100010));
wire t0_011000100, t0_011000101;
mixer mix_t0_01100011 (.a(t0_011000110), .b(t0_011000111), .y(t0_01100011));
wire t0_011000110, t0_011000111;
mixer mix_t0_011001 (.a(t0_0110010), .b(t0_0110011), .y(t0_011001));
wire t0_0110010, t0_0110011;
mixer mix_t0_0110010 (.a(t0_01100100), .b(t0_01100101), .y(t0_0110010));
wire t0_01100100, t0_01100101;
mixer mix_t0_01100100 (.a(t0_011001000), .b(t0_011001001), .y(t0_01100100));
wire t0_011001000, t0_011001001;
mixer mix_t0_01100101 (.a(t0_011001010), .b(t0_011001011), .y(t0_01100101));
wire t0_011001010, t0_011001011;
mixer mix_t0_0110011 (.a(t0_01100110), .b(t0_01100111), .y(t0_0110011));
wire t0_01100110, t0_01100111;
mixer mix_t0_01100110 (.a(t0_011001100), .b(t0_011001101), .y(t0_01100110));
wire t0_011001100, t0_011001101;
mixer mix_t0_01100111 (.a(t0_011001110), .b(t0_011001111), .y(t0_01100111));
wire t0_011001110, t0_011001111;
mixer mix_t0_01101 (.a(t0_011010), .b(t0_011011), .y(t0_01101));
wire t0_011010, t0_011011;
mixer mix_t0_011010 (.a(t0_0110100), .b(t0_0110101), .y(t0_011010));
wire t0_0110100, t0_0110101;
mixer mix_t0_0110100 (.a(t0_01101000), .b(t0_01101001), .y(t0_0110100));
wire t0_01101000, t0_01101001;
mixer mix_t0_01101000 (.a(t0_011010000), .b(t0_011010001), .y(t0_01101000));
wire t0_011010000, t0_011010001;
mixer mix_t0_01101001 (.a(t0_011010010), .b(t0_011010011), .y(t0_01101001));
wire t0_011010010, t0_011010011;
mixer mix_t0_0110101 (.a(t0_01101010), .b(t0_01101011), .y(t0_0110101));
wire t0_01101010, t0_01101011;
mixer mix_t0_01101010 (.a(t0_011010100), .b(t0_011010101), .y(t0_01101010));
wire t0_011010100, t0_011010101;
mixer mix_t0_01101011 (.a(t0_011010110), .b(t0_011010111), .y(t0_01101011));
wire t0_011010110, t0_011010111;
mixer mix_t0_011011 (.a(t0_0110110), .b(t0_0110111), .y(t0_011011));
wire t0_0110110, t0_0110111;
mixer mix_t0_0110110 (.a(t0_01101100), .b(t0_01101101), .y(t0_0110110));
wire t0_01101100, t0_01101101;
mixer mix_t0_01101100 (.a(t0_011011000), .b(t0_011011001), .y(t0_01101100));
wire t0_011011000, t0_011011001;
mixer mix_t0_01101101 (.a(t0_011011010), .b(t0_011011011), .y(t0_01101101));
wire t0_011011010, t0_011011011;
mixer mix_t0_0110111 (.a(t0_01101110), .b(t0_01101111), .y(t0_0110111));
wire t0_01101110, t0_01101111;
mixer mix_t0_01101110 (.a(t0_011011100), .b(t0_011011101), .y(t0_01101110));
wire t0_011011100, t0_011011101;
mixer mix_t0_01101111 (.a(t0_011011110), .b(t0_011011111), .y(t0_01101111));
wire t0_011011110, t0_011011111;
mixer mix_t0_0111 (.a(t0_01110), .b(t0_01111), .y(t0_0111));
wire t0_01110, t0_01111;
mixer mix_t0_01110 (.a(t0_011100), .b(t0_011101), .y(t0_01110));
wire t0_011100, t0_011101;
mixer mix_t0_011100 (.a(t0_0111000), .b(t0_0111001), .y(t0_011100));
wire t0_0111000, t0_0111001;
mixer mix_t0_0111000 (.a(t0_01110000), .b(t0_01110001), .y(t0_0111000));
wire t0_01110000, t0_01110001;
mixer mix_t0_01110000 (.a(t0_011100000), .b(t0_011100001), .y(t0_01110000));
wire t0_011100000, t0_011100001;
mixer mix_t0_01110001 (.a(t0_011100010), .b(t0_011100011), .y(t0_01110001));
wire t0_011100010, t0_011100011;
mixer mix_t0_0111001 (.a(t0_01110010), .b(t0_01110011), .y(t0_0111001));
wire t0_01110010, t0_01110011;
mixer mix_t0_01110010 (.a(t0_011100100), .b(t0_011100101), .y(t0_01110010));
wire t0_011100100, t0_011100101;
mixer mix_t0_01110011 (.a(t0_011100110), .b(t0_011100111), .y(t0_01110011));
wire t0_011100110, t0_011100111;
mixer mix_t0_011101 (.a(t0_0111010), .b(t0_0111011), .y(t0_011101));
wire t0_0111010, t0_0111011;
mixer mix_t0_0111010 (.a(t0_01110100), .b(t0_01110101), .y(t0_0111010));
wire t0_01110100, t0_01110101;
mixer mix_t0_01110100 (.a(t0_011101000), .b(t0_011101001), .y(t0_01110100));
wire t0_011101000, t0_011101001;
mixer mix_t0_01110101 (.a(t0_011101010), .b(t0_011101011), .y(t0_01110101));
wire t0_011101010, t0_011101011;
mixer mix_t0_0111011 (.a(t0_01110110), .b(t0_01110111), .y(t0_0111011));
wire t0_01110110, t0_01110111;
mixer mix_t0_01110110 (.a(t0_011101100), .b(t0_011101101), .y(t0_01110110));
wire t0_011101100, t0_011101101;
mixer mix_t0_01110111 (.a(t0_011101110), .b(t0_011101111), .y(t0_01110111));
wire t0_011101110, t0_011101111;
mixer mix_t0_01111 (.a(t0_011110), .b(t0_011111), .y(t0_01111));
wire t0_011110, t0_011111;
mixer mix_t0_011110 (.a(t0_0111100), .b(t0_0111101), .y(t0_011110));
wire t0_0111100, t0_0111101;
mixer mix_t0_0111100 (.a(t0_01111000), .b(t0_01111001), .y(t0_0111100));
wire t0_01111000, t0_01111001;
mixer mix_t0_01111000 (.a(t0_011110000), .b(t0_011110001), .y(t0_01111000));
wire t0_011110000, t0_011110001;
mixer mix_t0_01111001 (.a(t0_011110010), .b(t0_011110011), .y(t0_01111001));
wire t0_011110010, t0_011110011;
mixer mix_t0_0111101 (.a(t0_01111010), .b(t0_01111011), .y(t0_0111101));
wire t0_01111010, t0_01111011;
mixer mix_t0_01111010 (.a(t0_011110100), .b(t0_011110101), .y(t0_01111010));
wire t0_011110100, t0_011110101;
mixer mix_t0_01111011 (.a(t0_011110110), .b(t0_011110111), .y(t0_01111011));
wire t0_011110110, t0_011110111;
mixer mix_t0_011111 (.a(t0_0111110), .b(t0_0111111), .y(t0_011111));
wire t0_0111110, t0_0111111;
mixer mix_t0_0111110 (.a(t0_01111100), .b(t0_01111101), .y(t0_0111110));
wire t0_01111100, t0_01111101;
mixer mix_t0_01111100 (.a(t0_011111000), .b(t0_011111001), .y(t0_01111100));
wire t0_011111000, t0_011111001;
mixer mix_t0_01111101 (.a(t0_011111010), .b(t0_011111011), .y(t0_01111101));
wire t0_011111010, t0_011111011;
mixer mix_t0_0111111 (.a(t0_01111110), .b(t0_01111111), .y(t0_0111111));
wire t0_01111110, t0_01111111;
mixer mix_t0_01111110 (.a(t0_011111100), .b(t0_011111101), .y(t0_01111110));
wire t0_011111100, t0_011111101;
mixer mix_t0_01111111 (.a(t0_011111110), .b(t0_011111111), .y(t0_01111111));
wire t0_011111110, t0_011111111;
mixer mix_t1_0 (.a(t1_00), .b(t1_01), .y(t1_0));
wire t1_00, t1_01;
mixer mix_t1_00 (.a(t1_000), .b(t1_001), .y(t1_00));
wire t1_000, t1_001;
mixer mix_t1_000 (.a(t1_0000), .b(t1_0001), .y(t1_000));
wire t1_0000, t1_0001;
mixer mix_t1_0000 (.a(t1_00000), .b(t1_00001), .y(t1_0000));
wire t1_00000, t1_00001;
mixer mix_t1_00000 (.a(t1_000000), .b(t1_000001), .y(t1_00000));
wire t1_000000, t1_000001;
mixer mix_t1_000000 (.a(t1_0000000), .b(t1_0000001), .y(t1_000000));
wire t1_0000000, t1_0000001;
mixer mix_t1_0000000 (.a(t1_00000000), .b(t1_00000001), .y(t1_0000000));
wire t1_00000000, t1_00000001;
mixer mix_t1_00000000 (.a(t1_000000000), .b(t1_000000001), .y(t1_00000000));
wire t1_000000000, t1_000000001;
mixer mix_t1_00000001 (.a(t1_000000010), .b(t1_000000011), .y(t1_00000001));
wire t1_000000010, t1_000000011;
mixer mix_t1_0000001 (.a(t1_00000010), .b(t1_00000011), .y(t1_0000001));
wire t1_00000010, t1_00000011;
mixer mix_t1_00000010 (.a(t1_000000100), .b(t1_000000101), .y(t1_00000010));
wire t1_000000100, t1_000000101;
mixer mix_t1_00000011 (.a(t1_000000110), .b(t1_000000111), .y(t1_00000011));
wire t1_000000110, t1_000000111;
mixer mix_t1_000001 (.a(t1_0000010), .b(t1_0000011), .y(t1_000001));
wire t1_0000010, t1_0000011;
mixer mix_t1_0000010 (.a(t1_00000100), .b(t1_00000101), .y(t1_0000010));
wire t1_00000100, t1_00000101;
mixer mix_t1_00000100 (.a(t1_000001000), .b(t1_000001001), .y(t1_00000100));
wire t1_000001000, t1_000001001;
mixer mix_t1_00000101 (.a(t1_000001010), .b(t1_000001011), .y(t1_00000101));
wire t1_000001010, t1_000001011;
mixer mix_t1_0000011 (.a(t1_00000110), .b(t1_00000111), .y(t1_0000011));
wire t1_00000110, t1_00000111;
mixer mix_t1_00000110 (.a(t1_000001100), .b(t1_000001101), .y(t1_00000110));
wire t1_000001100, t1_000001101;
mixer mix_t1_00000111 (.a(t1_000001110), .b(t1_000001111), .y(t1_00000111));
wire t1_000001110, t1_000001111;
mixer mix_t1_00001 (.a(t1_000010), .b(t1_000011), .y(t1_00001));
wire t1_000010, t1_000011;
mixer mix_t1_000010 (.a(t1_0000100), .b(t1_0000101), .y(t1_000010));
wire t1_0000100, t1_0000101;
mixer mix_t1_0000100 (.a(t1_00001000), .b(t1_00001001), .y(t1_0000100));
wire t1_00001000, t1_00001001;
mixer mix_t1_00001000 (.a(t1_000010000), .b(t1_000010001), .y(t1_00001000));
wire t1_000010000, t1_000010001;
mixer mix_t1_00001001 (.a(t1_000010010), .b(t1_000010011), .y(t1_00001001));
wire t1_000010010, t1_000010011;
mixer mix_t1_0000101 (.a(t1_00001010), .b(t1_00001011), .y(t1_0000101));
wire t1_00001010, t1_00001011;
mixer mix_t1_00001010 (.a(t1_000010100), .b(t1_000010101), .y(t1_00001010));
wire t1_000010100, t1_000010101;
mixer mix_t1_00001011 (.a(t1_000010110), .b(t1_000010111), .y(t1_00001011));
wire t1_000010110, t1_000010111;
mixer mix_t1_000011 (.a(t1_0000110), .b(t1_0000111), .y(t1_000011));
wire t1_0000110, t1_0000111;
mixer mix_t1_0000110 (.a(t1_00001100), .b(t1_00001101), .y(t1_0000110));
wire t1_00001100, t1_00001101;
mixer mix_t1_00001100 (.a(t1_000011000), .b(t1_000011001), .y(t1_00001100));
wire t1_000011000, t1_000011001;
mixer mix_t1_00001101 (.a(t1_000011010), .b(t1_000011011), .y(t1_00001101));
wire t1_000011010, t1_000011011;
mixer mix_t1_0000111 (.a(t1_00001110), .b(t1_00001111), .y(t1_0000111));
wire t1_00001110, t1_00001111;
mixer mix_t1_00001110 (.a(t1_000011100), .b(t1_000011101), .y(t1_00001110));
wire t1_000011100, t1_000011101;
mixer mix_t1_00001111 (.a(t1_000011110), .b(t1_000011111), .y(t1_00001111));
wire t1_000011110, t1_000011111;
mixer mix_t1_0001 (.a(t1_00010), .b(t1_00011), .y(t1_0001));
wire t1_00010, t1_00011;
mixer mix_t1_00010 (.a(t1_000100), .b(t1_000101), .y(t1_00010));
wire t1_000100, t1_000101;
mixer mix_t1_000100 (.a(t1_0001000), .b(t1_0001001), .y(t1_000100));
wire t1_0001000, t1_0001001;
mixer mix_t1_0001000 (.a(t1_00010000), .b(t1_00010001), .y(t1_0001000));
wire t1_00010000, t1_00010001;
mixer mix_t1_00010000 (.a(t1_000100000), .b(t1_000100001), .y(t1_00010000));
wire t1_000100000, t1_000100001;
mixer mix_t1_00010001 (.a(t1_000100010), .b(t1_000100011), .y(t1_00010001));
wire t1_000100010, t1_000100011;
mixer mix_t1_0001001 (.a(t1_00010010), .b(t1_00010011), .y(t1_0001001));
wire t1_00010010, t1_00010011;
mixer mix_t1_00010010 (.a(t1_000100100), .b(t1_000100101), .y(t1_00010010));
wire t1_000100100, t1_000100101;
mixer mix_t1_00010011 (.a(t1_000100110), .b(t1_000100111), .y(t1_00010011));
wire t1_000100110, t1_000100111;
mixer mix_t1_000101 (.a(t1_0001010), .b(t1_0001011), .y(t1_000101));
wire t1_0001010, t1_0001011;
mixer mix_t1_0001010 (.a(t1_00010100), .b(t1_00010101), .y(t1_0001010));
wire t1_00010100, t1_00010101;
mixer mix_t1_00010100 (.a(t1_000101000), .b(t1_000101001), .y(t1_00010100));
wire t1_000101000, t1_000101001;
mixer mix_t1_00010101 (.a(t1_000101010), .b(t1_000101011), .y(t1_00010101));
wire t1_000101010, t1_000101011;
mixer mix_t1_0001011 (.a(t1_00010110), .b(t1_00010111), .y(t1_0001011));
wire t1_00010110, t1_00010111;
mixer mix_t1_00010110 (.a(t1_000101100), .b(t1_000101101), .y(t1_00010110));
wire t1_000101100, t1_000101101;
mixer mix_t1_00010111 (.a(t1_000101110), .b(t1_000101111), .y(t1_00010111));
wire t1_000101110, t1_000101111;
mixer mix_t1_00011 (.a(t1_000110), .b(t1_000111), .y(t1_00011));
wire t1_000110, t1_000111;
mixer mix_t1_000110 (.a(t1_0001100), .b(t1_0001101), .y(t1_000110));
wire t1_0001100, t1_0001101;
mixer mix_t1_0001100 (.a(t1_00011000), .b(t1_00011001), .y(t1_0001100));
wire t1_00011000, t1_00011001;
mixer mix_t1_00011000 (.a(t1_000110000), .b(t1_000110001), .y(t1_00011000));
wire t1_000110000, t1_000110001;
mixer mix_t1_00011001 (.a(t1_000110010), .b(t1_000110011), .y(t1_00011001));
wire t1_000110010, t1_000110011;
mixer mix_t1_0001101 (.a(t1_00011010), .b(t1_00011011), .y(t1_0001101));
wire t1_00011010, t1_00011011;
mixer mix_t1_00011010 (.a(t1_000110100), .b(t1_000110101), .y(t1_00011010));
wire t1_000110100, t1_000110101;
mixer mix_t1_00011011 (.a(t1_000110110), .b(t1_000110111), .y(t1_00011011));
wire t1_000110110, t1_000110111;
mixer mix_t1_000111 (.a(t1_0001110), .b(t1_0001111), .y(t1_000111));
wire t1_0001110, t1_0001111;
mixer mix_t1_0001110 (.a(t1_00011100), .b(t1_00011101), .y(t1_0001110));
wire t1_00011100, t1_00011101;
mixer mix_t1_00011100 (.a(t1_000111000), .b(t1_000111001), .y(t1_00011100));
wire t1_000111000, t1_000111001;
mixer mix_t1_00011101 (.a(t1_000111010), .b(t1_000111011), .y(t1_00011101));
wire t1_000111010, t1_000111011;
mixer mix_t1_0001111 (.a(t1_00011110), .b(t1_00011111), .y(t1_0001111));
wire t1_00011110, t1_00011111;
mixer mix_t1_00011110 (.a(t1_000111100), .b(t1_000111101), .y(t1_00011110));
wire t1_000111100, t1_000111101;
mixer mix_t1_00011111 (.a(t1_000111110), .b(t1_000111111), .y(t1_00011111));
wire t1_000111110, t1_000111111;
mixer mix_t1_001 (.a(t1_0010), .b(t1_0011), .y(t1_001));
wire t1_0010, t1_0011;
mixer mix_t1_0010 (.a(t1_00100), .b(t1_00101), .y(t1_0010));
wire t1_00100, t1_00101;
mixer mix_t1_00100 (.a(t1_001000), .b(t1_001001), .y(t1_00100));
wire t1_001000, t1_001001;
mixer mix_t1_001000 (.a(t1_0010000), .b(t1_0010001), .y(t1_001000));
wire t1_0010000, t1_0010001;
mixer mix_t1_0010000 (.a(t1_00100000), .b(t1_00100001), .y(t1_0010000));
wire t1_00100000, t1_00100001;
mixer mix_t1_00100000 (.a(t1_001000000), .b(t1_001000001), .y(t1_00100000));
wire t1_001000000, t1_001000001;
mixer mix_t1_00100001 (.a(t1_001000010), .b(t1_001000011), .y(t1_00100001));
wire t1_001000010, t1_001000011;
mixer mix_t1_0010001 (.a(t1_00100010), .b(t1_00100011), .y(t1_0010001));
wire t1_00100010, t1_00100011;
mixer mix_t1_00100010 (.a(t1_001000100), .b(t1_001000101), .y(t1_00100010));
wire t1_001000100, t1_001000101;
mixer mix_t1_00100011 (.a(t1_001000110), .b(t1_001000111), .y(t1_00100011));
wire t1_001000110, t1_001000111;
mixer mix_t1_001001 (.a(t1_0010010), .b(t1_0010011), .y(t1_001001));
wire t1_0010010, t1_0010011;
mixer mix_t1_0010010 (.a(t1_00100100), .b(t1_00100101), .y(t1_0010010));
wire t1_00100100, t1_00100101;
mixer mix_t1_00100100 (.a(t1_001001000), .b(t1_001001001), .y(t1_00100100));
wire t1_001001000, t1_001001001;
mixer mix_t1_00100101 (.a(t1_001001010), .b(t1_001001011), .y(t1_00100101));
wire t1_001001010, t1_001001011;
mixer mix_t1_0010011 (.a(t1_00100110), .b(t1_00100111), .y(t1_0010011));
wire t1_00100110, t1_00100111;
mixer mix_t1_00100110 (.a(t1_001001100), .b(t1_001001101), .y(t1_00100110));
wire t1_001001100, t1_001001101;
mixer mix_t1_00100111 (.a(t1_001001110), .b(t1_001001111), .y(t1_00100111));
wire t1_001001110, t1_001001111;
mixer mix_t1_00101 (.a(t1_001010), .b(t1_001011), .y(t1_00101));
wire t1_001010, t1_001011;
mixer mix_t1_001010 (.a(t1_0010100), .b(t1_0010101), .y(t1_001010));
wire t1_0010100, t1_0010101;
mixer mix_t1_0010100 (.a(t1_00101000), .b(t1_00101001), .y(t1_0010100));
wire t1_00101000, t1_00101001;
mixer mix_t1_00101000 (.a(t1_001010000), .b(t1_001010001), .y(t1_00101000));
wire t1_001010000, t1_001010001;
mixer mix_t1_00101001 (.a(t1_001010010), .b(t1_001010011), .y(t1_00101001));
wire t1_001010010, t1_001010011;
mixer mix_t1_0010101 (.a(t1_00101010), .b(t1_00101011), .y(t1_0010101));
wire t1_00101010, t1_00101011;
mixer mix_t1_00101010 (.a(t1_001010100), .b(t1_001010101), .y(t1_00101010));
wire t1_001010100, t1_001010101;
mixer mix_t1_00101011 (.a(t1_001010110), .b(t1_001010111), .y(t1_00101011));
wire t1_001010110, t1_001010111;
mixer mix_t1_001011 (.a(t1_0010110), .b(t1_0010111), .y(t1_001011));
wire t1_0010110, t1_0010111;
mixer mix_t1_0010110 (.a(t1_00101100), .b(t1_00101101), .y(t1_0010110));
wire t1_00101100, t1_00101101;
mixer mix_t1_00101100 (.a(t1_001011000), .b(t1_001011001), .y(t1_00101100));
wire t1_001011000, t1_001011001;
mixer mix_t1_00101101 (.a(t1_001011010), .b(t1_001011011), .y(t1_00101101));
wire t1_001011010, t1_001011011;
mixer mix_t1_0010111 (.a(t1_00101110), .b(t1_00101111), .y(t1_0010111));
wire t1_00101110, t1_00101111;
mixer mix_t1_00101110 (.a(t1_001011100), .b(t1_001011101), .y(t1_00101110));
wire t1_001011100, t1_001011101;
mixer mix_t1_00101111 (.a(t1_001011110), .b(t1_001011111), .y(t1_00101111));
wire t1_001011110, t1_001011111;
mixer mix_t1_0011 (.a(t1_00110), .b(t1_00111), .y(t1_0011));
wire t1_00110, t1_00111;
mixer mix_t1_00110 (.a(t1_001100), .b(t1_001101), .y(t1_00110));
wire t1_001100, t1_001101;
mixer mix_t1_001100 (.a(t1_0011000), .b(t1_0011001), .y(t1_001100));
wire t1_0011000, t1_0011001;
mixer mix_t1_0011000 (.a(t1_00110000), .b(t1_00110001), .y(t1_0011000));
wire t1_00110000, t1_00110001;
mixer mix_t1_00110000 (.a(t1_001100000), .b(t1_001100001), .y(t1_00110000));
wire t1_001100000, t1_001100001;
mixer mix_t1_00110001 (.a(t1_001100010), .b(t1_001100011), .y(t1_00110001));
wire t1_001100010, t1_001100011;
mixer mix_t1_0011001 (.a(t1_00110010), .b(t1_00110011), .y(t1_0011001));
wire t1_00110010, t1_00110011;
mixer mix_t1_00110010 (.a(t1_001100100), .b(t1_001100101), .y(t1_00110010));
wire t1_001100100, t1_001100101;
mixer mix_t1_00110011 (.a(t1_001100110), .b(t1_001100111), .y(t1_00110011));
wire t1_001100110, t1_001100111;
mixer mix_t1_001101 (.a(t1_0011010), .b(t1_0011011), .y(t1_001101));
wire t1_0011010, t1_0011011;
mixer mix_t1_0011010 (.a(t1_00110100), .b(t1_00110101), .y(t1_0011010));
wire t1_00110100, t1_00110101;
mixer mix_t1_00110100 (.a(t1_001101000), .b(t1_001101001), .y(t1_00110100));
wire t1_001101000, t1_001101001;
mixer mix_t1_00110101 (.a(t1_001101010), .b(t1_001101011), .y(t1_00110101));
wire t1_001101010, t1_001101011;
mixer mix_t1_0011011 (.a(t1_00110110), .b(t1_00110111), .y(t1_0011011));
wire t1_00110110, t1_00110111;
mixer mix_t1_00110110 (.a(t1_001101100), .b(t1_001101101), .y(t1_00110110));
wire t1_001101100, t1_001101101;
mixer mix_t1_00110111 (.a(t1_001101110), .b(t1_001101111), .y(t1_00110111));
wire t1_001101110, t1_001101111;
mixer mix_t1_00111 (.a(t1_001110), .b(t1_001111), .y(t1_00111));
wire t1_001110, t1_001111;
mixer mix_t1_001110 (.a(t1_0011100), .b(t1_0011101), .y(t1_001110));
wire t1_0011100, t1_0011101;
mixer mix_t1_0011100 (.a(t1_00111000), .b(t1_00111001), .y(t1_0011100));
wire t1_00111000, t1_00111001;
mixer mix_t1_00111000 (.a(t1_001110000), .b(t1_001110001), .y(t1_00111000));
wire t1_001110000, t1_001110001;
mixer mix_t1_00111001 (.a(t1_001110010), .b(t1_001110011), .y(t1_00111001));
wire t1_001110010, t1_001110011;
mixer mix_t1_0011101 (.a(t1_00111010), .b(t1_00111011), .y(t1_0011101));
wire t1_00111010, t1_00111011;
mixer mix_t1_00111010 (.a(t1_001110100), .b(t1_001110101), .y(t1_00111010));
wire t1_001110100, t1_001110101;
mixer mix_t1_00111011 (.a(t1_001110110), .b(t1_001110111), .y(t1_00111011));
wire t1_001110110, t1_001110111;
mixer mix_t1_001111 (.a(t1_0011110), .b(t1_0011111), .y(t1_001111));
wire t1_0011110, t1_0011111;
mixer mix_t1_0011110 (.a(t1_00111100), .b(t1_00111101), .y(t1_0011110));
wire t1_00111100, t1_00111101;
mixer mix_t1_00111100 (.a(t1_001111000), .b(t1_001111001), .y(t1_00111100));
wire t1_001111000, t1_001111001;
mixer mix_t1_00111101 (.a(t1_001111010), .b(t1_001111011), .y(t1_00111101));
wire t1_001111010, t1_001111011;
mixer mix_t1_0011111 (.a(t1_00111110), .b(t1_00111111), .y(t1_0011111));
wire t1_00111110, t1_00111111;
mixer mix_t1_00111110 (.a(t1_001111100), .b(t1_001111101), .y(t1_00111110));
wire t1_001111100, t1_001111101;
mixer mix_t1_00111111 (.a(t1_001111110), .b(t1_001111111), .y(t1_00111111));
wire t1_001111110, t1_001111111;
mixer mix_t1_01 (.a(t1_010), .b(t1_011), .y(t1_01));
wire t1_010, t1_011;
mixer mix_t1_010 (.a(t1_0100), .b(t1_0101), .y(t1_010));
wire t1_0100, t1_0101;
mixer mix_t1_0100 (.a(t1_01000), .b(t1_01001), .y(t1_0100));
wire t1_01000, t1_01001;
mixer mix_t1_01000 (.a(t1_010000), .b(t1_010001), .y(t1_01000));
wire t1_010000, t1_010001;
mixer mix_t1_010000 (.a(t1_0100000), .b(t1_0100001), .y(t1_010000));
wire t1_0100000, t1_0100001;
mixer mix_t1_0100000 (.a(t1_01000000), .b(t1_01000001), .y(t1_0100000));
wire t1_01000000, t1_01000001;
mixer mix_t1_01000000 (.a(t1_010000000), .b(t1_010000001), .y(t1_01000000));
wire t1_010000000, t1_010000001;
mixer mix_t1_01000001 (.a(t1_010000010), .b(t1_010000011), .y(t1_01000001));
wire t1_010000010, t1_010000011;
mixer mix_t1_0100001 (.a(t1_01000010), .b(t1_01000011), .y(t1_0100001));
wire t1_01000010, t1_01000011;
mixer mix_t1_01000010 (.a(t1_010000100), .b(t1_010000101), .y(t1_01000010));
wire t1_010000100, t1_010000101;
mixer mix_t1_01000011 (.a(t1_010000110), .b(t1_010000111), .y(t1_01000011));
wire t1_010000110, t1_010000111;
mixer mix_t1_010001 (.a(t1_0100010), .b(t1_0100011), .y(t1_010001));
wire t1_0100010, t1_0100011;
mixer mix_t1_0100010 (.a(t1_01000100), .b(t1_01000101), .y(t1_0100010));
wire t1_01000100, t1_01000101;
mixer mix_t1_01000100 (.a(t1_010001000), .b(t1_010001001), .y(t1_01000100));
wire t1_010001000, t1_010001001;
mixer mix_t1_01000101 (.a(t1_010001010), .b(t1_010001011), .y(t1_01000101));
wire t1_010001010, t1_010001011;
mixer mix_t1_0100011 (.a(t1_01000110), .b(t1_01000111), .y(t1_0100011));
wire t1_01000110, t1_01000111;
mixer mix_t1_01000110 (.a(t1_010001100), .b(t1_010001101), .y(t1_01000110));
wire t1_010001100, t1_010001101;
mixer mix_t1_01000111 (.a(t1_010001110), .b(t1_010001111), .y(t1_01000111));
wire t1_010001110, t1_010001111;
mixer mix_t1_01001 (.a(t1_010010), .b(t1_010011), .y(t1_01001));
wire t1_010010, t1_010011;
mixer mix_t1_010010 (.a(t1_0100100), .b(t1_0100101), .y(t1_010010));
wire t1_0100100, t1_0100101;
mixer mix_t1_0100100 (.a(t1_01001000), .b(t1_01001001), .y(t1_0100100));
wire t1_01001000, t1_01001001;
mixer mix_t1_01001000 (.a(t1_010010000), .b(t1_010010001), .y(t1_01001000));
wire t1_010010000, t1_010010001;
mixer mix_t1_01001001 (.a(t1_010010010), .b(t1_010010011), .y(t1_01001001));
wire t1_010010010, t1_010010011;
mixer mix_t1_0100101 (.a(t1_01001010), .b(t1_01001011), .y(t1_0100101));
wire t1_01001010, t1_01001011;
mixer mix_t1_01001010 (.a(t1_010010100), .b(t1_010010101), .y(t1_01001010));
wire t1_010010100, t1_010010101;
mixer mix_t1_01001011 (.a(t1_010010110), .b(t1_010010111), .y(t1_01001011));
wire t1_010010110, t1_010010111;
mixer mix_t1_010011 (.a(t1_0100110), .b(t1_0100111), .y(t1_010011));
wire t1_0100110, t1_0100111;
mixer mix_t1_0100110 (.a(t1_01001100), .b(t1_01001101), .y(t1_0100110));
wire t1_01001100, t1_01001101;
mixer mix_t1_01001100 (.a(t1_010011000), .b(t1_010011001), .y(t1_01001100));
wire t1_010011000, t1_010011001;
mixer mix_t1_01001101 (.a(t1_010011010), .b(t1_010011011), .y(t1_01001101));
wire t1_010011010, t1_010011011;
mixer mix_t1_0100111 (.a(t1_01001110), .b(t1_01001111), .y(t1_0100111));
wire t1_01001110, t1_01001111;
mixer mix_t1_01001110 (.a(t1_010011100), .b(t1_010011101), .y(t1_01001110));
wire t1_010011100, t1_010011101;
mixer mix_t1_01001111 (.a(t1_010011110), .b(t1_010011111), .y(t1_01001111));
wire t1_010011110, t1_010011111;
mixer mix_t1_0101 (.a(t1_01010), .b(t1_01011), .y(t1_0101));
wire t1_01010, t1_01011;
mixer mix_t1_01010 (.a(t1_010100), .b(t1_010101), .y(t1_01010));
wire t1_010100, t1_010101;
mixer mix_t1_010100 (.a(t1_0101000), .b(t1_0101001), .y(t1_010100));
wire t1_0101000, t1_0101001;
mixer mix_t1_0101000 (.a(t1_01010000), .b(t1_01010001), .y(t1_0101000));
wire t1_01010000, t1_01010001;
mixer mix_t1_01010000 (.a(t1_010100000), .b(t1_010100001), .y(t1_01010000));
wire t1_010100000, t1_010100001;
mixer mix_t1_01010001 (.a(t1_010100010), .b(t1_010100011), .y(t1_01010001));
wire t1_010100010, t1_010100011;
mixer mix_t1_0101001 (.a(t1_01010010), .b(t1_01010011), .y(t1_0101001));
wire t1_01010010, t1_01010011;
mixer mix_t1_01010010 (.a(t1_010100100), .b(t1_010100101), .y(t1_01010010));
wire t1_010100100, t1_010100101;
mixer mix_t1_01010011 (.a(t1_010100110), .b(t1_010100111), .y(t1_01010011));
wire t1_010100110, t1_010100111;
mixer mix_t1_010101 (.a(t1_0101010), .b(t1_0101011), .y(t1_010101));
wire t1_0101010, t1_0101011;
mixer mix_t1_0101010 (.a(t1_01010100), .b(t1_01010101), .y(t1_0101010));
wire t1_01010100, t1_01010101;
mixer mix_t1_01010100 (.a(t1_010101000), .b(t1_010101001), .y(t1_01010100));
wire t1_010101000, t1_010101001;
mixer mix_t1_01010101 (.a(t1_010101010), .b(t1_010101011), .y(t1_01010101));
wire t1_010101010, t1_010101011;
mixer mix_t1_0101011 (.a(t1_01010110), .b(t1_01010111), .y(t1_0101011));
wire t1_01010110, t1_01010111;
mixer mix_t1_01010110 (.a(t1_010101100), .b(t1_010101101), .y(t1_01010110));
wire t1_010101100, t1_010101101;
mixer mix_t1_01010111 (.a(t1_010101110), .b(t1_010101111), .y(t1_01010111));
wire t1_010101110, t1_010101111;
mixer mix_t1_01011 (.a(t1_010110), .b(t1_010111), .y(t1_01011));
wire t1_010110, t1_010111;
mixer mix_t1_010110 (.a(t1_0101100), .b(t1_0101101), .y(t1_010110));
wire t1_0101100, t1_0101101;
mixer mix_t1_0101100 (.a(t1_01011000), .b(t1_01011001), .y(t1_0101100));
wire t1_01011000, t1_01011001;
mixer mix_t1_01011000 (.a(t1_010110000), .b(t1_010110001), .y(t1_01011000));
wire t1_010110000, t1_010110001;
mixer mix_t1_01011001 (.a(t1_010110010), .b(t1_010110011), .y(t1_01011001));
wire t1_010110010, t1_010110011;
mixer mix_t1_0101101 (.a(t1_01011010), .b(t1_01011011), .y(t1_0101101));
wire t1_01011010, t1_01011011;
mixer mix_t1_01011010 (.a(t1_010110100), .b(t1_010110101), .y(t1_01011010));
wire t1_010110100, t1_010110101;
mixer mix_t1_01011011 (.a(t1_010110110), .b(t1_010110111), .y(t1_01011011));
wire t1_010110110, t1_010110111;
mixer mix_t1_010111 (.a(t1_0101110), .b(t1_0101111), .y(t1_010111));
wire t1_0101110, t1_0101111;
mixer mix_t1_0101110 (.a(t1_01011100), .b(t1_01011101), .y(t1_0101110));
wire t1_01011100, t1_01011101;
mixer mix_t1_01011100 (.a(t1_010111000), .b(t1_010111001), .y(t1_01011100));
wire t1_010111000, t1_010111001;
mixer mix_t1_01011101 (.a(t1_010111010), .b(t1_010111011), .y(t1_01011101));
wire t1_010111010, t1_010111011;
mixer mix_t1_0101111 (.a(t1_01011110), .b(t1_01011111), .y(t1_0101111));
wire t1_01011110, t1_01011111;
mixer mix_t1_01011110 (.a(t1_010111100), .b(t1_010111101), .y(t1_01011110));
wire t1_010111100, t1_010111101;
mixer mix_t1_01011111 (.a(t1_010111110), .b(t1_010111111), .y(t1_01011111));
wire t1_010111110, t1_010111111;
mixer mix_t1_011 (.a(t1_0110), .b(t1_0111), .y(t1_011));
wire t1_0110, t1_0111;
mixer mix_t1_0110 (.a(t1_01100), .b(t1_01101), .y(t1_0110));
wire t1_01100, t1_01101;
mixer mix_t1_01100 (.a(t1_011000), .b(t1_011001), .y(t1_01100));
wire t1_011000, t1_011001;
mixer mix_t1_011000 (.a(t1_0110000), .b(t1_0110001), .y(t1_011000));
wire t1_0110000, t1_0110001;
mixer mix_t1_0110000 (.a(t1_01100000), .b(t1_01100001), .y(t1_0110000));
wire t1_01100000, t1_01100001;
mixer mix_t1_01100000 (.a(t1_011000000), .b(t1_011000001), .y(t1_01100000));
wire t1_011000000, t1_011000001;
mixer mix_t1_01100001 (.a(t1_011000010), .b(t1_011000011), .y(t1_01100001));
wire t1_011000010, t1_011000011;
mixer mix_t1_0110001 (.a(t1_01100010), .b(t1_01100011), .y(t1_0110001));
wire t1_01100010, t1_01100011;
mixer mix_t1_01100010 (.a(t1_011000100), .b(t1_011000101), .y(t1_01100010));
wire t1_011000100, t1_011000101;
mixer mix_t1_01100011 (.a(t1_011000110), .b(t1_011000111), .y(t1_01100011));
wire t1_011000110, t1_011000111;
mixer mix_t1_011001 (.a(t1_0110010), .b(t1_0110011), .y(t1_011001));
wire t1_0110010, t1_0110011;
mixer mix_t1_0110010 (.a(t1_01100100), .b(t1_01100101), .y(t1_0110010));
wire t1_01100100, t1_01100101;
mixer mix_t1_01100100 (.a(t1_011001000), .b(t1_011001001), .y(t1_01100100));
wire t1_011001000, t1_011001001;
mixer mix_t1_01100101 (.a(t1_011001010), .b(t1_011001011), .y(t1_01100101));
wire t1_011001010, t1_011001011;
mixer mix_t1_0110011 (.a(t1_01100110), .b(t1_01100111), .y(t1_0110011));
wire t1_01100110, t1_01100111;
mixer mix_t1_01100110 (.a(t1_011001100), .b(t1_011001101), .y(t1_01100110));
wire t1_011001100, t1_011001101;
mixer mix_t1_01100111 (.a(t1_011001110), .b(t1_011001111), .y(t1_01100111));
wire t1_011001110, t1_011001111;
mixer mix_t1_01101 (.a(t1_011010), .b(t1_011011), .y(t1_01101));
wire t1_011010, t1_011011;
mixer mix_t1_011010 (.a(t1_0110100), .b(t1_0110101), .y(t1_011010));
wire t1_0110100, t1_0110101;
mixer mix_t1_0110100 (.a(t1_01101000), .b(t1_01101001), .y(t1_0110100));
wire t1_01101000, t1_01101001;
mixer mix_t1_01101000 (.a(t1_011010000), .b(t1_011010001), .y(t1_01101000));
wire t1_011010000, t1_011010001;
mixer mix_t1_01101001 (.a(t1_011010010), .b(t1_011010011), .y(t1_01101001));
wire t1_011010010, t1_011010011;
mixer mix_t1_0110101 (.a(t1_01101010), .b(t1_01101011), .y(t1_0110101));
wire t1_01101010, t1_01101011;
mixer mix_t1_01101010 (.a(t1_011010100), .b(t1_011010101), .y(t1_01101010));
wire t1_011010100, t1_011010101;
mixer mix_t1_01101011 (.a(t1_011010110), .b(t1_011010111), .y(t1_01101011));
wire t1_011010110, t1_011010111;
mixer mix_t1_011011 (.a(t1_0110110), .b(t1_0110111), .y(t1_011011));
wire t1_0110110, t1_0110111;
mixer mix_t1_0110110 (.a(t1_01101100), .b(t1_01101101), .y(t1_0110110));
wire t1_01101100, t1_01101101;
mixer mix_t1_01101100 (.a(t1_011011000), .b(t1_011011001), .y(t1_01101100));
wire t1_011011000, t1_011011001;
mixer mix_t1_01101101 (.a(t1_011011010), .b(t1_011011011), .y(t1_01101101));
wire t1_011011010, t1_011011011;
mixer mix_t1_0110111 (.a(t1_01101110), .b(t1_01101111), .y(t1_0110111));
wire t1_01101110, t1_01101111;
mixer mix_t1_01101110 (.a(t1_011011100), .b(t1_011011101), .y(t1_01101110));
wire t1_011011100, t1_011011101;
mixer mix_t1_01101111 (.a(t1_011011110), .b(t1_011011111), .y(t1_01101111));
wire t1_011011110, t1_011011111;
mixer mix_t1_0111 (.a(t1_01110), .b(t1_01111), .y(t1_0111));
wire t1_01110, t1_01111;
mixer mix_t1_01110 (.a(t1_011100), .b(t1_011101), .y(t1_01110));
wire t1_011100, t1_011101;
mixer mix_t1_011100 (.a(t1_0111000), .b(t1_0111001), .y(t1_011100));
wire t1_0111000, t1_0111001;
mixer mix_t1_0111000 (.a(t1_01110000), .b(t1_01110001), .y(t1_0111000));
wire t1_01110000, t1_01110001;
mixer mix_t1_01110000 (.a(t1_011100000), .b(t1_011100001), .y(t1_01110000));
wire t1_011100000, t1_011100001;
mixer mix_t1_01110001 (.a(t1_011100010), .b(t1_011100011), .y(t1_01110001));
wire t1_011100010, t1_011100011;
mixer mix_t1_0111001 (.a(t1_01110010), .b(t1_01110011), .y(t1_0111001));
wire t1_01110010, t1_01110011;
mixer mix_t1_01110010 (.a(t1_011100100), .b(t1_011100101), .y(t1_01110010));
wire t1_011100100, t1_011100101;
mixer mix_t1_01110011 (.a(t1_011100110), .b(t1_011100111), .y(t1_01110011));
wire t1_011100110, t1_011100111;
mixer mix_t1_011101 (.a(t1_0111010), .b(t1_0111011), .y(t1_011101));
wire t1_0111010, t1_0111011;
mixer mix_t1_0111010 (.a(t1_01110100), .b(t1_01110101), .y(t1_0111010));
wire t1_01110100, t1_01110101;
mixer mix_t1_01110100 (.a(t1_011101000), .b(t1_011101001), .y(t1_01110100));
wire t1_011101000, t1_011101001;
mixer mix_t1_01110101 (.a(t1_011101010), .b(t1_011101011), .y(t1_01110101));
wire t1_011101010, t1_011101011;
mixer mix_t1_0111011 (.a(t1_01110110), .b(t1_01110111), .y(t1_0111011));
wire t1_01110110, t1_01110111;
mixer mix_t1_01110110 (.a(t1_011101100), .b(t1_011101101), .y(t1_01110110));
wire t1_011101100, t1_011101101;
mixer mix_t1_01110111 (.a(t1_011101110), .b(t1_011101111), .y(t1_01110111));
wire t1_011101110, t1_011101111;
mixer mix_t1_01111 (.a(t1_011110), .b(t1_011111), .y(t1_01111));
wire t1_011110, t1_011111;
mixer mix_t1_011110 (.a(t1_0111100), .b(t1_0111101), .y(t1_011110));
wire t1_0111100, t1_0111101;
mixer mix_t1_0111100 (.a(t1_01111000), .b(t1_01111001), .y(t1_0111100));
wire t1_01111000, t1_01111001;
mixer mix_t1_01111000 (.a(t1_011110000), .b(t1_011110001), .y(t1_01111000));
wire t1_011110000, t1_011110001;
mixer mix_t1_01111001 (.a(t1_011110010), .b(t1_011110011), .y(t1_01111001));
wire t1_011110010, t1_011110011;
mixer mix_t1_0111101 (.a(t1_01111010), .b(t1_01111011), .y(t1_0111101));
wire t1_01111010, t1_01111011;
mixer mix_t1_01111010 (.a(t1_011110100), .b(t1_011110101), .y(t1_01111010));
wire t1_011110100, t1_011110101;
mixer mix_t1_01111011 (.a(t1_011110110), .b(t1_011110111), .y(t1_01111011));
wire t1_011110110, t1_011110111;
mixer mix_t1_011111 (.a(t1_0111110), .b(t1_0111111), .y(t1_011111));
wire t1_0111110, t1_0111111;
mixer mix_t1_0111110 (.a(t1_01111100), .b(t1_01111101), .y(t1_0111110));
wire t1_01111100, t1_01111101;
mixer mix_t1_01111100 (.a(t1_011111000), .b(t1_011111001), .y(t1_01111100));
wire t1_011111000, t1_011111001;
mixer mix_t1_01111101 (.a(t1_011111010), .b(t1_011111011), .y(t1_01111101));
wire t1_011111010, t1_011111011;
mixer mix_t1_0111111 (.a(t1_01111110), .b(t1_01111111), .y(t1_0111111));
wire t1_01111110, t1_01111111;
mixer mix_t1_01111110 (.a(t1_011111100), .b(t1_011111101), .y(t1_01111110));
wire t1_011111100, t1_011111101;
mixer mix_t1_01111111 (.a(t1_011111110), .b(t1_011111111), .y(t1_01111111));
wire t1_011111110, t1_011111111;
mixer mix_t2_0 (.a(t2_00), .b(t2_01), .y(t2_0));
wire t2_00, t2_01;
mixer mix_t2_00 (.a(t2_000), .b(t2_001), .y(t2_00));
wire t2_000, t2_001;
mixer mix_t2_000 (.a(t2_0000), .b(t2_0001), .y(t2_000));
wire t2_0000, t2_0001;
mixer mix_t2_0000 (.a(t2_00000), .b(t2_00001), .y(t2_0000));
wire t2_00000, t2_00001;
mixer mix_t2_00000 (.a(t2_000000), .b(t2_000001), .y(t2_00000));
wire t2_000000, t2_000001;
mixer mix_t2_000000 (.a(t2_0000000), .b(t2_0000001), .y(t2_000000));
wire t2_0000000, t2_0000001;
mixer mix_t2_0000000 (.a(t2_00000000), .b(t2_00000001), .y(t2_0000000));
wire t2_00000000, t2_00000001;
mixer mix_t2_00000000 (.a(t2_000000000), .b(t2_000000001), .y(t2_00000000));
wire t2_000000000, t2_000000001;
mixer mix_t2_00000001 (.a(t2_000000010), .b(t2_000000011), .y(t2_00000001));
wire t2_000000010, t2_000000011;
mixer mix_t2_0000001 (.a(t2_00000010), .b(t2_00000011), .y(t2_0000001));
wire t2_00000010, t2_00000011;
mixer mix_t2_00000010 (.a(t2_000000100), .b(t2_000000101), .y(t2_00000010));
wire t2_000000100, t2_000000101;
mixer mix_t2_00000011 (.a(t2_000000110), .b(t2_000000111), .y(t2_00000011));
wire t2_000000110, t2_000000111;
mixer mix_t2_000001 (.a(t2_0000010), .b(t2_0000011), .y(t2_000001));
wire t2_0000010, t2_0000011;
mixer mix_t2_0000010 (.a(t2_00000100), .b(t2_00000101), .y(t2_0000010));
wire t2_00000100, t2_00000101;
mixer mix_t2_00000100 (.a(t2_000001000), .b(t2_000001001), .y(t2_00000100));
wire t2_000001000, t2_000001001;
mixer mix_t2_00000101 (.a(t2_000001010), .b(t2_000001011), .y(t2_00000101));
wire t2_000001010, t2_000001011;
mixer mix_t2_0000011 (.a(t2_00000110), .b(t2_00000111), .y(t2_0000011));
wire t2_00000110, t2_00000111;
mixer mix_t2_00000110 (.a(t2_000001100), .b(t2_000001101), .y(t2_00000110));
wire t2_000001100, t2_000001101;
mixer mix_t2_00000111 (.a(t2_000001110), .b(t2_000001111), .y(t2_00000111));
wire t2_000001110, t2_000001111;
mixer mix_t2_00001 (.a(t2_000010), .b(t2_000011), .y(t2_00001));
wire t2_000010, t2_000011;
mixer mix_t2_000010 (.a(t2_0000100), .b(t2_0000101), .y(t2_000010));
wire t2_0000100, t2_0000101;
mixer mix_t2_0000100 (.a(t2_00001000), .b(t2_00001001), .y(t2_0000100));
wire t2_00001000, t2_00001001;
mixer mix_t2_00001000 (.a(t2_000010000), .b(t2_000010001), .y(t2_00001000));
wire t2_000010000, t2_000010001;
mixer mix_t2_00001001 (.a(t2_000010010), .b(t2_000010011), .y(t2_00001001));
wire t2_000010010, t2_000010011;
mixer mix_t2_0000101 (.a(t2_00001010), .b(t2_00001011), .y(t2_0000101));
wire t2_00001010, t2_00001011;
mixer mix_t2_00001010 (.a(t2_000010100), .b(t2_000010101), .y(t2_00001010));
wire t2_000010100, t2_000010101;
mixer mix_t2_00001011 (.a(t2_000010110), .b(t2_000010111), .y(t2_00001011));
wire t2_000010110, t2_000010111;
mixer mix_t2_000011 (.a(t2_0000110), .b(t2_0000111), .y(t2_000011));
wire t2_0000110, t2_0000111;
mixer mix_t2_0000110 (.a(t2_00001100), .b(t2_00001101), .y(t2_0000110));
wire t2_00001100, t2_00001101;
mixer mix_t2_00001100 (.a(t2_000011000), .b(t2_000011001), .y(t2_00001100));
wire t2_000011000, t2_000011001;
mixer mix_t2_00001101 (.a(t2_000011010), .b(t2_000011011), .y(t2_00001101));
wire t2_000011010, t2_000011011;
mixer mix_t2_0000111 (.a(t2_00001110), .b(t2_00001111), .y(t2_0000111));
wire t2_00001110, t2_00001111;
mixer mix_t2_00001110 (.a(t2_000011100), .b(t2_000011101), .y(t2_00001110));
wire t2_000011100, t2_000011101;
mixer mix_t2_00001111 (.a(t2_000011110), .b(t2_000011111), .y(t2_00001111));
wire t2_000011110, t2_000011111;
mixer mix_t2_0001 (.a(t2_00010), .b(t2_00011), .y(t2_0001));
wire t2_00010, t2_00011;
mixer mix_t2_00010 (.a(t2_000100), .b(t2_000101), .y(t2_00010));
wire t2_000100, t2_000101;
mixer mix_t2_000100 (.a(t2_0001000), .b(t2_0001001), .y(t2_000100));
wire t2_0001000, t2_0001001;
mixer mix_t2_0001000 (.a(t2_00010000), .b(t2_00010001), .y(t2_0001000));
wire t2_00010000, t2_00010001;
mixer mix_t2_00010000 (.a(t2_000100000), .b(t2_000100001), .y(t2_00010000));
wire t2_000100000, t2_000100001;
mixer mix_t2_00010001 (.a(t2_000100010), .b(t2_000100011), .y(t2_00010001));
wire t2_000100010, t2_000100011;
mixer mix_t2_0001001 (.a(t2_00010010), .b(t2_00010011), .y(t2_0001001));
wire t2_00010010, t2_00010011;
mixer mix_t2_00010010 (.a(t2_000100100), .b(t2_000100101), .y(t2_00010010));
wire t2_000100100, t2_000100101;
mixer mix_t2_00010011 (.a(t2_000100110), .b(t2_000100111), .y(t2_00010011));
wire t2_000100110, t2_000100111;
mixer mix_t2_000101 (.a(t2_0001010), .b(t2_0001011), .y(t2_000101));
wire t2_0001010, t2_0001011;
mixer mix_t2_0001010 (.a(t2_00010100), .b(t2_00010101), .y(t2_0001010));
wire t2_00010100, t2_00010101;
mixer mix_t2_00010100 (.a(t2_000101000), .b(t2_000101001), .y(t2_00010100));
wire t2_000101000, t2_000101001;
mixer mix_t2_00010101 (.a(t2_000101010), .b(t2_000101011), .y(t2_00010101));
wire t2_000101010, t2_000101011;
mixer mix_t2_0001011 (.a(t2_00010110), .b(t2_00010111), .y(t2_0001011));
wire t2_00010110, t2_00010111;
mixer mix_t2_00010110 (.a(t2_000101100), .b(t2_000101101), .y(t2_00010110));
wire t2_000101100, t2_000101101;
mixer mix_t2_00010111 (.a(t2_000101110), .b(t2_000101111), .y(t2_00010111));
wire t2_000101110, t2_000101111;
mixer mix_t2_00011 (.a(t2_000110), .b(t2_000111), .y(t2_00011));
wire t2_000110, t2_000111;
mixer mix_t2_000110 (.a(t2_0001100), .b(t2_0001101), .y(t2_000110));
wire t2_0001100, t2_0001101;
mixer mix_t2_0001100 (.a(t2_00011000), .b(t2_00011001), .y(t2_0001100));
wire t2_00011000, t2_00011001;
mixer mix_t2_00011000 (.a(t2_000110000), .b(t2_000110001), .y(t2_00011000));
wire t2_000110000, t2_000110001;
mixer mix_t2_00011001 (.a(t2_000110010), .b(t2_000110011), .y(t2_00011001));
wire t2_000110010, t2_000110011;
mixer mix_t2_0001101 (.a(t2_00011010), .b(t2_00011011), .y(t2_0001101));
wire t2_00011010, t2_00011011;
mixer mix_t2_00011010 (.a(t2_000110100), .b(t2_000110101), .y(t2_00011010));
wire t2_000110100, t2_000110101;
mixer mix_t2_00011011 (.a(t2_000110110), .b(t2_000110111), .y(t2_00011011));
wire t2_000110110, t2_000110111;
mixer mix_t2_000111 (.a(t2_0001110), .b(t2_0001111), .y(t2_000111));
wire t2_0001110, t2_0001111;
mixer mix_t2_0001110 (.a(t2_00011100), .b(t2_00011101), .y(t2_0001110));
wire t2_00011100, t2_00011101;
mixer mix_t2_00011100 (.a(t2_000111000), .b(t2_000111001), .y(t2_00011100));
wire t2_000111000, t2_000111001;
mixer mix_t2_00011101 (.a(t2_000111010), .b(t2_000111011), .y(t2_00011101));
wire t2_000111010, t2_000111011;
mixer mix_t2_0001111 (.a(t2_00011110), .b(t2_00011111), .y(t2_0001111));
wire t2_00011110, t2_00011111;
mixer mix_t2_00011110 (.a(t2_000111100), .b(t2_000111101), .y(t2_00011110));
wire t2_000111100, t2_000111101;
mixer mix_t2_00011111 (.a(t2_000111110), .b(t2_000111111), .y(t2_00011111));
wire t2_000111110, t2_000111111;
mixer mix_t2_001 (.a(t2_0010), .b(t2_0011), .y(t2_001));
wire t2_0010, t2_0011;
mixer mix_t2_0010 (.a(t2_00100), .b(t2_00101), .y(t2_0010));
wire t2_00100, t2_00101;
mixer mix_t2_00100 (.a(t2_001000), .b(t2_001001), .y(t2_00100));
wire t2_001000, t2_001001;
mixer mix_t2_001000 (.a(t2_0010000), .b(t2_0010001), .y(t2_001000));
wire t2_0010000, t2_0010001;
mixer mix_t2_0010000 (.a(t2_00100000), .b(t2_00100001), .y(t2_0010000));
wire t2_00100000, t2_00100001;
mixer mix_t2_00100000 (.a(t2_001000000), .b(t2_001000001), .y(t2_00100000));
wire t2_001000000, t2_001000001;
mixer mix_t2_00100001 (.a(t2_001000010), .b(t2_001000011), .y(t2_00100001));
wire t2_001000010, t2_001000011;
mixer mix_t2_0010001 (.a(t2_00100010), .b(t2_00100011), .y(t2_0010001));
wire t2_00100010, t2_00100011;
mixer mix_t2_00100010 (.a(t2_001000100), .b(t2_001000101), .y(t2_00100010));
wire t2_001000100, t2_001000101;
mixer mix_t2_00100011 (.a(t2_001000110), .b(t2_001000111), .y(t2_00100011));
wire t2_001000110, t2_001000111;
mixer mix_t2_001001 (.a(t2_0010010), .b(t2_0010011), .y(t2_001001));
wire t2_0010010, t2_0010011;
mixer mix_t2_0010010 (.a(t2_00100100), .b(t2_00100101), .y(t2_0010010));
wire t2_00100100, t2_00100101;
mixer mix_t2_00100100 (.a(t2_001001000), .b(t2_001001001), .y(t2_00100100));
wire t2_001001000, t2_001001001;
mixer mix_t2_00100101 (.a(t2_001001010), .b(t2_001001011), .y(t2_00100101));
wire t2_001001010, t2_001001011;
mixer mix_t2_0010011 (.a(t2_00100110), .b(t2_00100111), .y(t2_0010011));
wire t2_00100110, t2_00100111;
mixer mix_t2_00100110 (.a(t2_001001100), .b(t2_001001101), .y(t2_00100110));
wire t2_001001100, t2_001001101;
mixer mix_t2_00100111 (.a(t2_001001110), .b(t2_001001111), .y(t2_00100111));
wire t2_001001110, t2_001001111;
mixer mix_t2_00101 (.a(t2_001010), .b(t2_001011), .y(t2_00101));
wire t2_001010, t2_001011;
mixer mix_t2_001010 (.a(t2_0010100), .b(t2_0010101), .y(t2_001010));
wire t2_0010100, t2_0010101;
mixer mix_t2_0010100 (.a(t2_00101000), .b(t2_00101001), .y(t2_0010100));
wire t2_00101000, t2_00101001;
mixer mix_t2_00101000 (.a(t2_001010000), .b(t2_001010001), .y(t2_00101000));
wire t2_001010000, t2_001010001;
mixer mix_t2_00101001 (.a(t2_001010010), .b(t2_001010011), .y(t2_00101001));
wire t2_001010010, t2_001010011;
mixer mix_t2_0010101 (.a(t2_00101010), .b(t2_00101011), .y(t2_0010101));
wire t2_00101010, t2_00101011;
mixer mix_t2_00101010 (.a(t2_001010100), .b(t2_001010101), .y(t2_00101010));
wire t2_001010100, t2_001010101;
mixer mix_t2_00101011 (.a(t2_001010110), .b(t2_001010111), .y(t2_00101011));
wire t2_001010110, t2_001010111;
mixer mix_t2_001011 (.a(t2_0010110), .b(t2_0010111), .y(t2_001011));
wire t2_0010110, t2_0010111;
mixer mix_t2_0010110 (.a(t2_00101100), .b(t2_00101101), .y(t2_0010110));
wire t2_00101100, t2_00101101;
mixer mix_t2_00101100 (.a(t2_001011000), .b(t2_001011001), .y(t2_00101100));
wire t2_001011000, t2_001011001;
mixer mix_t2_00101101 (.a(t2_001011010), .b(t2_001011011), .y(t2_00101101));
wire t2_001011010, t2_001011011;
mixer mix_t2_0010111 (.a(t2_00101110), .b(t2_00101111), .y(t2_0010111));
wire t2_00101110, t2_00101111;
mixer mix_t2_00101110 (.a(t2_001011100), .b(t2_001011101), .y(t2_00101110));
wire t2_001011100, t2_001011101;
mixer mix_t2_00101111 (.a(t2_001011110), .b(t2_001011111), .y(t2_00101111));
wire t2_001011110, t2_001011111;
mixer mix_t2_0011 (.a(t2_00110), .b(t2_00111), .y(t2_0011));
wire t2_00110, t2_00111;
mixer mix_t2_00110 (.a(t2_001100), .b(t2_001101), .y(t2_00110));
wire t2_001100, t2_001101;
mixer mix_t2_001100 (.a(t2_0011000), .b(t2_0011001), .y(t2_001100));
wire t2_0011000, t2_0011001;
mixer mix_t2_0011000 (.a(t2_00110000), .b(t2_00110001), .y(t2_0011000));
wire t2_00110000, t2_00110001;
mixer mix_t2_00110000 (.a(t2_001100000), .b(t2_001100001), .y(t2_00110000));
wire t2_001100000, t2_001100001;
mixer mix_t2_00110001 (.a(t2_001100010), .b(t2_001100011), .y(t2_00110001));
wire t2_001100010, t2_001100011;
mixer mix_t2_0011001 (.a(t2_00110010), .b(t2_00110011), .y(t2_0011001));
wire t2_00110010, t2_00110011;
mixer mix_t2_00110010 (.a(t2_001100100), .b(t2_001100101), .y(t2_00110010));
wire t2_001100100, t2_001100101;
mixer mix_t2_00110011 (.a(t2_001100110), .b(t2_001100111), .y(t2_00110011));
wire t2_001100110, t2_001100111;
mixer mix_t2_001101 (.a(t2_0011010), .b(t2_0011011), .y(t2_001101));
wire t2_0011010, t2_0011011;
mixer mix_t2_0011010 (.a(t2_00110100), .b(t2_00110101), .y(t2_0011010));
wire t2_00110100, t2_00110101;
mixer mix_t2_00110100 (.a(t2_001101000), .b(t2_001101001), .y(t2_00110100));
wire t2_001101000, t2_001101001;
mixer mix_t2_00110101 (.a(t2_001101010), .b(t2_001101011), .y(t2_00110101));
wire t2_001101010, t2_001101011;
mixer mix_t2_0011011 (.a(t2_00110110), .b(t2_00110111), .y(t2_0011011));
wire t2_00110110, t2_00110111;
mixer mix_t2_00110110 (.a(t2_001101100), .b(t2_001101101), .y(t2_00110110));
wire t2_001101100, t2_001101101;
mixer mix_t2_00110111 (.a(t2_001101110), .b(t2_001101111), .y(t2_00110111));
wire t2_001101110, t2_001101111;
mixer mix_t2_00111 (.a(t2_001110), .b(t2_001111), .y(t2_00111));
wire t2_001110, t2_001111;
mixer mix_t2_001110 (.a(t2_0011100), .b(t2_0011101), .y(t2_001110));
wire t2_0011100, t2_0011101;
mixer mix_t2_0011100 (.a(t2_00111000), .b(t2_00111001), .y(t2_0011100));
wire t2_00111000, t2_00111001;
mixer mix_t2_00111000 (.a(t2_001110000), .b(t2_001110001), .y(t2_00111000));
wire t2_001110000, t2_001110001;
mixer mix_t2_00111001 (.a(t2_001110010), .b(t2_001110011), .y(t2_00111001));
wire t2_001110010, t2_001110011;
mixer mix_t2_0011101 (.a(t2_00111010), .b(t2_00111011), .y(t2_0011101));
wire t2_00111010, t2_00111011;
mixer mix_t2_00111010 (.a(t2_001110100), .b(t2_001110101), .y(t2_00111010));
wire t2_001110100, t2_001110101;
mixer mix_t2_00111011 (.a(t2_001110110), .b(t2_001110111), .y(t2_00111011));
wire t2_001110110, t2_001110111;
mixer mix_t2_001111 (.a(t2_0011110), .b(t2_0011111), .y(t2_001111));
wire t2_0011110, t2_0011111;
mixer mix_t2_0011110 (.a(t2_00111100), .b(t2_00111101), .y(t2_0011110));
wire t2_00111100, t2_00111101;
mixer mix_t2_00111100 (.a(t2_001111000), .b(t2_001111001), .y(t2_00111100));
wire t2_001111000, t2_001111001;
mixer mix_t2_00111101 (.a(t2_001111010), .b(t2_001111011), .y(t2_00111101));
wire t2_001111010, t2_001111011;
mixer mix_t2_0011111 (.a(t2_00111110), .b(t2_00111111), .y(t2_0011111));
wire t2_00111110, t2_00111111;
mixer mix_t2_00111110 (.a(t2_001111100), .b(t2_001111101), .y(t2_00111110));
wire t2_001111100, t2_001111101;
mixer mix_t2_00111111 (.a(t2_001111110), .b(t2_001111111), .y(t2_00111111));
wire t2_001111110, t2_001111111;
mixer mix_t2_01 (.a(t2_010), .b(t2_011), .y(t2_01));
wire t2_010, t2_011;
mixer mix_t2_010 (.a(t2_0100), .b(t2_0101), .y(t2_010));
wire t2_0100, t2_0101;
mixer mix_t2_0100 (.a(t2_01000), .b(t2_01001), .y(t2_0100));
wire t2_01000, t2_01001;
mixer mix_t2_01000 (.a(t2_010000), .b(t2_010001), .y(t2_01000));
wire t2_010000, t2_010001;
mixer mix_t2_010000 (.a(t2_0100000), .b(t2_0100001), .y(t2_010000));
wire t2_0100000, t2_0100001;
mixer mix_t2_0100000 (.a(t2_01000000), .b(t2_01000001), .y(t2_0100000));
wire t2_01000000, t2_01000001;
mixer mix_t2_01000000 (.a(t2_010000000), .b(t2_010000001), .y(t2_01000000));
wire t2_010000000, t2_010000001;
mixer mix_t2_01000001 (.a(t2_010000010), .b(t2_010000011), .y(t2_01000001));
wire t2_010000010, t2_010000011;
mixer mix_t2_0100001 (.a(t2_01000010), .b(t2_01000011), .y(t2_0100001));
wire t2_01000010, t2_01000011;
mixer mix_t2_01000010 (.a(t2_010000100), .b(t2_010000101), .y(t2_01000010));
wire t2_010000100, t2_010000101;
mixer mix_t2_01000011 (.a(t2_010000110), .b(t2_010000111), .y(t2_01000011));
wire t2_010000110, t2_010000111;
mixer mix_t2_010001 (.a(t2_0100010), .b(t2_0100011), .y(t2_010001));
wire t2_0100010, t2_0100011;
mixer mix_t2_0100010 (.a(t2_01000100), .b(t2_01000101), .y(t2_0100010));
wire t2_01000100, t2_01000101;
mixer mix_t2_01000100 (.a(t2_010001000), .b(t2_010001001), .y(t2_01000100));
wire t2_010001000, t2_010001001;
mixer mix_t2_01000101 (.a(t2_010001010), .b(t2_010001011), .y(t2_01000101));
wire t2_010001010, t2_010001011;
mixer mix_t2_0100011 (.a(t2_01000110), .b(t2_01000111), .y(t2_0100011));
wire t2_01000110, t2_01000111;
mixer mix_t2_01000110 (.a(t2_010001100), .b(t2_010001101), .y(t2_01000110));
wire t2_010001100, t2_010001101;
mixer mix_t2_01000111 (.a(t2_010001110), .b(t2_010001111), .y(t2_01000111));
wire t2_010001110, t2_010001111;
mixer mix_t2_01001 (.a(t2_010010), .b(t2_010011), .y(t2_01001));
wire t2_010010, t2_010011;
mixer mix_t2_010010 (.a(t2_0100100), .b(t2_0100101), .y(t2_010010));
wire t2_0100100, t2_0100101;
mixer mix_t2_0100100 (.a(t2_01001000), .b(t2_01001001), .y(t2_0100100));
wire t2_01001000, t2_01001001;
mixer mix_t2_01001000 (.a(t2_010010000), .b(t2_010010001), .y(t2_01001000));
wire t2_010010000, t2_010010001;
mixer mix_t2_01001001 (.a(t2_010010010), .b(t2_010010011), .y(t2_01001001));
wire t2_010010010, t2_010010011;
mixer mix_t2_0100101 (.a(t2_01001010), .b(t2_01001011), .y(t2_0100101));
wire t2_01001010, t2_01001011;
mixer mix_t2_01001010 (.a(t2_010010100), .b(t2_010010101), .y(t2_01001010));
wire t2_010010100, t2_010010101;
mixer mix_t2_01001011 (.a(t2_010010110), .b(t2_010010111), .y(t2_01001011));
wire t2_010010110, t2_010010111;
mixer mix_t2_010011 (.a(t2_0100110), .b(t2_0100111), .y(t2_010011));
wire t2_0100110, t2_0100111;
mixer mix_t2_0100110 (.a(t2_01001100), .b(t2_01001101), .y(t2_0100110));
wire t2_01001100, t2_01001101;
mixer mix_t2_01001100 (.a(t2_010011000), .b(t2_010011001), .y(t2_01001100));
wire t2_010011000, t2_010011001;
mixer mix_t2_01001101 (.a(t2_010011010), .b(t2_010011011), .y(t2_01001101));
wire t2_010011010, t2_010011011;
mixer mix_t2_0100111 (.a(t2_01001110), .b(t2_01001111), .y(t2_0100111));
wire t2_01001110, t2_01001111;
mixer mix_t2_01001110 (.a(t2_010011100), .b(t2_010011101), .y(t2_01001110));
wire t2_010011100, t2_010011101;
mixer mix_t2_01001111 (.a(t2_010011110), .b(t2_010011111), .y(t2_01001111));
wire t2_010011110, t2_010011111;
mixer mix_t2_0101 (.a(t2_01010), .b(t2_01011), .y(t2_0101));
wire t2_01010, t2_01011;
mixer mix_t2_01010 (.a(t2_010100), .b(t2_010101), .y(t2_01010));
wire t2_010100, t2_010101;
mixer mix_t2_010100 (.a(t2_0101000), .b(t2_0101001), .y(t2_010100));
wire t2_0101000, t2_0101001;
mixer mix_t2_0101000 (.a(t2_01010000), .b(t2_01010001), .y(t2_0101000));
wire t2_01010000, t2_01010001;
mixer mix_t2_01010000 (.a(t2_010100000), .b(t2_010100001), .y(t2_01010000));
wire t2_010100000, t2_010100001;
mixer mix_t2_01010001 (.a(t2_010100010), .b(t2_010100011), .y(t2_01010001));
wire t2_010100010, t2_010100011;
mixer mix_t2_0101001 (.a(t2_01010010), .b(t2_01010011), .y(t2_0101001));
wire t2_01010010, t2_01010011;
mixer mix_t2_01010010 (.a(t2_010100100), .b(t2_010100101), .y(t2_01010010));
wire t2_010100100, t2_010100101;
mixer mix_t2_01010011 (.a(t2_010100110), .b(t2_010100111), .y(t2_01010011));
wire t2_010100110, t2_010100111;
mixer mix_t2_010101 (.a(t2_0101010), .b(t2_0101011), .y(t2_010101));
wire t2_0101010, t2_0101011;
mixer mix_t2_0101010 (.a(t2_01010100), .b(t2_01010101), .y(t2_0101010));
wire t2_01010100, t2_01010101;
mixer mix_t2_01010100 (.a(t2_010101000), .b(t2_010101001), .y(t2_01010100));
wire t2_010101000, t2_010101001;
mixer mix_t2_01010101 (.a(t2_010101010), .b(t2_010101011), .y(t2_01010101));
wire t2_010101010, t2_010101011;
mixer mix_t2_0101011 (.a(t2_01010110), .b(t2_01010111), .y(t2_0101011));
wire t2_01010110, t2_01010111;
mixer mix_t2_01010110 (.a(t2_010101100), .b(t2_010101101), .y(t2_01010110));
wire t2_010101100, t2_010101101;
mixer mix_t2_01010111 (.a(t2_010101110), .b(t2_010101111), .y(t2_01010111));
wire t2_010101110, t2_010101111;
mixer mix_t2_01011 (.a(t2_010110), .b(t2_010111), .y(t2_01011));
wire t2_010110, t2_010111;
mixer mix_t2_010110 (.a(t2_0101100), .b(t2_0101101), .y(t2_010110));
wire t2_0101100, t2_0101101;
mixer mix_t2_0101100 (.a(t2_01011000), .b(t2_01011001), .y(t2_0101100));
wire t2_01011000, t2_01011001;
mixer mix_t2_01011000 (.a(t2_010110000), .b(t2_010110001), .y(t2_01011000));
wire t2_010110000, t2_010110001;
mixer mix_t2_01011001 (.a(t2_010110010), .b(t2_010110011), .y(t2_01011001));
wire t2_010110010, t2_010110011;
mixer mix_t2_0101101 (.a(t2_01011010), .b(t2_01011011), .y(t2_0101101));
wire t2_01011010, t2_01011011;
mixer mix_t2_01011010 (.a(t2_010110100), .b(t2_010110101), .y(t2_01011010));
wire t2_010110100, t2_010110101;
mixer mix_t2_01011011 (.a(t2_010110110), .b(t2_010110111), .y(t2_01011011));
wire t2_010110110, t2_010110111;
mixer mix_t2_010111 (.a(t2_0101110), .b(t2_0101111), .y(t2_010111));
wire t2_0101110, t2_0101111;
mixer mix_t2_0101110 (.a(t2_01011100), .b(t2_01011101), .y(t2_0101110));
wire t2_01011100, t2_01011101;
mixer mix_t2_01011100 (.a(t2_010111000), .b(t2_010111001), .y(t2_01011100));
wire t2_010111000, t2_010111001;
mixer mix_t2_01011101 (.a(t2_010111010), .b(t2_010111011), .y(t2_01011101));
wire t2_010111010, t2_010111011;
mixer mix_t2_0101111 (.a(t2_01011110), .b(t2_01011111), .y(t2_0101111));
wire t2_01011110, t2_01011111;
mixer mix_t2_01011110 (.a(t2_010111100), .b(t2_010111101), .y(t2_01011110));
wire t2_010111100, t2_010111101;
mixer mix_t2_01011111 (.a(t2_010111110), .b(t2_010111111), .y(t2_01011111));
wire t2_010111110, t2_010111111;
mixer mix_t2_011 (.a(t2_0110), .b(t2_0111), .y(t2_011));
wire t2_0110, t2_0111;
mixer mix_t2_0110 (.a(t2_01100), .b(t2_01101), .y(t2_0110));
wire t2_01100, t2_01101;
mixer mix_t2_01100 (.a(t2_011000), .b(t2_011001), .y(t2_01100));
wire t2_011000, t2_011001;
mixer mix_t2_011000 (.a(t2_0110000), .b(t2_0110001), .y(t2_011000));
wire t2_0110000, t2_0110001;
mixer mix_t2_0110000 (.a(t2_01100000), .b(t2_01100001), .y(t2_0110000));
wire t2_01100000, t2_01100001;
mixer mix_t2_01100000 (.a(t2_011000000), .b(t2_011000001), .y(t2_01100000));
wire t2_011000000, t2_011000001;
mixer mix_t2_01100001 (.a(t2_011000010), .b(t2_011000011), .y(t2_01100001));
wire t2_011000010, t2_011000011;
mixer mix_t2_0110001 (.a(t2_01100010), .b(t2_01100011), .y(t2_0110001));
wire t2_01100010, t2_01100011;
mixer mix_t2_01100010 (.a(t2_011000100), .b(t2_011000101), .y(t2_01100010));
wire t2_011000100, t2_011000101;
mixer mix_t2_01100011 (.a(t2_011000110), .b(t2_011000111), .y(t2_01100011));
wire t2_011000110, t2_011000111;
mixer mix_t2_011001 (.a(t2_0110010), .b(t2_0110011), .y(t2_011001));
wire t2_0110010, t2_0110011;
mixer mix_t2_0110010 (.a(t2_01100100), .b(t2_01100101), .y(t2_0110010));
wire t2_01100100, t2_01100101;
mixer mix_t2_01100100 (.a(t2_011001000), .b(t2_011001001), .y(t2_01100100));
wire t2_011001000, t2_011001001;
mixer mix_t2_01100101 (.a(t2_011001010), .b(t2_011001011), .y(t2_01100101));
wire t2_011001010, t2_011001011;
mixer mix_t2_0110011 (.a(t2_01100110), .b(t2_01100111), .y(t2_0110011));
wire t2_01100110, t2_01100111;
mixer mix_t2_01100110 (.a(t2_011001100), .b(t2_011001101), .y(t2_01100110));
wire t2_011001100, t2_011001101;
mixer mix_t2_01100111 (.a(t2_011001110), .b(t2_011001111), .y(t2_01100111));
wire t2_011001110, t2_011001111;
mixer mix_t2_01101 (.a(t2_011010), .b(t2_011011), .y(t2_01101));
wire t2_011010, t2_011011;
mixer mix_t2_011010 (.a(t2_0110100), .b(t2_0110101), .y(t2_011010));
wire t2_0110100, t2_0110101;
mixer mix_t2_0110100 (.a(t2_01101000), .b(t2_01101001), .y(t2_0110100));
wire t2_01101000, t2_01101001;
mixer mix_t2_01101000 (.a(t2_011010000), .b(t2_011010001), .y(t2_01101000));
wire t2_011010000, t2_011010001;
mixer mix_t2_01101001 (.a(t2_011010010), .b(t2_011010011), .y(t2_01101001));
wire t2_011010010, t2_011010011;
mixer mix_t2_0110101 (.a(t2_01101010), .b(t2_01101011), .y(t2_0110101));
wire t2_01101010, t2_01101011;
mixer mix_t2_01101010 (.a(t2_011010100), .b(t2_011010101), .y(t2_01101010));
wire t2_011010100, t2_011010101;
mixer mix_t2_01101011 (.a(t2_011010110), .b(t2_011010111), .y(t2_01101011));
wire t2_011010110, t2_011010111;
mixer mix_t2_011011 (.a(t2_0110110), .b(t2_0110111), .y(t2_011011));
wire t2_0110110, t2_0110111;
mixer mix_t2_0110110 (.a(t2_01101100), .b(t2_01101101), .y(t2_0110110));
wire t2_01101100, t2_01101101;
mixer mix_t2_01101100 (.a(t2_011011000), .b(t2_011011001), .y(t2_01101100));
wire t2_011011000, t2_011011001;
mixer mix_t2_01101101 (.a(t2_011011010), .b(t2_011011011), .y(t2_01101101));
wire t2_011011010, t2_011011011;
mixer mix_t2_0110111 (.a(t2_01101110), .b(t2_01101111), .y(t2_0110111));
wire t2_01101110, t2_01101111;
mixer mix_t2_01101110 (.a(t2_011011100), .b(t2_011011101), .y(t2_01101110));
wire t2_011011100, t2_011011101;
mixer mix_t2_01101111 (.a(t2_011011110), .b(t2_011011111), .y(t2_01101111));
wire t2_011011110, t2_011011111;
mixer mix_t2_0111 (.a(t2_01110), .b(t2_01111), .y(t2_0111));
wire t2_01110, t2_01111;
mixer mix_t2_01110 (.a(t2_011100), .b(t2_011101), .y(t2_01110));
wire t2_011100, t2_011101;
mixer mix_t2_011100 (.a(t2_0111000), .b(t2_0111001), .y(t2_011100));
wire t2_0111000, t2_0111001;
mixer mix_t2_0111000 (.a(t2_01110000), .b(t2_01110001), .y(t2_0111000));
wire t2_01110000, t2_01110001;
mixer mix_t2_01110000 (.a(t2_011100000), .b(t2_011100001), .y(t2_01110000));
wire t2_011100000, t2_011100001;
mixer mix_t2_01110001 (.a(t2_011100010), .b(t2_011100011), .y(t2_01110001));
wire t2_011100010, t2_011100011;
mixer mix_t2_0111001 (.a(t2_01110010), .b(t2_01110011), .y(t2_0111001));
wire t2_01110010, t2_01110011;
mixer mix_t2_01110010 (.a(t2_011100100), .b(t2_011100101), .y(t2_01110010));
wire t2_011100100, t2_011100101;
mixer mix_t2_01110011 (.a(t2_011100110), .b(t2_011100111), .y(t2_01110011));
wire t2_011100110, t2_011100111;
mixer mix_t2_011101 (.a(t2_0111010), .b(t2_0111011), .y(t2_011101));
wire t2_0111010, t2_0111011;
mixer mix_t2_0111010 (.a(t2_01110100), .b(t2_01110101), .y(t2_0111010));
wire t2_01110100, t2_01110101;
mixer mix_t2_01110100 (.a(t2_011101000), .b(t2_011101001), .y(t2_01110100));
wire t2_011101000, t2_011101001;
mixer mix_t2_01110101 (.a(t2_011101010), .b(t2_011101011), .y(t2_01110101));
wire t2_011101010, t2_011101011;
mixer mix_t2_0111011 (.a(t2_01110110), .b(t2_01110111), .y(t2_0111011));
wire t2_01110110, t2_01110111;
mixer mix_t2_01110110 (.a(t2_011101100), .b(t2_011101101), .y(t2_01110110));
wire t2_011101100, t2_011101101;
mixer mix_t2_01110111 (.a(t2_011101110), .b(t2_011101111), .y(t2_01110111));
wire t2_011101110, t2_011101111;
mixer mix_t2_01111 (.a(t2_011110), .b(t2_011111), .y(t2_01111));
wire t2_011110, t2_011111;
mixer mix_t2_011110 (.a(t2_0111100), .b(t2_0111101), .y(t2_011110));
wire t2_0111100, t2_0111101;
mixer mix_t2_0111100 (.a(t2_01111000), .b(t2_01111001), .y(t2_0111100));
wire t2_01111000, t2_01111001;
mixer mix_t2_01111000 (.a(t2_011110000), .b(t2_011110001), .y(t2_01111000));
wire t2_011110000, t2_011110001;
mixer mix_t2_01111001 (.a(t2_011110010), .b(t2_011110011), .y(t2_01111001));
wire t2_011110010, t2_011110011;
mixer mix_t2_0111101 (.a(t2_01111010), .b(t2_01111011), .y(t2_0111101));
wire t2_01111010, t2_01111011;
mixer mix_t2_01111010 (.a(t2_011110100), .b(t2_011110101), .y(t2_01111010));
wire t2_011110100, t2_011110101;
mixer mix_t2_01111011 (.a(t2_011110110), .b(t2_011110111), .y(t2_01111011));
wire t2_011110110, t2_011110111;
mixer mix_t2_011111 (.a(t2_0111110), .b(t2_0111111), .y(t2_011111));
wire t2_0111110, t2_0111111;
mixer mix_t2_0111110 (.a(t2_01111100), .b(t2_01111101), .y(t2_0111110));
wire t2_01111100, t2_01111101;
mixer mix_t2_01111100 (.a(t2_011111000), .b(t2_011111001), .y(t2_01111100));
wire t2_011111000, t2_011111001;
mixer mix_t2_01111101 (.a(t2_011111010), .b(t2_011111011), .y(t2_01111101));
wire t2_011111010, t2_011111011;
mixer mix_t2_0111111 (.a(t2_01111110), .b(t2_01111111), .y(t2_0111111));
wire t2_01111110, t2_01111111;
mixer mix_t2_01111110 (.a(t2_011111100), .b(t2_011111101), .y(t2_01111110));
wire t2_011111100, t2_011111101;
mixer mix_t2_01111111 (.a(t2_011111110), .b(t2_011111111), .y(t2_01111111));
wire t2_011111110, t2_011111111;
mixer mix_t3_0 (.a(t3_00), .b(t3_01), .y(t3_0));
wire t3_00, t3_01;
mixer mix_t3_00 (.a(t3_000), .b(t3_001), .y(t3_00));
wire t3_000, t3_001;
mixer mix_t3_000 (.a(t3_0000), .b(t3_0001), .y(t3_000));
wire t3_0000, t3_0001;
mixer mix_t3_0000 (.a(t3_00000), .b(t3_00001), .y(t3_0000));
wire t3_00000, t3_00001;
mixer mix_t3_00000 (.a(t3_000000), .b(t3_000001), .y(t3_00000));
wire t3_000000, t3_000001;
mixer mix_t3_000000 (.a(t3_0000000), .b(t3_0000001), .y(t3_000000));
wire t3_0000000, t3_0000001;
mixer mix_t3_0000000 (.a(t3_00000000), .b(t3_00000001), .y(t3_0000000));
wire t3_00000000, t3_00000001;
mixer mix_t3_00000000 (.a(t3_000000000), .b(t3_000000001), .y(t3_00000000));
wire t3_000000000, t3_000000001;
mixer mix_t3_00000001 (.a(t3_000000010), .b(t3_000000011), .y(t3_00000001));
wire t3_000000010, t3_000000011;
mixer mix_t3_0000001 (.a(t3_00000010), .b(t3_00000011), .y(t3_0000001));
wire t3_00000010, t3_00000011;
mixer mix_t3_00000010 (.a(t3_000000100), .b(t3_000000101), .y(t3_00000010));
wire t3_000000100, t3_000000101;
mixer mix_t3_00000011 (.a(t3_000000110), .b(t3_000000111), .y(t3_00000011));
wire t3_000000110, t3_000000111;
mixer mix_t3_000001 (.a(t3_0000010), .b(t3_0000011), .y(t3_000001));
wire t3_0000010, t3_0000011;
mixer mix_t3_0000010 (.a(t3_00000100), .b(t3_00000101), .y(t3_0000010));
wire t3_00000100, t3_00000101;
mixer mix_t3_00000100 (.a(t3_000001000), .b(t3_000001001), .y(t3_00000100));
wire t3_000001000, t3_000001001;
mixer mix_t3_00000101 (.a(t3_000001010), .b(t3_000001011), .y(t3_00000101));
wire t3_000001010, t3_000001011;
mixer mix_t3_0000011 (.a(t3_00000110), .b(t3_00000111), .y(t3_0000011));
wire t3_00000110, t3_00000111;
mixer mix_t3_00000110 (.a(t3_000001100), .b(t3_000001101), .y(t3_00000110));
wire t3_000001100, t3_000001101;
mixer mix_t3_00000111 (.a(t3_000001110), .b(t3_000001111), .y(t3_00000111));
wire t3_000001110, t3_000001111;
mixer mix_t3_00001 (.a(t3_000010), .b(t3_000011), .y(t3_00001));
wire t3_000010, t3_000011;
mixer mix_t3_000010 (.a(t3_0000100), .b(t3_0000101), .y(t3_000010));
wire t3_0000100, t3_0000101;
mixer mix_t3_0000100 (.a(t3_00001000), .b(t3_00001001), .y(t3_0000100));
wire t3_00001000, t3_00001001;
mixer mix_t3_00001000 (.a(t3_000010000), .b(t3_000010001), .y(t3_00001000));
wire t3_000010000, t3_000010001;
mixer mix_t3_00001001 (.a(t3_000010010), .b(t3_000010011), .y(t3_00001001));
wire t3_000010010, t3_000010011;
mixer mix_t3_0000101 (.a(t3_00001010), .b(t3_00001011), .y(t3_0000101));
wire t3_00001010, t3_00001011;
mixer mix_t3_00001010 (.a(t3_000010100), .b(t3_000010101), .y(t3_00001010));
wire t3_000010100, t3_000010101;
mixer mix_t3_00001011 (.a(t3_000010110), .b(t3_000010111), .y(t3_00001011));
wire t3_000010110, t3_000010111;
mixer mix_t3_000011 (.a(t3_0000110), .b(t3_0000111), .y(t3_000011));
wire t3_0000110, t3_0000111;
mixer mix_t3_0000110 (.a(t3_00001100), .b(t3_00001101), .y(t3_0000110));
wire t3_00001100, t3_00001101;
mixer mix_t3_00001100 (.a(t3_000011000), .b(t3_000011001), .y(t3_00001100));
wire t3_000011000, t3_000011001;
mixer mix_t3_00001101 (.a(t3_000011010), .b(t3_000011011), .y(t3_00001101));
wire t3_000011010, t3_000011011;
mixer mix_t3_0000111 (.a(t3_00001110), .b(t3_00001111), .y(t3_0000111));
wire t3_00001110, t3_00001111;
mixer mix_t3_00001110 (.a(t3_000011100), .b(t3_000011101), .y(t3_00001110));
wire t3_000011100, t3_000011101;
mixer mix_t3_00001111 (.a(t3_000011110), .b(t3_000011111), .y(t3_00001111));
wire t3_000011110, t3_000011111;
mixer mix_t3_0001 (.a(t3_00010), .b(t3_00011), .y(t3_0001));
wire t3_00010, t3_00011;
mixer mix_t3_00010 (.a(t3_000100), .b(t3_000101), .y(t3_00010));
wire t3_000100, t3_000101;
mixer mix_t3_000100 (.a(t3_0001000), .b(t3_0001001), .y(t3_000100));
wire t3_0001000, t3_0001001;
mixer mix_t3_0001000 (.a(t3_00010000), .b(t3_00010001), .y(t3_0001000));
wire t3_00010000, t3_00010001;
mixer mix_t3_00010000 (.a(t3_000100000), .b(t3_000100001), .y(t3_00010000));
wire t3_000100000, t3_000100001;
mixer mix_t3_00010001 (.a(t3_000100010), .b(t3_000100011), .y(t3_00010001));
wire t3_000100010, t3_000100011;
mixer mix_t3_0001001 (.a(t3_00010010), .b(t3_00010011), .y(t3_0001001));
wire t3_00010010, t3_00010011;
mixer mix_t3_00010010 (.a(t3_000100100), .b(t3_000100101), .y(t3_00010010));
wire t3_000100100, t3_000100101;
mixer mix_t3_00010011 (.a(t3_000100110), .b(t3_000100111), .y(t3_00010011));
wire t3_000100110, t3_000100111;
mixer mix_t3_000101 (.a(t3_0001010), .b(t3_0001011), .y(t3_000101));
wire t3_0001010, t3_0001011;
mixer mix_t3_0001010 (.a(t3_00010100), .b(t3_00010101), .y(t3_0001010));
wire t3_00010100, t3_00010101;
mixer mix_t3_00010100 (.a(t3_000101000), .b(t3_000101001), .y(t3_00010100));
wire t3_000101000, t3_000101001;
mixer mix_t3_00010101 (.a(t3_000101010), .b(t3_000101011), .y(t3_00010101));
wire t3_000101010, t3_000101011;
mixer mix_t3_0001011 (.a(t3_00010110), .b(t3_00010111), .y(t3_0001011));
wire t3_00010110, t3_00010111;
mixer mix_t3_00010110 (.a(t3_000101100), .b(t3_000101101), .y(t3_00010110));
wire t3_000101100, t3_000101101;
mixer mix_t3_00010111 (.a(t3_000101110), .b(t3_000101111), .y(t3_00010111));
wire t3_000101110, t3_000101111;
mixer mix_t3_00011 (.a(t3_000110), .b(t3_000111), .y(t3_00011));
wire t3_000110, t3_000111;
mixer mix_t3_000110 (.a(t3_0001100), .b(t3_0001101), .y(t3_000110));
wire t3_0001100, t3_0001101;
mixer mix_t3_0001100 (.a(t3_00011000), .b(t3_00011001), .y(t3_0001100));
wire t3_00011000, t3_00011001;
mixer mix_t3_00011000 (.a(t3_000110000), .b(t3_000110001), .y(t3_00011000));
wire t3_000110000, t3_000110001;
mixer mix_t3_00011001 (.a(t3_000110010), .b(t3_000110011), .y(t3_00011001));
wire t3_000110010, t3_000110011;
mixer mix_t3_0001101 (.a(t3_00011010), .b(t3_00011011), .y(t3_0001101));
wire t3_00011010, t3_00011011;
mixer mix_t3_00011010 (.a(t3_000110100), .b(t3_000110101), .y(t3_00011010));
wire t3_000110100, t3_000110101;
mixer mix_t3_00011011 (.a(t3_000110110), .b(t3_000110111), .y(t3_00011011));
wire t3_000110110, t3_000110111;
mixer mix_t3_000111 (.a(t3_0001110), .b(t3_0001111), .y(t3_000111));
wire t3_0001110, t3_0001111;
mixer mix_t3_0001110 (.a(t3_00011100), .b(t3_00011101), .y(t3_0001110));
wire t3_00011100, t3_00011101;
mixer mix_t3_00011100 (.a(t3_000111000), .b(t3_000111001), .y(t3_00011100));
wire t3_000111000, t3_000111001;
mixer mix_t3_00011101 (.a(t3_000111010), .b(t3_000111011), .y(t3_00011101));
wire t3_000111010, t3_000111011;
mixer mix_t3_0001111 (.a(t3_00011110), .b(t3_00011111), .y(t3_0001111));
wire t3_00011110, t3_00011111;
mixer mix_t3_00011110 (.a(t3_000111100), .b(t3_000111101), .y(t3_00011110));
wire t3_000111100, t3_000111101;
mixer mix_t3_00011111 (.a(t3_000111110), .b(t3_000111111), .y(t3_00011111));
wire t3_000111110, t3_000111111;
mixer mix_t3_001 (.a(t3_0010), .b(t3_0011), .y(t3_001));
wire t3_0010, t3_0011;
mixer mix_t3_0010 (.a(t3_00100), .b(t3_00101), .y(t3_0010));
wire t3_00100, t3_00101;
mixer mix_t3_00100 (.a(t3_001000), .b(t3_001001), .y(t3_00100));
wire t3_001000, t3_001001;
mixer mix_t3_001000 (.a(t3_0010000), .b(t3_0010001), .y(t3_001000));
wire t3_0010000, t3_0010001;
mixer mix_t3_0010000 (.a(t3_00100000), .b(t3_00100001), .y(t3_0010000));
wire t3_00100000, t3_00100001;
mixer mix_t3_00100000 (.a(t3_001000000), .b(t3_001000001), .y(t3_00100000));
wire t3_001000000, t3_001000001;
mixer mix_t3_00100001 (.a(t3_001000010), .b(t3_001000011), .y(t3_00100001));
wire t3_001000010, t3_001000011;
mixer mix_t3_0010001 (.a(t3_00100010), .b(t3_00100011), .y(t3_0010001));
wire t3_00100010, t3_00100011;
mixer mix_t3_00100010 (.a(t3_001000100), .b(t3_001000101), .y(t3_00100010));
wire t3_001000100, t3_001000101;
mixer mix_t3_00100011 (.a(t3_001000110), .b(t3_001000111), .y(t3_00100011));
wire t3_001000110, t3_001000111;
mixer mix_t3_001001 (.a(t3_0010010), .b(t3_0010011), .y(t3_001001));
wire t3_0010010, t3_0010011;
mixer mix_t3_0010010 (.a(t3_00100100), .b(t3_00100101), .y(t3_0010010));
wire t3_00100100, t3_00100101;
mixer mix_t3_00100100 (.a(t3_001001000), .b(t3_001001001), .y(t3_00100100));
wire t3_001001000, t3_001001001;
mixer mix_t3_00100101 (.a(t3_001001010), .b(t3_001001011), .y(t3_00100101));
wire t3_001001010, t3_001001011;
mixer mix_t3_0010011 (.a(t3_00100110), .b(t3_00100111), .y(t3_0010011));
wire t3_00100110, t3_00100111;
mixer mix_t3_00100110 (.a(t3_001001100), .b(t3_001001101), .y(t3_00100110));
wire t3_001001100, t3_001001101;
mixer mix_t3_00100111 (.a(t3_001001110), .b(t3_001001111), .y(t3_00100111));
wire t3_001001110, t3_001001111;
mixer mix_t3_00101 (.a(t3_001010), .b(t3_001011), .y(t3_00101));
wire t3_001010, t3_001011;
mixer mix_t3_001010 (.a(t3_0010100), .b(t3_0010101), .y(t3_001010));
wire t3_0010100, t3_0010101;
mixer mix_t3_0010100 (.a(t3_00101000), .b(t3_00101001), .y(t3_0010100));
wire t3_00101000, t3_00101001;
mixer mix_t3_00101000 (.a(t3_001010000), .b(t3_001010001), .y(t3_00101000));
wire t3_001010000, t3_001010001;
mixer mix_t3_00101001 (.a(t3_001010010), .b(t3_001010011), .y(t3_00101001));
wire t3_001010010, t3_001010011;
mixer mix_t3_0010101 (.a(t3_00101010), .b(t3_00101011), .y(t3_0010101));
wire t3_00101010, t3_00101011;
mixer mix_t3_00101010 (.a(t3_001010100), .b(t3_001010101), .y(t3_00101010));
wire t3_001010100, t3_001010101;
mixer mix_t3_00101011 (.a(t3_001010110), .b(t3_001010111), .y(t3_00101011));
wire t3_001010110, t3_001010111;
mixer mix_t3_001011 (.a(t3_0010110), .b(t3_0010111), .y(t3_001011));
wire t3_0010110, t3_0010111;
mixer mix_t3_0010110 (.a(t3_00101100), .b(t3_00101101), .y(t3_0010110));
wire t3_00101100, t3_00101101;
mixer mix_t3_00101100 (.a(t3_001011000), .b(t3_001011001), .y(t3_00101100));
wire t3_001011000, t3_001011001;
mixer mix_t3_00101101 (.a(t3_001011010), .b(t3_001011011), .y(t3_00101101));
wire t3_001011010, t3_001011011;
mixer mix_t3_0010111 (.a(t3_00101110), .b(t3_00101111), .y(t3_0010111));
wire t3_00101110, t3_00101111;
mixer mix_t3_00101110 (.a(t3_001011100), .b(t3_001011101), .y(t3_00101110));
wire t3_001011100, t3_001011101;
mixer mix_t3_00101111 (.a(t3_001011110), .b(t3_001011111), .y(t3_00101111));
wire t3_001011110, t3_001011111;
mixer mix_t3_0011 (.a(t3_00110), .b(t3_00111), .y(t3_0011));
wire t3_00110, t3_00111;
mixer mix_t3_00110 (.a(t3_001100), .b(t3_001101), .y(t3_00110));
wire t3_001100, t3_001101;
mixer mix_t3_001100 (.a(t3_0011000), .b(t3_0011001), .y(t3_001100));
wire t3_0011000, t3_0011001;
mixer mix_t3_0011000 (.a(t3_00110000), .b(t3_00110001), .y(t3_0011000));
wire t3_00110000, t3_00110001;
mixer mix_t3_00110000 (.a(t3_001100000), .b(t3_001100001), .y(t3_00110000));
wire t3_001100000, t3_001100001;
mixer mix_t3_00110001 (.a(t3_001100010), .b(t3_001100011), .y(t3_00110001));
wire t3_001100010, t3_001100011;
mixer mix_t3_0011001 (.a(t3_00110010), .b(t3_00110011), .y(t3_0011001));
wire t3_00110010, t3_00110011;
mixer mix_t3_00110010 (.a(t3_001100100), .b(t3_001100101), .y(t3_00110010));
wire t3_001100100, t3_001100101;
mixer mix_t3_00110011 (.a(t3_001100110), .b(t3_001100111), .y(t3_00110011));
wire t3_001100110, t3_001100111;
mixer mix_t3_001101 (.a(t3_0011010), .b(t3_0011011), .y(t3_001101));
wire t3_0011010, t3_0011011;
mixer mix_t3_0011010 (.a(t3_00110100), .b(t3_00110101), .y(t3_0011010));
wire t3_00110100, t3_00110101;
mixer mix_t3_00110100 (.a(t3_001101000), .b(t3_001101001), .y(t3_00110100));
wire t3_001101000, t3_001101001;
mixer mix_t3_00110101 (.a(t3_001101010), .b(t3_001101011), .y(t3_00110101));
wire t3_001101010, t3_001101011;
mixer mix_t3_0011011 (.a(t3_00110110), .b(t3_00110111), .y(t3_0011011));
wire t3_00110110, t3_00110111;
mixer mix_t3_00110110 (.a(t3_001101100), .b(t3_001101101), .y(t3_00110110));
wire t3_001101100, t3_001101101;
mixer mix_t3_00110111 (.a(t3_001101110), .b(t3_001101111), .y(t3_00110111));
wire t3_001101110, t3_001101111;
mixer mix_t3_00111 (.a(t3_001110), .b(t3_001111), .y(t3_00111));
wire t3_001110, t3_001111;
mixer mix_t3_001110 (.a(t3_0011100), .b(t3_0011101), .y(t3_001110));
wire t3_0011100, t3_0011101;
mixer mix_t3_0011100 (.a(t3_00111000), .b(t3_00111001), .y(t3_0011100));
wire t3_00111000, t3_00111001;
mixer mix_t3_00111000 (.a(t3_001110000), .b(t3_001110001), .y(t3_00111000));
wire t3_001110000, t3_001110001;
mixer mix_t3_00111001 (.a(t3_001110010), .b(t3_001110011), .y(t3_00111001));
wire t3_001110010, t3_001110011;
mixer mix_t3_0011101 (.a(t3_00111010), .b(t3_00111011), .y(t3_0011101));
wire t3_00111010, t3_00111011;
mixer mix_t3_00111010 (.a(t3_001110100), .b(t3_001110101), .y(t3_00111010));
wire t3_001110100, t3_001110101;
mixer mix_t3_00111011 (.a(t3_001110110), .b(t3_001110111), .y(t3_00111011));
wire t3_001110110, t3_001110111;
mixer mix_t3_001111 (.a(t3_0011110), .b(t3_0011111), .y(t3_001111));
wire t3_0011110, t3_0011111;
mixer mix_t3_0011110 (.a(t3_00111100), .b(t3_00111101), .y(t3_0011110));
wire t3_00111100, t3_00111101;
mixer mix_t3_00111100 (.a(t3_001111000), .b(t3_001111001), .y(t3_00111100));
wire t3_001111000, t3_001111001;
mixer mix_t3_00111101 (.a(t3_001111010), .b(t3_001111011), .y(t3_00111101));
wire t3_001111010, t3_001111011;
mixer mix_t3_0011111 (.a(t3_00111110), .b(t3_00111111), .y(t3_0011111));
wire t3_00111110, t3_00111111;
mixer mix_t3_00111110 (.a(t3_001111100), .b(t3_001111101), .y(t3_00111110));
wire t3_001111100, t3_001111101;
mixer mix_t3_00111111 (.a(t3_001111110), .b(t3_001111111), .y(t3_00111111));
wire t3_001111110, t3_001111111;
mixer mix_t3_01 (.a(t3_010), .b(t3_011), .y(t3_01));
wire t3_010, t3_011;
mixer mix_t3_010 (.a(t3_0100), .b(t3_0101), .y(t3_010));
wire t3_0100, t3_0101;
mixer mix_t3_0100 (.a(t3_01000), .b(t3_01001), .y(t3_0100));
wire t3_01000, t3_01001;
mixer mix_t3_01000 (.a(t3_010000), .b(t3_010001), .y(t3_01000));
wire t3_010000, t3_010001;
mixer mix_t3_010000 (.a(t3_0100000), .b(t3_0100001), .y(t3_010000));
wire t3_0100000, t3_0100001;
mixer mix_t3_0100000 (.a(t3_01000000), .b(t3_01000001), .y(t3_0100000));
wire t3_01000000, t3_01000001;
mixer mix_t3_01000000 (.a(t3_010000000), .b(t3_010000001), .y(t3_01000000));
wire t3_010000000, t3_010000001;
mixer mix_t3_01000001 (.a(t3_010000010), .b(t3_010000011), .y(t3_01000001));
wire t3_010000010, t3_010000011;
mixer mix_t3_0100001 (.a(t3_01000010), .b(t3_01000011), .y(t3_0100001));
wire t3_01000010, t3_01000011;
mixer mix_t3_01000010 (.a(t3_010000100), .b(t3_010000101), .y(t3_01000010));
wire t3_010000100, t3_010000101;
mixer mix_t3_01000011 (.a(t3_010000110), .b(t3_010000111), .y(t3_01000011));
wire t3_010000110, t3_010000111;
mixer mix_t3_010001 (.a(t3_0100010), .b(t3_0100011), .y(t3_010001));
wire t3_0100010, t3_0100011;
mixer mix_t3_0100010 (.a(t3_01000100), .b(t3_01000101), .y(t3_0100010));
wire t3_01000100, t3_01000101;
mixer mix_t3_01000100 (.a(t3_010001000), .b(t3_010001001), .y(t3_01000100));
wire t3_010001000, t3_010001001;
mixer mix_t3_01000101 (.a(t3_010001010), .b(t3_010001011), .y(t3_01000101));
wire t3_010001010, t3_010001011;
mixer mix_t3_0100011 (.a(t3_01000110), .b(t3_01000111), .y(t3_0100011));
wire t3_01000110, t3_01000111;
mixer mix_t3_01000110 (.a(t3_010001100), .b(t3_010001101), .y(t3_01000110));
wire t3_010001100, t3_010001101;
mixer mix_t3_01000111 (.a(t3_010001110), .b(t3_010001111), .y(t3_01000111));
wire t3_010001110, t3_010001111;
mixer mix_t3_01001 (.a(t3_010010), .b(t3_010011), .y(t3_01001));
wire t3_010010, t3_010011;
mixer mix_t3_010010 (.a(t3_0100100), .b(t3_0100101), .y(t3_010010));
wire t3_0100100, t3_0100101;
mixer mix_t3_0100100 (.a(t3_01001000), .b(t3_01001001), .y(t3_0100100));
wire t3_01001000, t3_01001001;
mixer mix_t3_01001000 (.a(t3_010010000), .b(t3_010010001), .y(t3_01001000));
wire t3_010010000, t3_010010001;
mixer mix_t3_01001001 (.a(t3_010010010), .b(t3_010010011), .y(t3_01001001));
wire t3_010010010, t3_010010011;
mixer mix_t3_0100101 (.a(t3_01001010), .b(t3_01001011), .y(t3_0100101));
wire t3_01001010, t3_01001011;
mixer mix_t3_01001010 (.a(t3_010010100), .b(t3_010010101), .y(t3_01001010));
wire t3_010010100, t3_010010101;
mixer mix_t3_01001011 (.a(t3_010010110), .b(t3_010010111), .y(t3_01001011));
wire t3_010010110, t3_010010111;
mixer mix_t3_010011 (.a(t3_0100110), .b(t3_0100111), .y(t3_010011));
wire t3_0100110, t3_0100111;
mixer mix_t3_0100110 (.a(t3_01001100), .b(t3_01001101), .y(t3_0100110));
wire t3_01001100, t3_01001101;
mixer mix_t3_01001100 (.a(t3_010011000), .b(t3_010011001), .y(t3_01001100));
wire t3_010011000, t3_010011001;
mixer mix_t3_01001101 (.a(t3_010011010), .b(t3_010011011), .y(t3_01001101));
wire t3_010011010, t3_010011011;
mixer mix_t3_0100111 (.a(t3_01001110), .b(t3_01001111), .y(t3_0100111));
wire t3_01001110, t3_01001111;
mixer mix_t3_01001110 (.a(t3_010011100), .b(t3_010011101), .y(t3_01001110));
wire t3_010011100, t3_010011101;
mixer mix_t3_01001111 (.a(t3_010011110), .b(t3_010011111), .y(t3_01001111));
wire t3_010011110, t3_010011111;
mixer mix_t3_0101 (.a(t3_01010), .b(t3_01011), .y(t3_0101));
wire t3_01010, t3_01011;
mixer mix_t3_01010 (.a(t3_010100), .b(t3_010101), .y(t3_01010));
wire t3_010100, t3_010101;
mixer mix_t3_010100 (.a(t3_0101000), .b(t3_0101001), .y(t3_010100));
wire t3_0101000, t3_0101001;
mixer mix_t3_0101000 (.a(t3_01010000), .b(t3_01010001), .y(t3_0101000));
wire t3_01010000, t3_01010001;
mixer mix_t3_01010000 (.a(t3_010100000), .b(t3_010100001), .y(t3_01010000));
wire t3_010100000, t3_010100001;
mixer mix_t3_01010001 (.a(t3_010100010), .b(t3_010100011), .y(t3_01010001));
wire t3_010100010, t3_010100011;
mixer mix_t3_0101001 (.a(t3_01010010), .b(t3_01010011), .y(t3_0101001));
wire t3_01010010, t3_01010011;
mixer mix_t3_01010010 (.a(t3_010100100), .b(t3_010100101), .y(t3_01010010));
wire t3_010100100, t3_010100101;
mixer mix_t3_01010011 (.a(t3_010100110), .b(t3_010100111), .y(t3_01010011));
wire t3_010100110, t3_010100111;
mixer mix_t3_010101 (.a(t3_0101010), .b(t3_0101011), .y(t3_010101));
wire t3_0101010, t3_0101011;
mixer mix_t3_0101010 (.a(t3_01010100), .b(t3_01010101), .y(t3_0101010));
wire t3_01010100, t3_01010101;
mixer mix_t3_01010100 (.a(t3_010101000), .b(t3_010101001), .y(t3_01010100));
wire t3_010101000, t3_010101001;
mixer mix_t3_01010101 (.a(t3_010101010), .b(t3_010101011), .y(t3_01010101));
wire t3_010101010, t3_010101011;
mixer mix_t3_0101011 (.a(t3_01010110), .b(t3_01010111), .y(t3_0101011));
wire t3_01010110, t3_01010111;
mixer mix_t3_01010110 (.a(t3_010101100), .b(t3_010101101), .y(t3_01010110));
wire t3_010101100, t3_010101101;
mixer mix_t3_01010111 (.a(t3_010101110), .b(t3_010101111), .y(t3_01010111));
wire t3_010101110, t3_010101111;
mixer mix_t3_01011 (.a(t3_010110), .b(t3_010111), .y(t3_01011));
wire t3_010110, t3_010111;
mixer mix_t3_010110 (.a(t3_0101100), .b(t3_0101101), .y(t3_010110));
wire t3_0101100, t3_0101101;
mixer mix_t3_0101100 (.a(t3_01011000), .b(t3_01011001), .y(t3_0101100));
wire t3_01011000, t3_01011001;
mixer mix_t3_01011000 (.a(t3_010110000), .b(t3_010110001), .y(t3_01011000));
wire t3_010110000, t3_010110001;
mixer mix_t3_01011001 (.a(t3_010110010), .b(t3_010110011), .y(t3_01011001));
wire t3_010110010, t3_010110011;
mixer mix_t3_0101101 (.a(t3_01011010), .b(t3_01011011), .y(t3_0101101));
wire t3_01011010, t3_01011011;
mixer mix_t3_01011010 (.a(t3_010110100), .b(t3_010110101), .y(t3_01011010));
wire t3_010110100, t3_010110101;
mixer mix_t3_01011011 (.a(t3_010110110), .b(t3_010110111), .y(t3_01011011));
wire t3_010110110, t3_010110111;
mixer mix_t3_010111 (.a(t3_0101110), .b(t3_0101111), .y(t3_010111));
wire t3_0101110, t3_0101111;
mixer mix_t3_0101110 (.a(t3_01011100), .b(t3_01011101), .y(t3_0101110));
wire t3_01011100, t3_01011101;
mixer mix_t3_01011100 (.a(t3_010111000), .b(t3_010111001), .y(t3_01011100));
wire t3_010111000, t3_010111001;
mixer mix_t3_01011101 (.a(t3_010111010), .b(t3_010111011), .y(t3_01011101));
wire t3_010111010, t3_010111011;
mixer mix_t3_0101111 (.a(t3_01011110), .b(t3_01011111), .y(t3_0101111));
wire t3_01011110, t3_01011111;
mixer mix_t3_01011110 (.a(t3_010111100), .b(t3_010111101), .y(t3_01011110));
wire t3_010111100, t3_010111101;
mixer mix_t3_01011111 (.a(t3_010111110), .b(t3_010111111), .y(t3_01011111));
wire t3_010111110, t3_010111111;
mixer mix_t3_011 (.a(t3_0110), .b(t3_0111), .y(t3_011));
wire t3_0110, t3_0111;
mixer mix_t3_0110 (.a(t3_01100), .b(t3_01101), .y(t3_0110));
wire t3_01100, t3_01101;
mixer mix_t3_01100 (.a(t3_011000), .b(t3_011001), .y(t3_01100));
wire t3_011000, t3_011001;
mixer mix_t3_011000 (.a(t3_0110000), .b(t3_0110001), .y(t3_011000));
wire t3_0110000, t3_0110001;
mixer mix_t3_0110000 (.a(t3_01100000), .b(t3_01100001), .y(t3_0110000));
wire t3_01100000, t3_01100001;
mixer mix_t3_01100000 (.a(t3_011000000), .b(t3_011000001), .y(t3_01100000));
wire t3_011000000, t3_011000001;
mixer mix_t3_01100001 (.a(t3_011000010), .b(t3_011000011), .y(t3_01100001));
wire t3_011000010, t3_011000011;
mixer mix_t3_0110001 (.a(t3_01100010), .b(t3_01100011), .y(t3_0110001));
wire t3_01100010, t3_01100011;
mixer mix_t3_01100010 (.a(t3_011000100), .b(t3_011000101), .y(t3_01100010));
wire t3_011000100, t3_011000101;
mixer mix_t3_01100011 (.a(t3_011000110), .b(t3_011000111), .y(t3_01100011));
wire t3_011000110, t3_011000111;
mixer mix_t3_011001 (.a(t3_0110010), .b(t3_0110011), .y(t3_011001));
wire t3_0110010, t3_0110011;
mixer mix_t3_0110010 (.a(t3_01100100), .b(t3_01100101), .y(t3_0110010));
wire t3_01100100, t3_01100101;
mixer mix_t3_01100100 (.a(t3_011001000), .b(t3_011001001), .y(t3_01100100));
wire t3_011001000, t3_011001001;
mixer mix_t3_01100101 (.a(t3_011001010), .b(t3_011001011), .y(t3_01100101));
wire t3_011001010, t3_011001011;
mixer mix_t3_0110011 (.a(t3_01100110), .b(t3_01100111), .y(t3_0110011));
wire t3_01100110, t3_01100111;
mixer mix_t3_01100110 (.a(t3_011001100), .b(t3_011001101), .y(t3_01100110));
wire t3_011001100, t3_011001101;
mixer mix_t3_01100111 (.a(t3_011001110), .b(t3_011001111), .y(t3_01100111));
wire t3_011001110, t3_011001111;
mixer mix_t3_01101 (.a(t3_011010), .b(t3_011011), .y(t3_01101));
wire t3_011010, t3_011011;
mixer mix_t3_011010 (.a(t3_0110100), .b(t3_0110101), .y(t3_011010));
wire t3_0110100, t3_0110101;
mixer mix_t3_0110100 (.a(t3_01101000), .b(t3_01101001), .y(t3_0110100));
wire t3_01101000, t3_01101001;
mixer mix_t3_01101000 (.a(t3_011010000), .b(t3_011010001), .y(t3_01101000));
wire t3_011010000, t3_011010001;
mixer mix_t3_01101001 (.a(t3_011010010), .b(t3_011010011), .y(t3_01101001));
wire t3_011010010, t3_011010011;
mixer mix_t3_0110101 (.a(t3_01101010), .b(t3_01101011), .y(t3_0110101));
wire t3_01101010, t3_01101011;
mixer mix_t3_01101010 (.a(t3_011010100), .b(t3_011010101), .y(t3_01101010));
wire t3_011010100, t3_011010101;
mixer mix_t3_01101011 (.a(t3_011010110), .b(t3_011010111), .y(t3_01101011));
wire t3_011010110, t3_011010111;
mixer mix_t3_011011 (.a(t3_0110110), .b(t3_0110111), .y(t3_011011));
wire t3_0110110, t3_0110111;
mixer mix_t3_0110110 (.a(t3_01101100), .b(t3_01101101), .y(t3_0110110));
wire t3_01101100, t3_01101101;
mixer mix_t3_01101100 (.a(t3_011011000), .b(t3_011011001), .y(t3_01101100));
wire t3_011011000, t3_011011001;
mixer mix_t3_01101101 (.a(t3_011011010), .b(t3_011011011), .y(t3_01101101));
wire t3_011011010, t3_011011011;
mixer mix_t3_0110111 (.a(t3_01101110), .b(t3_01101111), .y(t3_0110111));
wire t3_01101110, t3_01101111;
mixer mix_t3_01101110 (.a(t3_011011100), .b(t3_011011101), .y(t3_01101110));
wire t3_011011100, t3_011011101;
mixer mix_t3_01101111 (.a(t3_011011110), .b(t3_011011111), .y(t3_01101111));
wire t3_011011110, t3_011011111;
mixer mix_t3_0111 (.a(t3_01110), .b(t3_01111), .y(t3_0111));
wire t3_01110, t3_01111;
mixer mix_t3_01110 (.a(t3_011100), .b(t3_011101), .y(t3_01110));
wire t3_011100, t3_011101;
mixer mix_t3_011100 (.a(t3_0111000), .b(t3_0111001), .y(t3_011100));
wire t3_0111000, t3_0111001;
mixer mix_t3_0111000 (.a(t3_01110000), .b(t3_01110001), .y(t3_0111000));
wire t3_01110000, t3_01110001;
mixer mix_t3_01110000 (.a(t3_011100000), .b(t3_011100001), .y(t3_01110000));
wire t3_011100000, t3_011100001;
mixer mix_t3_01110001 (.a(t3_011100010), .b(t3_011100011), .y(t3_01110001));
wire t3_011100010, t3_011100011;
mixer mix_t3_0111001 (.a(t3_01110010), .b(t3_01110011), .y(t3_0111001));
wire t3_01110010, t3_01110011;
mixer mix_t3_01110010 (.a(t3_011100100), .b(t3_011100101), .y(t3_01110010));
wire t3_011100100, t3_011100101;
mixer mix_t3_01110011 (.a(t3_011100110), .b(t3_011100111), .y(t3_01110011));
wire t3_011100110, t3_011100111;
mixer mix_t3_011101 (.a(t3_0111010), .b(t3_0111011), .y(t3_011101));
wire t3_0111010, t3_0111011;
mixer mix_t3_0111010 (.a(t3_01110100), .b(t3_01110101), .y(t3_0111010));
wire t3_01110100, t3_01110101;
mixer mix_t3_01110100 (.a(t3_011101000), .b(t3_011101001), .y(t3_01110100));
wire t3_011101000, t3_011101001;
mixer mix_t3_01110101 (.a(t3_011101010), .b(t3_011101011), .y(t3_01110101));
wire t3_011101010, t3_011101011;
mixer mix_t3_0111011 (.a(t3_01110110), .b(t3_01110111), .y(t3_0111011));
wire t3_01110110, t3_01110111;
mixer mix_t3_01110110 (.a(t3_011101100), .b(t3_011101101), .y(t3_01110110));
wire t3_011101100, t3_011101101;
mixer mix_t3_01110111 (.a(t3_011101110), .b(t3_011101111), .y(t3_01110111));
wire t3_011101110, t3_011101111;
mixer mix_t3_01111 (.a(t3_011110), .b(t3_011111), .y(t3_01111));
wire t3_011110, t3_011111;
mixer mix_t3_011110 (.a(t3_0111100), .b(t3_0111101), .y(t3_011110));
wire t3_0111100, t3_0111101;
mixer mix_t3_0111100 (.a(t3_01111000), .b(t3_01111001), .y(t3_0111100));
wire t3_01111000, t3_01111001;
mixer mix_t3_01111000 (.a(t3_011110000), .b(t3_011110001), .y(t3_01111000));
wire t3_011110000, t3_011110001;
mixer mix_t3_01111001 (.a(t3_011110010), .b(t3_011110011), .y(t3_01111001));
wire t3_011110010, t3_011110011;
mixer mix_t3_0111101 (.a(t3_01111010), .b(t3_01111011), .y(t3_0111101));
wire t3_01111010, t3_01111011;
mixer mix_t3_01111010 (.a(t3_011110100), .b(t3_011110101), .y(t3_01111010));
wire t3_011110100, t3_011110101;
mixer mix_t3_01111011 (.a(t3_011110110), .b(t3_011110111), .y(t3_01111011));
wire t3_011110110, t3_011110111;
mixer mix_t3_011111 (.a(t3_0111110), .b(t3_0111111), .y(t3_011111));
wire t3_0111110, t3_0111111;
mixer mix_t3_0111110 (.a(t3_01111100), .b(t3_01111101), .y(t3_0111110));
wire t3_01111100, t3_01111101;
mixer mix_t3_01111100 (.a(t3_011111000), .b(t3_011111001), .y(t3_01111100));
wire t3_011111000, t3_011111001;
mixer mix_t3_01111101 (.a(t3_011111010), .b(t3_011111011), .y(t3_01111101));
wire t3_011111010, t3_011111011;
mixer mix_t3_0111111 (.a(t3_01111110), .b(t3_01111111), .y(t3_0111111));
wire t3_01111110, t3_01111111;
mixer mix_t3_01111110 (.a(t3_011111100), .b(t3_011111101), .y(t3_01111110));
wire t3_011111100, t3_011111101;
mixer mix_t3_01111111 (.a(t3_011111110), .b(t3_011111111), .y(t3_01111111));
wire t3_011111110, t3_011111111;
mixer mix_t4_0 (.a(t4_00), .b(t4_01), .y(t4_0));
wire t4_00, t4_01;
mixer mix_t4_00 (.a(t4_000), .b(t4_001), .y(t4_00));
wire t4_000, t4_001;
mixer mix_t4_000 (.a(t4_0000), .b(t4_0001), .y(t4_000));
wire t4_0000, t4_0001;
mixer mix_t4_0000 (.a(t4_00000), .b(t4_00001), .y(t4_0000));
wire t4_00000, t4_00001;
mixer mix_t4_00000 (.a(t4_000000), .b(t4_000001), .y(t4_00000));
wire t4_000000, t4_000001;
mixer mix_t4_000000 (.a(t4_0000000), .b(t4_0000001), .y(t4_000000));
wire t4_0000000, t4_0000001;
mixer mix_t4_0000000 (.a(t4_00000000), .b(t4_00000001), .y(t4_0000000));
wire t4_00000000, t4_00000001;
mixer mix_t4_00000000 (.a(t4_000000000), .b(t4_000000001), .y(t4_00000000));
wire t4_000000000, t4_000000001;
mixer mix_t4_00000001 (.a(t4_000000010), .b(t4_000000011), .y(t4_00000001));
wire t4_000000010, t4_000000011;
mixer mix_t4_0000001 (.a(t4_00000010), .b(t4_00000011), .y(t4_0000001));
wire t4_00000010, t4_00000011;
mixer mix_t4_00000010 (.a(t4_000000100), .b(t4_000000101), .y(t4_00000010));
wire t4_000000100, t4_000000101;
mixer mix_t4_00000011 (.a(t4_000000110), .b(t4_000000111), .y(t4_00000011));
wire t4_000000110, t4_000000111;
mixer mix_t4_000001 (.a(t4_0000010), .b(t4_0000011), .y(t4_000001));
wire t4_0000010, t4_0000011;
mixer mix_t4_0000010 (.a(t4_00000100), .b(t4_00000101), .y(t4_0000010));
wire t4_00000100, t4_00000101;
mixer mix_t4_00000100 (.a(t4_000001000), .b(t4_000001001), .y(t4_00000100));
wire t4_000001000, t4_000001001;
mixer mix_t4_00000101 (.a(t4_000001010), .b(t4_000001011), .y(t4_00000101));
wire t4_000001010, t4_000001011;
mixer mix_t4_0000011 (.a(t4_00000110), .b(t4_00000111), .y(t4_0000011));
wire t4_00000110, t4_00000111;
mixer mix_t4_00000110 (.a(t4_000001100), .b(t4_000001101), .y(t4_00000110));
wire t4_000001100, t4_000001101;
mixer mix_t4_00000111 (.a(t4_000001110), .b(t4_000001111), .y(t4_00000111));
wire t4_000001110, t4_000001111;
mixer mix_t4_00001 (.a(t4_000010), .b(t4_000011), .y(t4_00001));
wire t4_000010, t4_000011;
mixer mix_t4_000010 (.a(t4_0000100), .b(t4_0000101), .y(t4_000010));
wire t4_0000100, t4_0000101;
mixer mix_t4_0000100 (.a(t4_00001000), .b(t4_00001001), .y(t4_0000100));
wire t4_00001000, t4_00001001;
mixer mix_t4_00001000 (.a(t4_000010000), .b(t4_000010001), .y(t4_00001000));
wire t4_000010000, t4_000010001;
mixer mix_t4_00001001 (.a(t4_000010010), .b(t4_000010011), .y(t4_00001001));
wire t4_000010010, t4_000010011;
mixer mix_t4_0000101 (.a(t4_00001010), .b(t4_00001011), .y(t4_0000101));
wire t4_00001010, t4_00001011;
mixer mix_t4_00001010 (.a(t4_000010100), .b(t4_000010101), .y(t4_00001010));
wire t4_000010100, t4_000010101;
mixer mix_t4_00001011 (.a(t4_000010110), .b(t4_000010111), .y(t4_00001011));
wire t4_000010110, t4_000010111;
mixer mix_t4_000011 (.a(t4_0000110), .b(t4_0000111), .y(t4_000011));
wire t4_0000110, t4_0000111;
mixer mix_t4_0000110 (.a(t4_00001100), .b(t4_00001101), .y(t4_0000110));
wire t4_00001100, t4_00001101;
mixer mix_t4_00001100 (.a(t4_000011000), .b(t4_000011001), .y(t4_00001100));
wire t4_000011000, t4_000011001;
mixer mix_t4_00001101 (.a(t4_000011010), .b(t4_000011011), .y(t4_00001101));
wire t4_000011010, t4_000011011;
mixer mix_t4_0000111 (.a(t4_00001110), .b(t4_00001111), .y(t4_0000111));
wire t4_00001110, t4_00001111;
mixer mix_t4_00001110 (.a(t4_000011100), .b(t4_000011101), .y(t4_00001110));
wire t4_000011100, t4_000011101;
mixer mix_t4_00001111 (.a(t4_000011110), .b(t4_000011111), .y(t4_00001111));
wire t4_000011110, t4_000011111;
mixer mix_t4_0001 (.a(t4_00010), .b(t4_00011), .y(t4_0001));
wire t4_00010, t4_00011;
mixer mix_t4_00010 (.a(t4_000100), .b(t4_000101), .y(t4_00010));
wire t4_000100, t4_000101;
mixer mix_t4_000100 (.a(t4_0001000), .b(t4_0001001), .y(t4_000100));
wire t4_0001000, t4_0001001;
mixer mix_t4_0001000 (.a(t4_00010000), .b(t4_00010001), .y(t4_0001000));
wire t4_00010000, t4_00010001;
mixer mix_t4_00010000 (.a(t4_000100000), .b(t4_000100001), .y(t4_00010000));
wire t4_000100000, t4_000100001;
mixer mix_t4_00010001 (.a(t4_000100010), .b(t4_000100011), .y(t4_00010001));
wire t4_000100010, t4_000100011;
mixer mix_t4_0001001 (.a(t4_00010010), .b(t4_00010011), .y(t4_0001001));
wire t4_00010010, t4_00010011;
mixer mix_t4_00010010 (.a(t4_000100100), .b(t4_000100101), .y(t4_00010010));
wire t4_000100100, t4_000100101;
mixer mix_t4_00010011 (.a(t4_000100110), .b(t4_000100111), .y(t4_00010011));
wire t4_000100110, t4_000100111;
mixer mix_t4_000101 (.a(t4_0001010), .b(t4_0001011), .y(t4_000101));
wire t4_0001010, t4_0001011;
mixer mix_t4_0001010 (.a(t4_00010100), .b(t4_00010101), .y(t4_0001010));
wire t4_00010100, t4_00010101;
mixer mix_t4_00010100 (.a(t4_000101000), .b(t4_000101001), .y(t4_00010100));
wire t4_000101000, t4_000101001;
mixer mix_t4_00010101 (.a(t4_000101010), .b(t4_000101011), .y(t4_00010101));
wire t4_000101010, t4_000101011;
mixer mix_t4_0001011 (.a(t4_00010110), .b(t4_00010111), .y(t4_0001011));
wire t4_00010110, t4_00010111;
mixer mix_t4_00010110 (.a(t4_000101100), .b(t4_000101101), .y(t4_00010110));
wire t4_000101100, t4_000101101;
mixer mix_t4_00010111 (.a(t4_000101110), .b(t4_000101111), .y(t4_00010111));
wire t4_000101110, t4_000101111;
mixer mix_t4_00011 (.a(t4_000110), .b(t4_000111), .y(t4_00011));
wire t4_000110, t4_000111;
mixer mix_t4_000110 (.a(t4_0001100), .b(t4_0001101), .y(t4_000110));
wire t4_0001100, t4_0001101;
mixer mix_t4_0001100 (.a(t4_00011000), .b(t4_00011001), .y(t4_0001100));
wire t4_00011000, t4_00011001;
mixer mix_t4_00011000 (.a(t4_000110000), .b(t4_000110001), .y(t4_00011000));
wire t4_000110000, t4_000110001;
mixer mix_t4_00011001 (.a(t4_000110010), .b(t4_000110011), .y(t4_00011001));
wire t4_000110010, t4_000110011;
mixer mix_t4_0001101 (.a(t4_00011010), .b(t4_00011011), .y(t4_0001101));
wire t4_00011010, t4_00011011;
mixer mix_t4_00011010 (.a(t4_000110100), .b(t4_000110101), .y(t4_00011010));
wire t4_000110100, t4_000110101;
mixer mix_t4_00011011 (.a(t4_000110110), .b(t4_000110111), .y(t4_00011011));
wire t4_000110110, t4_000110111;
mixer mix_t4_000111 (.a(t4_0001110), .b(t4_0001111), .y(t4_000111));
wire t4_0001110, t4_0001111;
mixer mix_t4_0001110 (.a(t4_00011100), .b(t4_00011101), .y(t4_0001110));
wire t4_00011100, t4_00011101;
mixer mix_t4_00011100 (.a(t4_000111000), .b(t4_000111001), .y(t4_00011100));
wire t4_000111000, t4_000111001;
mixer mix_t4_00011101 (.a(t4_000111010), .b(t4_000111011), .y(t4_00011101));
wire t4_000111010, t4_000111011;
mixer mix_t4_0001111 (.a(t4_00011110), .b(t4_00011111), .y(t4_0001111));
wire t4_00011110, t4_00011111;
mixer mix_t4_00011110 (.a(t4_000111100), .b(t4_000111101), .y(t4_00011110));
wire t4_000111100, t4_000111101;
mixer mix_t4_00011111 (.a(t4_000111110), .b(t4_000111111), .y(t4_00011111));
wire t4_000111110, t4_000111111;
mixer mix_t4_001 (.a(t4_0010), .b(t4_0011), .y(t4_001));
wire t4_0010, t4_0011;
mixer mix_t4_0010 (.a(t4_00100), .b(t4_00101), .y(t4_0010));
wire t4_00100, t4_00101;
mixer mix_t4_00100 (.a(t4_001000), .b(t4_001001), .y(t4_00100));
wire t4_001000, t4_001001;
mixer mix_t4_001000 (.a(t4_0010000), .b(t4_0010001), .y(t4_001000));
wire t4_0010000, t4_0010001;
mixer mix_t4_0010000 (.a(t4_00100000), .b(t4_00100001), .y(t4_0010000));
wire t4_00100000, t4_00100001;
mixer mix_t4_00100000 (.a(t4_001000000), .b(t4_001000001), .y(t4_00100000));
wire t4_001000000, t4_001000001;
mixer mix_t4_00100001 (.a(t4_001000010), .b(t4_001000011), .y(t4_00100001));
wire t4_001000010, t4_001000011;
mixer mix_t4_0010001 (.a(t4_00100010), .b(t4_00100011), .y(t4_0010001));
wire t4_00100010, t4_00100011;
mixer mix_t4_00100010 (.a(t4_001000100), .b(t4_001000101), .y(t4_00100010));
wire t4_001000100, t4_001000101;
mixer mix_t4_00100011 (.a(t4_001000110), .b(t4_001000111), .y(t4_00100011));
wire t4_001000110, t4_001000111;
mixer mix_t4_001001 (.a(t4_0010010), .b(t4_0010011), .y(t4_001001));
wire t4_0010010, t4_0010011;
mixer mix_t4_0010010 (.a(t4_00100100), .b(t4_00100101), .y(t4_0010010));
wire t4_00100100, t4_00100101;
mixer mix_t4_00100100 (.a(t4_001001000), .b(t4_001001001), .y(t4_00100100));
wire t4_001001000, t4_001001001;
mixer mix_t4_00100101 (.a(t4_001001010), .b(t4_001001011), .y(t4_00100101));
wire t4_001001010, t4_001001011;
mixer mix_t4_0010011 (.a(t4_00100110), .b(t4_00100111), .y(t4_0010011));
wire t4_00100110, t4_00100111;
mixer mix_t4_00100110 (.a(t4_001001100), .b(t4_001001101), .y(t4_00100110));
wire t4_001001100, t4_001001101;
mixer mix_t4_00100111 (.a(t4_001001110), .b(t4_001001111), .y(t4_00100111));
wire t4_001001110, t4_001001111;
mixer mix_t4_00101 (.a(t4_001010), .b(t4_001011), .y(t4_00101));
wire t4_001010, t4_001011;
mixer mix_t4_001010 (.a(t4_0010100), .b(t4_0010101), .y(t4_001010));
wire t4_0010100, t4_0010101;
mixer mix_t4_0010100 (.a(t4_00101000), .b(t4_00101001), .y(t4_0010100));
wire t4_00101000, t4_00101001;
mixer mix_t4_00101000 (.a(t4_001010000), .b(t4_001010001), .y(t4_00101000));
wire t4_001010000, t4_001010001;
mixer mix_t4_00101001 (.a(t4_001010010), .b(t4_001010011), .y(t4_00101001));
wire t4_001010010, t4_001010011;
mixer mix_t4_0010101 (.a(t4_00101010), .b(t4_00101011), .y(t4_0010101));
wire t4_00101010, t4_00101011;
mixer mix_t4_00101010 (.a(t4_001010100), .b(t4_001010101), .y(t4_00101010));
wire t4_001010100, t4_001010101;
mixer mix_t4_00101011 (.a(t4_001010110), .b(t4_001010111), .y(t4_00101011));
wire t4_001010110, t4_001010111;
mixer mix_t4_001011 (.a(t4_0010110), .b(t4_0010111), .y(t4_001011));
wire t4_0010110, t4_0010111;
mixer mix_t4_0010110 (.a(t4_00101100), .b(t4_00101101), .y(t4_0010110));
wire t4_00101100, t4_00101101;
mixer mix_t4_00101100 (.a(t4_001011000), .b(t4_001011001), .y(t4_00101100));
wire t4_001011000, t4_001011001;
mixer mix_t4_00101101 (.a(t4_001011010), .b(t4_001011011), .y(t4_00101101));
wire t4_001011010, t4_001011011;
mixer mix_t4_0010111 (.a(t4_00101110), .b(t4_00101111), .y(t4_0010111));
wire t4_00101110, t4_00101111;
mixer mix_t4_00101110 (.a(t4_001011100), .b(t4_001011101), .y(t4_00101110));
wire t4_001011100, t4_001011101;
mixer mix_t4_00101111 (.a(t4_001011110), .b(t4_001011111), .y(t4_00101111));
wire t4_001011110, t4_001011111;
mixer mix_t4_0011 (.a(t4_00110), .b(t4_00111), .y(t4_0011));
wire t4_00110, t4_00111;
mixer mix_t4_00110 (.a(t4_001100), .b(t4_001101), .y(t4_00110));
wire t4_001100, t4_001101;
mixer mix_t4_001100 (.a(t4_0011000), .b(t4_0011001), .y(t4_001100));
wire t4_0011000, t4_0011001;
mixer mix_t4_0011000 (.a(t4_00110000), .b(t4_00110001), .y(t4_0011000));
wire t4_00110000, t4_00110001;
mixer mix_t4_00110000 (.a(t4_001100000), .b(t4_001100001), .y(t4_00110000));
wire t4_001100000, t4_001100001;
mixer mix_t4_00110001 (.a(t4_001100010), .b(t4_001100011), .y(t4_00110001));
wire t4_001100010, t4_001100011;
mixer mix_t4_0011001 (.a(t4_00110010), .b(t4_00110011), .y(t4_0011001));
wire t4_00110010, t4_00110011;
mixer mix_t4_00110010 (.a(t4_001100100), .b(t4_001100101), .y(t4_00110010));
wire t4_001100100, t4_001100101;
mixer mix_t4_00110011 (.a(t4_001100110), .b(t4_001100111), .y(t4_00110011));
wire t4_001100110, t4_001100111;
mixer mix_t4_001101 (.a(t4_0011010), .b(t4_0011011), .y(t4_001101));
wire t4_0011010, t4_0011011;
mixer mix_t4_0011010 (.a(t4_00110100), .b(t4_00110101), .y(t4_0011010));
wire t4_00110100, t4_00110101;
mixer mix_t4_00110100 (.a(t4_001101000), .b(t4_001101001), .y(t4_00110100));
wire t4_001101000, t4_001101001;
mixer mix_t4_00110101 (.a(t4_001101010), .b(t4_001101011), .y(t4_00110101));
wire t4_001101010, t4_001101011;
mixer mix_t4_0011011 (.a(t4_00110110), .b(t4_00110111), .y(t4_0011011));
wire t4_00110110, t4_00110111;
mixer mix_t4_00110110 (.a(t4_001101100), .b(t4_001101101), .y(t4_00110110));
wire t4_001101100, t4_001101101;
mixer mix_t4_00110111 (.a(t4_001101110), .b(t4_001101111), .y(t4_00110111));
wire t4_001101110, t4_001101111;
mixer mix_t4_00111 (.a(t4_001110), .b(t4_001111), .y(t4_00111));
wire t4_001110, t4_001111;
mixer mix_t4_001110 (.a(t4_0011100), .b(t4_0011101), .y(t4_001110));
wire t4_0011100, t4_0011101;
mixer mix_t4_0011100 (.a(t4_00111000), .b(t4_00111001), .y(t4_0011100));
wire t4_00111000, t4_00111001;
mixer mix_t4_00111000 (.a(t4_001110000), .b(t4_001110001), .y(t4_00111000));
wire t4_001110000, t4_001110001;
mixer mix_t4_00111001 (.a(t4_001110010), .b(t4_001110011), .y(t4_00111001));
wire t4_001110010, t4_001110011;
mixer mix_t4_0011101 (.a(t4_00111010), .b(t4_00111011), .y(t4_0011101));
wire t4_00111010, t4_00111011;
mixer mix_t4_00111010 (.a(t4_001110100), .b(t4_001110101), .y(t4_00111010));
wire t4_001110100, t4_001110101;
mixer mix_t4_00111011 (.a(t4_001110110), .b(t4_001110111), .y(t4_00111011));
wire t4_001110110, t4_001110111;
mixer mix_t4_001111 (.a(t4_0011110), .b(t4_0011111), .y(t4_001111));
wire t4_0011110, t4_0011111;
mixer mix_t4_0011110 (.a(t4_00111100), .b(t4_00111101), .y(t4_0011110));
wire t4_00111100, t4_00111101;
mixer mix_t4_00111100 (.a(t4_001111000), .b(t4_001111001), .y(t4_00111100));
wire t4_001111000, t4_001111001;
mixer mix_t4_00111101 (.a(t4_001111010), .b(t4_001111011), .y(t4_00111101));
wire t4_001111010, t4_001111011;
mixer mix_t4_0011111 (.a(t4_00111110), .b(t4_00111111), .y(t4_0011111));
wire t4_00111110, t4_00111111;
mixer mix_t4_00111110 (.a(t4_001111100), .b(t4_001111101), .y(t4_00111110));
wire t4_001111100, t4_001111101;
mixer mix_t4_00111111 (.a(t4_001111110), .b(t4_001111111), .y(t4_00111111));
wire t4_001111110, t4_001111111;
mixer mix_t4_01 (.a(t4_010), .b(t4_011), .y(t4_01));
wire t4_010, t4_011;
mixer mix_t4_010 (.a(t4_0100), .b(t4_0101), .y(t4_010));
wire t4_0100, t4_0101;
mixer mix_t4_0100 (.a(t4_01000), .b(t4_01001), .y(t4_0100));
wire t4_01000, t4_01001;
mixer mix_t4_01000 (.a(t4_010000), .b(t4_010001), .y(t4_01000));
wire t4_010000, t4_010001;
mixer mix_t4_010000 (.a(t4_0100000), .b(t4_0100001), .y(t4_010000));
wire t4_0100000, t4_0100001;
mixer mix_t4_0100000 (.a(t4_01000000), .b(t4_01000001), .y(t4_0100000));
wire t4_01000000, t4_01000001;
mixer mix_t4_01000000 (.a(t4_010000000), .b(t4_010000001), .y(t4_01000000));
wire t4_010000000, t4_010000001;
mixer mix_t4_01000001 (.a(t4_010000010), .b(t4_010000011), .y(t4_01000001));
wire t4_010000010, t4_010000011;
mixer mix_t4_0100001 (.a(t4_01000010), .b(t4_01000011), .y(t4_0100001));
wire t4_01000010, t4_01000011;
mixer mix_t4_01000010 (.a(t4_010000100), .b(t4_010000101), .y(t4_01000010));
wire t4_010000100, t4_010000101;
mixer mix_t4_01000011 (.a(t4_010000110), .b(t4_010000111), .y(t4_01000011));
wire t4_010000110, t4_010000111;
mixer mix_t4_010001 (.a(t4_0100010), .b(t4_0100011), .y(t4_010001));
wire t4_0100010, t4_0100011;
mixer mix_t4_0100010 (.a(t4_01000100), .b(t4_01000101), .y(t4_0100010));
wire t4_01000100, t4_01000101;
mixer mix_t4_01000100 (.a(t4_010001000), .b(t4_010001001), .y(t4_01000100));
wire t4_010001000, t4_010001001;
mixer mix_t4_01000101 (.a(t4_010001010), .b(t4_010001011), .y(t4_01000101));
wire t4_010001010, t4_010001011;
mixer mix_t4_0100011 (.a(t4_01000110), .b(t4_01000111), .y(t4_0100011));
wire t4_01000110, t4_01000111;
mixer mix_t4_01000110 (.a(t4_010001100), .b(t4_010001101), .y(t4_01000110));
wire t4_010001100, t4_010001101;
mixer mix_t4_01000111 (.a(t4_010001110), .b(t4_010001111), .y(t4_01000111));
wire t4_010001110, t4_010001111;
mixer mix_t4_01001 (.a(t4_010010), .b(t4_010011), .y(t4_01001));
wire t4_010010, t4_010011;
mixer mix_t4_010010 (.a(t4_0100100), .b(t4_0100101), .y(t4_010010));
wire t4_0100100, t4_0100101;
mixer mix_t4_0100100 (.a(t4_01001000), .b(t4_01001001), .y(t4_0100100));
wire t4_01001000, t4_01001001;
mixer mix_t4_01001000 (.a(t4_010010000), .b(t4_010010001), .y(t4_01001000));
wire t4_010010000, t4_010010001;
mixer mix_t4_01001001 (.a(t4_010010010), .b(t4_010010011), .y(t4_01001001));
wire t4_010010010, t4_010010011;
mixer mix_t4_0100101 (.a(t4_01001010), .b(t4_01001011), .y(t4_0100101));
wire t4_01001010, t4_01001011;
mixer mix_t4_01001010 (.a(t4_010010100), .b(t4_010010101), .y(t4_01001010));
wire t4_010010100, t4_010010101;
mixer mix_t4_01001011 (.a(t4_010010110), .b(t4_010010111), .y(t4_01001011));
wire t4_010010110, t4_010010111;
mixer mix_t4_010011 (.a(t4_0100110), .b(t4_0100111), .y(t4_010011));
wire t4_0100110, t4_0100111;
mixer mix_t4_0100110 (.a(t4_01001100), .b(t4_01001101), .y(t4_0100110));
wire t4_01001100, t4_01001101;
mixer mix_t4_01001100 (.a(t4_010011000), .b(t4_010011001), .y(t4_01001100));
wire t4_010011000, t4_010011001;
mixer mix_t4_01001101 (.a(t4_010011010), .b(t4_010011011), .y(t4_01001101));
wire t4_010011010, t4_010011011;
mixer mix_t4_0100111 (.a(t4_01001110), .b(t4_01001111), .y(t4_0100111));
wire t4_01001110, t4_01001111;
mixer mix_t4_01001110 (.a(t4_010011100), .b(t4_010011101), .y(t4_01001110));
wire t4_010011100, t4_010011101;
mixer mix_t4_01001111 (.a(t4_010011110), .b(t4_010011111), .y(t4_01001111));
wire t4_010011110, t4_010011111;
mixer mix_t4_0101 (.a(t4_01010), .b(t4_01011), .y(t4_0101));
wire t4_01010, t4_01011;
mixer mix_t4_01010 (.a(t4_010100), .b(t4_010101), .y(t4_01010));
wire t4_010100, t4_010101;
mixer mix_t4_010100 (.a(t4_0101000), .b(t4_0101001), .y(t4_010100));
wire t4_0101000, t4_0101001;
mixer mix_t4_0101000 (.a(t4_01010000), .b(t4_01010001), .y(t4_0101000));
wire t4_01010000, t4_01010001;
mixer mix_t4_01010000 (.a(t4_010100000), .b(t4_010100001), .y(t4_01010000));
wire t4_010100000, t4_010100001;
mixer mix_t4_01010001 (.a(t4_010100010), .b(t4_010100011), .y(t4_01010001));
wire t4_010100010, t4_010100011;
mixer mix_t4_0101001 (.a(t4_01010010), .b(t4_01010011), .y(t4_0101001));
wire t4_01010010, t4_01010011;
mixer mix_t4_01010010 (.a(t4_010100100), .b(t4_010100101), .y(t4_01010010));
wire t4_010100100, t4_010100101;
mixer mix_t4_01010011 (.a(t4_010100110), .b(t4_010100111), .y(t4_01010011));
wire t4_010100110, t4_010100111;
mixer mix_t4_010101 (.a(t4_0101010), .b(t4_0101011), .y(t4_010101));
wire t4_0101010, t4_0101011;
mixer mix_t4_0101010 (.a(t4_01010100), .b(t4_01010101), .y(t4_0101010));
wire t4_01010100, t4_01010101;
mixer mix_t4_01010100 (.a(t4_010101000), .b(t4_010101001), .y(t4_01010100));
wire t4_010101000, t4_010101001;
mixer mix_t4_01010101 (.a(t4_010101010), .b(t4_010101011), .y(t4_01010101));
wire t4_010101010, t4_010101011;
mixer mix_t4_0101011 (.a(t4_01010110), .b(t4_01010111), .y(t4_0101011));
wire t4_01010110, t4_01010111;
mixer mix_t4_01010110 (.a(t4_010101100), .b(t4_010101101), .y(t4_01010110));
wire t4_010101100, t4_010101101;
mixer mix_t4_01010111 (.a(t4_010101110), .b(t4_010101111), .y(t4_01010111));
wire t4_010101110, t4_010101111;
mixer mix_t4_01011 (.a(t4_010110), .b(t4_010111), .y(t4_01011));
wire t4_010110, t4_010111;
mixer mix_t4_010110 (.a(t4_0101100), .b(t4_0101101), .y(t4_010110));
wire t4_0101100, t4_0101101;
mixer mix_t4_0101100 (.a(t4_01011000), .b(t4_01011001), .y(t4_0101100));
wire t4_01011000, t4_01011001;
mixer mix_t4_01011000 (.a(t4_010110000), .b(t4_010110001), .y(t4_01011000));
wire t4_010110000, t4_010110001;
mixer mix_t4_01011001 (.a(t4_010110010), .b(t4_010110011), .y(t4_01011001));
wire t4_010110010, t4_010110011;
mixer mix_t4_0101101 (.a(t4_01011010), .b(t4_01011011), .y(t4_0101101));
wire t4_01011010, t4_01011011;
mixer mix_t4_01011010 (.a(t4_010110100), .b(t4_010110101), .y(t4_01011010));
wire t4_010110100, t4_010110101;
mixer mix_t4_01011011 (.a(t4_010110110), .b(t4_010110111), .y(t4_01011011));
wire t4_010110110, t4_010110111;
mixer mix_t4_010111 (.a(t4_0101110), .b(t4_0101111), .y(t4_010111));
wire t4_0101110, t4_0101111;
mixer mix_t4_0101110 (.a(t4_01011100), .b(t4_01011101), .y(t4_0101110));
wire t4_01011100, t4_01011101;
mixer mix_t4_01011100 (.a(t4_010111000), .b(t4_010111001), .y(t4_01011100));
wire t4_010111000, t4_010111001;
mixer mix_t4_01011101 (.a(t4_010111010), .b(t4_010111011), .y(t4_01011101));
wire t4_010111010, t4_010111011;
mixer mix_t4_0101111 (.a(t4_01011110), .b(t4_01011111), .y(t4_0101111));
wire t4_01011110, t4_01011111;
mixer mix_t4_01011110 (.a(t4_010111100), .b(t4_010111101), .y(t4_01011110));
wire t4_010111100, t4_010111101;
mixer mix_t4_01011111 (.a(t4_010111110), .b(t4_010111111), .y(t4_01011111));
wire t4_010111110, t4_010111111;
mixer mix_t4_011 (.a(t4_0110), .b(t4_0111), .y(t4_011));
wire t4_0110, t4_0111;
mixer mix_t4_0110 (.a(t4_01100), .b(t4_01101), .y(t4_0110));
wire t4_01100, t4_01101;
mixer mix_t4_01100 (.a(t4_011000), .b(t4_011001), .y(t4_01100));
wire t4_011000, t4_011001;
mixer mix_t4_011000 (.a(t4_0110000), .b(t4_0110001), .y(t4_011000));
wire t4_0110000, t4_0110001;
mixer mix_t4_0110000 (.a(t4_01100000), .b(t4_01100001), .y(t4_0110000));
wire t4_01100000, t4_01100001;
mixer mix_t4_01100000 (.a(t4_011000000), .b(t4_011000001), .y(t4_01100000));
wire t4_011000000, t4_011000001;
mixer mix_t4_01100001 (.a(t4_011000010), .b(t4_011000011), .y(t4_01100001));
wire t4_011000010, t4_011000011;
mixer mix_t4_0110001 (.a(t4_01100010), .b(t4_01100011), .y(t4_0110001));
wire t4_01100010, t4_01100011;
mixer mix_t4_01100010 (.a(t4_011000100), .b(t4_011000101), .y(t4_01100010));
wire t4_011000100, t4_011000101;
mixer mix_t4_01100011 (.a(t4_011000110), .b(t4_011000111), .y(t4_01100011));
wire t4_011000110, t4_011000111;
mixer mix_t4_011001 (.a(t4_0110010), .b(t4_0110011), .y(t4_011001));
wire t4_0110010, t4_0110011;
mixer mix_t4_0110010 (.a(t4_01100100), .b(t4_01100101), .y(t4_0110010));
wire t4_01100100, t4_01100101;
mixer mix_t4_01100100 (.a(t4_011001000), .b(t4_011001001), .y(t4_01100100));
wire t4_011001000, t4_011001001;
mixer mix_t4_01100101 (.a(t4_011001010), .b(t4_011001011), .y(t4_01100101));
wire t4_011001010, t4_011001011;
mixer mix_t4_0110011 (.a(t4_01100110), .b(t4_01100111), .y(t4_0110011));
wire t4_01100110, t4_01100111;
mixer mix_t4_01100110 (.a(t4_011001100), .b(t4_011001101), .y(t4_01100110));
wire t4_011001100, t4_011001101;
mixer mix_t4_01100111 (.a(t4_011001110), .b(t4_011001111), .y(t4_01100111));
wire t4_011001110, t4_011001111;
mixer mix_t4_01101 (.a(t4_011010), .b(t4_011011), .y(t4_01101));
wire t4_011010, t4_011011;
mixer mix_t4_011010 (.a(t4_0110100), .b(t4_0110101), .y(t4_011010));
wire t4_0110100, t4_0110101;
mixer mix_t4_0110100 (.a(t4_01101000), .b(t4_01101001), .y(t4_0110100));
wire t4_01101000, t4_01101001;
mixer mix_t4_01101000 (.a(t4_011010000), .b(t4_011010001), .y(t4_01101000));
wire t4_011010000, t4_011010001;
mixer mix_t4_01101001 (.a(t4_011010010), .b(t4_011010011), .y(t4_01101001));
wire t4_011010010, t4_011010011;
mixer mix_t4_0110101 (.a(t4_01101010), .b(t4_01101011), .y(t4_0110101));
wire t4_01101010, t4_01101011;
mixer mix_t4_01101010 (.a(t4_011010100), .b(t4_011010101), .y(t4_01101010));
wire t4_011010100, t4_011010101;
mixer mix_t4_01101011 (.a(t4_011010110), .b(t4_011010111), .y(t4_01101011));
wire t4_011010110, t4_011010111;
mixer mix_t4_011011 (.a(t4_0110110), .b(t4_0110111), .y(t4_011011));
wire t4_0110110, t4_0110111;
mixer mix_t4_0110110 (.a(t4_01101100), .b(t4_01101101), .y(t4_0110110));
wire t4_01101100, t4_01101101;
mixer mix_t4_01101100 (.a(t4_011011000), .b(t4_011011001), .y(t4_01101100));
wire t4_011011000, t4_011011001;
mixer mix_t4_01101101 (.a(t4_011011010), .b(t4_011011011), .y(t4_01101101));
wire t4_011011010, t4_011011011;
mixer mix_t4_0110111 (.a(t4_01101110), .b(t4_01101111), .y(t4_0110111));
wire t4_01101110, t4_01101111;
mixer mix_t4_01101110 (.a(t4_011011100), .b(t4_011011101), .y(t4_01101110));
wire t4_011011100, t4_011011101;
mixer mix_t4_01101111 (.a(t4_011011110), .b(t4_011011111), .y(t4_01101111));
wire t4_011011110, t4_011011111;
mixer mix_t4_0111 (.a(t4_01110), .b(t4_01111), .y(t4_0111));
wire t4_01110, t4_01111;
mixer mix_t4_01110 (.a(t4_011100), .b(t4_011101), .y(t4_01110));
wire t4_011100, t4_011101;
mixer mix_t4_011100 (.a(t4_0111000), .b(t4_0111001), .y(t4_011100));
wire t4_0111000, t4_0111001;
mixer mix_t4_0111000 (.a(t4_01110000), .b(t4_01110001), .y(t4_0111000));
wire t4_01110000, t4_01110001;
mixer mix_t4_01110000 (.a(t4_011100000), .b(t4_011100001), .y(t4_01110000));
wire t4_011100000, t4_011100001;
mixer mix_t4_01110001 (.a(t4_011100010), .b(t4_011100011), .y(t4_01110001));
wire t4_011100010, t4_011100011;
mixer mix_t4_0111001 (.a(t4_01110010), .b(t4_01110011), .y(t4_0111001));
wire t4_01110010, t4_01110011;
mixer mix_t4_01110010 (.a(t4_011100100), .b(t4_011100101), .y(t4_01110010));
wire t4_011100100, t4_011100101;
mixer mix_t4_01110011 (.a(t4_011100110), .b(t4_011100111), .y(t4_01110011));
wire t4_011100110, t4_011100111;
mixer mix_t4_011101 (.a(t4_0111010), .b(t4_0111011), .y(t4_011101));
wire t4_0111010, t4_0111011;
mixer mix_t4_0111010 (.a(t4_01110100), .b(t4_01110101), .y(t4_0111010));
wire t4_01110100, t4_01110101;
mixer mix_t4_01110100 (.a(t4_011101000), .b(t4_011101001), .y(t4_01110100));
wire t4_011101000, t4_011101001;
mixer mix_t4_01110101 (.a(t4_011101010), .b(t4_011101011), .y(t4_01110101));
wire t4_011101010, t4_011101011;
mixer mix_t4_0111011 (.a(t4_01110110), .b(t4_01110111), .y(t4_0111011));
wire t4_01110110, t4_01110111;
mixer mix_t4_01110110 (.a(t4_011101100), .b(t4_011101101), .y(t4_01110110));
wire t4_011101100, t4_011101101;
mixer mix_t4_01110111 (.a(t4_011101110), .b(t4_011101111), .y(t4_01110111));
wire t4_011101110, t4_011101111;
mixer mix_t4_01111 (.a(t4_011110), .b(t4_011111), .y(t4_01111));
wire t4_011110, t4_011111;
mixer mix_t4_011110 (.a(t4_0111100), .b(t4_0111101), .y(t4_011110));
wire t4_0111100, t4_0111101;
mixer mix_t4_0111100 (.a(t4_01111000), .b(t4_01111001), .y(t4_0111100));
wire t4_01111000, t4_01111001;
mixer mix_t4_01111000 (.a(t4_011110000), .b(t4_011110001), .y(t4_01111000));
wire t4_011110000, t4_011110001;
mixer mix_t4_01111001 (.a(t4_011110010), .b(t4_011110011), .y(t4_01111001));
wire t4_011110010, t4_011110011;
mixer mix_t4_0111101 (.a(t4_01111010), .b(t4_01111011), .y(t4_0111101));
wire t4_01111010, t4_01111011;
mixer mix_t4_01111010 (.a(t4_011110100), .b(t4_011110101), .y(t4_01111010));
wire t4_011110100, t4_011110101;
mixer mix_t4_01111011 (.a(t4_011110110), .b(t4_011110111), .y(t4_01111011));
wire t4_011110110, t4_011110111;
mixer mix_t4_011111 (.a(t4_0111110), .b(t4_0111111), .y(t4_011111));
wire t4_0111110, t4_0111111;
mixer mix_t4_0111110 (.a(t4_01111100), .b(t4_01111101), .y(t4_0111110));
wire t4_01111100, t4_01111101;
mixer mix_t4_01111100 (.a(t4_011111000), .b(t4_011111001), .y(t4_01111100));
wire t4_011111000, t4_011111001;
mixer mix_t4_01111101 (.a(t4_011111010), .b(t4_011111011), .y(t4_01111101));
wire t4_011111010, t4_011111011;
mixer mix_t4_0111111 (.a(t4_01111110), .b(t4_01111111), .y(t4_0111111));
wire t4_01111110, t4_01111111;
mixer mix_t4_01111110 (.a(t4_011111100), .b(t4_011111101), .y(t4_01111110));
wire t4_011111100, t4_011111101;
mixer mix_t4_01111111 (.a(t4_011111110), .b(t4_011111111), .y(t4_01111111));
wire t4_011111110, t4_011111111;
mixer mix_t5_0 (.a(t5_00), .b(t5_01), .y(t5_0));
wire t5_00, t5_01;
mixer mix_t5_00 (.a(t5_000), .b(t5_001), .y(t5_00));
wire t5_000, t5_001;
mixer mix_t5_000 (.a(t5_0000), .b(t5_0001), .y(t5_000));
wire t5_0000, t5_0001;
mixer mix_t5_0000 (.a(t5_00000), .b(t5_00001), .y(t5_0000));
wire t5_00000, t5_00001;
mixer mix_t5_00000 (.a(t5_000000), .b(t5_000001), .y(t5_00000));
wire t5_000000, t5_000001;
mixer mix_t5_000000 (.a(t5_0000000), .b(t5_0000001), .y(t5_000000));
wire t5_0000000, t5_0000001;
mixer mix_t5_0000000 (.a(t5_00000000), .b(t5_00000001), .y(t5_0000000));
wire t5_00000000, t5_00000001;
mixer mix_t5_00000000 (.a(t5_000000000), .b(t5_000000001), .y(t5_00000000));
wire t5_000000000, t5_000000001;
mixer mix_t5_00000001 (.a(t5_000000010), .b(t5_000000011), .y(t5_00000001));
wire t5_000000010, t5_000000011;
mixer mix_t5_0000001 (.a(t5_00000010), .b(t5_00000011), .y(t5_0000001));
wire t5_00000010, t5_00000011;
mixer mix_t5_00000010 (.a(t5_000000100), .b(t5_000000101), .y(t5_00000010));
wire t5_000000100, t5_000000101;
mixer mix_t5_00000011 (.a(t5_000000110), .b(t5_000000111), .y(t5_00000011));
wire t5_000000110, t5_000000111;
mixer mix_t5_000001 (.a(t5_0000010), .b(t5_0000011), .y(t5_000001));
wire t5_0000010, t5_0000011;
mixer mix_t5_0000010 (.a(t5_00000100), .b(t5_00000101), .y(t5_0000010));
wire t5_00000100, t5_00000101;
mixer mix_t5_00000100 (.a(t5_000001000), .b(t5_000001001), .y(t5_00000100));
wire t5_000001000, t5_000001001;
mixer mix_t5_00000101 (.a(t5_000001010), .b(t5_000001011), .y(t5_00000101));
wire t5_000001010, t5_000001011;
mixer mix_t5_0000011 (.a(t5_00000110), .b(t5_00000111), .y(t5_0000011));
wire t5_00000110, t5_00000111;
mixer mix_t5_00000110 (.a(t5_000001100), .b(t5_000001101), .y(t5_00000110));
wire t5_000001100, t5_000001101;
mixer mix_t5_00000111 (.a(t5_000001110), .b(t5_000001111), .y(t5_00000111));
wire t5_000001110, t5_000001111;
mixer mix_t5_00001 (.a(t5_000010), .b(t5_000011), .y(t5_00001));
wire t5_000010, t5_000011;
mixer mix_t5_000010 (.a(t5_0000100), .b(t5_0000101), .y(t5_000010));
wire t5_0000100, t5_0000101;
mixer mix_t5_0000100 (.a(t5_00001000), .b(t5_00001001), .y(t5_0000100));
wire t5_00001000, t5_00001001;
mixer mix_t5_00001000 (.a(t5_000010000), .b(t5_000010001), .y(t5_00001000));
wire t5_000010000, t5_000010001;
mixer mix_t5_00001001 (.a(t5_000010010), .b(t5_000010011), .y(t5_00001001));
wire t5_000010010, t5_000010011;
mixer mix_t5_0000101 (.a(t5_00001010), .b(t5_00001011), .y(t5_0000101));
wire t5_00001010, t5_00001011;
mixer mix_t5_00001010 (.a(t5_000010100), .b(t5_000010101), .y(t5_00001010));
wire t5_000010100, t5_000010101;
mixer mix_t5_00001011 (.a(t5_000010110), .b(t5_000010111), .y(t5_00001011));
wire t5_000010110, t5_000010111;
mixer mix_t5_000011 (.a(t5_0000110), .b(t5_0000111), .y(t5_000011));
wire t5_0000110, t5_0000111;
mixer mix_t5_0000110 (.a(t5_00001100), .b(t5_00001101), .y(t5_0000110));
wire t5_00001100, t5_00001101;
mixer mix_t5_00001100 (.a(t5_000011000), .b(t5_000011001), .y(t5_00001100));
wire t5_000011000, t5_000011001;
mixer mix_t5_00001101 (.a(t5_000011010), .b(t5_000011011), .y(t5_00001101));
wire t5_000011010, t5_000011011;
mixer mix_t5_0000111 (.a(t5_00001110), .b(t5_00001111), .y(t5_0000111));
wire t5_00001110, t5_00001111;
mixer mix_t5_00001110 (.a(t5_000011100), .b(t5_000011101), .y(t5_00001110));
wire t5_000011100, t5_000011101;
mixer mix_t5_00001111 (.a(t5_000011110), .b(t5_000011111), .y(t5_00001111));
wire t5_000011110, t5_000011111;
mixer mix_t5_0001 (.a(t5_00010), .b(t5_00011), .y(t5_0001));
wire t5_00010, t5_00011;
mixer mix_t5_00010 (.a(t5_000100), .b(t5_000101), .y(t5_00010));
wire t5_000100, t5_000101;
mixer mix_t5_000100 (.a(t5_0001000), .b(t5_0001001), .y(t5_000100));
wire t5_0001000, t5_0001001;
mixer mix_t5_0001000 (.a(t5_00010000), .b(t5_00010001), .y(t5_0001000));
wire t5_00010000, t5_00010001;
mixer mix_t5_00010000 (.a(t5_000100000), .b(t5_000100001), .y(t5_00010000));
wire t5_000100000, t5_000100001;
mixer mix_t5_00010001 (.a(t5_000100010), .b(t5_000100011), .y(t5_00010001));
wire t5_000100010, t5_000100011;
mixer mix_t5_0001001 (.a(t5_00010010), .b(t5_00010011), .y(t5_0001001));
wire t5_00010010, t5_00010011;
mixer mix_t5_00010010 (.a(t5_000100100), .b(t5_000100101), .y(t5_00010010));
wire t5_000100100, t5_000100101;
mixer mix_t5_00010011 (.a(t5_000100110), .b(t5_000100111), .y(t5_00010011));
wire t5_000100110, t5_000100111;
mixer mix_t5_000101 (.a(t5_0001010), .b(t5_0001011), .y(t5_000101));
wire t5_0001010, t5_0001011;
mixer mix_t5_0001010 (.a(t5_00010100), .b(t5_00010101), .y(t5_0001010));
wire t5_00010100, t5_00010101;
mixer mix_t5_00010100 (.a(t5_000101000), .b(t5_000101001), .y(t5_00010100));
wire t5_000101000, t5_000101001;
mixer mix_t5_00010101 (.a(t5_000101010), .b(t5_000101011), .y(t5_00010101));
wire t5_000101010, t5_000101011;
mixer mix_t5_0001011 (.a(t5_00010110), .b(t5_00010111), .y(t5_0001011));
wire t5_00010110, t5_00010111;
mixer mix_t5_00010110 (.a(t5_000101100), .b(t5_000101101), .y(t5_00010110));
wire t5_000101100, t5_000101101;
mixer mix_t5_00010111 (.a(t5_000101110), .b(t5_000101111), .y(t5_00010111));
wire t5_000101110, t5_000101111;
mixer mix_t5_00011 (.a(t5_000110), .b(t5_000111), .y(t5_00011));
wire t5_000110, t5_000111;
mixer mix_t5_000110 (.a(t5_0001100), .b(t5_0001101), .y(t5_000110));
wire t5_0001100, t5_0001101;
mixer mix_t5_0001100 (.a(t5_00011000), .b(t5_00011001), .y(t5_0001100));
wire t5_00011000, t5_00011001;
mixer mix_t5_00011000 (.a(t5_000110000), .b(t5_000110001), .y(t5_00011000));
wire t5_000110000, t5_000110001;
mixer mix_t5_00011001 (.a(t5_000110010), .b(t5_000110011), .y(t5_00011001));
wire t5_000110010, t5_000110011;
mixer mix_t5_0001101 (.a(t5_00011010), .b(t5_00011011), .y(t5_0001101));
wire t5_00011010, t5_00011011;
mixer mix_t5_00011010 (.a(t5_000110100), .b(t5_000110101), .y(t5_00011010));
wire t5_000110100, t5_000110101;
mixer mix_t5_00011011 (.a(t5_000110110), .b(t5_000110111), .y(t5_00011011));
wire t5_000110110, t5_000110111;
mixer mix_t5_000111 (.a(t5_0001110), .b(t5_0001111), .y(t5_000111));
wire t5_0001110, t5_0001111;
mixer mix_t5_0001110 (.a(t5_00011100), .b(t5_00011101), .y(t5_0001110));
wire t5_00011100, t5_00011101;
mixer mix_t5_00011100 (.a(t5_000111000), .b(t5_000111001), .y(t5_00011100));
wire t5_000111000, t5_000111001;
mixer mix_t5_00011101 (.a(t5_000111010), .b(t5_000111011), .y(t5_00011101));
wire t5_000111010, t5_000111011;
mixer mix_t5_0001111 (.a(t5_00011110), .b(t5_00011111), .y(t5_0001111));
wire t5_00011110, t5_00011111;
mixer mix_t5_00011110 (.a(t5_000111100), .b(t5_000111101), .y(t5_00011110));
wire t5_000111100, t5_000111101;
mixer mix_t5_00011111 (.a(t5_000111110), .b(t5_000111111), .y(t5_00011111));
wire t5_000111110, t5_000111111;
mixer mix_t5_001 (.a(t5_0010), .b(t5_0011), .y(t5_001));
wire t5_0010, t5_0011;
mixer mix_t5_0010 (.a(t5_00100), .b(t5_00101), .y(t5_0010));
wire t5_00100, t5_00101;
mixer mix_t5_00100 (.a(t5_001000), .b(t5_001001), .y(t5_00100));
wire t5_001000, t5_001001;
mixer mix_t5_001000 (.a(t5_0010000), .b(t5_0010001), .y(t5_001000));
wire t5_0010000, t5_0010001;
mixer mix_t5_0010000 (.a(t5_00100000), .b(t5_00100001), .y(t5_0010000));
wire t5_00100000, t5_00100001;
mixer mix_t5_00100000 (.a(t5_001000000), .b(t5_001000001), .y(t5_00100000));
wire t5_001000000, t5_001000001;
mixer mix_t5_00100001 (.a(t5_001000010), .b(t5_001000011), .y(t5_00100001));
wire t5_001000010, t5_001000011;
mixer mix_t5_0010001 (.a(t5_00100010), .b(t5_00100011), .y(t5_0010001));
wire t5_00100010, t5_00100011;
mixer mix_t5_00100010 (.a(t5_001000100), .b(t5_001000101), .y(t5_00100010));
wire t5_001000100, t5_001000101;
mixer mix_t5_00100011 (.a(t5_001000110), .b(t5_001000111), .y(t5_00100011));
wire t5_001000110, t5_001000111;
mixer mix_t5_001001 (.a(t5_0010010), .b(t5_0010011), .y(t5_001001));
wire t5_0010010, t5_0010011;
mixer mix_t5_0010010 (.a(t5_00100100), .b(t5_00100101), .y(t5_0010010));
wire t5_00100100, t5_00100101;
mixer mix_t5_00100100 (.a(t5_001001000), .b(t5_001001001), .y(t5_00100100));
wire t5_001001000, t5_001001001;
mixer mix_t5_00100101 (.a(t5_001001010), .b(t5_001001011), .y(t5_00100101));
wire t5_001001010, t5_001001011;
mixer mix_t5_0010011 (.a(t5_00100110), .b(t5_00100111), .y(t5_0010011));
wire t5_00100110, t5_00100111;
mixer mix_t5_00100110 (.a(t5_001001100), .b(t5_001001101), .y(t5_00100110));
wire t5_001001100, t5_001001101;
mixer mix_t5_00100111 (.a(t5_001001110), .b(t5_001001111), .y(t5_00100111));
wire t5_001001110, t5_001001111;
mixer mix_t5_00101 (.a(t5_001010), .b(t5_001011), .y(t5_00101));
wire t5_001010, t5_001011;
mixer mix_t5_001010 (.a(t5_0010100), .b(t5_0010101), .y(t5_001010));
wire t5_0010100, t5_0010101;
mixer mix_t5_0010100 (.a(t5_00101000), .b(t5_00101001), .y(t5_0010100));
wire t5_00101000, t5_00101001;
mixer mix_t5_00101000 (.a(t5_001010000), .b(t5_001010001), .y(t5_00101000));
wire t5_001010000, t5_001010001;
mixer mix_t5_00101001 (.a(t5_001010010), .b(t5_001010011), .y(t5_00101001));
wire t5_001010010, t5_001010011;
mixer mix_t5_0010101 (.a(t5_00101010), .b(t5_00101011), .y(t5_0010101));
wire t5_00101010, t5_00101011;
mixer mix_t5_00101010 (.a(t5_001010100), .b(t5_001010101), .y(t5_00101010));
wire t5_001010100, t5_001010101;
mixer mix_t5_00101011 (.a(t5_001010110), .b(t5_001010111), .y(t5_00101011));
wire t5_001010110, t5_001010111;
mixer mix_t5_001011 (.a(t5_0010110), .b(t5_0010111), .y(t5_001011));
wire t5_0010110, t5_0010111;
mixer mix_t5_0010110 (.a(t5_00101100), .b(t5_00101101), .y(t5_0010110));
wire t5_00101100, t5_00101101;
mixer mix_t5_00101100 (.a(t5_001011000), .b(t5_001011001), .y(t5_00101100));
wire t5_001011000, t5_001011001;
mixer mix_t5_00101101 (.a(t5_001011010), .b(t5_001011011), .y(t5_00101101));
wire t5_001011010, t5_001011011;
mixer mix_t5_0010111 (.a(t5_00101110), .b(t5_00101111), .y(t5_0010111));
wire t5_00101110, t5_00101111;
mixer mix_t5_00101110 (.a(t5_001011100), .b(t5_001011101), .y(t5_00101110));
wire t5_001011100, t5_001011101;
mixer mix_t5_00101111 (.a(t5_001011110), .b(t5_001011111), .y(t5_00101111));
wire t5_001011110, t5_001011111;
mixer mix_t5_0011 (.a(t5_00110), .b(t5_00111), .y(t5_0011));
wire t5_00110, t5_00111;
mixer mix_t5_00110 (.a(t5_001100), .b(t5_001101), .y(t5_00110));
wire t5_001100, t5_001101;
mixer mix_t5_001100 (.a(t5_0011000), .b(t5_0011001), .y(t5_001100));
wire t5_0011000, t5_0011001;
mixer mix_t5_0011000 (.a(t5_00110000), .b(t5_00110001), .y(t5_0011000));
wire t5_00110000, t5_00110001;
mixer mix_t5_00110000 (.a(t5_001100000), .b(t5_001100001), .y(t5_00110000));
wire t5_001100000, t5_001100001;
mixer mix_t5_00110001 (.a(t5_001100010), .b(t5_001100011), .y(t5_00110001));
wire t5_001100010, t5_001100011;
mixer mix_t5_0011001 (.a(t5_00110010), .b(t5_00110011), .y(t5_0011001));
wire t5_00110010, t5_00110011;
mixer mix_t5_00110010 (.a(t5_001100100), .b(t5_001100101), .y(t5_00110010));
wire t5_001100100, t5_001100101;
mixer mix_t5_00110011 (.a(t5_001100110), .b(t5_001100111), .y(t5_00110011));
wire t5_001100110, t5_001100111;
mixer mix_t5_001101 (.a(t5_0011010), .b(t5_0011011), .y(t5_001101));
wire t5_0011010, t5_0011011;
mixer mix_t5_0011010 (.a(t5_00110100), .b(t5_00110101), .y(t5_0011010));
wire t5_00110100, t5_00110101;
mixer mix_t5_00110100 (.a(t5_001101000), .b(t5_001101001), .y(t5_00110100));
wire t5_001101000, t5_001101001;
mixer mix_t5_00110101 (.a(t5_001101010), .b(t5_001101011), .y(t5_00110101));
wire t5_001101010, t5_001101011;
mixer mix_t5_0011011 (.a(t5_00110110), .b(t5_00110111), .y(t5_0011011));
wire t5_00110110, t5_00110111;
mixer mix_t5_00110110 (.a(t5_001101100), .b(t5_001101101), .y(t5_00110110));
wire t5_001101100, t5_001101101;
mixer mix_t5_00110111 (.a(t5_001101110), .b(t5_001101111), .y(t5_00110111));
wire t5_001101110, t5_001101111;
mixer mix_t5_00111 (.a(t5_001110), .b(t5_001111), .y(t5_00111));
wire t5_001110, t5_001111;
mixer mix_t5_001110 (.a(t5_0011100), .b(t5_0011101), .y(t5_001110));
wire t5_0011100, t5_0011101;
mixer mix_t5_0011100 (.a(t5_00111000), .b(t5_00111001), .y(t5_0011100));
wire t5_00111000, t5_00111001;
mixer mix_t5_00111000 (.a(t5_001110000), .b(t5_001110001), .y(t5_00111000));
wire t5_001110000, t5_001110001;
mixer mix_t5_00111001 (.a(t5_001110010), .b(t5_001110011), .y(t5_00111001));
wire t5_001110010, t5_001110011;
mixer mix_t5_0011101 (.a(t5_00111010), .b(t5_00111011), .y(t5_0011101));
wire t5_00111010, t5_00111011;
mixer mix_t5_00111010 (.a(t5_001110100), .b(t5_001110101), .y(t5_00111010));
wire t5_001110100, t5_001110101;
mixer mix_t5_00111011 (.a(t5_001110110), .b(t5_001110111), .y(t5_00111011));
wire t5_001110110, t5_001110111;
mixer mix_t5_001111 (.a(t5_0011110), .b(t5_0011111), .y(t5_001111));
wire t5_0011110, t5_0011111;
mixer mix_t5_0011110 (.a(t5_00111100), .b(t5_00111101), .y(t5_0011110));
wire t5_00111100, t5_00111101;
mixer mix_t5_00111100 (.a(t5_001111000), .b(t5_001111001), .y(t5_00111100));
wire t5_001111000, t5_001111001;
mixer mix_t5_00111101 (.a(t5_001111010), .b(t5_001111011), .y(t5_00111101));
wire t5_001111010, t5_001111011;
mixer mix_t5_0011111 (.a(t5_00111110), .b(t5_00111111), .y(t5_0011111));
wire t5_00111110, t5_00111111;
mixer mix_t5_00111110 (.a(t5_001111100), .b(t5_001111101), .y(t5_00111110));
wire t5_001111100, t5_001111101;
mixer mix_t5_00111111 (.a(t5_001111110), .b(t5_001111111), .y(t5_00111111));
wire t5_001111110, t5_001111111;
mixer mix_t5_01 (.a(t5_010), .b(t5_011), .y(t5_01));
wire t5_010, t5_011;
mixer mix_t5_010 (.a(t5_0100), .b(t5_0101), .y(t5_010));
wire t5_0100, t5_0101;
mixer mix_t5_0100 (.a(t5_01000), .b(t5_01001), .y(t5_0100));
wire t5_01000, t5_01001;
mixer mix_t5_01000 (.a(t5_010000), .b(t5_010001), .y(t5_01000));
wire t5_010000, t5_010001;
mixer mix_t5_010000 (.a(t5_0100000), .b(t5_0100001), .y(t5_010000));
wire t5_0100000, t5_0100001;
mixer mix_t5_0100000 (.a(t5_01000000), .b(t5_01000001), .y(t5_0100000));
wire t5_01000000, t5_01000001;
mixer mix_t5_01000000 (.a(t5_010000000), .b(t5_010000001), .y(t5_01000000));
wire t5_010000000, t5_010000001;
mixer mix_t5_01000001 (.a(t5_010000010), .b(t5_010000011), .y(t5_01000001));
wire t5_010000010, t5_010000011;
mixer mix_t5_0100001 (.a(t5_01000010), .b(t5_01000011), .y(t5_0100001));
wire t5_01000010, t5_01000011;
mixer mix_t5_01000010 (.a(t5_010000100), .b(t5_010000101), .y(t5_01000010));
wire t5_010000100, t5_010000101;
mixer mix_t5_01000011 (.a(t5_010000110), .b(t5_010000111), .y(t5_01000011));
wire t5_010000110, t5_010000111;
mixer mix_t5_010001 (.a(t5_0100010), .b(t5_0100011), .y(t5_010001));
wire t5_0100010, t5_0100011;
mixer mix_t5_0100010 (.a(t5_01000100), .b(t5_01000101), .y(t5_0100010));
wire t5_01000100, t5_01000101;
mixer mix_t5_01000100 (.a(t5_010001000), .b(t5_010001001), .y(t5_01000100));
wire t5_010001000, t5_010001001;
mixer mix_t5_01000101 (.a(t5_010001010), .b(t5_010001011), .y(t5_01000101));
wire t5_010001010, t5_010001011;
mixer mix_t5_0100011 (.a(t5_01000110), .b(t5_01000111), .y(t5_0100011));
wire t5_01000110, t5_01000111;
mixer mix_t5_01000110 (.a(t5_010001100), .b(t5_010001101), .y(t5_01000110));
wire t5_010001100, t5_010001101;
mixer mix_t5_01000111 (.a(t5_010001110), .b(t5_010001111), .y(t5_01000111));
wire t5_010001110, t5_010001111;
mixer mix_t5_01001 (.a(t5_010010), .b(t5_010011), .y(t5_01001));
wire t5_010010, t5_010011;
mixer mix_t5_010010 (.a(t5_0100100), .b(t5_0100101), .y(t5_010010));
wire t5_0100100, t5_0100101;
mixer mix_t5_0100100 (.a(t5_01001000), .b(t5_01001001), .y(t5_0100100));
wire t5_01001000, t5_01001001;
mixer mix_t5_01001000 (.a(t5_010010000), .b(t5_010010001), .y(t5_01001000));
wire t5_010010000, t5_010010001;
mixer mix_t5_01001001 (.a(t5_010010010), .b(t5_010010011), .y(t5_01001001));
wire t5_010010010, t5_010010011;
mixer mix_t5_0100101 (.a(t5_01001010), .b(t5_01001011), .y(t5_0100101));
wire t5_01001010, t5_01001011;
mixer mix_t5_01001010 (.a(t5_010010100), .b(t5_010010101), .y(t5_01001010));
wire t5_010010100, t5_010010101;
mixer mix_t5_01001011 (.a(t5_010010110), .b(t5_010010111), .y(t5_01001011));
wire t5_010010110, t5_010010111;
mixer mix_t5_010011 (.a(t5_0100110), .b(t5_0100111), .y(t5_010011));
wire t5_0100110, t5_0100111;
mixer mix_t5_0100110 (.a(t5_01001100), .b(t5_01001101), .y(t5_0100110));
wire t5_01001100, t5_01001101;
mixer mix_t5_01001100 (.a(t5_010011000), .b(t5_010011001), .y(t5_01001100));
wire t5_010011000, t5_010011001;
mixer mix_t5_01001101 (.a(t5_010011010), .b(t5_010011011), .y(t5_01001101));
wire t5_010011010, t5_010011011;
mixer mix_t5_0100111 (.a(t5_01001110), .b(t5_01001111), .y(t5_0100111));
wire t5_01001110, t5_01001111;
mixer mix_t5_01001110 (.a(t5_010011100), .b(t5_010011101), .y(t5_01001110));
wire t5_010011100, t5_010011101;
mixer mix_t5_01001111 (.a(t5_010011110), .b(t5_010011111), .y(t5_01001111));
wire t5_010011110, t5_010011111;
mixer mix_t5_0101 (.a(t5_01010), .b(t5_01011), .y(t5_0101));
wire t5_01010, t5_01011;
mixer mix_t5_01010 (.a(t5_010100), .b(t5_010101), .y(t5_01010));
wire t5_010100, t5_010101;
mixer mix_t5_010100 (.a(t5_0101000), .b(t5_0101001), .y(t5_010100));
wire t5_0101000, t5_0101001;
mixer mix_t5_0101000 (.a(t5_01010000), .b(t5_01010001), .y(t5_0101000));
wire t5_01010000, t5_01010001;
mixer mix_t5_01010000 (.a(t5_010100000), .b(t5_010100001), .y(t5_01010000));
wire t5_010100000, t5_010100001;
mixer mix_t5_01010001 (.a(t5_010100010), .b(t5_010100011), .y(t5_01010001));
wire t5_010100010, t5_010100011;
mixer mix_t5_0101001 (.a(t5_01010010), .b(t5_01010011), .y(t5_0101001));
wire t5_01010010, t5_01010011;
mixer mix_t5_01010010 (.a(t5_010100100), .b(t5_010100101), .y(t5_01010010));
wire t5_010100100, t5_010100101;
mixer mix_t5_01010011 (.a(t5_010100110), .b(t5_010100111), .y(t5_01010011));
wire t5_010100110, t5_010100111;
mixer mix_t5_010101 (.a(t5_0101010), .b(t5_0101011), .y(t5_010101));
wire t5_0101010, t5_0101011;
mixer mix_t5_0101010 (.a(t5_01010100), .b(t5_01010101), .y(t5_0101010));
wire t5_01010100, t5_01010101;
mixer mix_t5_01010100 (.a(t5_010101000), .b(t5_010101001), .y(t5_01010100));
wire t5_010101000, t5_010101001;
mixer mix_t5_01010101 (.a(t5_010101010), .b(t5_010101011), .y(t5_01010101));
wire t5_010101010, t5_010101011;
mixer mix_t5_0101011 (.a(t5_01010110), .b(t5_01010111), .y(t5_0101011));
wire t5_01010110, t5_01010111;
mixer mix_t5_01010110 (.a(t5_010101100), .b(t5_010101101), .y(t5_01010110));
wire t5_010101100, t5_010101101;
mixer mix_t5_01010111 (.a(t5_010101110), .b(t5_010101111), .y(t5_01010111));
wire t5_010101110, t5_010101111;
mixer mix_t5_01011 (.a(t5_010110), .b(t5_010111), .y(t5_01011));
wire t5_010110, t5_010111;
mixer mix_t5_010110 (.a(t5_0101100), .b(t5_0101101), .y(t5_010110));
wire t5_0101100, t5_0101101;
mixer mix_t5_0101100 (.a(t5_01011000), .b(t5_01011001), .y(t5_0101100));
wire t5_01011000, t5_01011001;
mixer mix_t5_01011000 (.a(t5_010110000), .b(t5_010110001), .y(t5_01011000));
wire t5_010110000, t5_010110001;
mixer mix_t5_01011001 (.a(t5_010110010), .b(t5_010110011), .y(t5_01011001));
wire t5_010110010, t5_010110011;
mixer mix_t5_0101101 (.a(t5_01011010), .b(t5_01011011), .y(t5_0101101));
wire t5_01011010, t5_01011011;
mixer mix_t5_01011010 (.a(t5_010110100), .b(t5_010110101), .y(t5_01011010));
wire t5_010110100, t5_010110101;
mixer mix_t5_01011011 (.a(t5_010110110), .b(t5_010110111), .y(t5_01011011));
wire t5_010110110, t5_010110111;
mixer mix_t5_010111 (.a(t5_0101110), .b(t5_0101111), .y(t5_010111));
wire t5_0101110, t5_0101111;
mixer mix_t5_0101110 (.a(t5_01011100), .b(t5_01011101), .y(t5_0101110));
wire t5_01011100, t5_01011101;
mixer mix_t5_01011100 (.a(t5_010111000), .b(t5_010111001), .y(t5_01011100));
wire t5_010111000, t5_010111001;
mixer mix_t5_01011101 (.a(t5_010111010), .b(t5_010111011), .y(t5_01011101));
wire t5_010111010, t5_010111011;
mixer mix_t5_0101111 (.a(t5_01011110), .b(t5_01011111), .y(t5_0101111));
wire t5_01011110, t5_01011111;
mixer mix_t5_01011110 (.a(t5_010111100), .b(t5_010111101), .y(t5_01011110));
wire t5_010111100, t5_010111101;
mixer mix_t5_01011111 (.a(t5_010111110), .b(t5_010111111), .y(t5_01011111));
wire t5_010111110, t5_010111111;
mixer mix_t5_011 (.a(t5_0110), .b(t5_0111), .y(t5_011));
wire t5_0110, t5_0111;
mixer mix_t5_0110 (.a(t5_01100), .b(t5_01101), .y(t5_0110));
wire t5_01100, t5_01101;
mixer mix_t5_01100 (.a(t5_011000), .b(t5_011001), .y(t5_01100));
wire t5_011000, t5_011001;
mixer mix_t5_011000 (.a(t5_0110000), .b(t5_0110001), .y(t5_011000));
wire t5_0110000, t5_0110001;
mixer mix_t5_0110000 (.a(t5_01100000), .b(t5_01100001), .y(t5_0110000));
wire t5_01100000, t5_01100001;
mixer mix_t5_01100000 (.a(t5_011000000), .b(t5_011000001), .y(t5_01100000));
wire t5_011000000, t5_011000001;
mixer mix_t5_01100001 (.a(t5_011000010), .b(t5_011000011), .y(t5_01100001));
wire t5_011000010, t5_011000011;
mixer mix_t5_0110001 (.a(t5_01100010), .b(t5_01100011), .y(t5_0110001));
wire t5_01100010, t5_01100011;
mixer mix_t5_01100010 (.a(t5_011000100), .b(t5_011000101), .y(t5_01100010));
wire t5_011000100, t5_011000101;
mixer mix_t5_01100011 (.a(t5_011000110), .b(t5_011000111), .y(t5_01100011));
wire t5_011000110, t5_011000111;
mixer mix_t5_011001 (.a(t5_0110010), .b(t5_0110011), .y(t5_011001));
wire t5_0110010, t5_0110011;
mixer mix_t5_0110010 (.a(t5_01100100), .b(t5_01100101), .y(t5_0110010));
wire t5_01100100, t5_01100101;
mixer mix_t5_01100100 (.a(t5_011001000), .b(t5_011001001), .y(t5_01100100));
wire t5_011001000, t5_011001001;
mixer mix_t5_01100101 (.a(t5_011001010), .b(t5_011001011), .y(t5_01100101));
wire t5_011001010, t5_011001011;
mixer mix_t5_0110011 (.a(t5_01100110), .b(t5_01100111), .y(t5_0110011));
wire t5_01100110, t5_01100111;
mixer mix_t5_01100110 (.a(t5_011001100), .b(t5_011001101), .y(t5_01100110));
wire t5_011001100, t5_011001101;
mixer mix_t5_01100111 (.a(t5_011001110), .b(t5_011001111), .y(t5_01100111));
wire t5_011001110, t5_011001111;
mixer mix_t5_01101 (.a(t5_011010), .b(t5_011011), .y(t5_01101));
wire t5_011010, t5_011011;
mixer mix_t5_011010 (.a(t5_0110100), .b(t5_0110101), .y(t5_011010));
wire t5_0110100, t5_0110101;
mixer mix_t5_0110100 (.a(t5_01101000), .b(t5_01101001), .y(t5_0110100));
wire t5_01101000, t5_01101001;
mixer mix_t5_01101000 (.a(t5_011010000), .b(t5_011010001), .y(t5_01101000));
wire t5_011010000, t5_011010001;
mixer mix_t5_01101001 (.a(t5_011010010), .b(t5_011010011), .y(t5_01101001));
wire t5_011010010, t5_011010011;
mixer mix_t5_0110101 (.a(t5_01101010), .b(t5_01101011), .y(t5_0110101));
wire t5_01101010, t5_01101011;
mixer mix_t5_01101010 (.a(t5_011010100), .b(t5_011010101), .y(t5_01101010));
wire t5_011010100, t5_011010101;
mixer mix_t5_01101011 (.a(t5_011010110), .b(t5_011010111), .y(t5_01101011));
wire t5_011010110, t5_011010111;
mixer mix_t5_011011 (.a(t5_0110110), .b(t5_0110111), .y(t5_011011));
wire t5_0110110, t5_0110111;
mixer mix_t5_0110110 (.a(t5_01101100), .b(t5_01101101), .y(t5_0110110));
wire t5_01101100, t5_01101101;
mixer mix_t5_01101100 (.a(t5_011011000), .b(t5_011011001), .y(t5_01101100));
wire t5_011011000, t5_011011001;
mixer mix_t5_01101101 (.a(t5_011011010), .b(t5_011011011), .y(t5_01101101));
wire t5_011011010, t5_011011011;
mixer mix_t5_0110111 (.a(t5_01101110), .b(t5_01101111), .y(t5_0110111));
wire t5_01101110, t5_01101111;
mixer mix_t5_01101110 (.a(t5_011011100), .b(t5_011011101), .y(t5_01101110));
wire t5_011011100, t5_011011101;
mixer mix_t5_01101111 (.a(t5_011011110), .b(t5_011011111), .y(t5_01101111));
wire t5_011011110, t5_011011111;
mixer mix_t5_0111 (.a(t5_01110), .b(t5_01111), .y(t5_0111));
wire t5_01110, t5_01111;
mixer mix_t5_01110 (.a(t5_011100), .b(t5_011101), .y(t5_01110));
wire t5_011100, t5_011101;
mixer mix_t5_011100 (.a(t5_0111000), .b(t5_0111001), .y(t5_011100));
wire t5_0111000, t5_0111001;
mixer mix_t5_0111000 (.a(t5_01110000), .b(t5_01110001), .y(t5_0111000));
wire t5_01110000, t5_01110001;
mixer mix_t5_01110000 (.a(t5_011100000), .b(t5_011100001), .y(t5_01110000));
wire t5_011100000, t5_011100001;
mixer mix_t5_01110001 (.a(t5_011100010), .b(t5_011100011), .y(t5_01110001));
wire t5_011100010, t5_011100011;
mixer mix_t5_0111001 (.a(t5_01110010), .b(t5_01110011), .y(t5_0111001));
wire t5_01110010, t5_01110011;
mixer mix_t5_01110010 (.a(t5_011100100), .b(t5_011100101), .y(t5_01110010));
wire t5_011100100, t5_011100101;
mixer mix_t5_01110011 (.a(t5_011100110), .b(t5_011100111), .y(t5_01110011));
wire t5_011100110, t5_011100111;
mixer mix_t5_011101 (.a(t5_0111010), .b(t5_0111011), .y(t5_011101));
wire t5_0111010, t5_0111011;
mixer mix_t5_0111010 (.a(t5_01110100), .b(t5_01110101), .y(t5_0111010));
wire t5_01110100, t5_01110101;
mixer mix_t5_01110100 (.a(t5_011101000), .b(t5_011101001), .y(t5_01110100));
wire t5_011101000, t5_011101001;
mixer mix_t5_01110101 (.a(t5_011101010), .b(t5_011101011), .y(t5_01110101));
wire t5_011101010, t5_011101011;
mixer mix_t5_0111011 (.a(t5_01110110), .b(t5_01110111), .y(t5_0111011));
wire t5_01110110, t5_01110111;
mixer mix_t5_01110110 (.a(t5_011101100), .b(t5_011101101), .y(t5_01110110));
wire t5_011101100, t5_011101101;
mixer mix_t5_01110111 (.a(t5_011101110), .b(t5_011101111), .y(t5_01110111));
wire t5_011101110, t5_011101111;
mixer mix_t5_01111 (.a(t5_011110), .b(t5_011111), .y(t5_01111));
wire t5_011110, t5_011111;
mixer mix_t5_011110 (.a(t5_0111100), .b(t5_0111101), .y(t5_011110));
wire t5_0111100, t5_0111101;
mixer mix_t5_0111100 (.a(t5_01111000), .b(t5_01111001), .y(t5_0111100));
wire t5_01111000, t5_01111001;
mixer mix_t5_01111000 (.a(t5_011110000), .b(t5_011110001), .y(t5_01111000));
wire t5_011110000, t5_011110001;
mixer mix_t5_01111001 (.a(t5_011110010), .b(t5_011110011), .y(t5_01111001));
wire t5_011110010, t5_011110011;
mixer mix_t5_0111101 (.a(t5_01111010), .b(t5_01111011), .y(t5_0111101));
wire t5_01111010, t5_01111011;
mixer mix_t5_01111010 (.a(t5_011110100), .b(t5_011110101), .y(t5_01111010));
wire t5_011110100, t5_011110101;
mixer mix_t5_01111011 (.a(t5_011110110), .b(t5_011110111), .y(t5_01111011));
wire t5_011110110, t5_011110111;
mixer mix_t5_011111 (.a(t5_0111110), .b(t5_0111111), .y(t5_011111));
wire t5_0111110, t5_0111111;
mixer mix_t5_0111110 (.a(t5_01111100), .b(t5_01111101), .y(t5_0111110));
wire t5_01111100, t5_01111101;
mixer mix_t5_01111100 (.a(t5_011111000), .b(t5_011111001), .y(t5_01111100));
wire t5_011111000, t5_011111001;
mixer mix_t5_01111101 (.a(t5_011111010), .b(t5_011111011), .y(t5_01111101));
wire t5_011111010, t5_011111011;
mixer mix_t5_0111111 (.a(t5_01111110), .b(t5_01111111), .y(t5_0111111));
wire t5_01111110, t5_01111111;
mixer mix_t5_01111110 (.a(t5_011111100), .b(t5_011111101), .y(t5_01111110));
wire t5_011111100, t5_011111101;
mixer mix_t5_01111111 (.a(t5_011111110), .b(t5_011111111), .y(t5_01111111));
wire t5_011111110, t5_011111111;
mixer mix_t6_0 (.a(t6_00), .b(t6_01), .y(t6_0));
wire t6_00, t6_01;
mixer mix_t6_00 (.a(t6_000), .b(t6_001), .y(t6_00));
wire t6_000, t6_001;
mixer mix_t6_000 (.a(t6_0000), .b(t6_0001), .y(t6_000));
wire t6_0000, t6_0001;
mixer mix_t6_0000 (.a(t6_00000), .b(t6_00001), .y(t6_0000));
wire t6_00000, t6_00001;
mixer mix_t6_00000 (.a(t6_000000), .b(t6_000001), .y(t6_00000));
wire t6_000000, t6_000001;
mixer mix_t6_000000 (.a(t6_0000000), .b(t6_0000001), .y(t6_000000));
wire t6_0000000, t6_0000001;
mixer mix_t6_0000000 (.a(t6_00000000), .b(t6_00000001), .y(t6_0000000));
wire t6_00000000, t6_00000001;
mixer mix_t6_00000000 (.a(t6_000000000), .b(t6_000000001), .y(t6_00000000));
wire t6_000000000, t6_000000001;
mixer mix_t6_00000001 (.a(t6_000000010), .b(t6_000000011), .y(t6_00000001));
wire t6_000000010, t6_000000011;
mixer mix_t6_0000001 (.a(t6_00000010), .b(t6_00000011), .y(t6_0000001));
wire t6_00000010, t6_00000011;
mixer mix_t6_00000010 (.a(t6_000000100), .b(t6_000000101), .y(t6_00000010));
wire t6_000000100, t6_000000101;
mixer mix_t6_00000011 (.a(t6_000000110), .b(t6_000000111), .y(t6_00000011));
wire t6_000000110, t6_000000111;
mixer mix_t6_000001 (.a(t6_0000010), .b(t6_0000011), .y(t6_000001));
wire t6_0000010, t6_0000011;
mixer mix_t6_0000010 (.a(t6_00000100), .b(t6_00000101), .y(t6_0000010));
wire t6_00000100, t6_00000101;
mixer mix_t6_00000100 (.a(t6_000001000), .b(t6_000001001), .y(t6_00000100));
wire t6_000001000, t6_000001001;
mixer mix_t6_00000101 (.a(t6_000001010), .b(t6_000001011), .y(t6_00000101));
wire t6_000001010, t6_000001011;
mixer mix_t6_0000011 (.a(t6_00000110), .b(t6_00000111), .y(t6_0000011));
wire t6_00000110, t6_00000111;
mixer mix_t6_00000110 (.a(t6_000001100), .b(t6_000001101), .y(t6_00000110));
wire t6_000001100, t6_000001101;
mixer mix_t6_00000111 (.a(t6_000001110), .b(t6_000001111), .y(t6_00000111));
wire t6_000001110, t6_000001111;
mixer mix_t6_00001 (.a(t6_000010), .b(t6_000011), .y(t6_00001));
wire t6_000010, t6_000011;
mixer mix_t6_000010 (.a(t6_0000100), .b(t6_0000101), .y(t6_000010));
wire t6_0000100, t6_0000101;
mixer mix_t6_0000100 (.a(t6_00001000), .b(t6_00001001), .y(t6_0000100));
wire t6_00001000, t6_00001001;
mixer mix_t6_00001000 (.a(t6_000010000), .b(t6_000010001), .y(t6_00001000));
wire t6_000010000, t6_000010001;
mixer mix_t6_00001001 (.a(t6_000010010), .b(t6_000010011), .y(t6_00001001));
wire t6_000010010, t6_000010011;
mixer mix_t6_0000101 (.a(t6_00001010), .b(t6_00001011), .y(t6_0000101));
wire t6_00001010, t6_00001011;
mixer mix_t6_00001010 (.a(t6_000010100), .b(t6_000010101), .y(t6_00001010));
wire t6_000010100, t6_000010101;
mixer mix_t6_00001011 (.a(t6_000010110), .b(t6_000010111), .y(t6_00001011));
wire t6_000010110, t6_000010111;
mixer mix_t6_000011 (.a(t6_0000110), .b(t6_0000111), .y(t6_000011));
wire t6_0000110, t6_0000111;
mixer mix_t6_0000110 (.a(t6_00001100), .b(t6_00001101), .y(t6_0000110));
wire t6_00001100, t6_00001101;
mixer mix_t6_00001100 (.a(t6_000011000), .b(t6_000011001), .y(t6_00001100));
wire t6_000011000, t6_000011001;
mixer mix_t6_00001101 (.a(t6_000011010), .b(t6_000011011), .y(t6_00001101));
wire t6_000011010, t6_000011011;
mixer mix_t6_0000111 (.a(t6_00001110), .b(t6_00001111), .y(t6_0000111));
wire t6_00001110, t6_00001111;
mixer mix_t6_00001110 (.a(t6_000011100), .b(t6_000011101), .y(t6_00001110));
wire t6_000011100, t6_000011101;
mixer mix_t6_00001111 (.a(t6_000011110), .b(t6_000011111), .y(t6_00001111));
wire t6_000011110, t6_000011111;
mixer mix_t6_0001 (.a(t6_00010), .b(t6_00011), .y(t6_0001));
wire t6_00010, t6_00011;
mixer mix_t6_00010 (.a(t6_000100), .b(t6_000101), .y(t6_00010));
wire t6_000100, t6_000101;
mixer mix_t6_000100 (.a(t6_0001000), .b(t6_0001001), .y(t6_000100));
wire t6_0001000, t6_0001001;
mixer mix_t6_0001000 (.a(t6_00010000), .b(t6_00010001), .y(t6_0001000));
wire t6_00010000, t6_00010001;
mixer mix_t6_00010000 (.a(t6_000100000), .b(t6_000100001), .y(t6_00010000));
wire t6_000100000, t6_000100001;
mixer mix_t6_00010001 (.a(t6_000100010), .b(t6_000100011), .y(t6_00010001));
wire t6_000100010, t6_000100011;
mixer mix_t6_0001001 (.a(t6_00010010), .b(t6_00010011), .y(t6_0001001));
wire t6_00010010, t6_00010011;
mixer mix_t6_00010010 (.a(t6_000100100), .b(t6_000100101), .y(t6_00010010));
wire t6_000100100, t6_000100101;
mixer mix_t6_00010011 (.a(t6_000100110), .b(t6_000100111), .y(t6_00010011));
wire t6_000100110, t6_000100111;
mixer mix_t6_000101 (.a(t6_0001010), .b(t6_0001011), .y(t6_000101));
wire t6_0001010, t6_0001011;
mixer mix_t6_0001010 (.a(t6_00010100), .b(t6_00010101), .y(t6_0001010));
wire t6_00010100, t6_00010101;
mixer mix_t6_00010100 (.a(t6_000101000), .b(t6_000101001), .y(t6_00010100));
wire t6_000101000, t6_000101001;
mixer mix_t6_00010101 (.a(t6_000101010), .b(t6_000101011), .y(t6_00010101));
wire t6_000101010, t6_000101011;
mixer mix_t6_0001011 (.a(t6_00010110), .b(t6_00010111), .y(t6_0001011));
wire t6_00010110, t6_00010111;
mixer mix_t6_00010110 (.a(t6_000101100), .b(t6_000101101), .y(t6_00010110));
wire t6_000101100, t6_000101101;
mixer mix_t6_00010111 (.a(t6_000101110), .b(t6_000101111), .y(t6_00010111));
wire t6_000101110, t6_000101111;
mixer mix_t6_00011 (.a(t6_000110), .b(t6_000111), .y(t6_00011));
wire t6_000110, t6_000111;
mixer mix_t6_000110 (.a(t6_0001100), .b(t6_0001101), .y(t6_000110));
wire t6_0001100, t6_0001101;
mixer mix_t6_0001100 (.a(t6_00011000), .b(t6_00011001), .y(t6_0001100));
wire t6_00011000, t6_00011001;
mixer mix_t6_00011000 (.a(t6_000110000), .b(t6_000110001), .y(t6_00011000));
wire t6_000110000, t6_000110001;
mixer mix_t6_00011001 (.a(t6_000110010), .b(t6_000110011), .y(t6_00011001));
wire t6_000110010, t6_000110011;
mixer mix_t6_0001101 (.a(t6_00011010), .b(t6_00011011), .y(t6_0001101));
wire t6_00011010, t6_00011011;
mixer mix_t6_00011010 (.a(t6_000110100), .b(t6_000110101), .y(t6_00011010));
wire t6_000110100, t6_000110101;
mixer mix_t6_00011011 (.a(t6_000110110), .b(t6_000110111), .y(t6_00011011));
wire t6_000110110, t6_000110111;
mixer mix_t6_000111 (.a(t6_0001110), .b(t6_0001111), .y(t6_000111));
wire t6_0001110, t6_0001111;
mixer mix_t6_0001110 (.a(t6_00011100), .b(t6_00011101), .y(t6_0001110));
wire t6_00011100, t6_00011101;
mixer mix_t6_00011100 (.a(t6_000111000), .b(t6_000111001), .y(t6_00011100));
wire t6_000111000, t6_000111001;
mixer mix_t6_00011101 (.a(t6_000111010), .b(t6_000111011), .y(t6_00011101));
wire t6_000111010, t6_000111011;
mixer mix_t6_0001111 (.a(t6_00011110), .b(t6_00011111), .y(t6_0001111));
wire t6_00011110, t6_00011111;
mixer mix_t6_00011110 (.a(t6_000111100), .b(t6_000111101), .y(t6_00011110));
wire t6_000111100, t6_000111101;
mixer mix_t6_00011111 (.a(t6_000111110), .b(t6_000111111), .y(t6_00011111));
wire t6_000111110, t6_000111111;
mixer mix_t6_001 (.a(t6_0010), .b(t6_0011), .y(t6_001));
wire t6_0010, t6_0011;
mixer mix_t6_0010 (.a(t6_00100), .b(t6_00101), .y(t6_0010));
wire t6_00100, t6_00101;
mixer mix_t6_00100 (.a(t6_001000), .b(t6_001001), .y(t6_00100));
wire t6_001000, t6_001001;
mixer mix_t6_001000 (.a(t6_0010000), .b(t6_0010001), .y(t6_001000));
wire t6_0010000, t6_0010001;
mixer mix_t6_0010000 (.a(t6_00100000), .b(t6_00100001), .y(t6_0010000));
wire t6_00100000, t6_00100001;
mixer mix_t6_00100000 (.a(t6_001000000), .b(t6_001000001), .y(t6_00100000));
wire t6_001000000, t6_001000001;
mixer mix_t6_00100001 (.a(t6_001000010), .b(t6_001000011), .y(t6_00100001));
wire t6_001000010, t6_001000011;
mixer mix_t6_0010001 (.a(t6_00100010), .b(t6_00100011), .y(t6_0010001));
wire t6_00100010, t6_00100011;
mixer mix_t6_00100010 (.a(t6_001000100), .b(t6_001000101), .y(t6_00100010));
wire t6_001000100, t6_001000101;
mixer mix_t6_00100011 (.a(t6_001000110), .b(t6_001000111), .y(t6_00100011));
wire t6_001000110, t6_001000111;
mixer mix_t6_001001 (.a(t6_0010010), .b(t6_0010011), .y(t6_001001));
wire t6_0010010, t6_0010011;
mixer mix_t6_0010010 (.a(t6_00100100), .b(t6_00100101), .y(t6_0010010));
wire t6_00100100, t6_00100101;
mixer mix_t6_00100100 (.a(t6_001001000), .b(t6_001001001), .y(t6_00100100));
wire t6_001001000, t6_001001001;
mixer mix_t6_00100101 (.a(t6_001001010), .b(t6_001001011), .y(t6_00100101));
wire t6_001001010, t6_001001011;
mixer mix_t6_0010011 (.a(t6_00100110), .b(t6_00100111), .y(t6_0010011));
wire t6_00100110, t6_00100111;
mixer mix_t6_00100110 (.a(t6_001001100), .b(t6_001001101), .y(t6_00100110));
wire t6_001001100, t6_001001101;
mixer mix_t6_00100111 (.a(t6_001001110), .b(t6_001001111), .y(t6_00100111));
wire t6_001001110, t6_001001111;
mixer mix_t6_00101 (.a(t6_001010), .b(t6_001011), .y(t6_00101));
wire t6_001010, t6_001011;
mixer mix_t6_001010 (.a(t6_0010100), .b(t6_0010101), .y(t6_001010));
wire t6_0010100, t6_0010101;
mixer mix_t6_0010100 (.a(t6_00101000), .b(t6_00101001), .y(t6_0010100));
wire t6_00101000, t6_00101001;
mixer mix_t6_00101000 (.a(t6_001010000), .b(t6_001010001), .y(t6_00101000));
wire t6_001010000, t6_001010001;
mixer mix_t6_00101001 (.a(t6_001010010), .b(t6_001010011), .y(t6_00101001));
wire t6_001010010, t6_001010011;
mixer mix_t6_0010101 (.a(t6_00101010), .b(t6_00101011), .y(t6_0010101));
wire t6_00101010, t6_00101011;
mixer mix_t6_00101010 (.a(t6_001010100), .b(t6_001010101), .y(t6_00101010));
wire t6_001010100, t6_001010101;
mixer mix_t6_00101011 (.a(t6_001010110), .b(t6_001010111), .y(t6_00101011));
wire t6_001010110, t6_001010111;
mixer mix_t6_001011 (.a(t6_0010110), .b(t6_0010111), .y(t6_001011));
wire t6_0010110, t6_0010111;
mixer mix_t6_0010110 (.a(t6_00101100), .b(t6_00101101), .y(t6_0010110));
wire t6_00101100, t6_00101101;
mixer mix_t6_00101100 (.a(t6_001011000), .b(t6_001011001), .y(t6_00101100));
wire t6_001011000, t6_001011001;
mixer mix_t6_00101101 (.a(t6_001011010), .b(t6_001011011), .y(t6_00101101));
wire t6_001011010, t6_001011011;
mixer mix_t6_0010111 (.a(t6_00101110), .b(t6_00101111), .y(t6_0010111));
wire t6_00101110, t6_00101111;
mixer mix_t6_00101110 (.a(t6_001011100), .b(t6_001011101), .y(t6_00101110));
wire t6_001011100, t6_001011101;
mixer mix_t6_00101111 (.a(t6_001011110), .b(t6_001011111), .y(t6_00101111));
wire t6_001011110, t6_001011111;
mixer mix_t6_0011 (.a(t6_00110), .b(t6_00111), .y(t6_0011));
wire t6_00110, t6_00111;
mixer mix_t6_00110 (.a(t6_001100), .b(t6_001101), .y(t6_00110));
wire t6_001100, t6_001101;
mixer mix_t6_001100 (.a(t6_0011000), .b(t6_0011001), .y(t6_001100));
wire t6_0011000, t6_0011001;
mixer mix_t6_0011000 (.a(t6_00110000), .b(t6_00110001), .y(t6_0011000));
wire t6_00110000, t6_00110001;
mixer mix_t6_00110000 (.a(t6_001100000), .b(t6_001100001), .y(t6_00110000));
wire t6_001100000, t6_001100001;
mixer mix_t6_00110001 (.a(t6_001100010), .b(t6_001100011), .y(t6_00110001));
wire t6_001100010, t6_001100011;
mixer mix_t6_0011001 (.a(t6_00110010), .b(t6_00110011), .y(t6_0011001));
wire t6_00110010, t6_00110011;
mixer mix_t6_00110010 (.a(t6_001100100), .b(t6_001100101), .y(t6_00110010));
wire t6_001100100, t6_001100101;
mixer mix_t6_00110011 (.a(t6_001100110), .b(t6_001100111), .y(t6_00110011));
wire t6_001100110, t6_001100111;
mixer mix_t6_001101 (.a(t6_0011010), .b(t6_0011011), .y(t6_001101));
wire t6_0011010, t6_0011011;
mixer mix_t6_0011010 (.a(t6_00110100), .b(t6_00110101), .y(t6_0011010));
wire t6_00110100, t6_00110101;
mixer mix_t6_00110100 (.a(t6_001101000), .b(t6_001101001), .y(t6_00110100));
wire t6_001101000, t6_001101001;
mixer mix_t6_00110101 (.a(t6_001101010), .b(t6_001101011), .y(t6_00110101));
wire t6_001101010, t6_001101011;
mixer mix_t6_0011011 (.a(t6_00110110), .b(t6_00110111), .y(t6_0011011));
wire t6_00110110, t6_00110111;
mixer mix_t6_00110110 (.a(t6_001101100), .b(t6_001101101), .y(t6_00110110));
wire t6_001101100, t6_001101101;
mixer mix_t6_00110111 (.a(t6_001101110), .b(t6_001101111), .y(t6_00110111));
wire t6_001101110, t6_001101111;
mixer mix_t6_00111 (.a(t6_001110), .b(t6_001111), .y(t6_00111));
wire t6_001110, t6_001111;
mixer mix_t6_001110 (.a(t6_0011100), .b(t6_0011101), .y(t6_001110));
wire t6_0011100, t6_0011101;
mixer mix_t6_0011100 (.a(t6_00111000), .b(t6_00111001), .y(t6_0011100));
wire t6_00111000, t6_00111001;
mixer mix_t6_00111000 (.a(t6_001110000), .b(t6_001110001), .y(t6_00111000));
wire t6_001110000, t6_001110001;
mixer mix_t6_00111001 (.a(t6_001110010), .b(t6_001110011), .y(t6_00111001));
wire t6_001110010, t6_001110011;
mixer mix_t6_0011101 (.a(t6_00111010), .b(t6_00111011), .y(t6_0011101));
wire t6_00111010, t6_00111011;
mixer mix_t6_00111010 (.a(t6_001110100), .b(t6_001110101), .y(t6_00111010));
wire t6_001110100, t6_001110101;
mixer mix_t6_00111011 (.a(t6_001110110), .b(t6_001110111), .y(t6_00111011));
wire t6_001110110, t6_001110111;
mixer mix_t6_001111 (.a(t6_0011110), .b(t6_0011111), .y(t6_001111));
wire t6_0011110, t6_0011111;
mixer mix_t6_0011110 (.a(t6_00111100), .b(t6_00111101), .y(t6_0011110));
wire t6_00111100, t6_00111101;
mixer mix_t6_00111100 (.a(t6_001111000), .b(t6_001111001), .y(t6_00111100));
wire t6_001111000, t6_001111001;
mixer mix_t6_00111101 (.a(t6_001111010), .b(t6_001111011), .y(t6_00111101));
wire t6_001111010, t6_001111011;
mixer mix_t6_0011111 (.a(t6_00111110), .b(t6_00111111), .y(t6_0011111));
wire t6_00111110, t6_00111111;
mixer mix_t6_00111110 (.a(t6_001111100), .b(t6_001111101), .y(t6_00111110));
wire t6_001111100, t6_001111101;
mixer mix_t6_00111111 (.a(t6_001111110), .b(t6_001111111), .y(t6_00111111));
wire t6_001111110, t6_001111111;
mixer mix_t6_01 (.a(t6_010), .b(t6_011), .y(t6_01));
wire t6_010, t6_011;
mixer mix_t6_010 (.a(t6_0100), .b(t6_0101), .y(t6_010));
wire t6_0100, t6_0101;
mixer mix_t6_0100 (.a(t6_01000), .b(t6_01001), .y(t6_0100));
wire t6_01000, t6_01001;
mixer mix_t6_01000 (.a(t6_010000), .b(t6_010001), .y(t6_01000));
wire t6_010000, t6_010001;
mixer mix_t6_010000 (.a(t6_0100000), .b(t6_0100001), .y(t6_010000));
wire t6_0100000, t6_0100001;
mixer mix_t6_0100000 (.a(t6_01000000), .b(t6_01000001), .y(t6_0100000));
wire t6_01000000, t6_01000001;
mixer mix_t6_01000000 (.a(t6_010000000), .b(t6_010000001), .y(t6_01000000));
wire t6_010000000, t6_010000001;
mixer mix_t6_01000001 (.a(t6_010000010), .b(t6_010000011), .y(t6_01000001));
wire t6_010000010, t6_010000011;
mixer mix_t6_0100001 (.a(t6_01000010), .b(t6_01000011), .y(t6_0100001));
wire t6_01000010, t6_01000011;
mixer mix_t6_01000010 (.a(t6_010000100), .b(t6_010000101), .y(t6_01000010));
wire t6_010000100, t6_010000101;
mixer mix_t6_01000011 (.a(t6_010000110), .b(t6_010000111), .y(t6_01000011));
wire t6_010000110, t6_010000111;
mixer mix_t6_010001 (.a(t6_0100010), .b(t6_0100011), .y(t6_010001));
wire t6_0100010, t6_0100011;
mixer mix_t6_0100010 (.a(t6_01000100), .b(t6_01000101), .y(t6_0100010));
wire t6_01000100, t6_01000101;
mixer mix_t6_01000100 (.a(t6_010001000), .b(t6_010001001), .y(t6_01000100));
wire t6_010001000, t6_010001001;
mixer mix_t6_01000101 (.a(t6_010001010), .b(t6_010001011), .y(t6_01000101));
wire t6_010001010, t6_010001011;
mixer mix_t6_0100011 (.a(t6_01000110), .b(t6_01000111), .y(t6_0100011));
wire t6_01000110, t6_01000111;
mixer mix_t6_01000110 (.a(t6_010001100), .b(t6_010001101), .y(t6_01000110));
wire t6_010001100, t6_010001101;
mixer mix_t6_01000111 (.a(t6_010001110), .b(t6_010001111), .y(t6_01000111));
wire t6_010001110, t6_010001111;
mixer mix_t6_01001 (.a(t6_010010), .b(t6_010011), .y(t6_01001));
wire t6_010010, t6_010011;
mixer mix_t6_010010 (.a(t6_0100100), .b(t6_0100101), .y(t6_010010));
wire t6_0100100, t6_0100101;
mixer mix_t6_0100100 (.a(t6_01001000), .b(t6_01001001), .y(t6_0100100));
wire t6_01001000, t6_01001001;
mixer mix_t6_01001000 (.a(t6_010010000), .b(t6_010010001), .y(t6_01001000));
wire t6_010010000, t6_010010001;
mixer mix_t6_01001001 (.a(t6_010010010), .b(t6_010010011), .y(t6_01001001));
wire t6_010010010, t6_010010011;
mixer mix_t6_0100101 (.a(t6_01001010), .b(t6_01001011), .y(t6_0100101));
wire t6_01001010, t6_01001011;
mixer mix_t6_01001010 (.a(t6_010010100), .b(t6_010010101), .y(t6_01001010));
wire t6_010010100, t6_010010101;
mixer mix_t6_01001011 (.a(t6_010010110), .b(t6_010010111), .y(t6_01001011));
wire t6_010010110, t6_010010111;
mixer mix_t6_010011 (.a(t6_0100110), .b(t6_0100111), .y(t6_010011));
wire t6_0100110, t6_0100111;
mixer mix_t6_0100110 (.a(t6_01001100), .b(t6_01001101), .y(t6_0100110));
wire t6_01001100, t6_01001101;
mixer mix_t6_01001100 (.a(t6_010011000), .b(t6_010011001), .y(t6_01001100));
wire t6_010011000, t6_010011001;
mixer mix_t6_01001101 (.a(t6_010011010), .b(t6_010011011), .y(t6_01001101));
wire t6_010011010, t6_010011011;
mixer mix_t6_0100111 (.a(t6_01001110), .b(t6_01001111), .y(t6_0100111));
wire t6_01001110, t6_01001111;
mixer mix_t6_01001110 (.a(t6_010011100), .b(t6_010011101), .y(t6_01001110));
wire t6_010011100, t6_010011101;
mixer mix_t6_01001111 (.a(t6_010011110), .b(t6_010011111), .y(t6_01001111));
wire t6_010011110, t6_010011111;
mixer mix_t6_0101 (.a(t6_01010), .b(t6_01011), .y(t6_0101));
wire t6_01010, t6_01011;
mixer mix_t6_01010 (.a(t6_010100), .b(t6_010101), .y(t6_01010));
wire t6_010100, t6_010101;
mixer mix_t6_010100 (.a(t6_0101000), .b(t6_0101001), .y(t6_010100));
wire t6_0101000, t6_0101001;
mixer mix_t6_0101000 (.a(t6_01010000), .b(t6_01010001), .y(t6_0101000));
wire t6_01010000, t6_01010001;
mixer mix_t6_01010000 (.a(t6_010100000), .b(t6_010100001), .y(t6_01010000));
wire t6_010100000, t6_010100001;
mixer mix_t6_01010001 (.a(t6_010100010), .b(t6_010100011), .y(t6_01010001));
wire t6_010100010, t6_010100011;
mixer mix_t6_0101001 (.a(t6_01010010), .b(t6_01010011), .y(t6_0101001));
wire t6_01010010, t6_01010011;
mixer mix_t6_01010010 (.a(t6_010100100), .b(t6_010100101), .y(t6_01010010));
wire t6_010100100, t6_010100101;
mixer mix_t6_01010011 (.a(t6_010100110), .b(t6_010100111), .y(t6_01010011));
wire t6_010100110, t6_010100111;
mixer mix_t6_010101 (.a(t6_0101010), .b(t6_0101011), .y(t6_010101));
wire t6_0101010, t6_0101011;
mixer mix_t6_0101010 (.a(t6_01010100), .b(t6_01010101), .y(t6_0101010));
wire t6_01010100, t6_01010101;
mixer mix_t6_01010100 (.a(t6_010101000), .b(t6_010101001), .y(t6_01010100));
wire t6_010101000, t6_010101001;
mixer mix_t6_01010101 (.a(t6_010101010), .b(t6_010101011), .y(t6_01010101));
wire t6_010101010, t6_010101011;
mixer mix_t6_0101011 (.a(t6_01010110), .b(t6_01010111), .y(t6_0101011));
wire t6_01010110, t6_01010111;
mixer mix_t6_01010110 (.a(t6_010101100), .b(t6_010101101), .y(t6_01010110));
wire t6_010101100, t6_010101101;
mixer mix_t6_01010111 (.a(t6_010101110), .b(t6_010101111), .y(t6_01010111));
wire t6_010101110, t6_010101111;
mixer mix_t6_01011 (.a(t6_010110), .b(t6_010111), .y(t6_01011));
wire t6_010110, t6_010111;
mixer mix_t6_010110 (.a(t6_0101100), .b(t6_0101101), .y(t6_010110));
wire t6_0101100, t6_0101101;
mixer mix_t6_0101100 (.a(t6_01011000), .b(t6_01011001), .y(t6_0101100));
wire t6_01011000, t6_01011001;
mixer mix_t6_01011000 (.a(t6_010110000), .b(t6_010110001), .y(t6_01011000));
wire t6_010110000, t6_010110001;
mixer mix_t6_01011001 (.a(t6_010110010), .b(t6_010110011), .y(t6_01011001));
wire t6_010110010, t6_010110011;
mixer mix_t6_0101101 (.a(t6_01011010), .b(t6_01011011), .y(t6_0101101));
wire t6_01011010, t6_01011011;
mixer mix_t6_01011010 (.a(t6_010110100), .b(t6_010110101), .y(t6_01011010));
wire t6_010110100, t6_010110101;
mixer mix_t6_01011011 (.a(t6_010110110), .b(t6_010110111), .y(t6_01011011));
wire t6_010110110, t6_010110111;
mixer mix_t6_010111 (.a(t6_0101110), .b(t6_0101111), .y(t6_010111));
wire t6_0101110, t6_0101111;
mixer mix_t6_0101110 (.a(t6_01011100), .b(t6_01011101), .y(t6_0101110));
wire t6_01011100, t6_01011101;
mixer mix_t6_01011100 (.a(t6_010111000), .b(t6_010111001), .y(t6_01011100));
wire t6_010111000, t6_010111001;
mixer mix_t6_01011101 (.a(t6_010111010), .b(t6_010111011), .y(t6_01011101));
wire t6_010111010, t6_010111011;
mixer mix_t6_0101111 (.a(t6_01011110), .b(t6_01011111), .y(t6_0101111));
wire t6_01011110, t6_01011111;
mixer mix_t6_01011110 (.a(t6_010111100), .b(t6_010111101), .y(t6_01011110));
wire t6_010111100, t6_010111101;
mixer mix_t6_01011111 (.a(t6_010111110), .b(t6_010111111), .y(t6_01011111));
wire t6_010111110, t6_010111111;
mixer mix_t6_011 (.a(t6_0110), .b(t6_0111), .y(t6_011));
wire t6_0110, t6_0111;
mixer mix_t6_0110 (.a(t6_01100), .b(t6_01101), .y(t6_0110));
wire t6_01100, t6_01101;
mixer mix_t6_01100 (.a(t6_011000), .b(t6_011001), .y(t6_01100));
wire t6_011000, t6_011001;
mixer mix_t6_011000 (.a(t6_0110000), .b(t6_0110001), .y(t6_011000));
wire t6_0110000, t6_0110001;
mixer mix_t6_0110000 (.a(t6_01100000), .b(t6_01100001), .y(t6_0110000));
wire t6_01100000, t6_01100001;
mixer mix_t6_01100000 (.a(t6_011000000), .b(t6_011000001), .y(t6_01100000));
wire t6_011000000, t6_011000001;
mixer mix_t6_01100001 (.a(t6_011000010), .b(t6_011000011), .y(t6_01100001));
wire t6_011000010, t6_011000011;
mixer mix_t6_0110001 (.a(t6_01100010), .b(t6_01100011), .y(t6_0110001));
wire t6_01100010, t6_01100011;
mixer mix_t6_01100010 (.a(t6_011000100), .b(t6_011000101), .y(t6_01100010));
wire t6_011000100, t6_011000101;
mixer mix_t6_01100011 (.a(t6_011000110), .b(t6_011000111), .y(t6_01100011));
wire t6_011000110, t6_011000111;
mixer mix_t6_011001 (.a(t6_0110010), .b(t6_0110011), .y(t6_011001));
wire t6_0110010, t6_0110011;
mixer mix_t6_0110010 (.a(t6_01100100), .b(t6_01100101), .y(t6_0110010));
wire t6_01100100, t6_01100101;
mixer mix_t6_01100100 (.a(t6_011001000), .b(t6_011001001), .y(t6_01100100));
wire t6_011001000, t6_011001001;
mixer mix_t6_01100101 (.a(t6_011001010), .b(t6_011001011), .y(t6_01100101));
wire t6_011001010, t6_011001011;
mixer mix_t6_0110011 (.a(t6_01100110), .b(t6_01100111), .y(t6_0110011));
wire t6_01100110, t6_01100111;
mixer mix_t6_01100110 (.a(t6_011001100), .b(t6_011001101), .y(t6_01100110));
wire t6_011001100, t6_011001101;
mixer mix_t6_01100111 (.a(t6_011001110), .b(t6_011001111), .y(t6_01100111));
wire t6_011001110, t6_011001111;
mixer mix_t6_01101 (.a(t6_011010), .b(t6_011011), .y(t6_01101));
wire t6_011010, t6_011011;
mixer mix_t6_011010 (.a(t6_0110100), .b(t6_0110101), .y(t6_011010));
wire t6_0110100, t6_0110101;
mixer mix_t6_0110100 (.a(t6_01101000), .b(t6_01101001), .y(t6_0110100));
wire t6_01101000, t6_01101001;
mixer mix_t6_01101000 (.a(t6_011010000), .b(t6_011010001), .y(t6_01101000));
wire t6_011010000, t6_011010001;
mixer mix_t6_01101001 (.a(t6_011010010), .b(t6_011010011), .y(t6_01101001));
wire t6_011010010, t6_011010011;
mixer mix_t6_0110101 (.a(t6_01101010), .b(t6_01101011), .y(t6_0110101));
wire t6_01101010, t6_01101011;
mixer mix_t6_01101010 (.a(t6_011010100), .b(t6_011010101), .y(t6_01101010));
wire t6_011010100, t6_011010101;
mixer mix_t6_01101011 (.a(t6_011010110), .b(t6_011010111), .y(t6_01101011));
wire t6_011010110, t6_011010111;
mixer mix_t6_011011 (.a(t6_0110110), .b(t6_0110111), .y(t6_011011));
wire t6_0110110, t6_0110111;
mixer mix_t6_0110110 (.a(t6_01101100), .b(t6_01101101), .y(t6_0110110));
wire t6_01101100, t6_01101101;
mixer mix_t6_01101100 (.a(t6_011011000), .b(t6_011011001), .y(t6_01101100));
wire t6_011011000, t6_011011001;
mixer mix_t6_01101101 (.a(t6_011011010), .b(t6_011011011), .y(t6_01101101));
wire t6_011011010, t6_011011011;
mixer mix_t6_0110111 (.a(t6_01101110), .b(t6_01101111), .y(t6_0110111));
wire t6_01101110, t6_01101111;
mixer mix_t6_01101110 (.a(t6_011011100), .b(t6_011011101), .y(t6_01101110));
wire t6_011011100, t6_011011101;
mixer mix_t6_01101111 (.a(t6_011011110), .b(t6_011011111), .y(t6_01101111));
wire t6_011011110, t6_011011111;
mixer mix_t6_0111 (.a(t6_01110), .b(t6_01111), .y(t6_0111));
wire t6_01110, t6_01111;
mixer mix_t6_01110 (.a(t6_011100), .b(t6_011101), .y(t6_01110));
wire t6_011100, t6_011101;
mixer mix_t6_011100 (.a(t6_0111000), .b(t6_0111001), .y(t6_011100));
wire t6_0111000, t6_0111001;
mixer mix_t6_0111000 (.a(t6_01110000), .b(t6_01110001), .y(t6_0111000));
wire t6_01110000, t6_01110001;
mixer mix_t6_01110000 (.a(t6_011100000), .b(t6_011100001), .y(t6_01110000));
wire t6_011100000, t6_011100001;
mixer mix_t6_01110001 (.a(t6_011100010), .b(t6_011100011), .y(t6_01110001));
wire t6_011100010, t6_011100011;
mixer mix_t6_0111001 (.a(t6_01110010), .b(t6_01110011), .y(t6_0111001));
wire t6_01110010, t6_01110011;
mixer mix_t6_01110010 (.a(t6_011100100), .b(t6_011100101), .y(t6_01110010));
wire t6_011100100, t6_011100101;
mixer mix_t6_01110011 (.a(t6_011100110), .b(t6_011100111), .y(t6_01110011));
wire t6_011100110, t6_011100111;
mixer mix_t6_011101 (.a(t6_0111010), .b(t6_0111011), .y(t6_011101));
wire t6_0111010, t6_0111011;
mixer mix_t6_0111010 (.a(t6_01110100), .b(t6_01110101), .y(t6_0111010));
wire t6_01110100, t6_01110101;
mixer mix_t6_01110100 (.a(t6_011101000), .b(t6_011101001), .y(t6_01110100));
wire t6_011101000, t6_011101001;
mixer mix_t6_01110101 (.a(t6_011101010), .b(t6_011101011), .y(t6_01110101));
wire t6_011101010, t6_011101011;
mixer mix_t6_0111011 (.a(t6_01110110), .b(t6_01110111), .y(t6_0111011));
wire t6_01110110, t6_01110111;
mixer mix_t6_01110110 (.a(t6_011101100), .b(t6_011101101), .y(t6_01110110));
wire t6_011101100, t6_011101101;
mixer mix_t6_01110111 (.a(t6_011101110), .b(t6_011101111), .y(t6_01110111));
wire t6_011101110, t6_011101111;
mixer mix_t6_01111 (.a(t6_011110), .b(t6_011111), .y(t6_01111));
wire t6_011110, t6_011111;
mixer mix_t6_011110 (.a(t6_0111100), .b(t6_0111101), .y(t6_011110));
wire t6_0111100, t6_0111101;
mixer mix_t6_0111100 (.a(t6_01111000), .b(t6_01111001), .y(t6_0111100));
wire t6_01111000, t6_01111001;
mixer mix_t6_01111000 (.a(t6_011110000), .b(t6_011110001), .y(t6_01111000));
wire t6_011110000, t6_011110001;
mixer mix_t6_01111001 (.a(t6_011110010), .b(t6_011110011), .y(t6_01111001));
wire t6_011110010, t6_011110011;
mixer mix_t6_0111101 (.a(t6_01111010), .b(t6_01111011), .y(t6_0111101));
wire t6_01111010, t6_01111011;
mixer mix_t6_01111010 (.a(t6_011110100), .b(t6_011110101), .y(t6_01111010));
wire t6_011110100, t6_011110101;
mixer mix_t6_01111011 (.a(t6_011110110), .b(t6_011110111), .y(t6_01111011));
wire t6_011110110, t6_011110111;
mixer mix_t6_011111 (.a(t6_0111110), .b(t6_0111111), .y(t6_011111));
wire t6_0111110, t6_0111111;
mixer mix_t6_0111110 (.a(t6_01111100), .b(t6_01111101), .y(t6_0111110));
wire t6_01111100, t6_01111101;
mixer mix_t6_01111100 (.a(t6_011111000), .b(t6_011111001), .y(t6_01111100));
wire t6_011111000, t6_011111001;
mixer mix_t6_01111101 (.a(t6_011111010), .b(t6_011111011), .y(t6_01111101));
wire t6_011111010, t6_011111011;
mixer mix_t6_0111111 (.a(t6_01111110), .b(t6_01111111), .y(t6_0111111));
wire t6_01111110, t6_01111111;
mixer mix_t6_01111110 (.a(t6_011111100), .b(t6_011111101), .y(t6_01111110));
wire t6_011111100, t6_011111101;
mixer mix_t6_01111111 (.a(t6_011111110), .b(t6_011111111), .y(t6_01111111));
wire t6_011111110, t6_011111111;
mixer mix_t7_0 (.a(t7_00), .b(t7_01), .y(t7_0));
wire t7_00, t7_01;
mixer mix_t7_00 (.a(t7_000), .b(t7_001), .y(t7_00));
wire t7_000, t7_001;
mixer mix_t7_000 (.a(t7_0000), .b(t7_0001), .y(t7_000));
wire t7_0000, t7_0001;
mixer mix_t7_0000 (.a(t7_00000), .b(t7_00001), .y(t7_0000));
wire t7_00000, t7_00001;
mixer mix_t7_00000 (.a(t7_000000), .b(t7_000001), .y(t7_00000));
wire t7_000000, t7_000001;
mixer mix_t7_000000 (.a(t7_0000000), .b(t7_0000001), .y(t7_000000));
wire t7_0000000, t7_0000001;
mixer mix_t7_0000000 (.a(t7_00000000), .b(t7_00000001), .y(t7_0000000));
wire t7_00000000, t7_00000001;
mixer mix_t7_00000000 (.a(t7_000000000), .b(t7_000000001), .y(t7_00000000));
wire t7_000000000, t7_000000001;
mixer mix_t7_00000001 (.a(t7_000000010), .b(t7_000000011), .y(t7_00000001));
wire t7_000000010, t7_000000011;
mixer mix_t7_0000001 (.a(t7_00000010), .b(t7_00000011), .y(t7_0000001));
wire t7_00000010, t7_00000011;
mixer mix_t7_00000010 (.a(t7_000000100), .b(t7_000000101), .y(t7_00000010));
wire t7_000000100, t7_000000101;
mixer mix_t7_00000011 (.a(t7_000000110), .b(t7_000000111), .y(t7_00000011));
wire t7_000000110, t7_000000111;
mixer mix_t7_000001 (.a(t7_0000010), .b(t7_0000011), .y(t7_000001));
wire t7_0000010, t7_0000011;
mixer mix_t7_0000010 (.a(t7_00000100), .b(t7_00000101), .y(t7_0000010));
wire t7_00000100, t7_00000101;
mixer mix_t7_00000100 (.a(t7_000001000), .b(t7_000001001), .y(t7_00000100));
wire t7_000001000, t7_000001001;
mixer mix_t7_00000101 (.a(t7_000001010), .b(t7_000001011), .y(t7_00000101));
wire t7_000001010, t7_000001011;
mixer mix_t7_0000011 (.a(t7_00000110), .b(t7_00000111), .y(t7_0000011));
wire t7_00000110, t7_00000111;
mixer mix_t7_00000110 (.a(t7_000001100), .b(t7_000001101), .y(t7_00000110));
wire t7_000001100, t7_000001101;
mixer mix_t7_00000111 (.a(t7_000001110), .b(t7_000001111), .y(t7_00000111));
wire t7_000001110, t7_000001111;
mixer mix_t7_00001 (.a(t7_000010), .b(t7_000011), .y(t7_00001));
wire t7_000010, t7_000011;
mixer mix_t7_000010 (.a(t7_0000100), .b(t7_0000101), .y(t7_000010));
wire t7_0000100, t7_0000101;
mixer mix_t7_0000100 (.a(t7_00001000), .b(t7_00001001), .y(t7_0000100));
wire t7_00001000, t7_00001001;
mixer mix_t7_00001000 (.a(t7_000010000), .b(t7_000010001), .y(t7_00001000));
wire t7_000010000, t7_000010001;
mixer mix_t7_00001001 (.a(t7_000010010), .b(t7_000010011), .y(t7_00001001));
wire t7_000010010, t7_000010011;
mixer mix_t7_0000101 (.a(t7_00001010), .b(t7_00001011), .y(t7_0000101));
wire t7_00001010, t7_00001011;
mixer mix_t7_00001010 (.a(t7_000010100), .b(t7_000010101), .y(t7_00001010));
wire t7_000010100, t7_000010101;
mixer mix_t7_00001011 (.a(t7_000010110), .b(t7_000010111), .y(t7_00001011));
wire t7_000010110, t7_000010111;
mixer mix_t7_000011 (.a(t7_0000110), .b(t7_0000111), .y(t7_000011));
wire t7_0000110, t7_0000111;
mixer mix_t7_0000110 (.a(t7_00001100), .b(t7_00001101), .y(t7_0000110));
wire t7_00001100, t7_00001101;
mixer mix_t7_00001100 (.a(t7_000011000), .b(t7_000011001), .y(t7_00001100));
wire t7_000011000, t7_000011001;
mixer mix_t7_00001101 (.a(t7_000011010), .b(t7_000011011), .y(t7_00001101));
wire t7_000011010, t7_000011011;
mixer mix_t7_0000111 (.a(t7_00001110), .b(t7_00001111), .y(t7_0000111));
wire t7_00001110, t7_00001111;
mixer mix_t7_00001110 (.a(t7_000011100), .b(t7_000011101), .y(t7_00001110));
wire t7_000011100, t7_000011101;
mixer mix_t7_00001111 (.a(t7_000011110), .b(t7_000011111), .y(t7_00001111));
wire t7_000011110, t7_000011111;
mixer mix_t7_0001 (.a(t7_00010), .b(t7_00011), .y(t7_0001));
wire t7_00010, t7_00011;
mixer mix_t7_00010 (.a(t7_000100), .b(t7_000101), .y(t7_00010));
wire t7_000100, t7_000101;
mixer mix_t7_000100 (.a(t7_0001000), .b(t7_0001001), .y(t7_000100));
wire t7_0001000, t7_0001001;
mixer mix_t7_0001000 (.a(t7_00010000), .b(t7_00010001), .y(t7_0001000));
wire t7_00010000, t7_00010001;
mixer mix_t7_00010000 (.a(t7_000100000), .b(t7_000100001), .y(t7_00010000));
wire t7_000100000, t7_000100001;
mixer mix_t7_00010001 (.a(t7_000100010), .b(t7_000100011), .y(t7_00010001));
wire t7_000100010, t7_000100011;
mixer mix_t7_0001001 (.a(t7_00010010), .b(t7_00010011), .y(t7_0001001));
wire t7_00010010, t7_00010011;
mixer mix_t7_00010010 (.a(t7_000100100), .b(t7_000100101), .y(t7_00010010));
wire t7_000100100, t7_000100101;
mixer mix_t7_00010011 (.a(t7_000100110), .b(t7_000100111), .y(t7_00010011));
wire t7_000100110, t7_000100111;
mixer mix_t7_000101 (.a(t7_0001010), .b(t7_0001011), .y(t7_000101));
wire t7_0001010, t7_0001011;
mixer mix_t7_0001010 (.a(t7_00010100), .b(t7_00010101), .y(t7_0001010));
wire t7_00010100, t7_00010101;
mixer mix_t7_00010100 (.a(t7_000101000), .b(t7_000101001), .y(t7_00010100));
wire t7_000101000, t7_000101001;
mixer mix_t7_00010101 (.a(t7_000101010), .b(t7_000101011), .y(t7_00010101));
wire t7_000101010, t7_000101011;
mixer mix_t7_0001011 (.a(t7_00010110), .b(t7_00010111), .y(t7_0001011));
wire t7_00010110, t7_00010111;
mixer mix_t7_00010110 (.a(t7_000101100), .b(t7_000101101), .y(t7_00010110));
wire t7_000101100, t7_000101101;
mixer mix_t7_00010111 (.a(t7_000101110), .b(t7_000101111), .y(t7_00010111));
wire t7_000101110, t7_000101111;
mixer mix_t7_00011 (.a(t7_000110), .b(t7_000111), .y(t7_00011));
wire t7_000110, t7_000111;
mixer mix_t7_000110 (.a(t7_0001100), .b(t7_0001101), .y(t7_000110));
wire t7_0001100, t7_0001101;
mixer mix_t7_0001100 (.a(t7_00011000), .b(t7_00011001), .y(t7_0001100));
wire t7_00011000, t7_00011001;
mixer mix_t7_00011000 (.a(t7_000110000), .b(t7_000110001), .y(t7_00011000));
wire t7_000110000, t7_000110001;
mixer mix_t7_00011001 (.a(t7_000110010), .b(t7_000110011), .y(t7_00011001));
wire t7_000110010, t7_000110011;
mixer mix_t7_0001101 (.a(t7_00011010), .b(t7_00011011), .y(t7_0001101));
wire t7_00011010, t7_00011011;
mixer mix_t7_00011010 (.a(t7_000110100), .b(t7_000110101), .y(t7_00011010));
wire t7_000110100, t7_000110101;
mixer mix_t7_00011011 (.a(t7_000110110), .b(t7_000110111), .y(t7_00011011));
wire t7_000110110, t7_000110111;
mixer mix_t7_000111 (.a(t7_0001110), .b(t7_0001111), .y(t7_000111));
wire t7_0001110, t7_0001111;
mixer mix_t7_0001110 (.a(t7_00011100), .b(t7_00011101), .y(t7_0001110));
wire t7_00011100, t7_00011101;
mixer mix_t7_00011100 (.a(t7_000111000), .b(t7_000111001), .y(t7_00011100));
wire t7_000111000, t7_000111001;
mixer mix_t7_00011101 (.a(t7_000111010), .b(t7_000111011), .y(t7_00011101));
wire t7_000111010, t7_000111011;
mixer mix_t7_0001111 (.a(t7_00011110), .b(t7_00011111), .y(t7_0001111));
wire t7_00011110, t7_00011111;
mixer mix_t7_00011110 (.a(t7_000111100), .b(t7_000111101), .y(t7_00011110));
wire t7_000111100, t7_000111101;
mixer mix_t7_00011111 (.a(t7_000111110), .b(t7_000111111), .y(t7_00011111));
wire t7_000111110, t7_000111111;
mixer mix_t7_001 (.a(t7_0010), .b(t7_0011), .y(t7_001));
wire t7_0010, t7_0011;
mixer mix_t7_0010 (.a(t7_00100), .b(t7_00101), .y(t7_0010));
wire t7_00100, t7_00101;
mixer mix_t7_00100 (.a(t7_001000), .b(t7_001001), .y(t7_00100));
wire t7_001000, t7_001001;
mixer mix_t7_001000 (.a(t7_0010000), .b(t7_0010001), .y(t7_001000));
wire t7_0010000, t7_0010001;
mixer mix_t7_0010000 (.a(t7_00100000), .b(t7_00100001), .y(t7_0010000));
wire t7_00100000, t7_00100001;
mixer mix_t7_00100000 (.a(t7_001000000), .b(t7_001000001), .y(t7_00100000));
wire t7_001000000, t7_001000001;
mixer mix_t7_00100001 (.a(t7_001000010), .b(t7_001000011), .y(t7_00100001));
wire t7_001000010, t7_001000011;
mixer mix_t7_0010001 (.a(t7_00100010), .b(t7_00100011), .y(t7_0010001));
wire t7_00100010, t7_00100011;
mixer mix_t7_00100010 (.a(t7_001000100), .b(t7_001000101), .y(t7_00100010));
wire t7_001000100, t7_001000101;
mixer mix_t7_00100011 (.a(t7_001000110), .b(t7_001000111), .y(t7_00100011));
wire t7_001000110, t7_001000111;
mixer mix_t7_001001 (.a(t7_0010010), .b(t7_0010011), .y(t7_001001));
wire t7_0010010, t7_0010011;
mixer mix_t7_0010010 (.a(t7_00100100), .b(t7_00100101), .y(t7_0010010));
wire t7_00100100, t7_00100101;
mixer mix_t7_00100100 (.a(t7_001001000), .b(t7_001001001), .y(t7_00100100));
wire t7_001001000, t7_001001001;
mixer mix_t7_00100101 (.a(t7_001001010), .b(t7_001001011), .y(t7_00100101));
wire t7_001001010, t7_001001011;
mixer mix_t7_0010011 (.a(t7_00100110), .b(t7_00100111), .y(t7_0010011));
wire t7_00100110, t7_00100111;
mixer mix_t7_00100110 (.a(t7_001001100), .b(t7_001001101), .y(t7_00100110));
wire t7_001001100, t7_001001101;
mixer mix_t7_00100111 (.a(t7_001001110), .b(t7_001001111), .y(t7_00100111));
wire t7_001001110, t7_001001111;
mixer mix_t7_00101 (.a(t7_001010), .b(t7_001011), .y(t7_00101));
wire t7_001010, t7_001011;
mixer mix_t7_001010 (.a(t7_0010100), .b(t7_0010101), .y(t7_001010));
wire t7_0010100, t7_0010101;
mixer mix_t7_0010100 (.a(t7_00101000), .b(t7_00101001), .y(t7_0010100));
wire t7_00101000, t7_00101001;
mixer mix_t7_00101000 (.a(t7_001010000), .b(t7_001010001), .y(t7_00101000));
wire t7_001010000, t7_001010001;
mixer mix_t7_00101001 (.a(t7_001010010), .b(t7_001010011), .y(t7_00101001));
wire t7_001010010, t7_001010011;
mixer mix_t7_0010101 (.a(t7_00101010), .b(t7_00101011), .y(t7_0010101));
wire t7_00101010, t7_00101011;
mixer mix_t7_00101010 (.a(t7_001010100), .b(t7_001010101), .y(t7_00101010));
wire t7_001010100, t7_001010101;
mixer mix_t7_00101011 (.a(t7_001010110), .b(t7_001010111), .y(t7_00101011));
wire t7_001010110, t7_001010111;
mixer mix_t7_001011 (.a(t7_0010110), .b(t7_0010111), .y(t7_001011));
wire t7_0010110, t7_0010111;
mixer mix_t7_0010110 (.a(t7_00101100), .b(t7_00101101), .y(t7_0010110));
wire t7_00101100, t7_00101101;
mixer mix_t7_00101100 (.a(t7_001011000), .b(t7_001011001), .y(t7_00101100));
wire t7_001011000, t7_001011001;
mixer mix_t7_00101101 (.a(t7_001011010), .b(t7_001011011), .y(t7_00101101));
wire t7_001011010, t7_001011011;
mixer mix_t7_0010111 (.a(t7_00101110), .b(t7_00101111), .y(t7_0010111));
wire t7_00101110, t7_00101111;
mixer mix_t7_00101110 (.a(t7_001011100), .b(t7_001011101), .y(t7_00101110));
wire t7_001011100, t7_001011101;
mixer mix_t7_00101111 (.a(t7_001011110), .b(t7_001011111), .y(t7_00101111));
wire t7_001011110, t7_001011111;
mixer mix_t7_0011 (.a(t7_00110), .b(t7_00111), .y(t7_0011));
wire t7_00110, t7_00111;
mixer mix_t7_00110 (.a(t7_001100), .b(t7_001101), .y(t7_00110));
wire t7_001100, t7_001101;
mixer mix_t7_001100 (.a(t7_0011000), .b(t7_0011001), .y(t7_001100));
wire t7_0011000, t7_0011001;
mixer mix_t7_0011000 (.a(t7_00110000), .b(t7_00110001), .y(t7_0011000));
wire t7_00110000, t7_00110001;
mixer mix_t7_00110000 (.a(t7_001100000), .b(t7_001100001), .y(t7_00110000));
wire t7_001100000, t7_001100001;
mixer mix_t7_00110001 (.a(t7_001100010), .b(t7_001100011), .y(t7_00110001));
wire t7_001100010, t7_001100011;
mixer mix_t7_0011001 (.a(t7_00110010), .b(t7_00110011), .y(t7_0011001));
wire t7_00110010, t7_00110011;
mixer mix_t7_00110010 (.a(t7_001100100), .b(t7_001100101), .y(t7_00110010));
wire t7_001100100, t7_001100101;
mixer mix_t7_00110011 (.a(t7_001100110), .b(t7_001100111), .y(t7_00110011));
wire t7_001100110, t7_001100111;
mixer mix_t7_001101 (.a(t7_0011010), .b(t7_0011011), .y(t7_001101));
wire t7_0011010, t7_0011011;
mixer mix_t7_0011010 (.a(t7_00110100), .b(t7_00110101), .y(t7_0011010));
wire t7_00110100, t7_00110101;
mixer mix_t7_00110100 (.a(t7_001101000), .b(t7_001101001), .y(t7_00110100));
wire t7_001101000, t7_001101001;
mixer mix_t7_00110101 (.a(t7_001101010), .b(t7_001101011), .y(t7_00110101));
wire t7_001101010, t7_001101011;
mixer mix_t7_0011011 (.a(t7_00110110), .b(t7_00110111), .y(t7_0011011));
wire t7_00110110, t7_00110111;
mixer mix_t7_00110110 (.a(t7_001101100), .b(t7_001101101), .y(t7_00110110));
wire t7_001101100, t7_001101101;
mixer mix_t7_00110111 (.a(t7_001101110), .b(t7_001101111), .y(t7_00110111));
wire t7_001101110, t7_001101111;
mixer mix_t7_00111 (.a(t7_001110), .b(t7_001111), .y(t7_00111));
wire t7_001110, t7_001111;
mixer mix_t7_001110 (.a(t7_0011100), .b(t7_0011101), .y(t7_001110));
wire t7_0011100, t7_0011101;
mixer mix_t7_0011100 (.a(t7_00111000), .b(t7_00111001), .y(t7_0011100));
wire t7_00111000, t7_00111001;
mixer mix_t7_00111000 (.a(t7_001110000), .b(t7_001110001), .y(t7_00111000));
wire t7_001110000, t7_001110001;
mixer mix_t7_00111001 (.a(t7_001110010), .b(t7_001110011), .y(t7_00111001));
wire t7_001110010, t7_001110011;
mixer mix_t7_0011101 (.a(t7_00111010), .b(t7_00111011), .y(t7_0011101));
wire t7_00111010, t7_00111011;
mixer mix_t7_00111010 (.a(t7_001110100), .b(t7_001110101), .y(t7_00111010));
wire t7_001110100, t7_001110101;
mixer mix_t7_00111011 (.a(t7_001110110), .b(t7_001110111), .y(t7_00111011));
wire t7_001110110, t7_001110111;
mixer mix_t7_001111 (.a(t7_0011110), .b(t7_0011111), .y(t7_001111));
wire t7_0011110, t7_0011111;
mixer mix_t7_0011110 (.a(t7_00111100), .b(t7_00111101), .y(t7_0011110));
wire t7_00111100, t7_00111101;
mixer mix_t7_00111100 (.a(t7_001111000), .b(t7_001111001), .y(t7_00111100));
wire t7_001111000, t7_001111001;
mixer mix_t7_00111101 (.a(t7_001111010), .b(t7_001111011), .y(t7_00111101));
wire t7_001111010, t7_001111011;
mixer mix_t7_0011111 (.a(t7_00111110), .b(t7_00111111), .y(t7_0011111));
wire t7_00111110, t7_00111111;
mixer mix_t7_00111110 (.a(t7_001111100), .b(t7_001111101), .y(t7_00111110));
wire t7_001111100, t7_001111101;
mixer mix_t7_00111111 (.a(t7_001111110), .b(t7_001111111), .y(t7_00111111));
wire t7_001111110, t7_001111111;
mixer mix_t7_01 (.a(t7_010), .b(t7_011), .y(t7_01));
wire t7_010, t7_011;
mixer mix_t7_010 (.a(t7_0100), .b(t7_0101), .y(t7_010));
wire t7_0100, t7_0101;
mixer mix_t7_0100 (.a(t7_01000), .b(t7_01001), .y(t7_0100));
wire t7_01000, t7_01001;
mixer mix_t7_01000 (.a(t7_010000), .b(t7_010001), .y(t7_01000));
wire t7_010000, t7_010001;
mixer mix_t7_010000 (.a(t7_0100000), .b(t7_0100001), .y(t7_010000));
wire t7_0100000, t7_0100001;
mixer mix_t7_0100000 (.a(t7_01000000), .b(t7_01000001), .y(t7_0100000));
wire t7_01000000, t7_01000001;
mixer mix_t7_01000000 (.a(t7_010000000), .b(t7_010000001), .y(t7_01000000));
wire t7_010000000, t7_010000001;
mixer mix_t7_01000001 (.a(t7_010000010), .b(t7_010000011), .y(t7_01000001));
wire t7_010000010, t7_010000011;
mixer mix_t7_0100001 (.a(t7_01000010), .b(t7_01000011), .y(t7_0100001));
wire t7_01000010, t7_01000011;
mixer mix_t7_01000010 (.a(t7_010000100), .b(t7_010000101), .y(t7_01000010));
wire t7_010000100, t7_010000101;
mixer mix_t7_01000011 (.a(t7_010000110), .b(t7_010000111), .y(t7_01000011));
wire t7_010000110, t7_010000111;
mixer mix_t7_010001 (.a(t7_0100010), .b(t7_0100011), .y(t7_010001));
wire t7_0100010, t7_0100011;
mixer mix_t7_0100010 (.a(t7_01000100), .b(t7_01000101), .y(t7_0100010));
wire t7_01000100, t7_01000101;
mixer mix_t7_01000100 (.a(t7_010001000), .b(t7_010001001), .y(t7_01000100));
wire t7_010001000, t7_010001001;
mixer mix_t7_01000101 (.a(t7_010001010), .b(t7_010001011), .y(t7_01000101));
wire t7_010001010, t7_010001011;
mixer mix_t7_0100011 (.a(t7_01000110), .b(t7_01000111), .y(t7_0100011));
wire t7_01000110, t7_01000111;
mixer mix_t7_01000110 (.a(t7_010001100), .b(t7_010001101), .y(t7_01000110));
wire t7_010001100, t7_010001101;
mixer mix_t7_01000111 (.a(t7_010001110), .b(t7_010001111), .y(t7_01000111));
wire t7_010001110, t7_010001111;
mixer mix_t7_01001 (.a(t7_010010), .b(t7_010011), .y(t7_01001));
wire t7_010010, t7_010011;
mixer mix_t7_010010 (.a(t7_0100100), .b(t7_0100101), .y(t7_010010));
wire t7_0100100, t7_0100101;
mixer mix_t7_0100100 (.a(t7_01001000), .b(t7_01001001), .y(t7_0100100));
wire t7_01001000, t7_01001001;
mixer mix_t7_01001000 (.a(t7_010010000), .b(t7_010010001), .y(t7_01001000));
wire t7_010010000, t7_010010001;
mixer mix_t7_01001001 (.a(t7_010010010), .b(t7_010010011), .y(t7_01001001));
wire t7_010010010, t7_010010011;
mixer mix_t7_0100101 (.a(t7_01001010), .b(t7_01001011), .y(t7_0100101));
wire t7_01001010, t7_01001011;
mixer mix_t7_01001010 (.a(t7_010010100), .b(t7_010010101), .y(t7_01001010));
wire t7_010010100, t7_010010101;
mixer mix_t7_01001011 (.a(t7_010010110), .b(t7_010010111), .y(t7_01001011));
wire t7_010010110, t7_010010111;
mixer mix_t7_010011 (.a(t7_0100110), .b(t7_0100111), .y(t7_010011));
wire t7_0100110, t7_0100111;
mixer mix_t7_0100110 (.a(t7_01001100), .b(t7_01001101), .y(t7_0100110));
wire t7_01001100, t7_01001101;
mixer mix_t7_01001100 (.a(t7_010011000), .b(t7_010011001), .y(t7_01001100));
wire t7_010011000, t7_010011001;
mixer mix_t7_01001101 (.a(t7_010011010), .b(t7_010011011), .y(t7_01001101));
wire t7_010011010, t7_010011011;
mixer mix_t7_0100111 (.a(t7_01001110), .b(t7_01001111), .y(t7_0100111));
wire t7_01001110, t7_01001111;
mixer mix_t7_01001110 (.a(t7_010011100), .b(t7_010011101), .y(t7_01001110));
wire t7_010011100, t7_010011101;
mixer mix_t7_01001111 (.a(t7_010011110), .b(t7_010011111), .y(t7_01001111));
wire t7_010011110, t7_010011111;
mixer mix_t7_0101 (.a(t7_01010), .b(t7_01011), .y(t7_0101));
wire t7_01010, t7_01011;
mixer mix_t7_01010 (.a(t7_010100), .b(t7_010101), .y(t7_01010));
wire t7_010100, t7_010101;
mixer mix_t7_010100 (.a(t7_0101000), .b(t7_0101001), .y(t7_010100));
wire t7_0101000, t7_0101001;
mixer mix_t7_0101000 (.a(t7_01010000), .b(t7_01010001), .y(t7_0101000));
wire t7_01010000, t7_01010001;
mixer mix_t7_01010000 (.a(t7_010100000), .b(t7_010100001), .y(t7_01010000));
wire t7_010100000, t7_010100001;
mixer mix_t7_01010001 (.a(t7_010100010), .b(t7_010100011), .y(t7_01010001));
wire t7_010100010, t7_010100011;
mixer mix_t7_0101001 (.a(t7_01010010), .b(t7_01010011), .y(t7_0101001));
wire t7_01010010, t7_01010011;
mixer mix_t7_01010010 (.a(t7_010100100), .b(t7_010100101), .y(t7_01010010));
wire t7_010100100, t7_010100101;
mixer mix_t7_01010011 (.a(t7_010100110), .b(t7_010100111), .y(t7_01010011));
wire t7_010100110, t7_010100111;
mixer mix_t7_010101 (.a(t7_0101010), .b(t7_0101011), .y(t7_010101));
wire t7_0101010, t7_0101011;
mixer mix_t7_0101010 (.a(t7_01010100), .b(t7_01010101), .y(t7_0101010));
wire t7_01010100, t7_01010101;
mixer mix_t7_01010100 (.a(t7_010101000), .b(t7_010101001), .y(t7_01010100));
wire t7_010101000, t7_010101001;
mixer mix_t7_01010101 (.a(t7_010101010), .b(t7_010101011), .y(t7_01010101));
wire t7_010101010, t7_010101011;
mixer mix_t7_0101011 (.a(t7_01010110), .b(t7_01010111), .y(t7_0101011));
wire t7_01010110, t7_01010111;
mixer mix_t7_01010110 (.a(t7_010101100), .b(t7_010101101), .y(t7_01010110));
wire t7_010101100, t7_010101101;
mixer mix_t7_01010111 (.a(t7_010101110), .b(t7_010101111), .y(t7_01010111));
wire t7_010101110, t7_010101111;
mixer mix_t7_01011 (.a(t7_010110), .b(t7_010111), .y(t7_01011));
wire t7_010110, t7_010111;
mixer mix_t7_010110 (.a(t7_0101100), .b(t7_0101101), .y(t7_010110));
wire t7_0101100, t7_0101101;
mixer mix_t7_0101100 (.a(t7_01011000), .b(t7_01011001), .y(t7_0101100));
wire t7_01011000, t7_01011001;
mixer mix_t7_01011000 (.a(t7_010110000), .b(t7_010110001), .y(t7_01011000));
wire t7_010110000, t7_010110001;
mixer mix_t7_01011001 (.a(t7_010110010), .b(t7_010110011), .y(t7_01011001));
wire t7_010110010, t7_010110011;
mixer mix_t7_0101101 (.a(t7_01011010), .b(t7_01011011), .y(t7_0101101));
wire t7_01011010, t7_01011011;
mixer mix_t7_01011010 (.a(t7_010110100), .b(t7_010110101), .y(t7_01011010));
wire t7_010110100, t7_010110101;
mixer mix_t7_01011011 (.a(t7_010110110), .b(t7_010110111), .y(t7_01011011));
wire t7_010110110, t7_010110111;
mixer mix_t7_010111 (.a(t7_0101110), .b(t7_0101111), .y(t7_010111));
wire t7_0101110, t7_0101111;
mixer mix_t7_0101110 (.a(t7_01011100), .b(t7_01011101), .y(t7_0101110));
wire t7_01011100, t7_01011101;
mixer mix_t7_01011100 (.a(t7_010111000), .b(t7_010111001), .y(t7_01011100));
wire t7_010111000, t7_010111001;
mixer mix_t7_01011101 (.a(t7_010111010), .b(t7_010111011), .y(t7_01011101));
wire t7_010111010, t7_010111011;
mixer mix_t7_0101111 (.a(t7_01011110), .b(t7_01011111), .y(t7_0101111));
wire t7_01011110, t7_01011111;
mixer mix_t7_01011110 (.a(t7_010111100), .b(t7_010111101), .y(t7_01011110));
wire t7_010111100, t7_010111101;
mixer mix_t7_01011111 (.a(t7_010111110), .b(t7_010111111), .y(t7_01011111));
wire t7_010111110, t7_010111111;
mixer mix_t7_011 (.a(t7_0110), .b(t7_0111), .y(t7_011));
wire t7_0110, t7_0111;
mixer mix_t7_0110 (.a(t7_01100), .b(t7_01101), .y(t7_0110));
wire t7_01100, t7_01101;
mixer mix_t7_01100 (.a(t7_011000), .b(t7_011001), .y(t7_01100));
wire t7_011000, t7_011001;
mixer mix_t7_011000 (.a(t7_0110000), .b(t7_0110001), .y(t7_011000));
wire t7_0110000, t7_0110001;
mixer mix_t7_0110000 (.a(t7_01100000), .b(t7_01100001), .y(t7_0110000));
wire t7_01100000, t7_01100001;
mixer mix_t7_01100000 (.a(t7_011000000), .b(t7_011000001), .y(t7_01100000));
wire t7_011000000, t7_011000001;
mixer mix_t7_01100001 (.a(t7_011000010), .b(t7_011000011), .y(t7_01100001));
wire t7_011000010, t7_011000011;
mixer mix_t7_0110001 (.a(t7_01100010), .b(t7_01100011), .y(t7_0110001));
wire t7_01100010, t7_01100011;
mixer mix_t7_01100010 (.a(t7_011000100), .b(t7_011000101), .y(t7_01100010));
wire t7_011000100, t7_011000101;
mixer mix_t7_01100011 (.a(t7_011000110), .b(t7_011000111), .y(t7_01100011));
wire t7_011000110, t7_011000111;
mixer mix_t7_011001 (.a(t7_0110010), .b(t7_0110011), .y(t7_011001));
wire t7_0110010, t7_0110011;
mixer mix_t7_0110010 (.a(t7_01100100), .b(t7_01100101), .y(t7_0110010));
wire t7_01100100, t7_01100101;
mixer mix_t7_01100100 (.a(t7_011001000), .b(t7_011001001), .y(t7_01100100));
wire t7_011001000, t7_011001001;
mixer mix_t7_01100101 (.a(t7_011001010), .b(t7_011001011), .y(t7_01100101));
wire t7_011001010, t7_011001011;
mixer mix_t7_0110011 (.a(t7_01100110), .b(t7_01100111), .y(t7_0110011));
wire t7_01100110, t7_01100111;
mixer mix_t7_01100110 (.a(t7_011001100), .b(t7_011001101), .y(t7_01100110));
wire t7_011001100, t7_011001101;
mixer mix_t7_01100111 (.a(t7_011001110), .b(t7_011001111), .y(t7_01100111));
wire t7_011001110, t7_011001111;
mixer mix_t7_01101 (.a(t7_011010), .b(t7_011011), .y(t7_01101));
wire t7_011010, t7_011011;
mixer mix_t7_011010 (.a(t7_0110100), .b(t7_0110101), .y(t7_011010));
wire t7_0110100, t7_0110101;
mixer mix_t7_0110100 (.a(t7_01101000), .b(t7_01101001), .y(t7_0110100));
wire t7_01101000, t7_01101001;
mixer mix_t7_01101000 (.a(t7_011010000), .b(t7_011010001), .y(t7_01101000));
wire t7_011010000, t7_011010001;
mixer mix_t7_01101001 (.a(t7_011010010), .b(t7_011010011), .y(t7_01101001));
wire t7_011010010, t7_011010011;
mixer mix_t7_0110101 (.a(t7_01101010), .b(t7_01101011), .y(t7_0110101));
wire t7_01101010, t7_01101011;
mixer mix_t7_01101010 (.a(t7_011010100), .b(t7_011010101), .y(t7_01101010));
wire t7_011010100, t7_011010101;
mixer mix_t7_01101011 (.a(t7_011010110), .b(t7_011010111), .y(t7_01101011));
wire t7_011010110, t7_011010111;
mixer mix_t7_011011 (.a(t7_0110110), .b(t7_0110111), .y(t7_011011));
wire t7_0110110, t7_0110111;
mixer mix_t7_0110110 (.a(t7_01101100), .b(t7_01101101), .y(t7_0110110));
wire t7_01101100, t7_01101101;
mixer mix_t7_01101100 (.a(t7_011011000), .b(t7_011011001), .y(t7_01101100));
wire t7_011011000, t7_011011001;
mixer mix_t7_01101101 (.a(t7_011011010), .b(t7_011011011), .y(t7_01101101));
wire t7_011011010, t7_011011011;
mixer mix_t7_0110111 (.a(t7_01101110), .b(t7_01101111), .y(t7_0110111));
wire t7_01101110, t7_01101111;
mixer mix_t7_01101110 (.a(t7_011011100), .b(t7_011011101), .y(t7_01101110));
wire t7_011011100, t7_011011101;
mixer mix_t7_01101111 (.a(t7_011011110), .b(t7_011011111), .y(t7_01101111));
wire t7_011011110, t7_011011111;
mixer mix_t7_0111 (.a(t7_01110), .b(t7_01111), .y(t7_0111));
wire t7_01110, t7_01111;
mixer mix_t7_01110 (.a(t7_011100), .b(t7_011101), .y(t7_01110));
wire t7_011100, t7_011101;
mixer mix_t7_011100 (.a(t7_0111000), .b(t7_0111001), .y(t7_011100));
wire t7_0111000, t7_0111001;
mixer mix_t7_0111000 (.a(t7_01110000), .b(t7_01110001), .y(t7_0111000));
wire t7_01110000, t7_01110001;
mixer mix_t7_01110000 (.a(t7_011100000), .b(t7_011100001), .y(t7_01110000));
wire t7_011100000, t7_011100001;
mixer mix_t7_01110001 (.a(t7_011100010), .b(t7_011100011), .y(t7_01110001));
wire t7_011100010, t7_011100011;
mixer mix_t7_0111001 (.a(t7_01110010), .b(t7_01110011), .y(t7_0111001));
wire t7_01110010, t7_01110011;
mixer mix_t7_01110010 (.a(t7_011100100), .b(t7_011100101), .y(t7_01110010));
wire t7_011100100, t7_011100101;
mixer mix_t7_01110011 (.a(t7_011100110), .b(t7_011100111), .y(t7_01110011));
wire t7_011100110, t7_011100111;
mixer mix_t7_011101 (.a(t7_0111010), .b(t7_0111011), .y(t7_011101));
wire t7_0111010, t7_0111011;
mixer mix_t7_0111010 (.a(t7_01110100), .b(t7_01110101), .y(t7_0111010));
wire t7_01110100, t7_01110101;
mixer mix_t7_01110100 (.a(t7_011101000), .b(t7_011101001), .y(t7_01110100));
wire t7_011101000, t7_011101001;
mixer mix_t7_01110101 (.a(t7_011101010), .b(t7_011101011), .y(t7_01110101));
wire t7_011101010, t7_011101011;
mixer mix_t7_0111011 (.a(t7_01110110), .b(t7_01110111), .y(t7_0111011));
wire t7_01110110, t7_01110111;
mixer mix_t7_01110110 (.a(t7_011101100), .b(t7_011101101), .y(t7_01110110));
wire t7_011101100, t7_011101101;
mixer mix_t7_01110111 (.a(t7_011101110), .b(t7_011101111), .y(t7_01110111));
wire t7_011101110, t7_011101111;
mixer mix_t7_01111 (.a(t7_011110), .b(t7_011111), .y(t7_01111));
wire t7_011110, t7_011111;
mixer mix_t7_011110 (.a(t7_0111100), .b(t7_0111101), .y(t7_011110));
wire t7_0111100, t7_0111101;
mixer mix_t7_0111100 (.a(t7_01111000), .b(t7_01111001), .y(t7_0111100));
wire t7_01111000, t7_01111001;
mixer mix_t7_01111000 (.a(t7_011110000), .b(t7_011110001), .y(t7_01111000));
wire t7_011110000, t7_011110001;
mixer mix_t7_01111001 (.a(t7_011110010), .b(t7_011110011), .y(t7_01111001));
wire t7_011110010, t7_011110011;
mixer mix_t7_0111101 (.a(t7_01111010), .b(t7_01111011), .y(t7_0111101));
wire t7_01111010, t7_01111011;
mixer mix_t7_01111010 (.a(t7_011110100), .b(t7_011110101), .y(t7_01111010));
wire t7_011110100, t7_011110101;
mixer mix_t7_01111011 (.a(t7_011110110), .b(t7_011110111), .y(t7_01111011));
wire t7_011110110, t7_011110111;
mixer mix_t7_011111 (.a(t7_0111110), .b(t7_0111111), .y(t7_011111));
wire t7_0111110, t7_0111111;
mixer mix_t7_0111110 (.a(t7_01111100), .b(t7_01111101), .y(t7_0111110));
wire t7_01111100, t7_01111101;
mixer mix_t7_01111100 (.a(t7_011111000), .b(t7_011111001), .y(t7_01111100));
wire t7_011111000, t7_011111001;
mixer mix_t7_01111101 (.a(t7_011111010), .b(t7_011111011), .y(t7_01111101));
wire t7_011111010, t7_011111011;
mixer mix_t7_0111111 (.a(t7_01111110), .b(t7_01111111), .y(t7_0111111));
wire t7_01111110, t7_01111111;
mixer mix_t7_01111110 (.a(t7_011111100), .b(t7_011111101), .y(t7_01111110));
wire t7_011111100, t7_011111101;
mixer mix_t7_01111111 (.a(t7_011111110), .b(t7_011111111), .y(t7_01111111));
wire t7_011111110, t7_011111111;
wire t0_0;
assign out_0 = t0_0;
wire t1_0;
assign out_1 = t1_0;
wire t2_0;
assign out_2 = t2_0;
wire t3_0;
assign out_3 = t3_0;
wire t4_0;
assign out_4 = t4_0;
wire t5_0;
assign out_5 = t5_0;
wire t6_0;
assign out_6 = t6_0;
wire t7_0;
assign out_7 = t7_0;
assign input_0 = t0_000000000;
assign input_1 = t0_000000001;
assign input_2 = t0_000000010;
assign input_3 = t0_000000011;
assign input_4 = t0_000000100;
assign input_5 = t0_000000101;
assign input_6 = t0_000000110;
assign input_7 = t0_000000111;
assign input_8 = t0_000001000;
assign input_9 = t0_000001001;
assign input_10 = t0_000001010;
assign input_11 = t0_000001011;
assign input_12 = t0_000001100;
assign input_13 = t0_000001101;
assign input_14 = t0_000001110;
assign input_15 = t0_000001111;
assign input_16 = t0_000010000;
assign input_17 = t0_000010001;
assign input_18 = t0_000010010;
assign input_19 = t0_000010011;
assign input_20 = t0_000010100;
assign input_21 = t0_000010101;
assign input_22 = t0_000010110;
assign input_23 = t0_000010111;
assign input_24 = t0_000011000;
assign input_25 = t0_000011001;
assign input_26 = t0_000011010;
assign input_27 = t0_000011011;
assign input_28 = t0_000011100;
assign input_29 = t0_000011101;
assign input_30 = t0_000011110;
assign input_31 = t0_000011111;
assign input_32 = t0_000100000;
assign input_33 = t0_000100001;
assign input_34 = t0_000100010;
assign input_35 = t0_000100011;
assign input_36 = t0_000100100;
assign input_37 = t0_000100101;
assign input_38 = t0_000100110;
assign input_39 = t0_000100111;
assign input_40 = t0_000101000;
assign input_41 = t0_000101001;
assign input_42 = t0_000101010;
assign input_43 = t0_000101011;
assign input_44 = t0_000101100;
assign input_45 = t0_000101101;
assign input_46 = t0_000101110;
assign input_47 = t0_000101111;
assign input_48 = t0_000110000;
assign input_49 = t0_000110001;
assign input_50 = t0_000110010;
assign input_51 = t0_000110011;
assign input_52 = t0_000110100;
assign input_53 = t0_000110101;
assign input_54 = t0_000110110;
assign input_55 = t0_000110111;
assign input_56 = t0_000111000;
assign input_57 = t0_000111001;
assign input_58 = t0_000111010;
assign input_59 = t0_000111011;
assign input_60 = t0_000111100;
assign input_61 = t0_000111101;
assign input_62 = t0_000111110;
assign input_63 = t0_000111111;
assign input_64 = t0_001000000;
assign input_65 = t0_001000001;
assign input_66 = t0_001000010;
assign input_67 = t0_001000011;
assign input_68 = t0_001000100;
assign input_69 = t0_001000101;
assign input_70 = t0_001000110;
assign input_71 = t0_001000111;
assign input_72 = t0_001001000;
assign input_73 = t0_001001001;
assign input_74 = t0_001001010;
assign input_75 = t0_001001011;
assign input_76 = t0_001001100;
assign input_77 = t0_001001101;
assign input_78 = t0_001001110;
assign input_79 = t0_001001111;
assign input_80 = t0_001010000;
assign input_81 = t0_001010001;
assign input_82 = t0_001010010;
assign input_83 = t0_001010011;
assign input_84 = t0_001010100;
assign input_85 = t0_001010101;
assign input_86 = t0_001010110;
assign input_87 = t0_001010111;
assign input_88 = t0_001011000;
assign input_89 = t0_001011001;
assign input_90 = t0_001011010;
assign input_91 = t0_001011011;
assign input_92 = t0_001011100;
assign input_93 = t0_001011101;
assign input_94 = t0_001011110;
assign input_95 = t0_001011111;
assign input_96 = t0_001100000;
assign input_97 = t0_001100001;
assign input_98 = t0_001100010;
assign input_99 = t0_001100011;
assign input_100 = t0_001100100;
assign input_101 = t0_001100101;
assign input_102 = t0_001100110;
assign input_103 = t0_001100111;
assign input_104 = t0_001101000;
assign input_105 = t0_001101001;
assign input_106 = t0_001101010;
assign input_107 = t0_001101011;
assign input_108 = t0_001101100;
assign input_109 = t0_001101101;
assign input_110 = t0_001101110;
assign input_111 = t0_001101111;
assign input_112 = t0_001110000;
assign input_113 = t0_001110001;
assign input_114 = t0_001110010;
assign input_115 = t0_001110011;
assign input_116 = t0_001110100;
assign input_117 = t0_001110101;
assign input_118 = t0_001110110;
assign input_119 = t0_001110111;
assign input_120 = t0_001111000;
assign input_121 = t0_001111001;
assign input_122 = t0_001111010;
assign input_123 = t0_001111011;
assign input_124 = t0_001111100;
assign input_125 = t0_001111101;
assign input_126 = t0_001111110;
assign input_127 = t0_001111111;
assign input_128 = t0_010000000;
assign input_129 = t0_010000001;
assign input_130 = t0_010000010;
assign input_131 = t0_010000011;
assign input_132 = t0_010000100;
assign input_133 = t0_010000101;
assign input_134 = t0_010000110;
assign input_135 = t0_010000111;
assign input_136 = t0_010001000;
assign input_137 = t0_010001001;
assign input_138 = t0_010001010;
assign input_139 = t0_010001011;
assign input_140 = t0_010001100;
assign input_141 = t0_010001101;
assign input_142 = t0_010001110;
assign input_143 = t0_010001111;
assign input_144 = t0_010010000;
assign input_145 = t0_010010001;
assign input_146 = t0_010010010;
assign input_147 = t0_010010011;
assign input_148 = t0_010010100;
assign input_149 = t0_010010101;
assign input_150 = t0_010010110;
assign input_151 = t0_010010111;
assign input_152 = t0_010011000;
assign input_153 = t0_010011001;
assign input_154 = t0_010011010;
assign input_155 = t0_010011011;
assign input_156 = t0_010011100;
assign input_157 = t0_010011101;
assign input_158 = t0_010011110;
assign input_159 = t0_010011111;
assign input_160 = t0_010100000;
assign input_161 = t0_010100001;
assign input_162 = t0_010100010;
assign input_163 = t0_010100011;
assign input_164 = t0_010100100;
assign input_165 = t0_010100101;
assign input_166 = t0_010100110;
assign input_167 = t0_010100111;
assign input_168 = t0_010101000;
assign input_169 = t0_010101001;
assign input_170 = t0_010101010;
assign input_171 = t0_010101011;
assign input_172 = t0_010101100;
assign input_173 = t0_010101101;
assign input_174 = t0_010101110;
assign input_175 = t0_010101111;
assign input_176 = t0_010110000;
assign input_177 = t0_010110001;
assign input_178 = t0_010110010;
assign input_179 = t0_010110011;
assign input_180 = t0_010110100;
assign input_181 = t0_010110101;
assign input_182 = t0_010110110;
assign input_183 = t0_010110111;
assign input_184 = t0_010111000;
assign input_185 = t0_010111001;
assign input_186 = t0_010111010;
assign input_187 = t0_010111011;
assign input_188 = t0_010111100;
assign input_189 = t0_010111101;
assign input_190 = t0_010111110;
assign input_191 = t0_010111111;
assign input_192 = t0_011000000;
assign input_193 = t0_011000001;
assign input_194 = t0_011000010;
assign input_195 = t0_011000011;
assign input_196 = t0_011000100;
assign input_197 = t0_011000101;
assign input_198 = t0_011000110;
assign input_199 = t0_011000111;
assign input_200 = t0_011001000;
assign input_201 = t0_011001001;
assign input_202 = t0_011001010;
assign input_203 = t0_011001011;
assign input_204 = t0_011001100;
assign input_205 = t0_011001101;
assign input_206 = t0_011001110;
assign input_207 = t0_011001111;
assign input_208 = t0_011010000;
assign input_209 = t0_011010001;
assign input_210 = t0_011010010;
assign input_211 = t0_011010011;
assign input_212 = t0_011010100;
assign input_213 = t0_011010101;
assign input_214 = t0_011010110;
assign input_215 = t0_011010111;
assign input_216 = t0_011011000;
assign input_217 = t0_011011001;
assign input_218 = t0_011011010;
assign input_219 = t0_011011011;
assign input_220 = t0_011011100;
assign input_221 = t0_011011101;
assign input_222 = t0_011011110;
assign input_223 = t0_011011111;
assign input_224 = t0_011100000;
assign input_225 = t0_011100001;
assign input_226 = t0_011100010;
assign input_227 = t0_011100011;
assign input_228 = t0_011100100;
assign input_229 = t0_011100101;
assign input_230 = t0_011100110;
assign input_231 = t0_011100111;
assign input_232 = t0_011101000;
assign input_233 = t0_011101001;
assign input_234 = t0_011101010;
assign input_235 = t0_011101011;
assign input_236 = t0_011101100;
assign input_237 = t0_011101101;
assign input_238 = t0_011101110;
assign input_239 = t0_011101111;
assign input_240 = t0_011110000;
assign input_241 = t0_011110001;
assign input_242 = t0_011110010;
assign input_243 = t0_011110011;
assign input_244 = t0_011110100;
assign input_245 = t0_011110101;
assign input_246 = t0_011110110;
assign input_247 = t0_011110111;
assign input_248 = t0_011111000;
assign input_249 = t0_011111001;
assign input_250 = t0_011111010;
assign input_251 = t0_011111011;
assign input_252 = t0_011111100;
assign input_253 = t0_011111101;
assign input_254 = t0_011111110;
assign input_255 = t0_011111111;
assign input_256 = t1_000000000;
assign input_257 = t1_000000001;
assign input_258 = t1_000000010;
assign input_259 = t1_000000011;
assign input_260 = t1_000000100;
assign input_261 = t1_000000101;
assign input_262 = t1_000000110;
assign input_263 = t1_000000111;
assign input_264 = t1_000001000;
assign input_265 = t1_000001001;
assign input_266 = t1_000001010;
assign input_267 = t1_000001011;
assign input_268 = t1_000001100;
assign input_269 = t1_000001101;
assign input_270 = t1_000001110;
assign input_271 = t1_000001111;
assign input_272 = t1_000010000;
assign input_273 = t1_000010001;
assign input_274 = t1_000010010;
assign input_275 = t1_000010011;
assign input_276 = t1_000010100;
assign input_277 = t1_000010101;
assign input_278 = t1_000010110;
assign input_279 = t1_000010111;
assign input_280 = t1_000011000;
assign input_281 = t1_000011001;
assign input_282 = t1_000011010;
assign input_283 = t1_000011011;
assign input_284 = t1_000011100;
assign input_285 = t1_000011101;
assign input_286 = t1_000011110;
assign input_287 = t1_000011111;
assign input_288 = t1_000100000;
assign input_289 = t1_000100001;
assign input_290 = t1_000100010;
assign input_291 = t1_000100011;
assign input_292 = t1_000100100;
assign input_293 = t1_000100101;
assign input_294 = t1_000100110;
assign input_295 = t1_000100111;
assign input_296 = t1_000101000;
assign input_297 = t1_000101001;
assign input_298 = t1_000101010;
assign input_299 = t1_000101011;
assign input_300 = t1_000101100;
assign input_301 = t1_000101101;
assign input_302 = t1_000101110;
assign input_303 = t1_000101111;
assign input_304 = t1_000110000;
assign input_305 = t1_000110001;
assign input_306 = t1_000110010;
assign input_307 = t1_000110011;
assign input_308 = t1_000110100;
assign input_309 = t1_000110101;
assign input_310 = t1_000110110;
assign input_311 = t1_000110111;
assign input_312 = t1_000111000;
assign input_313 = t1_000111001;
assign input_314 = t1_000111010;
assign input_315 = t1_000111011;
assign input_316 = t1_000111100;
assign input_317 = t1_000111101;
assign input_318 = t1_000111110;
assign input_319 = t1_000111111;
assign input_320 = t1_001000000;
assign input_321 = t1_001000001;
assign input_322 = t1_001000010;
assign input_323 = t1_001000011;
assign input_324 = t1_001000100;
assign input_325 = t1_001000101;
assign input_326 = t1_001000110;
assign input_327 = t1_001000111;
assign input_328 = t1_001001000;
assign input_329 = t1_001001001;
assign input_330 = t1_001001010;
assign input_331 = t1_001001011;
assign input_332 = t1_001001100;
assign input_333 = t1_001001101;
assign input_334 = t1_001001110;
assign input_335 = t1_001001111;
assign input_336 = t1_001010000;
assign input_337 = t1_001010001;
assign input_338 = t1_001010010;
assign input_339 = t1_001010011;
assign input_340 = t1_001010100;
assign input_341 = t1_001010101;
assign input_342 = t1_001010110;
assign input_343 = t1_001010111;
assign input_344 = t1_001011000;
assign input_345 = t1_001011001;
assign input_346 = t1_001011010;
assign input_347 = t1_001011011;
assign input_348 = t1_001011100;
assign input_349 = t1_001011101;
assign input_350 = t1_001011110;
assign input_351 = t1_001011111;
assign input_352 = t1_001100000;
assign input_353 = t1_001100001;
assign input_354 = t1_001100010;
assign input_355 = t1_001100011;
assign input_356 = t1_001100100;
assign input_357 = t1_001100101;
assign input_358 = t1_001100110;
assign input_359 = t1_001100111;
assign input_360 = t1_001101000;
assign input_361 = t1_001101001;
assign input_362 = t1_001101010;
assign input_363 = t1_001101011;
assign input_364 = t1_001101100;
assign input_365 = t1_001101101;
assign input_366 = t1_001101110;
assign input_367 = t1_001101111;
assign input_368 = t1_001110000;
assign input_369 = t1_001110001;
assign input_370 = t1_001110010;
assign input_371 = t1_001110011;
assign input_372 = t1_001110100;
assign input_373 = t1_001110101;
assign input_374 = t1_001110110;
assign input_375 = t1_001110111;
assign input_376 = t1_001111000;
assign input_377 = t1_001111001;
assign input_378 = t1_001111010;
assign input_379 = t1_001111011;
assign input_380 = t1_001111100;
assign input_381 = t1_001111101;
assign input_382 = t1_001111110;
assign input_383 = t1_001111111;
assign input_384 = t1_010000000;
assign input_385 = t1_010000001;
assign input_386 = t1_010000010;
assign input_387 = t1_010000011;
assign input_388 = t1_010000100;
assign input_389 = t1_010000101;
assign input_390 = t1_010000110;
assign input_391 = t1_010000111;
assign input_392 = t1_010001000;
assign input_393 = t1_010001001;
assign input_394 = t1_010001010;
assign input_395 = t1_010001011;
assign input_396 = t1_010001100;
assign input_397 = t1_010001101;
assign input_398 = t1_010001110;
assign input_399 = t1_010001111;
assign input_400 = t1_010010000;
assign input_401 = t1_010010001;
assign input_402 = t1_010010010;
assign input_403 = t1_010010011;
assign input_404 = t1_010010100;
assign input_405 = t1_010010101;
assign input_406 = t1_010010110;
assign input_407 = t1_010010111;
assign input_408 = t1_010011000;
assign input_409 = t1_010011001;
assign input_410 = t1_010011010;
assign input_411 = t1_010011011;
assign input_412 = t1_010011100;
assign input_413 = t1_010011101;
assign input_414 = t1_010011110;
assign input_415 = t1_010011111;
assign input_416 = t1_010100000;
assign input_417 = t1_010100001;
assign input_418 = t1_010100010;
assign input_419 = t1_010100011;
assign input_420 = t1_010100100;
assign input_421 = t1_010100101;
assign input_422 = t1_010100110;
assign input_423 = t1_010100111;
assign input_424 = t1_010101000;
assign input_425 = t1_010101001;
assign input_426 = t1_010101010;
assign input_427 = t1_010101011;
assign input_428 = t1_010101100;
assign input_429 = t1_010101101;
assign input_430 = t1_010101110;
assign input_431 = t1_010101111;
assign input_432 = t1_010110000;
assign input_433 = t1_010110001;
assign input_434 = t1_010110010;
assign input_435 = t1_010110011;
assign input_436 = t1_010110100;
assign input_437 = t1_010110101;
assign input_438 = t1_010110110;
assign input_439 = t1_010110111;
assign input_440 = t1_010111000;
assign input_441 = t1_010111001;
assign input_442 = t1_010111010;
assign input_443 = t1_010111011;
assign input_444 = t1_010111100;
assign input_445 = t1_010111101;
assign input_446 = t1_010111110;
assign input_447 = t1_010111111;
assign input_448 = t1_011000000;
assign input_449 = t1_011000001;
assign input_450 = t1_011000010;
assign input_451 = t1_011000011;
assign input_452 = t1_011000100;
assign input_453 = t1_011000101;
assign input_454 = t1_011000110;
assign input_455 = t1_011000111;
assign input_456 = t1_011001000;
assign input_457 = t1_011001001;
assign input_458 = t1_011001010;
assign input_459 = t1_011001011;
assign input_460 = t1_011001100;
assign input_461 = t1_011001101;
assign input_462 = t1_011001110;
assign input_463 = t1_011001111;
assign input_464 = t1_011010000;
assign input_465 = t1_011010001;
assign input_466 = t1_011010010;
assign input_467 = t1_011010011;
assign input_468 = t1_011010100;
assign input_469 = t1_011010101;
assign input_470 = t1_011010110;
assign input_471 = t1_011010111;
assign input_472 = t1_011011000;
assign input_473 = t1_011011001;
assign input_474 = t1_011011010;
assign input_475 = t1_011011011;
assign input_476 = t1_011011100;
assign input_477 = t1_011011101;
assign input_478 = t1_011011110;
assign input_479 = t1_011011111;
assign input_480 = t1_011100000;
assign input_481 = t1_011100001;
assign input_482 = t1_011100010;
assign input_483 = t1_011100011;
assign input_484 = t1_011100100;
assign input_485 = t1_011100101;
assign input_486 = t1_011100110;
assign input_487 = t1_011100111;
assign input_488 = t1_011101000;
assign input_489 = t1_011101001;
assign input_490 = t1_011101010;
assign input_491 = t1_011101011;
assign input_492 = t1_011101100;
assign input_493 = t1_011101101;
assign input_494 = t1_011101110;
assign input_495 = t1_011101111;
assign input_496 = t1_011110000;
assign input_497 = t1_011110001;
assign input_498 = t1_011110010;
assign input_499 = t1_011110011;
assign input_500 = t1_011110100;
assign input_501 = t1_011110101;
assign input_502 = t1_011110110;
assign input_503 = t1_011110111;
assign input_504 = t1_011111000;
assign input_505 = t1_011111001;
assign input_506 = t1_011111010;
assign input_507 = t1_011111011;
assign input_508 = t1_011111100;
assign input_509 = t1_011111101;
assign input_510 = t1_011111110;
assign input_511 = t1_011111111;
assign input_512 = t2_000000000;
assign input_513 = t2_000000001;
assign input_514 = t2_000000010;
assign input_515 = t2_000000011;
assign input_516 = t2_000000100;
assign input_517 = t2_000000101;
assign input_518 = t2_000000110;
assign input_519 = t2_000000111;
assign input_520 = t2_000001000;
assign input_521 = t2_000001001;
assign input_522 = t2_000001010;
assign input_523 = t2_000001011;
assign input_524 = t2_000001100;
assign input_525 = t2_000001101;
assign input_526 = t2_000001110;
assign input_527 = t2_000001111;
assign input_528 = t2_000010000;
assign input_529 = t2_000010001;
assign input_530 = t2_000010010;
assign input_531 = t2_000010011;
assign input_532 = t2_000010100;
assign input_533 = t2_000010101;
assign input_534 = t2_000010110;
assign input_535 = t2_000010111;
assign input_536 = t2_000011000;
assign input_537 = t2_000011001;
assign input_538 = t2_000011010;
assign input_539 = t2_000011011;
assign input_540 = t2_000011100;
assign input_541 = t2_000011101;
assign input_542 = t2_000011110;
assign input_543 = t2_000011111;
assign input_544 = t2_000100000;
assign input_545 = t2_000100001;
assign input_546 = t2_000100010;
assign input_547 = t2_000100011;
assign input_548 = t2_000100100;
assign input_549 = t2_000100101;
assign input_550 = t2_000100110;
assign input_551 = t2_000100111;
assign input_552 = t2_000101000;
assign input_553 = t2_000101001;
assign input_554 = t2_000101010;
assign input_555 = t2_000101011;
assign input_556 = t2_000101100;
assign input_557 = t2_000101101;
assign input_558 = t2_000101110;
assign input_559 = t2_000101111;
assign input_560 = t2_000110000;
assign input_561 = t2_000110001;
assign input_562 = t2_000110010;
assign input_563 = t2_000110011;
assign input_564 = t2_000110100;
assign input_565 = t2_000110101;
assign input_566 = t2_000110110;
assign input_567 = t2_000110111;
assign input_568 = t2_000111000;
assign input_569 = t2_000111001;
assign input_570 = t2_000111010;
assign input_571 = t2_000111011;
assign input_572 = t2_000111100;
assign input_573 = t2_000111101;
assign input_574 = t2_000111110;
assign input_575 = t2_000111111;
assign input_576 = t2_001000000;
assign input_577 = t2_001000001;
assign input_578 = t2_001000010;
assign input_579 = t2_001000011;
assign input_580 = t2_001000100;
assign input_581 = t2_001000101;
assign input_582 = t2_001000110;
assign input_583 = t2_001000111;
assign input_584 = t2_001001000;
assign input_585 = t2_001001001;
assign input_586 = t2_001001010;
assign input_587 = t2_001001011;
assign input_588 = t2_001001100;
assign input_589 = t2_001001101;
assign input_590 = t2_001001110;
assign input_591 = t2_001001111;
assign input_592 = t2_001010000;
assign input_593 = t2_001010001;
assign input_594 = t2_001010010;
assign input_595 = t2_001010011;
assign input_596 = t2_001010100;
assign input_597 = t2_001010101;
assign input_598 = t2_001010110;
assign input_599 = t2_001010111;
assign input_600 = t2_001011000;
assign input_601 = t2_001011001;
assign input_602 = t2_001011010;
assign input_603 = t2_001011011;
assign input_604 = t2_001011100;
assign input_605 = t2_001011101;
assign input_606 = t2_001011110;
assign input_607 = t2_001011111;
assign input_608 = t2_001100000;
assign input_609 = t2_001100001;
assign input_610 = t2_001100010;
assign input_611 = t2_001100011;
assign input_612 = t2_001100100;
assign input_613 = t2_001100101;
assign input_614 = t2_001100110;
assign input_615 = t2_001100111;
assign input_616 = t2_001101000;
assign input_617 = t2_001101001;
assign input_618 = t2_001101010;
assign input_619 = t2_001101011;
assign input_620 = t2_001101100;
assign input_621 = t2_001101101;
assign input_622 = t2_001101110;
assign input_623 = t2_001101111;
assign input_624 = t2_001110000;
assign input_625 = t2_001110001;
assign input_626 = t2_001110010;
assign input_627 = t2_001110011;
assign input_628 = t2_001110100;
assign input_629 = t2_001110101;
assign input_630 = t2_001110110;
assign input_631 = t2_001110111;
assign input_632 = t2_001111000;
assign input_633 = t2_001111001;
assign input_634 = t2_001111010;
assign input_635 = t2_001111011;
assign input_636 = t2_001111100;
assign input_637 = t2_001111101;
assign input_638 = t2_001111110;
assign input_639 = t2_001111111;
assign input_640 = t2_010000000;
assign input_641 = t2_010000001;
assign input_642 = t2_010000010;
assign input_643 = t2_010000011;
assign input_644 = t2_010000100;
assign input_645 = t2_010000101;
assign input_646 = t2_010000110;
assign input_647 = t2_010000111;
assign input_648 = t2_010001000;
assign input_649 = t2_010001001;
assign input_650 = t2_010001010;
assign input_651 = t2_010001011;
assign input_652 = t2_010001100;
assign input_653 = t2_010001101;
assign input_654 = t2_010001110;
assign input_655 = t2_010001111;
assign input_656 = t2_010010000;
assign input_657 = t2_010010001;
assign input_658 = t2_010010010;
assign input_659 = t2_010010011;
assign input_660 = t2_010010100;
assign input_661 = t2_010010101;
assign input_662 = t2_010010110;
assign input_663 = t2_010010111;
assign input_664 = t2_010011000;
assign input_665 = t2_010011001;
assign input_666 = t2_010011010;
assign input_667 = t2_010011011;
assign input_668 = t2_010011100;
assign input_669 = t2_010011101;
assign input_670 = t2_010011110;
assign input_671 = t2_010011111;
assign input_672 = t2_010100000;
assign input_673 = t2_010100001;
assign input_674 = t2_010100010;
assign input_675 = t2_010100011;
assign input_676 = t2_010100100;
assign input_677 = t2_010100101;
assign input_678 = t2_010100110;
assign input_679 = t2_010100111;
assign input_680 = t2_010101000;
assign input_681 = t2_010101001;
assign input_682 = t2_010101010;
assign input_683 = t2_010101011;
assign input_684 = t2_010101100;
assign input_685 = t2_010101101;
assign input_686 = t2_010101110;
assign input_687 = t2_010101111;
assign input_688 = t2_010110000;
assign input_689 = t2_010110001;
assign input_690 = t2_010110010;
assign input_691 = t2_010110011;
assign input_692 = t2_010110100;
assign input_693 = t2_010110101;
assign input_694 = t2_010110110;
assign input_695 = t2_010110111;
assign input_696 = t2_010111000;
assign input_697 = t2_010111001;
assign input_698 = t2_010111010;
assign input_699 = t2_010111011;
assign input_700 = t2_010111100;
assign input_701 = t2_010111101;
assign input_702 = t2_010111110;
assign input_703 = t2_010111111;
assign input_704 = t2_011000000;
assign input_705 = t2_011000001;
assign input_706 = t2_011000010;
assign input_707 = t2_011000011;
assign input_708 = t2_011000100;
assign input_709 = t2_011000101;
assign input_710 = t2_011000110;
assign input_711 = t2_011000111;
assign input_712 = t2_011001000;
assign input_713 = t2_011001001;
assign input_714 = t2_011001010;
assign input_715 = t2_011001011;
assign input_716 = t2_011001100;
assign input_717 = t2_011001101;
assign input_718 = t2_011001110;
assign input_719 = t2_011001111;
assign input_720 = t2_011010000;
assign input_721 = t2_011010001;
assign input_722 = t2_011010010;
assign input_723 = t2_011010011;
assign input_724 = t2_011010100;
assign input_725 = t2_011010101;
assign input_726 = t2_011010110;
assign input_727 = t2_011010111;
assign input_728 = t2_011011000;
assign input_729 = t2_011011001;
assign input_730 = t2_011011010;
assign input_731 = t2_011011011;
assign input_732 = t2_011011100;
assign input_733 = t2_011011101;
assign input_734 = t2_011011110;
assign input_735 = t2_011011111;
assign input_736 = t2_011100000;
assign input_737 = t2_011100001;
assign input_738 = t2_011100010;
assign input_739 = t2_011100011;
assign input_740 = t2_011100100;
assign input_741 = t2_011100101;
assign input_742 = t2_011100110;
assign input_743 = t2_011100111;
assign input_744 = t2_011101000;
assign input_745 = t2_011101001;
assign input_746 = t2_011101010;
assign input_747 = t2_011101011;
assign input_748 = t2_011101100;
assign input_749 = t2_011101101;
assign input_750 = t2_011101110;
assign input_751 = t2_011101111;
assign input_752 = t2_011110000;
assign input_753 = t2_011110001;
assign input_754 = t2_011110010;
assign input_755 = t2_011110011;
assign input_756 = t2_011110100;
assign input_757 = t2_011110101;
assign input_758 = t2_011110110;
assign input_759 = t2_011110111;
assign input_760 = t2_011111000;
assign input_761 = t2_011111001;
assign input_762 = t2_011111010;
assign input_763 = t2_011111011;
assign input_764 = t2_011111100;
assign input_765 = t2_011111101;
assign input_766 = t2_011111110;
assign input_767 = t2_011111111;
assign input_768 = t3_000000000;
assign input_769 = t3_000000001;
assign input_770 = t3_000000010;
assign input_771 = t3_000000011;
assign input_772 = t3_000000100;
assign input_773 = t3_000000101;
assign input_774 = t3_000000110;
assign input_775 = t3_000000111;
assign input_776 = t3_000001000;
assign input_777 = t3_000001001;
assign input_778 = t3_000001010;
assign input_779 = t3_000001011;
assign input_780 = t3_000001100;
assign input_781 = t3_000001101;
assign input_782 = t3_000001110;
assign input_783 = t3_000001111;
assign input_784 = t3_000010000;
assign input_785 = t3_000010001;
assign input_786 = t3_000010010;
assign input_787 = t3_000010011;
assign input_788 = t3_000010100;
assign input_789 = t3_000010101;
assign input_790 = t3_000010110;
assign input_791 = t3_000010111;
assign input_792 = t3_000011000;
assign input_793 = t3_000011001;
assign input_794 = t3_000011010;
assign input_795 = t3_000011011;
assign input_796 = t3_000011100;
assign input_797 = t3_000011101;
assign input_798 = t3_000011110;
assign input_799 = t3_000011111;
assign input_800 = t3_000100000;
assign input_801 = t3_000100001;
assign input_802 = t3_000100010;
assign input_803 = t3_000100011;
assign input_804 = t3_000100100;
assign input_805 = t3_000100101;
assign input_806 = t3_000100110;
assign input_807 = t3_000100111;
assign input_808 = t3_000101000;
assign input_809 = t3_000101001;
assign input_810 = t3_000101010;
assign input_811 = t3_000101011;
assign input_812 = t3_000101100;
assign input_813 = t3_000101101;
assign input_814 = t3_000101110;
assign input_815 = t3_000101111;
assign input_816 = t3_000110000;
assign input_817 = t3_000110001;
assign input_818 = t3_000110010;
assign input_819 = t3_000110011;
assign input_820 = t3_000110100;
assign input_821 = t3_000110101;
assign input_822 = t3_000110110;
assign input_823 = t3_000110111;
assign input_824 = t3_000111000;
assign input_825 = t3_000111001;
assign input_826 = t3_000111010;
assign input_827 = t3_000111011;
assign input_828 = t3_000111100;
assign input_829 = t3_000111101;
assign input_830 = t3_000111110;
assign input_831 = t3_000111111;
assign input_832 = t3_001000000;
assign input_833 = t3_001000001;
assign input_834 = t3_001000010;
assign input_835 = t3_001000011;
assign input_836 = t3_001000100;
assign input_837 = t3_001000101;
assign input_838 = t3_001000110;
assign input_839 = t3_001000111;
assign input_840 = t3_001001000;
assign input_841 = t3_001001001;
assign input_842 = t3_001001010;
assign input_843 = t3_001001011;
assign input_844 = t3_001001100;
assign input_845 = t3_001001101;
assign input_846 = t3_001001110;
assign input_847 = t3_001001111;
assign input_848 = t3_001010000;
assign input_849 = t3_001010001;
assign input_850 = t3_001010010;
assign input_851 = t3_001010011;
assign input_852 = t3_001010100;
assign input_853 = t3_001010101;
assign input_854 = t3_001010110;
assign input_855 = t3_001010111;
assign input_856 = t3_001011000;
assign input_857 = t3_001011001;
assign input_858 = t3_001011010;
assign input_859 = t3_001011011;
assign input_860 = t3_001011100;
assign input_861 = t3_001011101;
assign input_862 = t3_001011110;
assign input_863 = t3_001011111;
assign input_864 = t3_001100000;
assign input_865 = t3_001100001;
assign input_866 = t3_001100010;
assign input_867 = t3_001100011;
assign input_868 = t3_001100100;
assign input_869 = t3_001100101;
assign input_870 = t3_001100110;
assign input_871 = t3_001100111;
assign input_872 = t3_001101000;
assign input_873 = t3_001101001;
assign input_874 = t3_001101010;
assign input_875 = t3_001101011;
assign input_876 = t3_001101100;
assign input_877 = t3_001101101;
assign input_878 = t3_001101110;
assign input_879 = t3_001101111;
assign input_880 = t3_001110000;
assign input_881 = t3_001110001;
assign input_882 = t3_001110010;
assign input_883 = t3_001110011;
assign input_884 = t3_001110100;
assign input_885 = t3_001110101;
assign input_886 = t3_001110110;
assign input_887 = t3_001110111;
assign input_888 = t3_001111000;
assign input_889 = t3_001111001;
assign input_890 = t3_001111010;
assign input_891 = t3_001111011;
assign input_892 = t3_001111100;
assign input_893 = t3_001111101;
assign input_894 = t3_001111110;
assign input_895 = t3_001111111;
assign input_896 = t3_010000000;
assign input_897 = t3_010000001;
assign input_898 = t3_010000010;
assign input_899 = t3_010000011;
assign input_900 = t3_010000100;
assign input_901 = t3_010000101;
assign input_902 = t3_010000110;
assign input_903 = t3_010000111;
assign input_904 = t3_010001000;
assign input_905 = t3_010001001;
assign input_906 = t3_010001010;
assign input_907 = t3_010001011;
assign input_908 = t3_010001100;
assign input_909 = t3_010001101;
assign input_910 = t3_010001110;
assign input_911 = t3_010001111;
assign input_912 = t3_010010000;
assign input_913 = t3_010010001;
assign input_914 = t3_010010010;
assign input_915 = t3_010010011;
assign input_916 = t3_010010100;
assign input_917 = t3_010010101;
assign input_918 = t3_010010110;
assign input_919 = t3_010010111;
assign input_920 = t3_010011000;
assign input_921 = t3_010011001;
assign input_922 = t3_010011010;
assign input_923 = t3_010011011;
assign input_924 = t3_010011100;
assign input_925 = t3_010011101;
assign input_926 = t3_010011110;
assign input_927 = t3_010011111;
assign input_928 = t3_010100000;
assign input_929 = t3_010100001;
assign input_930 = t3_010100010;
assign input_931 = t3_010100011;
assign input_932 = t3_010100100;
assign input_933 = t3_010100101;
assign input_934 = t3_010100110;
assign input_935 = t3_010100111;
assign input_936 = t3_010101000;
assign input_937 = t3_010101001;
assign input_938 = t3_010101010;
assign input_939 = t3_010101011;
assign input_940 = t3_010101100;
assign input_941 = t3_010101101;
assign input_942 = t3_010101110;
assign input_943 = t3_010101111;
assign input_944 = t3_010110000;
assign input_945 = t3_010110001;
assign input_946 = t3_010110010;
assign input_947 = t3_010110011;
assign input_948 = t3_010110100;
assign input_949 = t3_010110101;
assign input_950 = t3_010110110;
assign input_951 = t3_010110111;
assign input_952 = t3_010111000;
assign input_953 = t3_010111001;
assign input_954 = t3_010111010;
assign input_955 = t3_010111011;
assign input_956 = t3_010111100;
assign input_957 = t3_010111101;
assign input_958 = t3_010111110;
assign input_959 = t3_010111111;
assign input_960 = t3_011000000;
assign input_961 = t3_011000001;
assign input_962 = t3_011000010;
assign input_963 = t3_011000011;
assign input_964 = t3_011000100;
assign input_965 = t3_011000101;
assign input_966 = t3_011000110;
assign input_967 = t3_011000111;
assign input_968 = t3_011001000;
assign input_969 = t3_011001001;
assign input_970 = t3_011001010;
assign input_971 = t3_011001011;
assign input_972 = t3_011001100;
assign input_973 = t3_011001101;
assign input_974 = t3_011001110;
assign input_975 = t3_011001111;
assign input_976 = t3_011010000;
assign input_977 = t3_011010001;
assign input_978 = t3_011010010;
assign input_979 = t3_011010011;
assign input_980 = t3_011010100;
assign input_981 = t3_011010101;
assign input_982 = t3_011010110;
assign input_983 = t3_011010111;
assign input_984 = t3_011011000;
assign input_985 = t3_011011001;
assign input_986 = t3_011011010;
assign input_987 = t3_011011011;
assign input_988 = t3_011011100;
assign input_989 = t3_011011101;
assign input_990 = t3_011011110;
assign input_991 = t3_011011111;
assign input_992 = t3_011100000;
assign input_993 = t3_011100001;
assign input_994 = t3_011100010;
assign input_995 = t3_011100011;
assign input_996 = t3_011100100;
assign input_997 = t3_011100101;
assign input_998 = t3_011100110;
assign input_999 = t3_011100111;
assign input_1000 = t3_011101000;
assign input_1001 = t3_011101001;
assign input_1002 = t3_011101010;
assign input_1003 = t3_011101011;
assign input_1004 = t3_011101100;
assign input_1005 = t3_011101101;
assign input_1006 = t3_011101110;
assign input_1007 = t3_011101111;
assign input_1008 = t3_011110000;
assign input_1009 = t3_011110001;
assign input_1010 = t3_011110010;
assign input_1011 = t3_011110011;
assign input_1012 = t3_011110100;
assign input_1013 = t3_011110101;
assign input_1014 = t3_011110110;
assign input_1015 = t3_011110111;
assign input_1016 = t3_011111000;
assign input_1017 = t3_011111001;
assign input_1018 = t3_011111010;
assign input_1019 = t3_011111011;
assign input_1020 = t3_011111100;
assign input_1021 = t3_011111101;
assign input_1022 = t3_011111110;
assign input_1023 = t3_011111111;
assign input_1024 = t4_000000000;
assign input_1025 = t4_000000001;
assign input_1026 = t4_000000010;
assign input_1027 = t4_000000011;
assign input_1028 = t4_000000100;
assign input_1029 = t4_000000101;
assign input_1030 = t4_000000110;
assign input_1031 = t4_000000111;
assign input_1032 = t4_000001000;
assign input_1033 = t4_000001001;
assign input_1034 = t4_000001010;
assign input_1035 = t4_000001011;
assign input_1036 = t4_000001100;
assign input_1037 = t4_000001101;
assign input_1038 = t4_000001110;
assign input_1039 = t4_000001111;
assign input_1040 = t4_000010000;
assign input_1041 = t4_000010001;
assign input_1042 = t4_000010010;
assign input_1043 = t4_000010011;
assign input_1044 = t4_000010100;
assign input_1045 = t4_000010101;
assign input_1046 = t4_000010110;
assign input_1047 = t4_000010111;
assign input_1048 = t4_000011000;
assign input_1049 = t4_000011001;
assign input_1050 = t4_000011010;
assign input_1051 = t4_000011011;
assign input_1052 = t4_000011100;
assign input_1053 = t4_000011101;
assign input_1054 = t4_000011110;
assign input_1055 = t4_000011111;
assign input_1056 = t4_000100000;
assign input_1057 = t4_000100001;
assign input_1058 = t4_000100010;
assign input_1059 = t4_000100011;
assign input_1060 = t4_000100100;
assign input_1061 = t4_000100101;
assign input_1062 = t4_000100110;
assign input_1063 = t4_000100111;
assign input_1064 = t4_000101000;
assign input_1065 = t4_000101001;
assign input_1066 = t4_000101010;
assign input_1067 = t4_000101011;
assign input_1068 = t4_000101100;
assign input_1069 = t4_000101101;
assign input_1070 = t4_000101110;
assign input_1071 = t4_000101111;
assign input_1072 = t4_000110000;
assign input_1073 = t4_000110001;
assign input_1074 = t4_000110010;
assign input_1075 = t4_000110011;
assign input_1076 = t4_000110100;
assign input_1077 = t4_000110101;
assign input_1078 = t4_000110110;
assign input_1079 = t4_000110111;
assign input_1080 = t4_000111000;
assign input_1081 = t4_000111001;
assign input_1082 = t4_000111010;
assign input_1083 = t4_000111011;
assign input_1084 = t4_000111100;
assign input_1085 = t4_000111101;
assign input_1086 = t4_000111110;
assign input_1087 = t4_000111111;
assign input_1088 = t4_001000000;
assign input_1089 = t4_001000001;
assign input_1090 = t4_001000010;
assign input_1091 = t4_001000011;
assign input_1092 = t4_001000100;
assign input_1093 = t4_001000101;
assign input_1094 = t4_001000110;
assign input_1095 = t4_001000111;
assign input_1096 = t4_001001000;
assign input_1097 = t4_001001001;
assign input_1098 = t4_001001010;
assign input_1099 = t4_001001011;
assign input_1100 = t4_001001100;
assign input_1101 = t4_001001101;
assign input_1102 = t4_001001110;
assign input_1103 = t4_001001111;
assign input_1104 = t4_001010000;
assign input_1105 = t4_001010001;
assign input_1106 = t4_001010010;
assign input_1107 = t4_001010011;
assign input_1108 = t4_001010100;
assign input_1109 = t4_001010101;
assign input_1110 = t4_001010110;
assign input_1111 = t4_001010111;
assign input_1112 = t4_001011000;
assign input_1113 = t4_001011001;
assign input_1114 = t4_001011010;
assign input_1115 = t4_001011011;
assign input_1116 = t4_001011100;
assign input_1117 = t4_001011101;
assign input_1118 = t4_001011110;
assign input_1119 = t4_001011111;
assign input_1120 = t4_001100000;
assign input_1121 = t4_001100001;
assign input_1122 = t4_001100010;
assign input_1123 = t4_001100011;
assign input_1124 = t4_001100100;
assign input_1125 = t4_001100101;
assign input_1126 = t4_001100110;
assign input_1127 = t4_001100111;
assign input_1128 = t4_001101000;
assign input_1129 = t4_001101001;
assign input_1130 = t4_001101010;
assign input_1131 = t4_001101011;
assign input_1132 = t4_001101100;
assign input_1133 = t4_001101101;
assign input_1134 = t4_001101110;
assign input_1135 = t4_001101111;
assign input_1136 = t4_001110000;
assign input_1137 = t4_001110001;
assign input_1138 = t4_001110010;
assign input_1139 = t4_001110011;
assign input_1140 = t4_001110100;
assign input_1141 = t4_001110101;
assign input_1142 = t4_001110110;
assign input_1143 = t4_001110111;
assign input_1144 = t4_001111000;
assign input_1145 = t4_001111001;
assign input_1146 = t4_001111010;
assign input_1147 = t4_001111011;
assign input_1148 = t4_001111100;
assign input_1149 = t4_001111101;
assign input_1150 = t4_001111110;
assign input_1151 = t4_001111111;
assign input_1152 = t4_010000000;
assign input_1153 = t4_010000001;
assign input_1154 = t4_010000010;
assign input_1155 = t4_010000011;
assign input_1156 = t4_010000100;
assign input_1157 = t4_010000101;
assign input_1158 = t4_010000110;
assign input_1159 = t4_010000111;
assign input_1160 = t4_010001000;
assign input_1161 = t4_010001001;
assign input_1162 = t4_010001010;
assign input_1163 = t4_010001011;
assign input_1164 = t4_010001100;
assign input_1165 = t4_010001101;
assign input_1166 = t4_010001110;
assign input_1167 = t4_010001111;
assign input_1168 = t4_010010000;
assign input_1169 = t4_010010001;
assign input_1170 = t4_010010010;
assign input_1171 = t4_010010011;
assign input_1172 = t4_010010100;
assign input_1173 = t4_010010101;
assign input_1174 = t4_010010110;
assign input_1175 = t4_010010111;
assign input_1176 = t4_010011000;
assign input_1177 = t4_010011001;
assign input_1178 = t4_010011010;
assign input_1179 = t4_010011011;
assign input_1180 = t4_010011100;
assign input_1181 = t4_010011101;
assign input_1182 = t4_010011110;
assign input_1183 = t4_010011111;
assign input_1184 = t4_010100000;
assign input_1185 = t4_010100001;
assign input_1186 = t4_010100010;
assign input_1187 = t4_010100011;
assign input_1188 = t4_010100100;
assign input_1189 = t4_010100101;
assign input_1190 = t4_010100110;
assign input_1191 = t4_010100111;
assign input_1192 = t4_010101000;
assign input_1193 = t4_010101001;
assign input_1194 = t4_010101010;
assign input_1195 = t4_010101011;
assign input_1196 = t4_010101100;
assign input_1197 = t4_010101101;
assign input_1198 = t4_010101110;
assign input_1199 = t4_010101111;
assign input_1200 = t4_010110000;
assign input_1201 = t4_010110001;
assign input_1202 = t4_010110010;
assign input_1203 = t4_010110011;
assign input_1204 = t4_010110100;
assign input_1205 = t4_010110101;
assign input_1206 = t4_010110110;
assign input_1207 = t4_010110111;
assign input_1208 = t4_010111000;
assign input_1209 = t4_010111001;
assign input_1210 = t4_010111010;
assign input_1211 = t4_010111011;
assign input_1212 = t4_010111100;
assign input_1213 = t4_010111101;
assign input_1214 = t4_010111110;
assign input_1215 = t4_010111111;
assign input_1216 = t4_011000000;
assign input_1217 = t4_011000001;
assign input_1218 = t4_011000010;
assign input_1219 = t4_011000011;
assign input_1220 = t4_011000100;
assign input_1221 = t4_011000101;
assign input_1222 = t4_011000110;
assign input_1223 = t4_011000111;
assign input_1224 = t4_011001000;
assign input_1225 = t4_011001001;
assign input_1226 = t4_011001010;
assign input_1227 = t4_011001011;
assign input_1228 = t4_011001100;
assign input_1229 = t4_011001101;
assign input_1230 = t4_011001110;
assign input_1231 = t4_011001111;
assign input_1232 = t4_011010000;
assign input_1233 = t4_011010001;
assign input_1234 = t4_011010010;
assign input_1235 = t4_011010011;
assign input_1236 = t4_011010100;
assign input_1237 = t4_011010101;
assign input_1238 = t4_011010110;
assign input_1239 = t4_011010111;
assign input_1240 = t4_011011000;
assign input_1241 = t4_011011001;
assign input_1242 = t4_011011010;
assign input_1243 = t4_011011011;
assign input_1244 = t4_011011100;
assign input_1245 = t4_011011101;
assign input_1246 = t4_011011110;
assign input_1247 = t4_011011111;
assign input_1248 = t4_011100000;
assign input_1249 = t4_011100001;
assign input_1250 = t4_011100010;
assign input_1251 = t4_011100011;
assign input_1252 = t4_011100100;
assign input_1253 = t4_011100101;
assign input_1254 = t4_011100110;
assign input_1255 = t4_011100111;
assign input_1256 = t4_011101000;
assign input_1257 = t4_011101001;
assign input_1258 = t4_011101010;
assign input_1259 = t4_011101011;
assign input_1260 = t4_011101100;
assign input_1261 = t4_011101101;
assign input_1262 = t4_011101110;
assign input_1263 = t4_011101111;
assign input_1264 = t4_011110000;
assign input_1265 = t4_011110001;
assign input_1266 = t4_011110010;
assign input_1267 = t4_011110011;
assign input_1268 = t4_011110100;
assign input_1269 = t4_011110101;
assign input_1270 = t4_011110110;
assign input_1271 = t4_011110111;
assign input_1272 = t4_011111000;
assign input_1273 = t4_011111001;
assign input_1274 = t4_011111010;
assign input_1275 = t4_011111011;
assign input_1276 = t4_011111100;
assign input_1277 = t4_011111101;
assign input_1278 = t4_011111110;
assign input_1279 = t4_011111111;
assign input_1280 = t5_000000000;
assign input_1281 = t5_000000001;
assign input_1282 = t5_000000010;
assign input_1283 = t5_000000011;
assign input_1284 = t5_000000100;
assign input_1285 = t5_000000101;
assign input_1286 = t5_000000110;
assign input_1287 = t5_000000111;
assign input_1288 = t5_000001000;
assign input_1289 = t5_000001001;
assign input_1290 = t5_000001010;
assign input_1291 = t5_000001011;
assign input_1292 = t5_000001100;
assign input_1293 = t5_000001101;
assign input_1294 = t5_000001110;
assign input_1295 = t5_000001111;
assign input_1296 = t5_000010000;
assign input_1297 = t5_000010001;
assign input_1298 = t5_000010010;
assign input_1299 = t5_000010011;
assign input_1300 = t5_000010100;
assign input_1301 = t5_000010101;
assign input_1302 = t5_000010110;
assign input_1303 = t5_000010111;
assign input_1304 = t5_000011000;
assign input_1305 = t5_000011001;
assign input_1306 = t5_000011010;
assign input_1307 = t5_000011011;
assign input_1308 = t5_000011100;
assign input_1309 = t5_000011101;
assign input_1310 = t5_000011110;
assign input_1311 = t5_000011111;
assign input_1312 = t5_000100000;
assign input_1313 = t5_000100001;
assign input_1314 = t5_000100010;
assign input_1315 = t5_000100011;
assign input_1316 = t5_000100100;
assign input_1317 = t5_000100101;
assign input_1318 = t5_000100110;
assign input_1319 = t5_000100111;
assign input_1320 = t5_000101000;
assign input_1321 = t5_000101001;
assign input_1322 = t5_000101010;
assign input_1323 = t5_000101011;
assign input_1324 = t5_000101100;
assign input_1325 = t5_000101101;
assign input_1326 = t5_000101110;
assign input_1327 = t5_000101111;
assign input_1328 = t5_000110000;
assign input_1329 = t5_000110001;
assign input_1330 = t5_000110010;
assign input_1331 = t5_000110011;
assign input_1332 = t5_000110100;
assign input_1333 = t5_000110101;
assign input_1334 = t5_000110110;
assign input_1335 = t5_000110111;
assign input_1336 = t5_000111000;
assign input_1337 = t5_000111001;
assign input_1338 = t5_000111010;
assign input_1339 = t5_000111011;
assign input_1340 = t5_000111100;
assign input_1341 = t5_000111101;
assign input_1342 = t5_000111110;
assign input_1343 = t5_000111111;
assign input_1344 = t5_001000000;
assign input_1345 = t5_001000001;
assign input_1346 = t5_001000010;
assign input_1347 = t5_001000011;
assign input_1348 = t5_001000100;
assign input_1349 = t5_001000101;
assign input_1350 = t5_001000110;
assign input_1351 = t5_001000111;
assign input_1352 = t5_001001000;
assign input_1353 = t5_001001001;
assign input_1354 = t5_001001010;
assign input_1355 = t5_001001011;
assign input_1356 = t5_001001100;
assign input_1357 = t5_001001101;
assign input_1358 = t5_001001110;
assign input_1359 = t5_001001111;
assign input_1360 = t5_001010000;
assign input_1361 = t5_001010001;
assign input_1362 = t5_001010010;
assign input_1363 = t5_001010011;
assign input_1364 = t5_001010100;
assign input_1365 = t5_001010101;
assign input_1366 = t5_001010110;
assign input_1367 = t5_001010111;
assign input_1368 = t5_001011000;
assign input_1369 = t5_001011001;
assign input_1370 = t5_001011010;
assign input_1371 = t5_001011011;
assign input_1372 = t5_001011100;
assign input_1373 = t5_001011101;
assign input_1374 = t5_001011110;
assign input_1375 = t5_001011111;
assign input_1376 = t5_001100000;
assign input_1377 = t5_001100001;
assign input_1378 = t5_001100010;
assign input_1379 = t5_001100011;
assign input_1380 = t5_001100100;
assign input_1381 = t5_001100101;
assign input_1382 = t5_001100110;
assign input_1383 = t5_001100111;
assign input_1384 = t5_001101000;
assign input_1385 = t5_001101001;
assign input_1386 = t5_001101010;
assign input_1387 = t5_001101011;
assign input_1388 = t5_001101100;
assign input_1389 = t5_001101101;
assign input_1390 = t5_001101110;
assign input_1391 = t5_001101111;
assign input_1392 = t5_001110000;
assign input_1393 = t5_001110001;
assign input_1394 = t5_001110010;
assign input_1395 = t5_001110011;
assign input_1396 = t5_001110100;
assign input_1397 = t5_001110101;
assign input_1398 = t5_001110110;
assign input_1399 = t5_001110111;
assign input_1400 = t5_001111000;
assign input_1401 = t5_001111001;
assign input_1402 = t5_001111010;
assign input_1403 = t5_001111011;
assign input_1404 = t5_001111100;
assign input_1405 = t5_001111101;
assign input_1406 = t5_001111110;
assign input_1407 = t5_001111111;
assign input_1408 = t5_010000000;
assign input_1409 = t5_010000001;
assign input_1410 = t5_010000010;
assign input_1411 = t5_010000011;
assign input_1412 = t5_010000100;
assign input_1413 = t5_010000101;
assign input_1414 = t5_010000110;
assign input_1415 = t5_010000111;
assign input_1416 = t5_010001000;
assign input_1417 = t5_010001001;
assign input_1418 = t5_010001010;
assign input_1419 = t5_010001011;
assign input_1420 = t5_010001100;
assign input_1421 = t5_010001101;
assign input_1422 = t5_010001110;
assign input_1423 = t5_010001111;
assign input_1424 = t5_010010000;
assign input_1425 = t5_010010001;
assign input_1426 = t5_010010010;
assign input_1427 = t5_010010011;
assign input_1428 = t5_010010100;
assign input_1429 = t5_010010101;
assign input_1430 = t5_010010110;
assign input_1431 = t5_010010111;
assign input_1432 = t5_010011000;
assign input_1433 = t5_010011001;
assign input_1434 = t5_010011010;
assign input_1435 = t5_010011011;
assign input_1436 = t5_010011100;
assign input_1437 = t5_010011101;
assign input_1438 = t5_010011110;
assign input_1439 = t5_010011111;
assign input_1440 = t5_010100000;
assign input_1441 = t5_010100001;
assign input_1442 = t5_010100010;
assign input_1443 = t5_010100011;
assign input_1444 = t5_010100100;
assign input_1445 = t5_010100101;
assign input_1446 = t5_010100110;
assign input_1447 = t5_010100111;
assign input_1448 = t5_010101000;
assign input_1449 = t5_010101001;
assign input_1450 = t5_010101010;
assign input_1451 = t5_010101011;
assign input_1452 = t5_010101100;
assign input_1453 = t5_010101101;
assign input_1454 = t5_010101110;
assign input_1455 = t5_010101111;
assign input_1456 = t5_010110000;
assign input_1457 = t5_010110001;
assign input_1458 = t5_010110010;
assign input_1459 = t5_010110011;
assign input_1460 = t5_010110100;
assign input_1461 = t5_010110101;
assign input_1462 = t5_010110110;
assign input_1463 = t5_010110111;
assign input_1464 = t5_010111000;
assign input_1465 = t5_010111001;
assign input_1466 = t5_010111010;
assign input_1467 = t5_010111011;
assign input_1468 = t5_010111100;
assign input_1469 = t5_010111101;
assign input_1470 = t5_010111110;
assign input_1471 = t5_010111111;
assign input_1472 = t5_011000000;
assign input_1473 = t5_011000001;
assign input_1474 = t5_011000010;
assign input_1475 = t5_011000011;
assign input_1476 = t5_011000100;
assign input_1477 = t5_011000101;
assign input_1478 = t5_011000110;
assign input_1479 = t5_011000111;
assign input_1480 = t5_011001000;
assign input_1481 = t5_011001001;
assign input_1482 = t5_011001010;
assign input_1483 = t5_011001011;
assign input_1484 = t5_011001100;
assign input_1485 = t5_011001101;
assign input_1486 = t5_011001110;
assign input_1487 = t5_011001111;
assign input_1488 = t5_011010000;
assign input_1489 = t5_011010001;
assign input_1490 = t5_011010010;
assign input_1491 = t5_011010011;
assign input_1492 = t5_011010100;
assign input_1493 = t5_011010101;
assign input_1494 = t5_011010110;
assign input_1495 = t5_011010111;
assign input_1496 = t5_011011000;
assign input_1497 = t5_011011001;
assign input_1498 = t5_011011010;
assign input_1499 = t5_011011011;
assign input_1500 = t5_011011100;
assign input_1501 = t5_011011101;
assign input_1502 = t5_011011110;
assign input_1503 = t5_011011111;
assign input_1504 = t5_011100000;
assign input_1505 = t5_011100001;
assign input_1506 = t5_011100010;
assign input_1507 = t5_011100011;
assign input_1508 = t5_011100100;
assign input_1509 = t5_011100101;
assign input_1510 = t5_011100110;
assign input_1511 = t5_011100111;
assign input_1512 = t5_011101000;
assign input_1513 = t5_011101001;
assign input_1514 = t5_011101010;
assign input_1515 = t5_011101011;
assign input_1516 = t5_011101100;
assign input_1517 = t5_011101101;
assign input_1518 = t5_011101110;
assign input_1519 = t5_011101111;
assign input_1520 = t5_011110000;
assign input_1521 = t5_011110001;
assign input_1522 = t5_011110010;
assign input_1523 = t5_011110011;
assign input_1524 = t5_011110100;
assign input_1525 = t5_011110101;
assign input_1526 = t5_011110110;
assign input_1527 = t5_011110111;
assign input_1528 = t5_011111000;
assign input_1529 = t5_011111001;
assign input_1530 = t5_011111010;
assign input_1531 = t5_011111011;
assign input_1532 = t5_011111100;
assign input_1533 = t5_011111101;
assign input_1534 = t5_011111110;
assign input_1535 = t5_011111111;
assign input_1536 = t6_000000000;
assign input_1537 = t6_000000001;
assign input_1538 = t6_000000010;
assign input_1539 = t6_000000011;
assign input_1540 = t6_000000100;
assign input_1541 = t6_000000101;
assign input_1542 = t6_000000110;
assign input_1543 = t6_000000111;
assign input_1544 = t6_000001000;
assign input_1545 = t6_000001001;
assign input_1546 = t6_000001010;
assign input_1547 = t6_000001011;
assign input_1548 = t6_000001100;
assign input_1549 = t6_000001101;
assign input_1550 = t6_000001110;
assign input_1551 = t6_000001111;
assign input_1552 = t6_000010000;
assign input_1553 = t6_000010001;
assign input_1554 = t6_000010010;
assign input_1555 = t6_000010011;
assign input_1556 = t6_000010100;
assign input_1557 = t6_000010101;
assign input_1558 = t6_000010110;
assign input_1559 = t6_000010111;
assign input_1560 = t6_000011000;
assign input_1561 = t6_000011001;
assign input_1562 = t6_000011010;
assign input_1563 = t6_000011011;
assign input_1564 = t6_000011100;
assign input_1565 = t6_000011101;
assign input_1566 = t6_000011110;
assign input_1567 = t6_000011111;
assign input_1568 = t6_000100000;
assign input_1569 = t6_000100001;
assign input_1570 = t6_000100010;
assign input_1571 = t6_000100011;
assign input_1572 = t6_000100100;
assign input_1573 = t6_000100101;
assign input_1574 = t6_000100110;
assign input_1575 = t6_000100111;
assign input_1576 = t6_000101000;
assign input_1577 = t6_000101001;
assign input_1578 = t6_000101010;
assign input_1579 = t6_000101011;
assign input_1580 = t6_000101100;
assign input_1581 = t6_000101101;
assign input_1582 = t6_000101110;
assign input_1583 = t6_000101111;
assign input_1584 = t6_000110000;
assign input_1585 = t6_000110001;
assign input_1586 = t6_000110010;
assign input_1587 = t6_000110011;
assign input_1588 = t6_000110100;
assign input_1589 = t6_000110101;
assign input_1590 = t6_000110110;
assign input_1591 = t6_000110111;
assign input_1592 = t6_000111000;
assign input_1593 = t6_000111001;
assign input_1594 = t6_000111010;
assign input_1595 = t6_000111011;
assign input_1596 = t6_000111100;
assign input_1597 = t6_000111101;
assign input_1598 = t6_000111110;
assign input_1599 = t6_000111111;
assign input_1600 = t6_001000000;
assign input_1601 = t6_001000001;
assign input_1602 = t6_001000010;
assign input_1603 = t6_001000011;
assign input_1604 = t6_001000100;
assign input_1605 = t6_001000101;
assign input_1606 = t6_001000110;
assign input_1607 = t6_001000111;
assign input_1608 = t6_001001000;
assign input_1609 = t6_001001001;
assign input_1610 = t6_001001010;
assign input_1611 = t6_001001011;
assign input_1612 = t6_001001100;
assign input_1613 = t6_001001101;
assign input_1614 = t6_001001110;
assign input_1615 = t6_001001111;
assign input_1616 = t6_001010000;
assign input_1617 = t6_001010001;
assign input_1618 = t6_001010010;
assign input_1619 = t6_001010011;
assign input_1620 = t6_001010100;
assign input_1621 = t6_001010101;
assign input_1622 = t6_001010110;
assign input_1623 = t6_001010111;
assign input_1624 = t6_001011000;
assign input_1625 = t6_001011001;
assign input_1626 = t6_001011010;
assign input_1627 = t6_001011011;
assign input_1628 = t6_001011100;
assign input_1629 = t6_001011101;
assign input_1630 = t6_001011110;
assign input_1631 = t6_001011111;
assign input_1632 = t6_001100000;
assign input_1633 = t6_001100001;
assign input_1634 = t6_001100010;
assign input_1635 = t6_001100011;
assign input_1636 = t6_001100100;
assign input_1637 = t6_001100101;
assign input_1638 = t6_001100110;
assign input_1639 = t6_001100111;
assign input_1640 = t6_001101000;
assign input_1641 = t6_001101001;
assign input_1642 = t6_001101010;
assign input_1643 = t6_001101011;
assign input_1644 = t6_001101100;
assign input_1645 = t6_001101101;
assign input_1646 = t6_001101110;
assign input_1647 = t6_001101111;
assign input_1648 = t6_001110000;
assign input_1649 = t6_001110001;
assign input_1650 = t6_001110010;
assign input_1651 = t6_001110011;
assign input_1652 = t6_001110100;
assign input_1653 = t6_001110101;
assign input_1654 = t6_001110110;
assign input_1655 = t6_001110111;
assign input_1656 = t6_001111000;
assign input_1657 = t6_001111001;
assign input_1658 = t6_001111010;
assign input_1659 = t6_001111011;
assign input_1660 = t6_001111100;
assign input_1661 = t6_001111101;
assign input_1662 = t6_001111110;
assign input_1663 = t6_001111111;
assign input_1664 = t6_010000000;
assign input_1665 = t6_010000001;
assign input_1666 = t6_010000010;
assign input_1667 = t6_010000011;
assign input_1668 = t6_010000100;
assign input_1669 = t6_010000101;
assign input_1670 = t6_010000110;
assign input_1671 = t6_010000111;
assign input_1672 = t6_010001000;
assign input_1673 = t6_010001001;
assign input_1674 = t6_010001010;
assign input_1675 = t6_010001011;
assign input_1676 = t6_010001100;
assign input_1677 = t6_010001101;
assign input_1678 = t6_010001110;
assign input_1679 = t6_010001111;
assign input_1680 = t6_010010000;
assign input_1681 = t6_010010001;
assign input_1682 = t6_010010010;
assign input_1683 = t6_010010011;
assign input_1684 = t6_010010100;
assign input_1685 = t6_010010101;
assign input_1686 = t6_010010110;
assign input_1687 = t6_010010111;
assign input_1688 = t6_010011000;
assign input_1689 = t6_010011001;
assign input_1690 = t6_010011010;
assign input_1691 = t6_010011011;
assign input_1692 = t6_010011100;
assign input_1693 = t6_010011101;
assign input_1694 = t6_010011110;
assign input_1695 = t6_010011111;
assign input_1696 = t6_010100000;
assign input_1697 = t6_010100001;
assign input_1698 = t6_010100010;
assign input_1699 = t6_010100011;
assign input_1700 = t6_010100100;
assign input_1701 = t6_010100101;
assign input_1702 = t6_010100110;
assign input_1703 = t6_010100111;
assign input_1704 = t6_010101000;
assign input_1705 = t6_010101001;
assign input_1706 = t6_010101010;
assign input_1707 = t6_010101011;
assign input_1708 = t6_010101100;
assign input_1709 = t6_010101101;
assign input_1710 = t6_010101110;
assign input_1711 = t6_010101111;
assign input_1712 = t6_010110000;
assign input_1713 = t6_010110001;
assign input_1714 = t6_010110010;
assign input_1715 = t6_010110011;
assign input_1716 = t6_010110100;
assign input_1717 = t6_010110101;
assign input_1718 = t6_010110110;
assign input_1719 = t6_010110111;
assign input_1720 = t6_010111000;
assign input_1721 = t6_010111001;
assign input_1722 = t6_010111010;
assign input_1723 = t6_010111011;
assign input_1724 = t6_010111100;
assign input_1725 = t6_010111101;
assign input_1726 = t6_010111110;
assign input_1727 = t6_010111111;
assign input_1728 = t6_011000000;
assign input_1729 = t6_011000001;
assign input_1730 = t6_011000010;
assign input_1731 = t6_011000011;
assign input_1732 = t6_011000100;
assign input_1733 = t6_011000101;
assign input_1734 = t6_011000110;
assign input_1735 = t6_011000111;
assign input_1736 = t6_011001000;
assign input_1737 = t6_011001001;
assign input_1738 = t6_011001010;
assign input_1739 = t6_011001011;
assign input_1740 = t6_011001100;
assign input_1741 = t6_011001101;
assign input_1742 = t6_011001110;
assign input_1743 = t6_011001111;
assign input_1744 = t6_011010000;
assign input_1745 = t6_011010001;
assign input_1746 = t6_011010010;
assign input_1747 = t6_011010011;
assign input_1748 = t6_011010100;
assign input_1749 = t6_011010101;
assign input_1750 = t6_011010110;
assign input_1751 = t6_011010111;
assign input_1752 = t6_011011000;
assign input_1753 = t6_011011001;
assign input_1754 = t6_011011010;
assign input_1755 = t6_011011011;
assign input_1756 = t6_011011100;
assign input_1757 = t6_011011101;
assign input_1758 = t6_011011110;
assign input_1759 = t6_011011111;
assign input_1760 = t6_011100000;
assign input_1761 = t6_011100001;
assign input_1762 = t6_011100010;
assign input_1763 = t6_011100011;
assign input_1764 = t6_011100100;
assign input_1765 = t6_011100101;
assign input_1766 = t6_011100110;
assign input_1767 = t6_011100111;
assign input_1768 = t6_011101000;
assign input_1769 = t6_011101001;
assign input_1770 = t6_011101010;
assign input_1771 = t6_011101011;
assign input_1772 = t6_011101100;
assign input_1773 = t6_011101101;
assign input_1774 = t6_011101110;
assign input_1775 = t6_011101111;
assign input_1776 = t6_011110000;
assign input_1777 = t6_011110001;
assign input_1778 = t6_011110010;
assign input_1779 = t6_011110011;
assign input_1780 = t6_011110100;
assign input_1781 = t6_011110101;
assign input_1782 = t6_011110110;
assign input_1783 = t6_011110111;
assign input_1784 = t6_011111000;
assign input_1785 = t6_011111001;
assign input_1786 = t6_011111010;
assign input_1787 = t6_011111011;
assign input_1788 = t6_011111100;
assign input_1789 = t6_011111101;
assign input_1790 = t6_011111110;
assign input_1791 = t6_011111111;
assign input_1792 = t7_000000000;
assign input_1793 = t7_000000001;
assign input_1794 = t7_000000010;
assign input_1795 = t7_000000011;
assign input_1796 = t7_000000100;
assign input_1797 = t7_000000101;
assign input_1798 = t7_000000110;
assign input_1799 = t7_000000111;
assign input_1800 = t7_000001000;
assign input_1801 = t7_000001001;
assign input_1802 = t7_000001010;
assign input_1803 = t7_000001011;
assign input_1804 = t7_000001100;
assign input_1805 = t7_000001101;
assign input_1806 = t7_000001110;
assign input_1807 = t7_000001111;
assign input_1808 = t7_000010000;
assign input_1809 = t7_000010001;
assign input_1810 = t7_000010010;
assign input_1811 = t7_000010011;
assign input_1812 = t7_000010100;
assign input_1813 = t7_000010101;
assign input_1814 = t7_000010110;
assign input_1815 = t7_000010111;
assign input_1816 = t7_000011000;
assign input_1817 = t7_000011001;
assign input_1818 = t7_000011010;
assign input_1819 = t7_000011011;
assign input_1820 = t7_000011100;
assign input_1821 = t7_000011101;
assign input_1822 = t7_000011110;
assign input_1823 = t7_000011111;
assign input_1824 = t7_000100000;
assign input_1825 = t7_000100001;
assign input_1826 = t7_000100010;
assign input_1827 = t7_000100011;
assign input_1828 = t7_000100100;
assign input_1829 = t7_000100101;
assign input_1830 = t7_000100110;
assign input_1831 = t7_000100111;
assign input_1832 = t7_000101000;
assign input_1833 = t7_000101001;
assign input_1834 = t7_000101010;
assign input_1835 = t7_000101011;
assign input_1836 = t7_000101100;
assign input_1837 = t7_000101101;
assign input_1838 = t7_000101110;
assign input_1839 = t7_000101111;
assign input_1840 = t7_000110000;
assign input_1841 = t7_000110001;
assign input_1842 = t7_000110010;
assign input_1843 = t7_000110011;
assign input_1844 = t7_000110100;
assign input_1845 = t7_000110101;
assign input_1846 = t7_000110110;
assign input_1847 = t7_000110111;
assign input_1848 = t7_000111000;
assign input_1849 = t7_000111001;
assign input_1850 = t7_000111010;
assign input_1851 = t7_000111011;
assign input_1852 = t7_000111100;
assign input_1853 = t7_000111101;
assign input_1854 = t7_000111110;
assign input_1855 = t7_000111111;
assign input_1856 = t7_001000000;
assign input_1857 = t7_001000001;
assign input_1858 = t7_001000010;
assign input_1859 = t7_001000011;
assign input_1860 = t7_001000100;
assign input_1861 = t7_001000101;
assign input_1862 = t7_001000110;
assign input_1863 = t7_001000111;
assign input_1864 = t7_001001000;
assign input_1865 = t7_001001001;
assign input_1866 = t7_001001010;
assign input_1867 = t7_001001011;
assign input_1868 = t7_001001100;
assign input_1869 = t7_001001101;
assign input_1870 = t7_001001110;
assign input_1871 = t7_001001111;
assign input_1872 = t7_001010000;
assign input_1873 = t7_001010001;
assign input_1874 = t7_001010010;
assign input_1875 = t7_001010011;
assign input_1876 = t7_001010100;
assign input_1877 = t7_001010101;
assign input_1878 = t7_001010110;
assign input_1879 = t7_001010111;
assign input_1880 = t7_001011000;
assign input_1881 = t7_001011001;
assign input_1882 = t7_001011010;
assign input_1883 = t7_001011011;
assign input_1884 = t7_001011100;
assign input_1885 = t7_001011101;
assign input_1886 = t7_001011110;
assign input_1887 = t7_001011111;
assign input_1888 = t7_001100000;
assign input_1889 = t7_001100001;
assign input_1890 = t7_001100010;
assign input_1891 = t7_001100011;
assign input_1892 = t7_001100100;
assign input_1893 = t7_001100101;
assign input_1894 = t7_001100110;
assign input_1895 = t7_001100111;
assign input_1896 = t7_001101000;
assign input_1897 = t7_001101001;
assign input_1898 = t7_001101010;
assign input_1899 = t7_001101011;
assign input_1900 = t7_001101100;
assign input_1901 = t7_001101101;
assign input_1902 = t7_001101110;
assign input_1903 = t7_001101111;
assign input_1904 = t7_001110000;
assign input_1905 = t7_001110001;
assign input_1906 = t7_001110010;
assign input_1907 = t7_001110011;
assign input_1908 = t7_001110100;
assign input_1909 = t7_001110101;
assign input_1910 = t7_001110110;
assign input_1911 = t7_001110111;
assign input_1912 = t7_001111000;
assign input_1913 = t7_001111001;
assign input_1914 = t7_001111010;
assign input_1915 = t7_001111011;
assign input_1916 = t7_001111100;
assign input_1917 = t7_001111101;
assign input_1918 = t7_001111110;
assign input_1919 = t7_001111111;
assign input_1920 = t7_010000000;
assign input_1921 = t7_010000001;
assign input_1922 = t7_010000010;
assign input_1923 = t7_010000011;
assign input_1924 = t7_010000100;
assign input_1925 = t7_010000101;
assign input_1926 = t7_010000110;
assign input_1927 = t7_010000111;
assign input_1928 = t7_010001000;
assign input_1929 = t7_010001001;
assign input_1930 = t7_010001010;
assign input_1931 = t7_010001011;
assign input_1932 = t7_010001100;
assign input_1933 = t7_010001101;
assign input_1934 = t7_010001110;
assign input_1935 = t7_010001111;
assign input_1936 = t7_010010000;
assign input_1937 = t7_010010001;
assign input_1938 = t7_010010010;
assign input_1939 = t7_010010011;
assign input_1940 = t7_010010100;
assign input_1941 = t7_010010101;
assign input_1942 = t7_010010110;
assign input_1943 = t7_010010111;
assign input_1944 = t7_010011000;
assign input_1945 = t7_010011001;
assign input_1946 = t7_010011010;
assign input_1947 = t7_010011011;
assign input_1948 = t7_010011100;
assign input_1949 = t7_010011101;
assign input_1950 = t7_010011110;
assign input_1951 = t7_010011111;
assign input_1952 = t7_010100000;
assign input_1953 = t7_010100001;
assign input_1954 = t7_010100010;
assign input_1955 = t7_010100011;
assign input_1956 = t7_010100100;
assign input_1957 = t7_010100101;
assign input_1958 = t7_010100110;
assign input_1959 = t7_010100111;
assign input_1960 = t7_010101000;
assign input_1961 = t7_010101001;
assign input_1962 = t7_010101010;
assign input_1963 = t7_010101011;
assign input_1964 = t7_010101100;
assign input_1965 = t7_010101101;
assign input_1966 = t7_010101110;
assign input_1967 = t7_010101111;
assign input_1968 = t7_010110000;
assign input_1969 = t7_010110001;
assign input_1970 = t7_010110010;
assign input_1971 = t7_010110011;
assign input_1972 = t7_010110100;
assign input_1973 = t7_010110101;
assign input_1974 = t7_010110110;
assign input_1975 = t7_010110111;
assign input_1976 = t7_010111000;
assign input_1977 = t7_010111001;
assign input_1978 = t7_010111010;
assign input_1979 = t7_010111011;
assign input_1980 = t7_010111100;
assign input_1981 = t7_010111101;
assign input_1982 = t7_010111110;
assign input_1983 = t7_010111111;
assign input_1984 = t7_011000000;
assign input_1985 = t7_011000001;
assign input_1986 = t7_011000010;
assign input_1987 = t7_011000011;
assign input_1988 = t7_011000100;
assign input_1989 = t7_011000101;
assign input_1990 = t7_011000110;
assign input_1991 = t7_011000111;
assign input_1992 = t7_011001000;
assign input_1993 = t7_011001001;
assign input_1994 = t7_011001010;
assign input_1995 = t7_011001011;
assign input_1996 = t7_011001100;
assign input_1997 = t7_011001101;
assign input_1998 = t7_011001110;
assign input_1999 = t7_011001111;
assign input_2000 = t7_011010000;
assign input_2001 = t7_011010001;
assign input_2002 = t7_011010010;
assign input_2003 = t7_011010011;
assign input_2004 = t7_011010100;
assign input_2005 = t7_011010101;
assign input_2006 = t7_011010110;
assign input_2007 = t7_011010111;
assign input_2008 = t7_011011000;
assign input_2009 = t7_011011001;
assign input_2010 = t7_011011010;
assign input_2011 = t7_011011011;
assign input_2012 = t7_011011100;
assign input_2013 = t7_011011101;
assign input_2014 = t7_011011110;
assign input_2015 = t7_011011111;
assign input_2016 = t7_011100000;
assign input_2017 = t7_011100001;
assign input_2018 = t7_011100010;
assign input_2019 = t7_011100011;
assign input_2020 = t7_011100100;
assign input_2021 = t7_011100101;
assign input_2022 = t7_011100110;
assign input_2023 = t7_011100111;
assign input_2024 = t7_011101000;
assign input_2025 = t7_011101001;
assign input_2026 = t7_011101010;
assign input_2027 = t7_011101011;
assign input_2028 = t7_011101100;
assign input_2029 = t7_011101101;
assign input_2030 = t7_011101110;
assign input_2031 = t7_011101111;
assign input_2032 = t7_011110000;
assign input_2033 = t7_011110001;
assign input_2034 = t7_011110010;
assign input_2035 = t7_011110011;
assign input_2036 = t7_011110100;
assign input_2037 = t7_011110101;
assign input_2038 = t7_011110110;
assign input_2039 = t7_011110111;
assign input_2040 = t7_011111000;
assign input_2041 = t7_011111001;
assign input_2042 = t7_011111010;
assign input_2043 = t7_011111011;
assign input_2044 = t7_011111100;
assign input_2045 = t7_011111101;
assign input_2046 = t7_011111110;
assign input_2047 = t7_011111111;
endmodule
