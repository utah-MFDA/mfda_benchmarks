module Planar_Synthetic_5(
input Source1,
input Source2,
output Out1
);
wire flow_switch4_1-Source1;
wire flow_switch4_1-Mixer1;
wire flow_switch4_1-Mixer2;
wire flow_switch4_2-flow_switch4_1;
wire flow_switch4_2-Mixer3;
wire flow_switch4_2-Mixer4;
wire flow_switch4_3-flow_switch4_2;
wire flow_switch4_3-Mixer5;
wire flow_switch4_3-Mixer6;
wire flow_switch4_4-flow_switch4_3;
wire flow_switch4_4-Mixer7;
wire flow_switch4_4-Mixer8;
wire flow_switch4_5-flow_switch4_4;
wire flow_switch4_5-Heater1;
wire flow_switch4_5-Heater2;
wire flow_switch4_6-flow_switch4_5;
wire flow_switch4_6-Filter1;
wire flow_switch4_6-Filter2;
wire flow_switch4_7-Source2;
wire flow_switch4_7-Mixer9;
wire flow_switch4_7-Mixer10;
wire flow_switch4_8-flow_switch4_7;
wire flow_switch4_8-Mixer11;
wire flow_switch4_8-Mixer12;
wire flow_switch4_9-flow_switch4_8;
wire flow_switch4_9-Mixer13;
wire flow_switch4_9-Mixer14;
wire flow_switch4_10-flow_switch4_9;
wire flow_switch4_10-Mixer15;
wire flow_switch4_10-Mixer16;
wire flow_switch4_11-flow_switch4_10;
wire flow_switch4_11-Heater3;
wire flow_switch4_11-Heater4;
wire flow_switch4_12-flow_switch4_11;
wire flow_switch4_12-Filter3;
wire flow_switch4_12-Filter4;
wire Heater5-flow_switch4_6;
wire Heater6-flow_switch4_12;
wire Filter5-Heater5;
wire Filter6-Heater6;
wire flow_switch3_1-Filter5;
wire flow_switch3_1-Filter6;
wire Mixer17-flow_switch3_1;
wire Filter7-Mixer17;
wire Out1-Filter7;
assign flow_switch4_1-Source1 = Source1;
assign flow_switch4_7-Source2 = Source2;
Mixer Mixer1(.port0(flow_switch4_1-Mixer1),.port1(None));
Mixer Mixer2(.port0(None),.port1(flow_switch4_1-Mixer2));
Mixer Mixer3(.port0(None),.port1(flow_switch4_2-Mixer3));
Mixer Mixer4(.port0(None),.port1(flow_switch4_2-Mixer4));
Mixer Mixer5(.port0(None),.port1(flow_switch4_3-Mixer5));
Mixer Mixer6(.port0(None),.port1(flow_switch4_3-Mixer6));
Mixer Mixer7(.port0(None),.port1(flow_switch4_4-Mixer7));
Mixer Mixer8(.port0(None),.port1(flow_switch4_4-Mixer8));
Mixer Mixer9(.port0(flow_switch4_7-Mixer9),.port1(None));
Mixer Mixer10(.port0(None),.port1(flow_switch4_7-Mixer10));
Mixer Mixer11(.port0(None),.port1(flow_switch4_8-Mixer11));
Mixer Mixer12(.port0(None),.port1(flow_switch4_8-Mixer12));
Mixer Mixer13(.port0(None),.port1(flow_switch4_9-Mixer13));
Mixer Mixer14(.port0(None),.port1(flow_switch4_9-Mixer14));
Mixer Mixer15(.port0(None),.port1(flow_switch4_10-Mixer15));
Mixer Mixer16(.port0(None),.port1(flow_switch4_10-Mixer16));
Mixer Mixer17(.port0(Filter7-Mixer17),.port1(Mixer17-flow_switch3_1));
Heater Heater1(.port0(flow_switch4_5-Heater1),.port1(None));
Heater Heater2(.port0(flow_switch4_5-Heater2),.port1(None));
Heater Heater3(.port0(flow_switch4_11-Heater3),.port1(None));
Heater Heater4(.port0(flow_switch4_11-Heater4),.port1(None));
Heater Heater5(.port0(Filter5-Heater5),.port1(Heater5-flow_switch4_6));
Heater Heater6(.port0(Heater6-flow_switch4_12),.port1(Filter6-Heater6));
Filter Filter1(.port0(flow_switch4_6-Filter1),.port1(None));
Filter Filter2(.port0(flow_switch4_6-Filter2),.port1(None));
Filter Filter3(.port0(flow_switch4_12-Filter3),.port1(None));
Filter Filter4(.port0(flow_switch4_12-Filter4),.port1(None));
Filter Filter5(.port0(flow_switch3_1-Filter5),.port1(Filter5-Heater5));
Filter Filter6(.port0(flow_switch3_1-Filter6),.port1(Filter6-Heater6));
Filter Filter7(.port0(Filter7-Mixer17),.port1(Out1-Filter7));
assign Out1 = Out1-Filter7;
Switch flow_switch4_1(.port0(flow_switch4_2-flow_switch4_1),.port1(flow_switch4_1-Source1),.port2(flow_switch4_1-Mixer1),.port3(flow_switch4_1-Mixer2));
Switch flow_switch4_2(.port0(flow_switch4_2-Mixer4),.port1(flow_switch4_3-flow_switch4_2),.port2(flow_switch4_2-flow_switch4_1),.port3(flow_switch4_2-Mixer3));
Switch flow_switch4_3(.port0(flow_switch4_3-Mixer6),.port1(flow_switch4_3-flow_switch4_2),.port2(flow_switch4_4-flow_switch4_3),.port3(flow_switch4_3-Mixer5));
Switch flow_switch4_4(.port0(flow_switch4_4-Mixer8),.port1(flow_switch4_5-flow_switch4_4),.port2(flow_switch4_4-flow_switch4_3),.port3(flow_switch4_4-Mixer7));
Switch flow_switch4_5(.port0(flow_switch4_5-Heater2),.port1(flow_switch4_5-flow_switch4_4),.port2(flow_switch4_6-flow_switch4_5),.port3(flow_switch4_5-Heater1));
Switch flow_switch4_6(.port0(flow_switch4_6-Filter2),.port1(flow_switch4_6-flow_switch4_5),.port2(Heater5-flow_switch4_6),.port3(flow_switch4_6-Filter1));
Switch flow_switch4_7(.port0(flow_switch4_7-Source2),.port1(flow_switch4_8-flow_switch4_7),.port2(flow_switch4_7-Mixer9),.port3(flow_switch4_7-Mixer10));
Switch flow_switch4_8(.port0(flow_switch4_8-Mixer12),.port1(flow_switch4_9-flow_switch4_8),.port2(flow_switch4_8-flow_switch4_7),.port3(flow_switch4_8-Mixer11));
Switch flow_switch4_9(.port0(flow_switch4_9-Mixer14),.port1(flow_switch4_9-flow_switch4_8),.port2(flow_switch4_10-flow_switch4_9),.port3(flow_switch4_9-Mixer13));
Switch flow_switch4_10(.port0(flow_switch4_10-Mixer16),.port1(flow_switch4_10-flow_switch4_9),.port2(flow_switch4_11-flow_switch4_10),.port3(flow_switch4_10-Mixer15));
Switch flow_switch4_11(.port0(flow_switch4_11-Heater4),.port1(flow_switch4_11-flow_switch4_10),.port2(flow_switch4_12-flow_switch4_11),.port3(flow_switch4_11-Heater3));
Switch flow_switch4_12(.port0(flow_switch4_12-Filter3),.port1(Heater6-flow_switch4_12),.port2(flow_switch4_12-Filter4),.port3(flow_switch4_12-flow_switch4_11));
Switch flow_switch3_1(.port0(None),.port1(Mixer17-flow_switch3_1),.port2(flow_switch3_1-Filter6),.port3(flow_switch3_1-Filter5));
endmodule
