module chain_mixer_32 (
output j32,input j0,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32,input k32
);
mixer m0(.a(in), .b(k0), .y(j1));
wire j1;
wire j2;
wire j3;
wire j4;
wire j5;
wire j6;
wire j7;
wire j8;
wire j9;
wire j10;
wire j11;
wire j12;
wire j13;
wire j14;
wire j15;
wire j16;
wire j17;
wire j18;
wire j19;
wire j20;
wire j21;
wire j22;
wire j23;
wire j24;
wire j25;
wire j26;
wire j27;
wire j28;
wire j29;
wire j30;
wire j31;
mixer m0(.a(j0), .b(k0), .y(j1));
mixer m1(.a(j1), .b(k1), .y(j2));
mixer m2(.a(j2), .b(k2), .y(j3));
mixer m3(.a(j3), .b(k3), .y(j4));
mixer m4(.a(j4), .b(k4), .y(j5));
mixer m5(.a(j5), .b(k5), .y(j6));
mixer m6(.a(j6), .b(k6), .y(j7));
mixer m7(.a(j7), .b(k7), .y(j8));
mixer m8(.a(j8), .b(k8), .y(j9));
mixer m9(.a(j9), .b(k9), .y(j10));
mixer m10(.a(j10), .b(k10), .y(j11));
mixer m11(.a(j11), .b(k11), .y(j12));
mixer m12(.a(j12), .b(k12), .y(j13));
mixer m13(.a(j13), .b(k13), .y(j14));
mixer m14(.a(j14), .b(k14), .y(j15));
mixer m15(.a(j15), .b(k15), .y(j16));
mixer m16(.a(j16), .b(k16), .y(j17));
mixer m17(.a(j17), .b(k17), .y(j18));
mixer m18(.a(j18), .b(k18), .y(j19));
mixer m19(.a(j19), .b(k19), .y(j20));
mixer m20(.a(j20), .b(k20), .y(j21));
mixer m21(.a(j21), .b(k21), .y(j22));
mixer m22(.a(j22), .b(k22), .y(j23));
mixer m23(.a(j23), .b(k23), .y(j24));
mixer m24(.a(j24), .b(k24), .y(j25));
mixer m25(.a(j25), .b(k25), .y(j26));
mixer m26(.a(j26), .b(k26), .y(j27));
mixer m27(.a(j27), .b(k27), .y(j28));
mixer m28(.a(j28), .b(k28), .y(j29));
mixer m29(.a(j29), .b(k29), .y(j30));
mixer m30(.a(j30), .b(k30), .y(j31));
mixer m31(.a(j31), .b(k31), .y(j32));
endmodule
