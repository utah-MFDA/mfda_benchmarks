module chain_128 (
inout k0, k128
);
wire {wires};
chamber ch0 (.in(k0), .out(k1)
chamber ch1 (.in(k1), .out(k2)
chamber ch2 (.in(k2), .out(k3)
chamber ch3 (.in(k3), .out(k4)
chamber ch4 (.in(k4), .out(k5)
chamber ch5 (.in(k5), .out(k6)
chamber ch6 (.in(k6), .out(k7)
chamber ch7 (.in(k7), .out(k8)
chamber ch8 (.in(k8), .out(k9)
chamber ch9 (.in(k9), .out(k10)
chamber ch10 (.in(k10), .out(k11)
chamber ch11 (.in(k11), .out(k12)
chamber ch12 (.in(k12), .out(k13)
chamber ch13 (.in(k13), .out(k14)
chamber ch14 (.in(k14), .out(k15)
chamber ch15 (.in(k15), .out(k16)
chamber ch16 (.in(k16), .out(k17)
chamber ch17 (.in(k17), .out(k18)
chamber ch18 (.in(k18), .out(k19)
chamber ch19 (.in(k19), .out(k20)
chamber ch20 (.in(k20), .out(k21)
chamber ch21 (.in(k21), .out(k22)
chamber ch22 (.in(k22), .out(k23)
chamber ch23 (.in(k23), .out(k24)
chamber ch24 (.in(k24), .out(k25)
chamber ch25 (.in(k25), .out(k26)
chamber ch26 (.in(k26), .out(k27)
chamber ch27 (.in(k27), .out(k28)
chamber ch28 (.in(k28), .out(k29)
chamber ch29 (.in(k29), .out(k30)
chamber ch30 (.in(k30), .out(k31)
chamber ch31 (.in(k31), .out(k32)
chamber ch32 (.in(k32), .out(k33)
chamber ch33 (.in(k33), .out(k34)
chamber ch34 (.in(k34), .out(k35)
chamber ch35 (.in(k35), .out(k36)
chamber ch36 (.in(k36), .out(k37)
chamber ch37 (.in(k37), .out(k38)
chamber ch38 (.in(k38), .out(k39)
chamber ch39 (.in(k39), .out(k40)
chamber ch40 (.in(k40), .out(k41)
chamber ch41 (.in(k41), .out(k42)
chamber ch42 (.in(k42), .out(k43)
chamber ch43 (.in(k43), .out(k44)
chamber ch44 (.in(k44), .out(k45)
chamber ch45 (.in(k45), .out(k46)
chamber ch46 (.in(k46), .out(k47)
chamber ch47 (.in(k47), .out(k48)
chamber ch48 (.in(k48), .out(k49)
chamber ch49 (.in(k49), .out(k50)
chamber ch50 (.in(k50), .out(k51)
chamber ch51 (.in(k51), .out(k52)
chamber ch52 (.in(k52), .out(k53)
chamber ch53 (.in(k53), .out(k54)
chamber ch54 (.in(k54), .out(k55)
chamber ch55 (.in(k55), .out(k56)
chamber ch56 (.in(k56), .out(k57)
chamber ch57 (.in(k57), .out(k58)
chamber ch58 (.in(k58), .out(k59)
chamber ch59 (.in(k59), .out(k60)
chamber ch60 (.in(k60), .out(k61)
chamber ch61 (.in(k61), .out(k62)
chamber ch62 (.in(k62), .out(k63)
chamber ch63 (.in(k63), .out(k64)
chamber ch64 (.in(k64), .out(k65)
chamber ch65 (.in(k65), .out(k66)
chamber ch66 (.in(k66), .out(k67)
chamber ch67 (.in(k67), .out(k68)
chamber ch68 (.in(k68), .out(k69)
chamber ch69 (.in(k69), .out(k70)
chamber ch70 (.in(k70), .out(k71)
chamber ch71 (.in(k71), .out(k72)
chamber ch72 (.in(k72), .out(k73)
chamber ch73 (.in(k73), .out(k74)
chamber ch74 (.in(k74), .out(k75)
chamber ch75 (.in(k75), .out(k76)
chamber ch76 (.in(k76), .out(k77)
chamber ch77 (.in(k77), .out(k78)
chamber ch78 (.in(k78), .out(k79)
chamber ch79 (.in(k79), .out(k80)
chamber ch80 (.in(k80), .out(k81)
chamber ch81 (.in(k81), .out(k82)
chamber ch82 (.in(k82), .out(k83)
chamber ch83 (.in(k83), .out(k84)
chamber ch84 (.in(k84), .out(k85)
chamber ch85 (.in(k85), .out(k86)
chamber ch86 (.in(k86), .out(k87)
chamber ch87 (.in(k87), .out(k88)
chamber ch88 (.in(k88), .out(k89)
chamber ch89 (.in(k89), .out(k90)
chamber ch90 (.in(k90), .out(k91)
chamber ch91 (.in(k91), .out(k92)
chamber ch92 (.in(k92), .out(k93)
chamber ch93 (.in(k93), .out(k94)
chamber ch94 (.in(k94), .out(k95)
chamber ch95 (.in(k95), .out(k96)
chamber ch96 (.in(k96), .out(k97)
chamber ch97 (.in(k97), .out(k98)
chamber ch98 (.in(k98), .out(k99)
chamber ch99 (.in(k99), .out(k100)
chamber ch100 (.in(k100), .out(k101)
chamber ch101 (.in(k101), .out(k102)
chamber ch102 (.in(k102), .out(k103)
chamber ch103 (.in(k103), .out(k104)
chamber ch104 (.in(k104), .out(k105)
chamber ch105 (.in(k105), .out(k106)
chamber ch106 (.in(k106), .out(k107)
chamber ch107 (.in(k107), .out(k108)
chamber ch108 (.in(k108), .out(k109)
chamber ch109 (.in(k109), .out(k110)
chamber ch110 (.in(k110), .out(k111)
chamber ch111 (.in(k111), .out(k112)
chamber ch112 (.in(k112), .out(k113)
chamber ch113 (.in(k113), .out(k114)
chamber ch114 (.in(k114), .out(k115)
chamber ch115 (.in(k115), .out(k116)
chamber ch116 (.in(k116), .out(k117)
chamber ch117 (.in(k117), .out(k118)
chamber ch118 (.in(k118), .out(k119)
chamber ch119 (.in(k119), .out(k120)
chamber ch120 (.in(k120), .out(k121)
chamber ch121 (.in(k121), .out(k122)
chamber ch122 (.in(k122), .out(k123)
chamber ch123 (.in(k123), .out(k124)
chamber ch124 (.in(k124), .out(k125)
chamber ch125 (.in(k125), .out(k126)
chamber ch126 (.in(k126), .out(k127)
chamber ch127 (.in(k127), .out(k128)
endmodule
