module fanout2_braid_16_32 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,output output_8,output output_9,output output_10,output output_11,output output_12,output output_13,output output_14,output output_15,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_9_0, output_9_1, output_8_0;
mixer gate_output_8_0(.a(output_9_0), .b(output_9_1), .y(output_8_0));
wire output_10_0, output_10_1, output_9_0;
mixer gate_output_9_0(.a(output_10_0), .b(output_10_1), .y(output_9_0));
wire output_11_0, output_11_1, output_10_0;
mixer gate_output_10_0(.a(output_11_0), .b(output_11_1), .y(output_10_0));
wire output_12_0, output_12_1, output_11_0;
mixer gate_output_11_0(.a(output_12_0), .b(output_12_1), .y(output_11_0));
wire output_13_0, output_13_1, output_12_0;
mixer gate_output_12_0(.a(output_13_0), .b(output_13_1), .y(output_12_0));
wire output_14_0, output_14_1, output_13_0;
mixer gate_output_13_0(.a(output_14_0), .b(output_14_1), .y(output_13_0));
wire output_15_0, output_15_1, output_14_0;
mixer gate_output_14_0(.a(output_15_0), .b(output_15_1), .y(output_14_0));
wire output_16_0, output_16_1, output_15_0;
mixer gate_output_15_0(.a(output_16_0), .b(output_16_1), .y(output_15_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_9_1, output_9_2, output_8_1;
mixer gate_output_8_1(.a(output_9_1), .b(output_9_2), .y(output_8_1));
wire output_10_1, output_10_2, output_9_1;
mixer gate_output_9_1(.a(output_10_1), .b(output_10_2), .y(output_9_1));
wire output_11_1, output_11_2, output_10_1;
mixer gate_output_10_1(.a(output_11_1), .b(output_11_2), .y(output_10_1));
wire output_12_1, output_12_2, output_11_1;
mixer gate_output_11_1(.a(output_12_1), .b(output_12_2), .y(output_11_1));
wire output_13_1, output_13_2, output_12_1;
mixer gate_output_12_1(.a(output_13_1), .b(output_13_2), .y(output_12_1));
wire output_14_1, output_14_2, output_13_1;
mixer gate_output_13_1(.a(output_14_1), .b(output_14_2), .y(output_13_1));
wire output_15_1, output_15_2, output_14_1;
mixer gate_output_14_1(.a(output_15_1), .b(output_15_2), .y(output_14_1));
wire output_16_1, output_16_2, output_15_1;
mixer gate_output_15_1(.a(output_16_1), .b(output_16_2), .y(output_15_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_9_2, output_9_3, output_8_2;
mixer gate_output_8_2(.a(output_9_2), .b(output_9_3), .y(output_8_2));
wire output_10_2, output_10_3, output_9_2;
mixer gate_output_9_2(.a(output_10_2), .b(output_10_3), .y(output_9_2));
wire output_11_2, output_11_3, output_10_2;
mixer gate_output_10_2(.a(output_11_2), .b(output_11_3), .y(output_10_2));
wire output_12_2, output_12_3, output_11_2;
mixer gate_output_11_2(.a(output_12_2), .b(output_12_3), .y(output_11_2));
wire output_13_2, output_13_3, output_12_2;
mixer gate_output_12_2(.a(output_13_2), .b(output_13_3), .y(output_12_2));
wire output_14_2, output_14_3, output_13_2;
mixer gate_output_13_2(.a(output_14_2), .b(output_14_3), .y(output_13_2));
wire output_15_2, output_15_3, output_14_2;
mixer gate_output_14_2(.a(output_15_2), .b(output_15_3), .y(output_14_2));
wire output_16_2, output_16_3, output_15_2;
mixer gate_output_15_2(.a(output_16_2), .b(output_16_3), .y(output_15_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_9_3, output_9_4, output_8_3;
mixer gate_output_8_3(.a(output_9_3), .b(output_9_4), .y(output_8_3));
wire output_10_3, output_10_4, output_9_3;
mixer gate_output_9_3(.a(output_10_3), .b(output_10_4), .y(output_9_3));
wire output_11_3, output_11_4, output_10_3;
mixer gate_output_10_3(.a(output_11_3), .b(output_11_4), .y(output_10_3));
wire output_12_3, output_12_4, output_11_3;
mixer gate_output_11_3(.a(output_12_3), .b(output_12_4), .y(output_11_3));
wire output_13_3, output_13_4, output_12_3;
mixer gate_output_12_3(.a(output_13_3), .b(output_13_4), .y(output_12_3));
wire output_14_3, output_14_4, output_13_3;
mixer gate_output_13_3(.a(output_14_3), .b(output_14_4), .y(output_13_3));
wire output_15_3, output_15_4, output_14_3;
mixer gate_output_14_3(.a(output_15_3), .b(output_15_4), .y(output_14_3));
wire output_16_3, output_16_4, output_15_3;
mixer gate_output_15_3(.a(output_16_3), .b(output_16_4), .y(output_15_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_9_4, output_9_5, output_8_4;
mixer gate_output_8_4(.a(output_9_4), .b(output_9_5), .y(output_8_4));
wire output_10_4, output_10_5, output_9_4;
mixer gate_output_9_4(.a(output_10_4), .b(output_10_5), .y(output_9_4));
wire output_11_4, output_11_5, output_10_4;
mixer gate_output_10_4(.a(output_11_4), .b(output_11_5), .y(output_10_4));
wire output_12_4, output_12_5, output_11_4;
mixer gate_output_11_4(.a(output_12_4), .b(output_12_5), .y(output_11_4));
wire output_13_4, output_13_5, output_12_4;
mixer gate_output_12_4(.a(output_13_4), .b(output_13_5), .y(output_12_4));
wire output_14_4, output_14_5, output_13_4;
mixer gate_output_13_4(.a(output_14_4), .b(output_14_5), .y(output_13_4));
wire output_15_4, output_15_5, output_14_4;
mixer gate_output_14_4(.a(output_15_4), .b(output_15_5), .y(output_14_4));
wire output_16_4, output_16_5, output_15_4;
mixer gate_output_15_4(.a(output_16_4), .b(output_16_5), .y(output_15_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_9_5, output_9_6, output_8_5;
mixer gate_output_8_5(.a(output_9_5), .b(output_9_6), .y(output_8_5));
wire output_10_5, output_10_6, output_9_5;
mixer gate_output_9_5(.a(output_10_5), .b(output_10_6), .y(output_9_5));
wire output_11_5, output_11_6, output_10_5;
mixer gate_output_10_5(.a(output_11_5), .b(output_11_6), .y(output_10_5));
wire output_12_5, output_12_6, output_11_5;
mixer gate_output_11_5(.a(output_12_5), .b(output_12_6), .y(output_11_5));
wire output_13_5, output_13_6, output_12_5;
mixer gate_output_12_5(.a(output_13_5), .b(output_13_6), .y(output_12_5));
wire output_14_5, output_14_6, output_13_5;
mixer gate_output_13_5(.a(output_14_5), .b(output_14_6), .y(output_13_5));
wire output_15_5, output_15_6, output_14_5;
mixer gate_output_14_5(.a(output_15_5), .b(output_15_6), .y(output_14_5));
wire output_16_5, output_16_6, output_15_5;
mixer gate_output_15_5(.a(output_16_5), .b(output_16_6), .y(output_15_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_9_6, output_9_7, output_8_6;
mixer gate_output_8_6(.a(output_9_6), .b(output_9_7), .y(output_8_6));
wire output_10_6, output_10_7, output_9_6;
mixer gate_output_9_6(.a(output_10_6), .b(output_10_7), .y(output_9_6));
wire output_11_6, output_11_7, output_10_6;
mixer gate_output_10_6(.a(output_11_6), .b(output_11_7), .y(output_10_6));
wire output_12_6, output_12_7, output_11_6;
mixer gate_output_11_6(.a(output_12_6), .b(output_12_7), .y(output_11_6));
wire output_13_6, output_13_7, output_12_6;
mixer gate_output_12_6(.a(output_13_6), .b(output_13_7), .y(output_12_6));
wire output_14_6, output_14_7, output_13_6;
mixer gate_output_13_6(.a(output_14_6), .b(output_14_7), .y(output_13_6));
wire output_15_6, output_15_7, output_14_6;
mixer gate_output_14_6(.a(output_15_6), .b(output_15_7), .y(output_14_6));
wire output_16_6, output_16_7, output_15_6;
mixer gate_output_15_6(.a(output_16_6), .b(output_16_7), .y(output_15_6));
wire output_1_7, output_1_8, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_8), .y(output_0_7));
wire output_2_7, output_2_8, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_8), .y(output_1_7));
wire output_3_7, output_3_8, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_8), .y(output_2_7));
wire output_4_7, output_4_8, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_8), .y(output_3_7));
wire output_5_7, output_5_8, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_8), .y(output_4_7));
wire output_6_7, output_6_8, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_8), .y(output_5_7));
wire output_7_7, output_7_8, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_8), .y(output_6_7));
wire output_8_7, output_8_8, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_8), .y(output_7_7));
wire output_9_7, output_9_8, output_8_7;
mixer gate_output_8_7(.a(output_9_7), .b(output_9_8), .y(output_8_7));
wire output_10_7, output_10_8, output_9_7;
mixer gate_output_9_7(.a(output_10_7), .b(output_10_8), .y(output_9_7));
wire output_11_7, output_11_8, output_10_7;
mixer gate_output_10_7(.a(output_11_7), .b(output_11_8), .y(output_10_7));
wire output_12_7, output_12_8, output_11_7;
mixer gate_output_11_7(.a(output_12_7), .b(output_12_8), .y(output_11_7));
wire output_13_7, output_13_8, output_12_7;
mixer gate_output_12_7(.a(output_13_7), .b(output_13_8), .y(output_12_7));
wire output_14_7, output_14_8, output_13_7;
mixer gate_output_13_7(.a(output_14_7), .b(output_14_8), .y(output_13_7));
wire output_15_7, output_15_8, output_14_7;
mixer gate_output_14_7(.a(output_15_7), .b(output_15_8), .y(output_14_7));
wire output_16_7, output_16_8, output_15_7;
mixer gate_output_15_7(.a(output_16_7), .b(output_16_8), .y(output_15_7));
wire output_1_8, output_1_9, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_9), .y(output_0_8));
wire output_2_8, output_2_9, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_9), .y(output_1_8));
wire output_3_8, output_3_9, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_9), .y(output_2_8));
wire output_4_8, output_4_9, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_9), .y(output_3_8));
wire output_5_8, output_5_9, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_9), .y(output_4_8));
wire output_6_8, output_6_9, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_9), .y(output_5_8));
wire output_7_8, output_7_9, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_9), .y(output_6_8));
wire output_8_8, output_8_9, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_9), .y(output_7_8));
wire output_9_8, output_9_9, output_8_8;
mixer gate_output_8_8(.a(output_9_8), .b(output_9_9), .y(output_8_8));
wire output_10_8, output_10_9, output_9_8;
mixer gate_output_9_8(.a(output_10_8), .b(output_10_9), .y(output_9_8));
wire output_11_8, output_11_9, output_10_8;
mixer gate_output_10_8(.a(output_11_8), .b(output_11_9), .y(output_10_8));
wire output_12_8, output_12_9, output_11_8;
mixer gate_output_11_8(.a(output_12_8), .b(output_12_9), .y(output_11_8));
wire output_13_8, output_13_9, output_12_8;
mixer gate_output_12_8(.a(output_13_8), .b(output_13_9), .y(output_12_8));
wire output_14_8, output_14_9, output_13_8;
mixer gate_output_13_8(.a(output_14_8), .b(output_14_9), .y(output_13_8));
wire output_15_8, output_15_9, output_14_8;
mixer gate_output_14_8(.a(output_15_8), .b(output_15_9), .y(output_14_8));
wire output_16_8, output_16_9, output_15_8;
mixer gate_output_15_8(.a(output_16_8), .b(output_16_9), .y(output_15_8));
wire output_1_9, output_1_10, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_10), .y(output_0_9));
wire output_2_9, output_2_10, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_10), .y(output_1_9));
wire output_3_9, output_3_10, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_10), .y(output_2_9));
wire output_4_9, output_4_10, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_10), .y(output_3_9));
wire output_5_9, output_5_10, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_10), .y(output_4_9));
wire output_6_9, output_6_10, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_10), .y(output_5_9));
wire output_7_9, output_7_10, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_10), .y(output_6_9));
wire output_8_9, output_8_10, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_10), .y(output_7_9));
wire output_9_9, output_9_10, output_8_9;
mixer gate_output_8_9(.a(output_9_9), .b(output_9_10), .y(output_8_9));
wire output_10_9, output_10_10, output_9_9;
mixer gate_output_9_9(.a(output_10_9), .b(output_10_10), .y(output_9_9));
wire output_11_9, output_11_10, output_10_9;
mixer gate_output_10_9(.a(output_11_9), .b(output_11_10), .y(output_10_9));
wire output_12_9, output_12_10, output_11_9;
mixer gate_output_11_9(.a(output_12_9), .b(output_12_10), .y(output_11_9));
wire output_13_9, output_13_10, output_12_9;
mixer gate_output_12_9(.a(output_13_9), .b(output_13_10), .y(output_12_9));
wire output_14_9, output_14_10, output_13_9;
mixer gate_output_13_9(.a(output_14_9), .b(output_14_10), .y(output_13_9));
wire output_15_9, output_15_10, output_14_9;
mixer gate_output_14_9(.a(output_15_9), .b(output_15_10), .y(output_14_9));
wire output_16_9, output_16_10, output_15_9;
mixer gate_output_15_9(.a(output_16_9), .b(output_16_10), .y(output_15_9));
wire output_1_10, output_1_11, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_11), .y(output_0_10));
wire output_2_10, output_2_11, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_11), .y(output_1_10));
wire output_3_10, output_3_11, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_11), .y(output_2_10));
wire output_4_10, output_4_11, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_11), .y(output_3_10));
wire output_5_10, output_5_11, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_11), .y(output_4_10));
wire output_6_10, output_6_11, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_11), .y(output_5_10));
wire output_7_10, output_7_11, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_11), .y(output_6_10));
wire output_8_10, output_8_11, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_11), .y(output_7_10));
wire output_9_10, output_9_11, output_8_10;
mixer gate_output_8_10(.a(output_9_10), .b(output_9_11), .y(output_8_10));
wire output_10_10, output_10_11, output_9_10;
mixer gate_output_9_10(.a(output_10_10), .b(output_10_11), .y(output_9_10));
wire output_11_10, output_11_11, output_10_10;
mixer gate_output_10_10(.a(output_11_10), .b(output_11_11), .y(output_10_10));
wire output_12_10, output_12_11, output_11_10;
mixer gate_output_11_10(.a(output_12_10), .b(output_12_11), .y(output_11_10));
wire output_13_10, output_13_11, output_12_10;
mixer gate_output_12_10(.a(output_13_10), .b(output_13_11), .y(output_12_10));
wire output_14_10, output_14_11, output_13_10;
mixer gate_output_13_10(.a(output_14_10), .b(output_14_11), .y(output_13_10));
wire output_15_10, output_15_11, output_14_10;
mixer gate_output_14_10(.a(output_15_10), .b(output_15_11), .y(output_14_10));
wire output_16_10, output_16_11, output_15_10;
mixer gate_output_15_10(.a(output_16_10), .b(output_16_11), .y(output_15_10));
wire output_1_11, output_1_12, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_12), .y(output_0_11));
wire output_2_11, output_2_12, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_12), .y(output_1_11));
wire output_3_11, output_3_12, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_12), .y(output_2_11));
wire output_4_11, output_4_12, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_12), .y(output_3_11));
wire output_5_11, output_5_12, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_12), .y(output_4_11));
wire output_6_11, output_6_12, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_12), .y(output_5_11));
wire output_7_11, output_7_12, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_12), .y(output_6_11));
wire output_8_11, output_8_12, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_12), .y(output_7_11));
wire output_9_11, output_9_12, output_8_11;
mixer gate_output_8_11(.a(output_9_11), .b(output_9_12), .y(output_8_11));
wire output_10_11, output_10_12, output_9_11;
mixer gate_output_9_11(.a(output_10_11), .b(output_10_12), .y(output_9_11));
wire output_11_11, output_11_12, output_10_11;
mixer gate_output_10_11(.a(output_11_11), .b(output_11_12), .y(output_10_11));
wire output_12_11, output_12_12, output_11_11;
mixer gate_output_11_11(.a(output_12_11), .b(output_12_12), .y(output_11_11));
wire output_13_11, output_13_12, output_12_11;
mixer gate_output_12_11(.a(output_13_11), .b(output_13_12), .y(output_12_11));
wire output_14_11, output_14_12, output_13_11;
mixer gate_output_13_11(.a(output_14_11), .b(output_14_12), .y(output_13_11));
wire output_15_11, output_15_12, output_14_11;
mixer gate_output_14_11(.a(output_15_11), .b(output_15_12), .y(output_14_11));
wire output_16_11, output_16_12, output_15_11;
mixer gate_output_15_11(.a(output_16_11), .b(output_16_12), .y(output_15_11));
wire output_1_12, output_1_13, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_13), .y(output_0_12));
wire output_2_12, output_2_13, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_13), .y(output_1_12));
wire output_3_12, output_3_13, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_13), .y(output_2_12));
wire output_4_12, output_4_13, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_13), .y(output_3_12));
wire output_5_12, output_5_13, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_13), .y(output_4_12));
wire output_6_12, output_6_13, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_13), .y(output_5_12));
wire output_7_12, output_7_13, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_13), .y(output_6_12));
wire output_8_12, output_8_13, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_13), .y(output_7_12));
wire output_9_12, output_9_13, output_8_12;
mixer gate_output_8_12(.a(output_9_12), .b(output_9_13), .y(output_8_12));
wire output_10_12, output_10_13, output_9_12;
mixer gate_output_9_12(.a(output_10_12), .b(output_10_13), .y(output_9_12));
wire output_11_12, output_11_13, output_10_12;
mixer gate_output_10_12(.a(output_11_12), .b(output_11_13), .y(output_10_12));
wire output_12_12, output_12_13, output_11_12;
mixer gate_output_11_12(.a(output_12_12), .b(output_12_13), .y(output_11_12));
wire output_13_12, output_13_13, output_12_12;
mixer gate_output_12_12(.a(output_13_12), .b(output_13_13), .y(output_12_12));
wire output_14_12, output_14_13, output_13_12;
mixer gate_output_13_12(.a(output_14_12), .b(output_14_13), .y(output_13_12));
wire output_15_12, output_15_13, output_14_12;
mixer gate_output_14_12(.a(output_15_12), .b(output_15_13), .y(output_14_12));
wire output_16_12, output_16_13, output_15_12;
mixer gate_output_15_12(.a(output_16_12), .b(output_16_13), .y(output_15_12));
wire output_1_13, output_1_14, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_14), .y(output_0_13));
wire output_2_13, output_2_14, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_14), .y(output_1_13));
wire output_3_13, output_3_14, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_14), .y(output_2_13));
wire output_4_13, output_4_14, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_14), .y(output_3_13));
wire output_5_13, output_5_14, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_14), .y(output_4_13));
wire output_6_13, output_6_14, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_14), .y(output_5_13));
wire output_7_13, output_7_14, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_14), .y(output_6_13));
wire output_8_13, output_8_14, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_14), .y(output_7_13));
wire output_9_13, output_9_14, output_8_13;
mixer gate_output_8_13(.a(output_9_13), .b(output_9_14), .y(output_8_13));
wire output_10_13, output_10_14, output_9_13;
mixer gate_output_9_13(.a(output_10_13), .b(output_10_14), .y(output_9_13));
wire output_11_13, output_11_14, output_10_13;
mixer gate_output_10_13(.a(output_11_13), .b(output_11_14), .y(output_10_13));
wire output_12_13, output_12_14, output_11_13;
mixer gate_output_11_13(.a(output_12_13), .b(output_12_14), .y(output_11_13));
wire output_13_13, output_13_14, output_12_13;
mixer gate_output_12_13(.a(output_13_13), .b(output_13_14), .y(output_12_13));
wire output_14_13, output_14_14, output_13_13;
mixer gate_output_13_13(.a(output_14_13), .b(output_14_14), .y(output_13_13));
wire output_15_13, output_15_14, output_14_13;
mixer gate_output_14_13(.a(output_15_13), .b(output_15_14), .y(output_14_13));
wire output_16_13, output_16_14, output_15_13;
mixer gate_output_15_13(.a(output_16_13), .b(output_16_14), .y(output_15_13));
wire output_1_14, output_1_15, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_15), .y(output_0_14));
wire output_2_14, output_2_15, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_15), .y(output_1_14));
wire output_3_14, output_3_15, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_15), .y(output_2_14));
wire output_4_14, output_4_15, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_15), .y(output_3_14));
wire output_5_14, output_5_15, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_15), .y(output_4_14));
wire output_6_14, output_6_15, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_15), .y(output_5_14));
wire output_7_14, output_7_15, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_15), .y(output_6_14));
wire output_8_14, output_8_15, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_15), .y(output_7_14));
wire output_9_14, output_9_15, output_8_14;
mixer gate_output_8_14(.a(output_9_14), .b(output_9_15), .y(output_8_14));
wire output_10_14, output_10_15, output_9_14;
mixer gate_output_9_14(.a(output_10_14), .b(output_10_15), .y(output_9_14));
wire output_11_14, output_11_15, output_10_14;
mixer gate_output_10_14(.a(output_11_14), .b(output_11_15), .y(output_10_14));
wire output_12_14, output_12_15, output_11_14;
mixer gate_output_11_14(.a(output_12_14), .b(output_12_15), .y(output_11_14));
wire output_13_14, output_13_15, output_12_14;
mixer gate_output_12_14(.a(output_13_14), .b(output_13_15), .y(output_12_14));
wire output_14_14, output_14_15, output_13_14;
mixer gate_output_13_14(.a(output_14_14), .b(output_14_15), .y(output_13_14));
wire output_15_14, output_15_15, output_14_14;
mixer gate_output_14_14(.a(output_15_14), .b(output_15_15), .y(output_14_14));
wire output_16_14, output_16_15, output_15_14;
mixer gate_output_15_14(.a(output_16_14), .b(output_16_15), .y(output_15_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
wire output_9_15, output_9_0, output_8_15;
mixer gate_output_8_15(.a(output_9_15), .b(output_9_0), .y(output_8_15));
wire output_10_15, output_10_0, output_9_15;
mixer gate_output_9_15(.a(output_10_15), .b(output_10_0), .y(output_9_15));
wire output_11_15, output_11_0, output_10_15;
mixer gate_output_10_15(.a(output_11_15), .b(output_11_0), .y(output_10_15));
wire output_12_15, output_12_0, output_11_15;
mixer gate_output_11_15(.a(output_12_15), .b(output_12_0), .y(output_11_15));
wire output_13_15, output_13_0, output_12_15;
mixer gate_output_12_15(.a(output_13_15), .b(output_13_0), .y(output_12_15));
wire output_14_15, output_14_0, output_13_15;
mixer gate_output_13_15(.a(output_14_15), .b(output_14_0), .y(output_13_15));
wire output_15_15, output_15_0, output_14_15;
mixer gate_output_14_15(.a(output_15_15), .b(output_15_0), .y(output_14_15));
wire output_16_15, output_16_0, output_15_15;
mixer gate_output_15_15(.a(output_16_15), .b(output_16_0), .y(output_15_15));
wire output_1_16, output_1_1, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_1), .y(output_0_16));
wire output_2_16, output_2_1, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_1), .y(output_1_16));
wire output_3_16, output_3_1, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_1), .y(output_2_16));
wire output_4_16, output_4_1, output_3_16;
mixer gate_output_3_16(.a(output_4_16), .b(output_4_1), .y(output_3_16));
wire output_5_16, output_5_1, output_4_16;
mixer gate_output_4_16(.a(output_5_16), .b(output_5_1), .y(output_4_16));
wire output_6_16, output_6_1, output_5_16;
mixer gate_output_5_16(.a(output_6_16), .b(output_6_1), .y(output_5_16));
wire output_7_16, output_7_1, output_6_16;
mixer gate_output_6_16(.a(output_7_16), .b(output_7_1), .y(output_6_16));
wire output_8_16, output_8_1, output_7_16;
mixer gate_output_7_16(.a(output_8_16), .b(output_8_1), .y(output_7_16));
wire output_9_16, output_9_1, output_8_16;
mixer gate_output_8_16(.a(output_9_16), .b(output_9_1), .y(output_8_16));
wire output_10_16, output_10_1, output_9_16;
mixer gate_output_9_16(.a(output_10_16), .b(output_10_1), .y(output_9_16));
wire output_11_16, output_11_1, output_10_16;
mixer gate_output_10_16(.a(output_11_16), .b(output_11_1), .y(output_10_16));
wire output_12_16, output_12_1, output_11_16;
mixer gate_output_11_16(.a(output_12_16), .b(output_12_1), .y(output_11_16));
wire output_13_16, output_13_1, output_12_16;
mixer gate_output_12_16(.a(output_13_16), .b(output_13_1), .y(output_12_16));
wire output_14_16, output_14_1, output_13_16;
mixer gate_output_13_16(.a(output_14_16), .b(output_14_1), .y(output_13_16));
wire output_15_16, output_15_1, output_14_16;
mixer gate_output_14_16(.a(output_15_16), .b(output_15_1), .y(output_14_16));
wire output_16_16, output_16_1, output_15_16;
mixer gate_output_15_16(.a(output_16_16), .b(output_16_1), .y(output_15_16));
wire output_1_17, output_1_2, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_2), .y(output_0_17));
wire output_2_17, output_2_2, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_2), .y(output_1_17));
wire output_3_17, output_3_2, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_2), .y(output_2_17));
wire output_4_17, output_4_2, output_3_17;
mixer gate_output_3_17(.a(output_4_17), .b(output_4_2), .y(output_3_17));
wire output_5_17, output_5_2, output_4_17;
mixer gate_output_4_17(.a(output_5_17), .b(output_5_2), .y(output_4_17));
wire output_6_17, output_6_2, output_5_17;
mixer gate_output_5_17(.a(output_6_17), .b(output_6_2), .y(output_5_17));
wire output_7_17, output_7_2, output_6_17;
mixer gate_output_6_17(.a(output_7_17), .b(output_7_2), .y(output_6_17));
wire output_8_17, output_8_2, output_7_17;
mixer gate_output_7_17(.a(output_8_17), .b(output_8_2), .y(output_7_17));
wire output_9_17, output_9_2, output_8_17;
mixer gate_output_8_17(.a(output_9_17), .b(output_9_2), .y(output_8_17));
wire output_10_17, output_10_2, output_9_17;
mixer gate_output_9_17(.a(output_10_17), .b(output_10_2), .y(output_9_17));
wire output_11_17, output_11_2, output_10_17;
mixer gate_output_10_17(.a(output_11_17), .b(output_11_2), .y(output_10_17));
wire output_12_17, output_12_2, output_11_17;
mixer gate_output_11_17(.a(output_12_17), .b(output_12_2), .y(output_11_17));
wire output_13_17, output_13_2, output_12_17;
mixer gate_output_12_17(.a(output_13_17), .b(output_13_2), .y(output_12_17));
wire output_14_17, output_14_2, output_13_17;
mixer gate_output_13_17(.a(output_14_17), .b(output_14_2), .y(output_13_17));
wire output_15_17, output_15_2, output_14_17;
mixer gate_output_14_17(.a(output_15_17), .b(output_15_2), .y(output_14_17));
wire output_16_17, output_16_2, output_15_17;
mixer gate_output_15_17(.a(output_16_17), .b(output_16_2), .y(output_15_17));
wire output_1_18, output_1_3, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_3), .y(output_0_18));
wire output_2_18, output_2_3, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_3), .y(output_1_18));
wire output_3_18, output_3_3, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_3), .y(output_2_18));
wire output_4_18, output_4_3, output_3_18;
mixer gate_output_3_18(.a(output_4_18), .b(output_4_3), .y(output_3_18));
wire output_5_18, output_5_3, output_4_18;
mixer gate_output_4_18(.a(output_5_18), .b(output_5_3), .y(output_4_18));
wire output_6_18, output_6_3, output_5_18;
mixer gate_output_5_18(.a(output_6_18), .b(output_6_3), .y(output_5_18));
wire output_7_18, output_7_3, output_6_18;
mixer gate_output_6_18(.a(output_7_18), .b(output_7_3), .y(output_6_18));
wire output_8_18, output_8_3, output_7_18;
mixer gate_output_7_18(.a(output_8_18), .b(output_8_3), .y(output_7_18));
wire output_9_18, output_9_3, output_8_18;
mixer gate_output_8_18(.a(output_9_18), .b(output_9_3), .y(output_8_18));
wire output_10_18, output_10_3, output_9_18;
mixer gate_output_9_18(.a(output_10_18), .b(output_10_3), .y(output_9_18));
wire output_11_18, output_11_3, output_10_18;
mixer gate_output_10_18(.a(output_11_18), .b(output_11_3), .y(output_10_18));
wire output_12_18, output_12_3, output_11_18;
mixer gate_output_11_18(.a(output_12_18), .b(output_12_3), .y(output_11_18));
wire output_13_18, output_13_3, output_12_18;
mixer gate_output_12_18(.a(output_13_18), .b(output_13_3), .y(output_12_18));
wire output_14_18, output_14_3, output_13_18;
mixer gate_output_13_18(.a(output_14_18), .b(output_14_3), .y(output_13_18));
wire output_15_18, output_15_3, output_14_18;
mixer gate_output_14_18(.a(output_15_18), .b(output_15_3), .y(output_14_18));
wire output_16_18, output_16_3, output_15_18;
mixer gate_output_15_18(.a(output_16_18), .b(output_16_3), .y(output_15_18));
wire output_1_19, output_1_4, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_4), .y(output_0_19));
wire output_2_19, output_2_4, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_4), .y(output_1_19));
wire output_3_19, output_3_4, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_4), .y(output_2_19));
wire output_4_19, output_4_4, output_3_19;
mixer gate_output_3_19(.a(output_4_19), .b(output_4_4), .y(output_3_19));
wire output_5_19, output_5_4, output_4_19;
mixer gate_output_4_19(.a(output_5_19), .b(output_5_4), .y(output_4_19));
wire output_6_19, output_6_4, output_5_19;
mixer gate_output_5_19(.a(output_6_19), .b(output_6_4), .y(output_5_19));
wire output_7_19, output_7_4, output_6_19;
mixer gate_output_6_19(.a(output_7_19), .b(output_7_4), .y(output_6_19));
wire output_8_19, output_8_4, output_7_19;
mixer gate_output_7_19(.a(output_8_19), .b(output_8_4), .y(output_7_19));
wire output_9_19, output_9_4, output_8_19;
mixer gate_output_8_19(.a(output_9_19), .b(output_9_4), .y(output_8_19));
wire output_10_19, output_10_4, output_9_19;
mixer gate_output_9_19(.a(output_10_19), .b(output_10_4), .y(output_9_19));
wire output_11_19, output_11_4, output_10_19;
mixer gate_output_10_19(.a(output_11_19), .b(output_11_4), .y(output_10_19));
wire output_12_19, output_12_4, output_11_19;
mixer gate_output_11_19(.a(output_12_19), .b(output_12_4), .y(output_11_19));
wire output_13_19, output_13_4, output_12_19;
mixer gate_output_12_19(.a(output_13_19), .b(output_13_4), .y(output_12_19));
wire output_14_19, output_14_4, output_13_19;
mixer gate_output_13_19(.a(output_14_19), .b(output_14_4), .y(output_13_19));
wire output_15_19, output_15_4, output_14_19;
mixer gate_output_14_19(.a(output_15_19), .b(output_15_4), .y(output_14_19));
wire output_16_19, output_16_4, output_15_19;
mixer gate_output_15_19(.a(output_16_19), .b(output_16_4), .y(output_15_19));
wire output_1_20, output_1_5, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_5), .y(output_0_20));
wire output_2_20, output_2_5, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_5), .y(output_1_20));
wire output_3_20, output_3_5, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_5), .y(output_2_20));
wire output_4_20, output_4_5, output_3_20;
mixer gate_output_3_20(.a(output_4_20), .b(output_4_5), .y(output_3_20));
wire output_5_20, output_5_5, output_4_20;
mixer gate_output_4_20(.a(output_5_20), .b(output_5_5), .y(output_4_20));
wire output_6_20, output_6_5, output_5_20;
mixer gate_output_5_20(.a(output_6_20), .b(output_6_5), .y(output_5_20));
wire output_7_20, output_7_5, output_6_20;
mixer gate_output_6_20(.a(output_7_20), .b(output_7_5), .y(output_6_20));
wire output_8_20, output_8_5, output_7_20;
mixer gate_output_7_20(.a(output_8_20), .b(output_8_5), .y(output_7_20));
wire output_9_20, output_9_5, output_8_20;
mixer gate_output_8_20(.a(output_9_20), .b(output_9_5), .y(output_8_20));
wire output_10_20, output_10_5, output_9_20;
mixer gate_output_9_20(.a(output_10_20), .b(output_10_5), .y(output_9_20));
wire output_11_20, output_11_5, output_10_20;
mixer gate_output_10_20(.a(output_11_20), .b(output_11_5), .y(output_10_20));
wire output_12_20, output_12_5, output_11_20;
mixer gate_output_11_20(.a(output_12_20), .b(output_12_5), .y(output_11_20));
wire output_13_20, output_13_5, output_12_20;
mixer gate_output_12_20(.a(output_13_20), .b(output_13_5), .y(output_12_20));
wire output_14_20, output_14_5, output_13_20;
mixer gate_output_13_20(.a(output_14_20), .b(output_14_5), .y(output_13_20));
wire output_15_20, output_15_5, output_14_20;
mixer gate_output_14_20(.a(output_15_20), .b(output_15_5), .y(output_14_20));
wire output_16_20, output_16_5, output_15_20;
mixer gate_output_15_20(.a(output_16_20), .b(output_16_5), .y(output_15_20));
wire output_1_21, output_1_6, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_6), .y(output_0_21));
wire output_2_21, output_2_6, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_6), .y(output_1_21));
wire output_3_21, output_3_6, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_6), .y(output_2_21));
wire output_4_21, output_4_6, output_3_21;
mixer gate_output_3_21(.a(output_4_21), .b(output_4_6), .y(output_3_21));
wire output_5_21, output_5_6, output_4_21;
mixer gate_output_4_21(.a(output_5_21), .b(output_5_6), .y(output_4_21));
wire output_6_21, output_6_6, output_5_21;
mixer gate_output_5_21(.a(output_6_21), .b(output_6_6), .y(output_5_21));
wire output_7_21, output_7_6, output_6_21;
mixer gate_output_6_21(.a(output_7_21), .b(output_7_6), .y(output_6_21));
wire output_8_21, output_8_6, output_7_21;
mixer gate_output_7_21(.a(output_8_21), .b(output_8_6), .y(output_7_21));
wire output_9_21, output_9_6, output_8_21;
mixer gate_output_8_21(.a(output_9_21), .b(output_9_6), .y(output_8_21));
wire output_10_21, output_10_6, output_9_21;
mixer gate_output_9_21(.a(output_10_21), .b(output_10_6), .y(output_9_21));
wire output_11_21, output_11_6, output_10_21;
mixer gate_output_10_21(.a(output_11_21), .b(output_11_6), .y(output_10_21));
wire output_12_21, output_12_6, output_11_21;
mixer gate_output_11_21(.a(output_12_21), .b(output_12_6), .y(output_11_21));
wire output_13_21, output_13_6, output_12_21;
mixer gate_output_12_21(.a(output_13_21), .b(output_13_6), .y(output_12_21));
wire output_14_21, output_14_6, output_13_21;
mixer gate_output_13_21(.a(output_14_21), .b(output_14_6), .y(output_13_21));
wire output_15_21, output_15_6, output_14_21;
mixer gate_output_14_21(.a(output_15_21), .b(output_15_6), .y(output_14_21));
wire output_16_21, output_16_6, output_15_21;
mixer gate_output_15_21(.a(output_16_21), .b(output_16_6), .y(output_15_21));
wire output_1_22, output_1_7, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_7), .y(output_0_22));
wire output_2_22, output_2_7, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_7), .y(output_1_22));
wire output_3_22, output_3_7, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_7), .y(output_2_22));
wire output_4_22, output_4_7, output_3_22;
mixer gate_output_3_22(.a(output_4_22), .b(output_4_7), .y(output_3_22));
wire output_5_22, output_5_7, output_4_22;
mixer gate_output_4_22(.a(output_5_22), .b(output_5_7), .y(output_4_22));
wire output_6_22, output_6_7, output_5_22;
mixer gate_output_5_22(.a(output_6_22), .b(output_6_7), .y(output_5_22));
wire output_7_22, output_7_7, output_6_22;
mixer gate_output_6_22(.a(output_7_22), .b(output_7_7), .y(output_6_22));
wire output_8_22, output_8_7, output_7_22;
mixer gate_output_7_22(.a(output_8_22), .b(output_8_7), .y(output_7_22));
wire output_9_22, output_9_7, output_8_22;
mixer gate_output_8_22(.a(output_9_22), .b(output_9_7), .y(output_8_22));
wire output_10_22, output_10_7, output_9_22;
mixer gate_output_9_22(.a(output_10_22), .b(output_10_7), .y(output_9_22));
wire output_11_22, output_11_7, output_10_22;
mixer gate_output_10_22(.a(output_11_22), .b(output_11_7), .y(output_10_22));
wire output_12_22, output_12_7, output_11_22;
mixer gate_output_11_22(.a(output_12_22), .b(output_12_7), .y(output_11_22));
wire output_13_22, output_13_7, output_12_22;
mixer gate_output_12_22(.a(output_13_22), .b(output_13_7), .y(output_12_22));
wire output_14_22, output_14_7, output_13_22;
mixer gate_output_13_22(.a(output_14_22), .b(output_14_7), .y(output_13_22));
wire output_15_22, output_15_7, output_14_22;
mixer gate_output_14_22(.a(output_15_22), .b(output_15_7), .y(output_14_22));
wire output_16_22, output_16_7, output_15_22;
mixer gate_output_15_22(.a(output_16_22), .b(output_16_7), .y(output_15_22));
wire output_1_23, output_1_8, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_8), .y(output_0_23));
wire output_2_23, output_2_8, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_8), .y(output_1_23));
wire output_3_23, output_3_8, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_8), .y(output_2_23));
wire output_4_23, output_4_8, output_3_23;
mixer gate_output_3_23(.a(output_4_23), .b(output_4_8), .y(output_3_23));
wire output_5_23, output_5_8, output_4_23;
mixer gate_output_4_23(.a(output_5_23), .b(output_5_8), .y(output_4_23));
wire output_6_23, output_6_8, output_5_23;
mixer gate_output_5_23(.a(output_6_23), .b(output_6_8), .y(output_5_23));
wire output_7_23, output_7_8, output_6_23;
mixer gate_output_6_23(.a(output_7_23), .b(output_7_8), .y(output_6_23));
wire output_8_23, output_8_8, output_7_23;
mixer gate_output_7_23(.a(output_8_23), .b(output_8_8), .y(output_7_23));
wire output_9_23, output_9_8, output_8_23;
mixer gate_output_8_23(.a(output_9_23), .b(output_9_8), .y(output_8_23));
wire output_10_23, output_10_8, output_9_23;
mixer gate_output_9_23(.a(output_10_23), .b(output_10_8), .y(output_9_23));
wire output_11_23, output_11_8, output_10_23;
mixer gate_output_10_23(.a(output_11_23), .b(output_11_8), .y(output_10_23));
wire output_12_23, output_12_8, output_11_23;
mixer gate_output_11_23(.a(output_12_23), .b(output_12_8), .y(output_11_23));
wire output_13_23, output_13_8, output_12_23;
mixer gate_output_12_23(.a(output_13_23), .b(output_13_8), .y(output_12_23));
wire output_14_23, output_14_8, output_13_23;
mixer gate_output_13_23(.a(output_14_23), .b(output_14_8), .y(output_13_23));
wire output_15_23, output_15_8, output_14_23;
mixer gate_output_14_23(.a(output_15_23), .b(output_15_8), .y(output_14_23));
wire output_16_23, output_16_8, output_15_23;
mixer gate_output_15_23(.a(output_16_23), .b(output_16_8), .y(output_15_23));
wire output_1_24, output_1_9, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_9), .y(output_0_24));
wire output_2_24, output_2_9, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_9), .y(output_1_24));
wire output_3_24, output_3_9, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_9), .y(output_2_24));
wire output_4_24, output_4_9, output_3_24;
mixer gate_output_3_24(.a(output_4_24), .b(output_4_9), .y(output_3_24));
wire output_5_24, output_5_9, output_4_24;
mixer gate_output_4_24(.a(output_5_24), .b(output_5_9), .y(output_4_24));
wire output_6_24, output_6_9, output_5_24;
mixer gate_output_5_24(.a(output_6_24), .b(output_6_9), .y(output_5_24));
wire output_7_24, output_7_9, output_6_24;
mixer gate_output_6_24(.a(output_7_24), .b(output_7_9), .y(output_6_24));
wire output_8_24, output_8_9, output_7_24;
mixer gate_output_7_24(.a(output_8_24), .b(output_8_9), .y(output_7_24));
wire output_9_24, output_9_9, output_8_24;
mixer gate_output_8_24(.a(output_9_24), .b(output_9_9), .y(output_8_24));
wire output_10_24, output_10_9, output_9_24;
mixer gate_output_9_24(.a(output_10_24), .b(output_10_9), .y(output_9_24));
wire output_11_24, output_11_9, output_10_24;
mixer gate_output_10_24(.a(output_11_24), .b(output_11_9), .y(output_10_24));
wire output_12_24, output_12_9, output_11_24;
mixer gate_output_11_24(.a(output_12_24), .b(output_12_9), .y(output_11_24));
wire output_13_24, output_13_9, output_12_24;
mixer gate_output_12_24(.a(output_13_24), .b(output_13_9), .y(output_12_24));
wire output_14_24, output_14_9, output_13_24;
mixer gate_output_13_24(.a(output_14_24), .b(output_14_9), .y(output_13_24));
wire output_15_24, output_15_9, output_14_24;
mixer gate_output_14_24(.a(output_15_24), .b(output_15_9), .y(output_14_24));
wire output_16_24, output_16_9, output_15_24;
mixer gate_output_15_24(.a(output_16_24), .b(output_16_9), .y(output_15_24));
wire output_1_25, output_1_10, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_10), .y(output_0_25));
wire output_2_25, output_2_10, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_10), .y(output_1_25));
wire output_3_25, output_3_10, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_10), .y(output_2_25));
wire output_4_25, output_4_10, output_3_25;
mixer gate_output_3_25(.a(output_4_25), .b(output_4_10), .y(output_3_25));
wire output_5_25, output_5_10, output_4_25;
mixer gate_output_4_25(.a(output_5_25), .b(output_5_10), .y(output_4_25));
wire output_6_25, output_6_10, output_5_25;
mixer gate_output_5_25(.a(output_6_25), .b(output_6_10), .y(output_5_25));
wire output_7_25, output_7_10, output_6_25;
mixer gate_output_6_25(.a(output_7_25), .b(output_7_10), .y(output_6_25));
wire output_8_25, output_8_10, output_7_25;
mixer gate_output_7_25(.a(output_8_25), .b(output_8_10), .y(output_7_25));
wire output_9_25, output_9_10, output_8_25;
mixer gate_output_8_25(.a(output_9_25), .b(output_9_10), .y(output_8_25));
wire output_10_25, output_10_10, output_9_25;
mixer gate_output_9_25(.a(output_10_25), .b(output_10_10), .y(output_9_25));
wire output_11_25, output_11_10, output_10_25;
mixer gate_output_10_25(.a(output_11_25), .b(output_11_10), .y(output_10_25));
wire output_12_25, output_12_10, output_11_25;
mixer gate_output_11_25(.a(output_12_25), .b(output_12_10), .y(output_11_25));
wire output_13_25, output_13_10, output_12_25;
mixer gate_output_12_25(.a(output_13_25), .b(output_13_10), .y(output_12_25));
wire output_14_25, output_14_10, output_13_25;
mixer gate_output_13_25(.a(output_14_25), .b(output_14_10), .y(output_13_25));
wire output_15_25, output_15_10, output_14_25;
mixer gate_output_14_25(.a(output_15_25), .b(output_15_10), .y(output_14_25));
wire output_16_25, output_16_10, output_15_25;
mixer gate_output_15_25(.a(output_16_25), .b(output_16_10), .y(output_15_25));
wire output_1_26, output_1_11, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_11), .y(output_0_26));
wire output_2_26, output_2_11, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_11), .y(output_1_26));
wire output_3_26, output_3_11, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_11), .y(output_2_26));
wire output_4_26, output_4_11, output_3_26;
mixer gate_output_3_26(.a(output_4_26), .b(output_4_11), .y(output_3_26));
wire output_5_26, output_5_11, output_4_26;
mixer gate_output_4_26(.a(output_5_26), .b(output_5_11), .y(output_4_26));
wire output_6_26, output_6_11, output_5_26;
mixer gate_output_5_26(.a(output_6_26), .b(output_6_11), .y(output_5_26));
wire output_7_26, output_7_11, output_6_26;
mixer gate_output_6_26(.a(output_7_26), .b(output_7_11), .y(output_6_26));
wire output_8_26, output_8_11, output_7_26;
mixer gate_output_7_26(.a(output_8_26), .b(output_8_11), .y(output_7_26));
wire output_9_26, output_9_11, output_8_26;
mixer gate_output_8_26(.a(output_9_26), .b(output_9_11), .y(output_8_26));
wire output_10_26, output_10_11, output_9_26;
mixer gate_output_9_26(.a(output_10_26), .b(output_10_11), .y(output_9_26));
wire output_11_26, output_11_11, output_10_26;
mixer gate_output_10_26(.a(output_11_26), .b(output_11_11), .y(output_10_26));
wire output_12_26, output_12_11, output_11_26;
mixer gate_output_11_26(.a(output_12_26), .b(output_12_11), .y(output_11_26));
wire output_13_26, output_13_11, output_12_26;
mixer gate_output_12_26(.a(output_13_26), .b(output_13_11), .y(output_12_26));
wire output_14_26, output_14_11, output_13_26;
mixer gate_output_13_26(.a(output_14_26), .b(output_14_11), .y(output_13_26));
wire output_15_26, output_15_11, output_14_26;
mixer gate_output_14_26(.a(output_15_26), .b(output_15_11), .y(output_14_26));
wire output_16_26, output_16_11, output_15_26;
mixer gate_output_15_26(.a(output_16_26), .b(output_16_11), .y(output_15_26));
wire output_1_27, output_1_12, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_12), .y(output_0_27));
wire output_2_27, output_2_12, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_12), .y(output_1_27));
wire output_3_27, output_3_12, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_12), .y(output_2_27));
wire output_4_27, output_4_12, output_3_27;
mixer gate_output_3_27(.a(output_4_27), .b(output_4_12), .y(output_3_27));
wire output_5_27, output_5_12, output_4_27;
mixer gate_output_4_27(.a(output_5_27), .b(output_5_12), .y(output_4_27));
wire output_6_27, output_6_12, output_5_27;
mixer gate_output_5_27(.a(output_6_27), .b(output_6_12), .y(output_5_27));
wire output_7_27, output_7_12, output_6_27;
mixer gate_output_6_27(.a(output_7_27), .b(output_7_12), .y(output_6_27));
wire output_8_27, output_8_12, output_7_27;
mixer gate_output_7_27(.a(output_8_27), .b(output_8_12), .y(output_7_27));
wire output_9_27, output_9_12, output_8_27;
mixer gate_output_8_27(.a(output_9_27), .b(output_9_12), .y(output_8_27));
wire output_10_27, output_10_12, output_9_27;
mixer gate_output_9_27(.a(output_10_27), .b(output_10_12), .y(output_9_27));
wire output_11_27, output_11_12, output_10_27;
mixer gate_output_10_27(.a(output_11_27), .b(output_11_12), .y(output_10_27));
wire output_12_27, output_12_12, output_11_27;
mixer gate_output_11_27(.a(output_12_27), .b(output_12_12), .y(output_11_27));
wire output_13_27, output_13_12, output_12_27;
mixer gate_output_12_27(.a(output_13_27), .b(output_13_12), .y(output_12_27));
wire output_14_27, output_14_12, output_13_27;
mixer gate_output_13_27(.a(output_14_27), .b(output_14_12), .y(output_13_27));
wire output_15_27, output_15_12, output_14_27;
mixer gate_output_14_27(.a(output_15_27), .b(output_15_12), .y(output_14_27));
wire output_16_27, output_16_12, output_15_27;
mixer gate_output_15_27(.a(output_16_27), .b(output_16_12), .y(output_15_27));
wire output_1_28, output_1_13, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_13), .y(output_0_28));
wire output_2_28, output_2_13, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_13), .y(output_1_28));
wire output_3_28, output_3_13, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_13), .y(output_2_28));
wire output_4_28, output_4_13, output_3_28;
mixer gate_output_3_28(.a(output_4_28), .b(output_4_13), .y(output_3_28));
wire output_5_28, output_5_13, output_4_28;
mixer gate_output_4_28(.a(output_5_28), .b(output_5_13), .y(output_4_28));
wire output_6_28, output_6_13, output_5_28;
mixer gate_output_5_28(.a(output_6_28), .b(output_6_13), .y(output_5_28));
wire output_7_28, output_7_13, output_6_28;
mixer gate_output_6_28(.a(output_7_28), .b(output_7_13), .y(output_6_28));
wire output_8_28, output_8_13, output_7_28;
mixer gate_output_7_28(.a(output_8_28), .b(output_8_13), .y(output_7_28));
wire output_9_28, output_9_13, output_8_28;
mixer gate_output_8_28(.a(output_9_28), .b(output_9_13), .y(output_8_28));
wire output_10_28, output_10_13, output_9_28;
mixer gate_output_9_28(.a(output_10_28), .b(output_10_13), .y(output_9_28));
wire output_11_28, output_11_13, output_10_28;
mixer gate_output_10_28(.a(output_11_28), .b(output_11_13), .y(output_10_28));
wire output_12_28, output_12_13, output_11_28;
mixer gate_output_11_28(.a(output_12_28), .b(output_12_13), .y(output_11_28));
wire output_13_28, output_13_13, output_12_28;
mixer gate_output_12_28(.a(output_13_28), .b(output_13_13), .y(output_12_28));
wire output_14_28, output_14_13, output_13_28;
mixer gate_output_13_28(.a(output_14_28), .b(output_14_13), .y(output_13_28));
wire output_15_28, output_15_13, output_14_28;
mixer gate_output_14_28(.a(output_15_28), .b(output_15_13), .y(output_14_28));
wire output_16_28, output_16_13, output_15_28;
mixer gate_output_15_28(.a(output_16_28), .b(output_16_13), .y(output_15_28));
wire output_1_29, output_1_14, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_14), .y(output_0_29));
wire output_2_29, output_2_14, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_14), .y(output_1_29));
wire output_3_29, output_3_14, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_14), .y(output_2_29));
wire output_4_29, output_4_14, output_3_29;
mixer gate_output_3_29(.a(output_4_29), .b(output_4_14), .y(output_3_29));
wire output_5_29, output_5_14, output_4_29;
mixer gate_output_4_29(.a(output_5_29), .b(output_5_14), .y(output_4_29));
wire output_6_29, output_6_14, output_5_29;
mixer gate_output_5_29(.a(output_6_29), .b(output_6_14), .y(output_5_29));
wire output_7_29, output_7_14, output_6_29;
mixer gate_output_6_29(.a(output_7_29), .b(output_7_14), .y(output_6_29));
wire output_8_29, output_8_14, output_7_29;
mixer gate_output_7_29(.a(output_8_29), .b(output_8_14), .y(output_7_29));
wire output_9_29, output_9_14, output_8_29;
mixer gate_output_8_29(.a(output_9_29), .b(output_9_14), .y(output_8_29));
wire output_10_29, output_10_14, output_9_29;
mixer gate_output_9_29(.a(output_10_29), .b(output_10_14), .y(output_9_29));
wire output_11_29, output_11_14, output_10_29;
mixer gate_output_10_29(.a(output_11_29), .b(output_11_14), .y(output_10_29));
wire output_12_29, output_12_14, output_11_29;
mixer gate_output_11_29(.a(output_12_29), .b(output_12_14), .y(output_11_29));
wire output_13_29, output_13_14, output_12_29;
mixer gate_output_12_29(.a(output_13_29), .b(output_13_14), .y(output_12_29));
wire output_14_29, output_14_14, output_13_29;
mixer gate_output_13_29(.a(output_14_29), .b(output_14_14), .y(output_13_29));
wire output_15_29, output_15_14, output_14_29;
mixer gate_output_14_29(.a(output_15_29), .b(output_15_14), .y(output_14_29));
wire output_16_29, output_16_14, output_15_29;
mixer gate_output_15_29(.a(output_16_29), .b(output_16_14), .y(output_15_29));
wire output_1_30, output_1_15, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_15), .y(output_0_30));
wire output_2_30, output_2_15, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_15), .y(output_1_30));
wire output_3_30, output_3_15, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_15), .y(output_2_30));
wire output_4_30, output_4_15, output_3_30;
mixer gate_output_3_30(.a(output_4_30), .b(output_4_15), .y(output_3_30));
wire output_5_30, output_5_15, output_4_30;
mixer gate_output_4_30(.a(output_5_30), .b(output_5_15), .y(output_4_30));
wire output_6_30, output_6_15, output_5_30;
mixer gate_output_5_30(.a(output_6_30), .b(output_6_15), .y(output_5_30));
wire output_7_30, output_7_15, output_6_30;
mixer gate_output_6_30(.a(output_7_30), .b(output_7_15), .y(output_6_30));
wire output_8_30, output_8_15, output_7_30;
mixer gate_output_7_30(.a(output_8_30), .b(output_8_15), .y(output_7_30));
wire output_9_30, output_9_15, output_8_30;
mixer gate_output_8_30(.a(output_9_30), .b(output_9_15), .y(output_8_30));
wire output_10_30, output_10_15, output_9_30;
mixer gate_output_9_30(.a(output_10_30), .b(output_10_15), .y(output_9_30));
wire output_11_30, output_11_15, output_10_30;
mixer gate_output_10_30(.a(output_11_30), .b(output_11_15), .y(output_10_30));
wire output_12_30, output_12_15, output_11_30;
mixer gate_output_11_30(.a(output_12_30), .b(output_12_15), .y(output_11_30));
wire output_13_30, output_13_15, output_12_30;
mixer gate_output_12_30(.a(output_13_30), .b(output_13_15), .y(output_12_30));
wire output_14_30, output_14_15, output_13_30;
mixer gate_output_13_30(.a(output_14_30), .b(output_14_15), .y(output_13_30));
wire output_15_30, output_15_15, output_14_30;
mixer gate_output_14_30(.a(output_15_30), .b(output_15_15), .y(output_14_30));
wire output_16_30, output_16_15, output_15_30;
mixer gate_output_15_30(.a(output_16_30), .b(output_16_15), .y(output_15_30));
wire output_1_31, output_1_0, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_0), .y(output_0_31));
wire output_2_31, output_2_0, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_0), .y(output_1_31));
wire output_3_31, output_3_0, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_0), .y(output_2_31));
wire output_4_31, output_4_0, output_3_31;
mixer gate_output_3_31(.a(output_4_31), .b(output_4_0), .y(output_3_31));
wire output_5_31, output_5_0, output_4_31;
mixer gate_output_4_31(.a(output_5_31), .b(output_5_0), .y(output_4_31));
wire output_6_31, output_6_0, output_5_31;
mixer gate_output_5_31(.a(output_6_31), .b(output_6_0), .y(output_5_31));
wire output_7_31, output_7_0, output_6_31;
mixer gate_output_6_31(.a(output_7_31), .b(output_7_0), .y(output_6_31));
wire output_8_31, output_8_0, output_7_31;
mixer gate_output_7_31(.a(output_8_31), .b(output_8_0), .y(output_7_31));
wire output_9_31, output_9_0, output_8_31;
mixer gate_output_8_31(.a(output_9_31), .b(output_9_0), .y(output_8_31));
wire output_10_31, output_10_0, output_9_31;
mixer gate_output_9_31(.a(output_10_31), .b(output_10_0), .y(output_9_31));
wire output_11_31, output_11_0, output_10_31;
mixer gate_output_10_31(.a(output_11_31), .b(output_11_0), .y(output_10_31));
wire output_12_31, output_12_0, output_11_31;
mixer gate_output_11_31(.a(output_12_31), .b(output_12_0), .y(output_11_31));
wire output_13_31, output_13_0, output_12_31;
mixer gate_output_12_31(.a(output_13_31), .b(output_13_0), .y(output_12_31));
wire output_14_31, output_14_0, output_13_31;
mixer gate_output_13_31(.a(output_14_31), .b(output_14_0), .y(output_13_31));
wire output_15_31, output_15_0, output_14_31;
mixer gate_output_14_31(.a(output_15_31), .b(output_15_0), .y(output_14_31));
wire output_16_31, output_16_0, output_15_31;
mixer gate_output_15_31(.a(output_16_31), .b(output_16_0), .y(output_15_31));
assign output_0 = output_0_0;
wire output_0_32;
assign output_0_32 = input_0;
assign output_1 = output_1_0;
wire output_1_32;
assign output_1_32 = input_1;
assign output_2 = output_2_0;
wire output_2_32;
assign output_2_32 = input_2;
assign output_3 = output_3_0;
wire output_3_32;
assign output_3_32 = input_3;
assign output_4 = output_4_0;
wire output_4_32;
assign output_4_32 = input_4;
assign output_5 = output_5_0;
wire output_5_32;
assign output_5_32 = input_5;
assign output_6 = output_6_0;
wire output_6_32;
assign output_6_32 = input_6;
assign output_7 = output_7_0;
wire output_7_32;
assign output_7_32 = input_7;
assign output_8 = output_8_0;
wire output_8_32;
assign output_8_32 = input_8;
assign output_9 = output_9_0;
wire output_9_32;
assign output_9_32 = input_9;
assign output_10 = output_10_0;
wire output_10_32;
assign output_10_32 = input_10;
assign output_11 = output_11_0;
wire output_11_32;
assign output_11_32 = input_11;
assign output_12 = output_12_0;
wire output_12_32;
assign output_12_32 = input_12;
assign output_13 = output_13_0;
wire output_13_32;
assign output_13_32 = input_13;
assign output_14 = output_14_0;
wire output_14_32;
assign output_14_32 = input_14;
assign output_15 = output_15_0;
wire output_15_32;
assign output_15_32 = input_15;
endmodule
