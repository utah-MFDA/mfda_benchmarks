module multiplexer_12 (
inout k_0_0,k_12_0,k_12_1,k_12_2,k_12_3,k_12_4,k_12_5,k_12_6,k_12_7,k_12_8,k_12_9,k_12_10,k_12_11,k_12_12,k_12_13,k_12_14,k_12_15,k_12_16,k_12_17,k_12_18,k_12_19,k_12_20,k_12_21,k_12_22,k_12_23,k_12_24,k_12_25,k_12_26,k_12_27,k_12_28,k_12_29,k_12_30,k_12_31,k_12_32,k_12_33,k_12_34,k_12_35,k_12_36,k_12_37,k_12_38,k_12_39,k_12_40,k_12_41,k_12_42,k_12_43,k_12_44,k_12_45,k_12_46,k_12_47,k_12_48,k_12_49,k_12_50,k_12_51,k_12_52,k_12_53,k_12_54,k_12_55,k_12_56,k_12_57,k_12_58,k_12_59,k_12_60,k_12_61,k_12_62,k_12_63,k_12_64,k_12_65,k_12_66,k_12_67,k_12_68,k_12_69,k_12_70,k_12_71,k_12_72,k_12_73,k_12_74,k_12_75,k_12_76,k_12_77,k_12_78,k_12_79,k_12_80,k_12_81,k_12_82,k_12_83,k_12_84,k_12_85,k_12_86,k_12_87,k_12_88,k_12_89,k_12_90,k_12_91,k_12_92,k_12_93,k_12_94,k_12_95,k_12_96,k_12_97,k_12_98,k_12_99,k_12_100,k_12_101,k_12_102,k_12_103,k_12_104,k_12_105,k_12_106,k_12_107,k_12_108,k_12_109,k_12_110,k_12_111,k_12_112,k_12_113,k_12_114,k_12_115,k_12_116,k_12_117,k_12_118,k_12_119,k_12_120,k_12_121,k_12_122,k_12_123,k_12_124,k_12_125,k_12_126,k_12_127,k_12_128,k_12_129,k_12_130,k_12_131,k_12_132,k_12_133,k_12_134,k_12_135,k_12_136,k_12_137,k_12_138,k_12_139,k_12_140,k_12_141,k_12_142,k_12_143,k_12_144,k_12_145,k_12_146,k_12_147,k_12_148,k_12_149,k_12_150,k_12_151,k_12_152,k_12_153,k_12_154,k_12_155,k_12_156,k_12_157,k_12_158,k_12_159,k_12_160,k_12_161,k_12_162,k_12_163,k_12_164,k_12_165,k_12_166,k_12_167,k_12_168,k_12_169,k_12_170,k_12_171,k_12_172,k_12_173,k_12_174,k_12_175,k_12_176,k_12_177,k_12_178,k_12_179,k_12_180,k_12_181,k_12_182,k_12_183,k_12_184,k_12_185,k_12_186,k_12_187,k_12_188,k_12_189,k_12_190,k_12_191,k_12_192,k_12_193,k_12_194,k_12_195,k_12_196,k_12_197,k_12_198,k_12_199,k_12_200,k_12_201,k_12_202,k_12_203,k_12_204,k_12_205,k_12_206,k_12_207,k_12_208,k_12_209,k_12_210,k_12_211,k_12_212,k_12_213,k_12_214,k_12_215,k_12_216,k_12_217,k_12_218,k_12_219,k_12_220,k_12_221,k_12_222,k_12_223,k_12_224,k_12_225,k_12_226,k_12_227,k_12_228,k_12_229,k_12_230,k_12_231,k_12_232,k_12_233,k_12_234,k_12_235,k_12_236,k_12_237,k_12_238,k_12_239,k_12_240,k_12_241,k_12_242,k_12_243,k_12_244,k_12_245,k_12_246,k_12_247,k_12_248,k_12_249,k_12_250,k_12_251,k_12_252,k_12_253,k_12_254,k_12_255,k_12_256,k_12_257,k_12_258,k_12_259,k_12_260,k_12_261,k_12_262,k_12_263,k_12_264,k_12_265,k_12_266,k_12_267,k_12_268,k_12_269,k_12_270,k_12_271,k_12_272,k_12_273,k_12_274,k_12_275,k_12_276,k_12_277,k_12_278,k_12_279,k_12_280,k_12_281,k_12_282,k_12_283,k_12_284,k_12_285,k_12_286,k_12_287,k_12_288,k_12_289,k_12_290,k_12_291,k_12_292,k_12_293,k_12_294,k_12_295,k_12_296,k_12_297,k_12_298,k_12_299,k_12_300,k_12_301,k_12_302,k_12_303,k_12_304,k_12_305,k_12_306,k_12_307,k_12_308,k_12_309,k_12_310,k_12_311,k_12_312,k_12_313,k_12_314,k_12_315,k_12_316,k_12_317,k_12_318,k_12_319,k_12_320,k_12_321,k_12_322,k_12_323,k_12_324,k_12_325,k_12_326,k_12_327,k_12_328,k_12_329,k_12_330,k_12_331,k_12_332,k_12_333,k_12_334,k_12_335,k_12_336,k_12_337,k_12_338,k_12_339,k_12_340,k_12_341,k_12_342,k_12_343,k_12_344,k_12_345,k_12_346,k_12_347,k_12_348,k_12_349,k_12_350,k_12_351,k_12_352,k_12_353,k_12_354,k_12_355,k_12_356,k_12_357,k_12_358,k_12_359,k_12_360,k_12_361,k_12_362,k_12_363,k_12_364,k_12_365,k_12_366,k_12_367,k_12_368,k_12_369,k_12_370,k_12_371,k_12_372,k_12_373,k_12_374,k_12_375,k_12_376,k_12_377,k_12_378,k_12_379,k_12_380,k_12_381,k_12_382,k_12_383,k_12_384,k_12_385,k_12_386,k_12_387,k_12_388,k_12_389,k_12_390,k_12_391,k_12_392,k_12_393,k_12_394,k_12_395,k_12_396,k_12_397,k_12_398,k_12_399,k_12_400,k_12_401,k_12_402,k_12_403,k_12_404,k_12_405,k_12_406,k_12_407,k_12_408,k_12_409,k_12_410,k_12_411,k_12_412,k_12_413,k_12_414,k_12_415,k_12_416,k_12_417,k_12_418,k_12_419,k_12_420,k_12_421,k_12_422,k_12_423,k_12_424,k_12_425,k_12_426,k_12_427,k_12_428,k_12_429,k_12_430,k_12_431,k_12_432,k_12_433,k_12_434,k_12_435,k_12_436,k_12_437,k_12_438,k_12_439,k_12_440,k_12_441,k_12_442,k_12_443,k_12_444,k_12_445,k_12_446,k_12_447,k_12_448,k_12_449,k_12_450,k_12_451,k_12_452,k_12_453,k_12_454,k_12_455,k_12_456,k_12_457,k_12_458,k_12_459,k_12_460,k_12_461,k_12_462,k_12_463,k_12_464,k_12_465,k_12_466,k_12_467,k_12_468,k_12_469,k_12_470,k_12_471,k_12_472,k_12_473,k_12_474,k_12_475,k_12_476,k_12_477,k_12_478,k_12_479,k_12_480,k_12_481,k_12_482,k_12_483,k_12_484,k_12_485,k_12_486,k_12_487,k_12_488,k_12_489,k_12_490,k_12_491,k_12_492,k_12_493,k_12_494,k_12_495,k_12_496,k_12_497,k_12_498,k_12_499,k_12_500,k_12_501,k_12_502,k_12_503,k_12_504,k_12_505,k_12_506,k_12_507,k_12_508,k_12_509,k_12_510,k_12_511,k_12_512,k_12_513,k_12_514,k_12_515,k_12_516,k_12_517,k_12_518,k_12_519,k_12_520,k_12_521,k_12_522,k_12_523,k_12_524,k_12_525,k_12_526,k_12_527,k_12_528,k_12_529,k_12_530,k_12_531,k_12_532,k_12_533,k_12_534,k_12_535,k_12_536,k_12_537,k_12_538,k_12_539,k_12_540,k_12_541,k_12_542,k_12_543,k_12_544,k_12_545,k_12_546,k_12_547,k_12_548,k_12_549,k_12_550,k_12_551,k_12_552,k_12_553,k_12_554,k_12_555,k_12_556,k_12_557,k_12_558,k_12_559,k_12_560,k_12_561,k_12_562,k_12_563,k_12_564,k_12_565,k_12_566,k_12_567,k_12_568,k_12_569,k_12_570,k_12_571,k_12_572,k_12_573,k_12_574,k_12_575,k_12_576,k_12_577,k_12_578,k_12_579,k_12_580,k_12_581,k_12_582,k_12_583,k_12_584,k_12_585,k_12_586,k_12_587,k_12_588,k_12_589,k_12_590,k_12_591,k_12_592,k_12_593,k_12_594,k_12_595,k_12_596,k_12_597,k_12_598,k_12_599,k_12_600,k_12_601,k_12_602,k_12_603,k_12_604,k_12_605,k_12_606,k_12_607,k_12_608,k_12_609,k_12_610,k_12_611,k_12_612,k_12_613,k_12_614,k_12_615,k_12_616,k_12_617,k_12_618,k_12_619,k_12_620,k_12_621,k_12_622,k_12_623,k_12_624,k_12_625,k_12_626,k_12_627,k_12_628,k_12_629,k_12_630,k_12_631,k_12_632,k_12_633,k_12_634,k_12_635,k_12_636,k_12_637,k_12_638,k_12_639,k_12_640,k_12_641,k_12_642,k_12_643,k_12_644,k_12_645,k_12_646,k_12_647,k_12_648,k_12_649,k_12_650,k_12_651,k_12_652,k_12_653,k_12_654,k_12_655,k_12_656,k_12_657,k_12_658,k_12_659,k_12_660,k_12_661,k_12_662,k_12_663,k_12_664,k_12_665,k_12_666,k_12_667,k_12_668,k_12_669,k_12_670,k_12_671,k_12_672,k_12_673,k_12_674,k_12_675,k_12_676,k_12_677,k_12_678,k_12_679,k_12_680,k_12_681,k_12_682,k_12_683,k_12_684,k_12_685,k_12_686,k_12_687,k_12_688,k_12_689,k_12_690,k_12_691,k_12_692,k_12_693,k_12_694,k_12_695,k_12_696,k_12_697,k_12_698,k_12_699,k_12_700,k_12_701,k_12_702,k_12_703,k_12_704,k_12_705,k_12_706,k_12_707,k_12_708,k_12_709,k_12_710,k_12_711,k_12_712,k_12_713,k_12_714,k_12_715,k_12_716,k_12_717,k_12_718,k_12_719,k_12_720,k_12_721,k_12_722,k_12_723,k_12_724,k_12_725,k_12_726,k_12_727,k_12_728,k_12_729,k_12_730,k_12_731,k_12_732,k_12_733,k_12_734,k_12_735,k_12_736,k_12_737,k_12_738,k_12_739,k_12_740,k_12_741,k_12_742,k_12_743,k_12_744,k_12_745,k_12_746,k_12_747,k_12_748,k_12_749,k_12_750,k_12_751,k_12_752,k_12_753,k_12_754,k_12_755,k_12_756,k_12_757,k_12_758,k_12_759,k_12_760,k_12_761,k_12_762,k_12_763,k_12_764,k_12_765,k_12_766,k_12_767,k_12_768,k_12_769,k_12_770,k_12_771,k_12_772,k_12_773,k_12_774,k_12_775,k_12_776,k_12_777,k_12_778,k_12_779,k_12_780,k_12_781,k_12_782,k_12_783,k_12_784,k_12_785,k_12_786,k_12_787,k_12_788,k_12_789,k_12_790,k_12_791,k_12_792,k_12_793,k_12_794,k_12_795,k_12_796,k_12_797,k_12_798,k_12_799,k_12_800,k_12_801,k_12_802,k_12_803,k_12_804,k_12_805,k_12_806,k_12_807,k_12_808,k_12_809,k_12_810,k_12_811,k_12_812,k_12_813,k_12_814,k_12_815,k_12_816,k_12_817,k_12_818,k_12_819,k_12_820,k_12_821,k_12_822,k_12_823,k_12_824,k_12_825,k_12_826,k_12_827,k_12_828,k_12_829,k_12_830,k_12_831,k_12_832,k_12_833,k_12_834,k_12_835,k_12_836,k_12_837,k_12_838,k_12_839,k_12_840,k_12_841,k_12_842,k_12_843,k_12_844,k_12_845,k_12_846,k_12_847,k_12_848,k_12_849,k_12_850,k_12_851,k_12_852,k_12_853,k_12_854,k_12_855,k_12_856,k_12_857,k_12_858,k_12_859,k_12_860,k_12_861,k_12_862,k_12_863,k_12_864,k_12_865,k_12_866,k_12_867,k_12_868,k_12_869,k_12_870,k_12_871,k_12_872,k_12_873,k_12_874,k_12_875,k_12_876,k_12_877,k_12_878,k_12_879,k_12_880,k_12_881,k_12_882,k_12_883,k_12_884,k_12_885,k_12_886,k_12_887,k_12_888,k_12_889,k_12_890,k_12_891,k_12_892,k_12_893,k_12_894,k_12_895,k_12_896,k_12_897,k_12_898,k_12_899,k_12_900,k_12_901,k_12_902,k_12_903,k_12_904,k_12_905,k_12_906,k_12_907,k_12_908,k_12_909,k_12_910,k_12_911,k_12_912,k_12_913,k_12_914,k_12_915,k_12_916,k_12_917,k_12_918,k_12_919,k_12_920,k_12_921,k_12_922,k_12_923,k_12_924,k_12_925,k_12_926,k_12_927,k_12_928,k_12_929,k_12_930,k_12_931,k_12_932,k_12_933,k_12_934,k_12_935,k_12_936,k_12_937,k_12_938,k_12_939,k_12_940,k_12_941,k_12_942,k_12_943,k_12_944,k_12_945,k_12_946,k_12_947,k_12_948,k_12_949,k_12_950,k_12_951,k_12_952,k_12_953,k_12_954,k_12_955,k_12_956,k_12_957,k_12_958,k_12_959,k_12_960,k_12_961,k_12_962,k_12_963,k_12_964,k_12_965,k_12_966,k_12_967,k_12_968,k_12_969,k_12_970,k_12_971,k_12_972,k_12_973,k_12_974,k_12_975,k_12_976,k_12_977,k_12_978,k_12_979,k_12_980,k_12_981,k_12_982,k_12_983,k_12_984,k_12_985,k_12_986,k_12_987,k_12_988,k_12_989,k_12_990,k_12_991,k_12_992,k_12_993,k_12_994,k_12_995,k_12_996,k_12_997,k_12_998,k_12_999,k_12_1000,k_12_1001,k_12_1002,k_12_1003,k_12_1004,k_12_1005,k_12_1006,k_12_1007,k_12_1008,k_12_1009,k_12_1010,k_12_1011,k_12_1012,k_12_1013,k_12_1014,k_12_1015,k_12_1016,k_12_1017,k_12_1018,k_12_1019,k_12_1020,k_12_1021,k_12_1022,k_12_1023,k_12_1024,k_12_1025,k_12_1026,k_12_1027,k_12_1028,k_12_1029,k_12_1030,k_12_1031,k_12_1032,k_12_1033,k_12_1034,k_12_1035,k_12_1036,k_12_1037,k_12_1038,k_12_1039,k_12_1040,k_12_1041,k_12_1042,k_12_1043,k_12_1044,k_12_1045,k_12_1046,k_12_1047,k_12_1048,k_12_1049,k_12_1050,k_12_1051,k_12_1052,k_12_1053,k_12_1054,k_12_1055,k_12_1056,k_12_1057,k_12_1058,k_12_1059,k_12_1060,k_12_1061,k_12_1062,k_12_1063,k_12_1064,k_12_1065,k_12_1066,k_12_1067,k_12_1068,k_12_1069,k_12_1070,k_12_1071,k_12_1072,k_12_1073,k_12_1074,k_12_1075,k_12_1076,k_12_1077,k_12_1078,k_12_1079,k_12_1080,k_12_1081,k_12_1082,k_12_1083,k_12_1084,k_12_1085,k_12_1086,k_12_1087,k_12_1088,k_12_1089,k_12_1090,k_12_1091,k_12_1092,k_12_1093,k_12_1094,k_12_1095,k_12_1096,k_12_1097,k_12_1098,k_12_1099,k_12_1100,k_12_1101,k_12_1102,k_12_1103,k_12_1104,k_12_1105,k_12_1106,k_12_1107,k_12_1108,k_12_1109,k_12_1110,k_12_1111,k_12_1112,k_12_1113,k_12_1114,k_12_1115,k_12_1116,k_12_1117,k_12_1118,k_12_1119,k_12_1120,k_12_1121,k_12_1122,k_12_1123,k_12_1124,k_12_1125,k_12_1126,k_12_1127,k_12_1128,k_12_1129,k_12_1130,k_12_1131,k_12_1132,k_12_1133,k_12_1134,k_12_1135,k_12_1136,k_12_1137,k_12_1138,k_12_1139,k_12_1140,k_12_1141,k_12_1142,k_12_1143,k_12_1144,k_12_1145,k_12_1146,k_12_1147,k_12_1148,k_12_1149,k_12_1150,k_12_1151,k_12_1152,k_12_1153,k_12_1154,k_12_1155,k_12_1156,k_12_1157,k_12_1158,k_12_1159,k_12_1160,k_12_1161,k_12_1162,k_12_1163,k_12_1164,k_12_1165,k_12_1166,k_12_1167,k_12_1168,k_12_1169,k_12_1170,k_12_1171,k_12_1172,k_12_1173,k_12_1174,k_12_1175,k_12_1176,k_12_1177,k_12_1178,k_12_1179,k_12_1180,k_12_1181,k_12_1182,k_12_1183,k_12_1184,k_12_1185,k_12_1186,k_12_1187,k_12_1188,k_12_1189,k_12_1190,k_12_1191,k_12_1192,k_12_1193,k_12_1194,k_12_1195,k_12_1196,k_12_1197,k_12_1198,k_12_1199,k_12_1200,k_12_1201,k_12_1202,k_12_1203,k_12_1204,k_12_1205,k_12_1206,k_12_1207,k_12_1208,k_12_1209,k_12_1210,k_12_1211,k_12_1212,k_12_1213,k_12_1214,k_12_1215,k_12_1216,k_12_1217,k_12_1218,k_12_1219,k_12_1220,k_12_1221,k_12_1222,k_12_1223,k_12_1224,k_12_1225,k_12_1226,k_12_1227,k_12_1228,k_12_1229,k_12_1230,k_12_1231,k_12_1232,k_12_1233,k_12_1234,k_12_1235,k_12_1236,k_12_1237,k_12_1238,k_12_1239,k_12_1240,k_12_1241,k_12_1242,k_12_1243,k_12_1244,k_12_1245,k_12_1246,k_12_1247,k_12_1248,k_12_1249,k_12_1250,k_12_1251,k_12_1252,k_12_1253,k_12_1254,k_12_1255,k_12_1256,k_12_1257,k_12_1258,k_12_1259,k_12_1260,k_12_1261,k_12_1262,k_12_1263,k_12_1264,k_12_1265,k_12_1266,k_12_1267,k_12_1268,k_12_1269,k_12_1270,k_12_1271,k_12_1272,k_12_1273,k_12_1274,k_12_1275,k_12_1276,k_12_1277,k_12_1278,k_12_1279,k_12_1280,k_12_1281,k_12_1282,k_12_1283,k_12_1284,k_12_1285,k_12_1286,k_12_1287,k_12_1288,k_12_1289,k_12_1290,k_12_1291,k_12_1292,k_12_1293,k_12_1294,k_12_1295,k_12_1296,k_12_1297,k_12_1298,k_12_1299,k_12_1300,k_12_1301,k_12_1302,k_12_1303,k_12_1304,k_12_1305,k_12_1306,k_12_1307,k_12_1308,k_12_1309,k_12_1310,k_12_1311,k_12_1312,k_12_1313,k_12_1314,k_12_1315,k_12_1316,k_12_1317,k_12_1318,k_12_1319,k_12_1320,k_12_1321,k_12_1322,k_12_1323,k_12_1324,k_12_1325,k_12_1326,k_12_1327,k_12_1328,k_12_1329,k_12_1330,k_12_1331,k_12_1332,k_12_1333,k_12_1334,k_12_1335,k_12_1336,k_12_1337,k_12_1338,k_12_1339,k_12_1340,k_12_1341,k_12_1342,k_12_1343,k_12_1344,k_12_1345,k_12_1346,k_12_1347,k_12_1348,k_12_1349,k_12_1350,k_12_1351,k_12_1352,k_12_1353,k_12_1354,k_12_1355,k_12_1356,k_12_1357,k_12_1358,k_12_1359,k_12_1360,k_12_1361,k_12_1362,k_12_1363,k_12_1364,k_12_1365,k_12_1366,k_12_1367,k_12_1368,k_12_1369,k_12_1370,k_12_1371,k_12_1372,k_12_1373,k_12_1374,k_12_1375,k_12_1376,k_12_1377,k_12_1378,k_12_1379,k_12_1380,k_12_1381,k_12_1382,k_12_1383,k_12_1384,k_12_1385,k_12_1386,k_12_1387,k_12_1388,k_12_1389,k_12_1390,k_12_1391,k_12_1392,k_12_1393,k_12_1394,k_12_1395,k_12_1396,k_12_1397,k_12_1398,k_12_1399,k_12_1400,k_12_1401,k_12_1402,k_12_1403,k_12_1404,k_12_1405,k_12_1406,k_12_1407,k_12_1408,k_12_1409,k_12_1410,k_12_1411,k_12_1412,k_12_1413,k_12_1414,k_12_1415,k_12_1416,k_12_1417,k_12_1418,k_12_1419,k_12_1420,k_12_1421,k_12_1422,k_12_1423,k_12_1424,k_12_1425,k_12_1426,k_12_1427,k_12_1428,k_12_1429,k_12_1430,k_12_1431,k_12_1432,k_12_1433,k_12_1434,k_12_1435,k_12_1436,k_12_1437,k_12_1438,k_12_1439,k_12_1440,k_12_1441,k_12_1442,k_12_1443,k_12_1444,k_12_1445,k_12_1446,k_12_1447,k_12_1448,k_12_1449,k_12_1450,k_12_1451,k_12_1452,k_12_1453,k_12_1454,k_12_1455,k_12_1456,k_12_1457,k_12_1458,k_12_1459,k_12_1460,k_12_1461,k_12_1462,k_12_1463,k_12_1464,k_12_1465,k_12_1466,k_12_1467,k_12_1468,k_12_1469,k_12_1470,k_12_1471,k_12_1472,k_12_1473,k_12_1474,k_12_1475,k_12_1476,k_12_1477,k_12_1478,k_12_1479,k_12_1480,k_12_1481,k_12_1482,k_12_1483,k_12_1484,k_12_1485,k_12_1486,k_12_1487,k_12_1488,k_12_1489,k_12_1490,k_12_1491,k_12_1492,k_12_1493,k_12_1494,k_12_1495,k_12_1496,k_12_1497,k_12_1498,k_12_1499,k_12_1500,k_12_1501,k_12_1502,k_12_1503,k_12_1504,k_12_1505,k_12_1506,k_12_1507,k_12_1508,k_12_1509,k_12_1510,k_12_1511,k_12_1512,k_12_1513,k_12_1514,k_12_1515,k_12_1516,k_12_1517,k_12_1518,k_12_1519,k_12_1520,k_12_1521,k_12_1522,k_12_1523,k_12_1524,k_12_1525,k_12_1526,k_12_1527,k_12_1528,k_12_1529,k_12_1530,k_12_1531,k_12_1532,k_12_1533,k_12_1534,k_12_1535,k_12_1536,k_12_1537,k_12_1538,k_12_1539,k_12_1540,k_12_1541,k_12_1542,k_12_1543,k_12_1544,k_12_1545,k_12_1546,k_12_1547,k_12_1548,k_12_1549,k_12_1550,k_12_1551,k_12_1552,k_12_1553,k_12_1554,k_12_1555,k_12_1556,k_12_1557,k_12_1558,k_12_1559,k_12_1560,k_12_1561,k_12_1562,k_12_1563,k_12_1564,k_12_1565,k_12_1566,k_12_1567,k_12_1568,k_12_1569,k_12_1570,k_12_1571,k_12_1572,k_12_1573,k_12_1574,k_12_1575,k_12_1576,k_12_1577,k_12_1578,k_12_1579,k_12_1580,k_12_1581,k_12_1582,k_12_1583,k_12_1584,k_12_1585,k_12_1586,k_12_1587,k_12_1588,k_12_1589,k_12_1590,k_12_1591,k_12_1592,k_12_1593,k_12_1594,k_12_1595,k_12_1596,k_12_1597,k_12_1598,k_12_1599,k_12_1600,k_12_1601,k_12_1602,k_12_1603,k_12_1604,k_12_1605,k_12_1606,k_12_1607,k_12_1608,k_12_1609,k_12_1610,k_12_1611,k_12_1612,k_12_1613,k_12_1614,k_12_1615,k_12_1616,k_12_1617,k_12_1618,k_12_1619,k_12_1620,k_12_1621,k_12_1622,k_12_1623,k_12_1624,k_12_1625,k_12_1626,k_12_1627,k_12_1628,k_12_1629,k_12_1630,k_12_1631,k_12_1632,k_12_1633,k_12_1634,k_12_1635,k_12_1636,k_12_1637,k_12_1638,k_12_1639,k_12_1640,k_12_1641,k_12_1642,k_12_1643,k_12_1644,k_12_1645,k_12_1646,k_12_1647,k_12_1648,k_12_1649,k_12_1650,k_12_1651,k_12_1652,k_12_1653,k_12_1654,k_12_1655,k_12_1656,k_12_1657,k_12_1658,k_12_1659,k_12_1660,k_12_1661,k_12_1662,k_12_1663,k_12_1664,k_12_1665,k_12_1666,k_12_1667,k_12_1668,k_12_1669,k_12_1670,k_12_1671,k_12_1672,k_12_1673,k_12_1674,k_12_1675,k_12_1676,k_12_1677,k_12_1678,k_12_1679,k_12_1680,k_12_1681,k_12_1682,k_12_1683,k_12_1684,k_12_1685,k_12_1686,k_12_1687,k_12_1688,k_12_1689,k_12_1690,k_12_1691,k_12_1692,k_12_1693,k_12_1694,k_12_1695,k_12_1696,k_12_1697,k_12_1698,k_12_1699,k_12_1700,k_12_1701,k_12_1702,k_12_1703,k_12_1704,k_12_1705,k_12_1706,k_12_1707,k_12_1708,k_12_1709,k_12_1710,k_12_1711,k_12_1712,k_12_1713,k_12_1714,k_12_1715,k_12_1716,k_12_1717,k_12_1718,k_12_1719,k_12_1720,k_12_1721,k_12_1722,k_12_1723,k_12_1724,k_12_1725,k_12_1726,k_12_1727,k_12_1728,k_12_1729,k_12_1730,k_12_1731,k_12_1732,k_12_1733,k_12_1734,k_12_1735,k_12_1736,k_12_1737,k_12_1738,k_12_1739,k_12_1740,k_12_1741,k_12_1742,k_12_1743,k_12_1744,k_12_1745,k_12_1746,k_12_1747,k_12_1748,k_12_1749,k_12_1750,k_12_1751,k_12_1752,k_12_1753,k_12_1754,k_12_1755,k_12_1756,k_12_1757,k_12_1758,k_12_1759,k_12_1760,k_12_1761,k_12_1762,k_12_1763,k_12_1764,k_12_1765,k_12_1766,k_12_1767,k_12_1768,k_12_1769,k_12_1770,k_12_1771,k_12_1772,k_12_1773,k_12_1774,k_12_1775,k_12_1776,k_12_1777,k_12_1778,k_12_1779,k_12_1780,k_12_1781,k_12_1782,k_12_1783,k_12_1784,k_12_1785,k_12_1786,k_12_1787,k_12_1788,k_12_1789,k_12_1790,k_12_1791,k_12_1792,k_12_1793,k_12_1794,k_12_1795,k_12_1796,k_12_1797,k_12_1798,k_12_1799,k_12_1800,k_12_1801,k_12_1802,k_12_1803,k_12_1804,k_12_1805,k_12_1806,k_12_1807,k_12_1808,k_12_1809,k_12_1810,k_12_1811,k_12_1812,k_12_1813,k_12_1814,k_12_1815,k_12_1816,k_12_1817,k_12_1818,k_12_1819,k_12_1820,k_12_1821,k_12_1822,k_12_1823,k_12_1824,k_12_1825,k_12_1826,k_12_1827,k_12_1828,k_12_1829,k_12_1830,k_12_1831,k_12_1832,k_12_1833,k_12_1834,k_12_1835,k_12_1836,k_12_1837,k_12_1838,k_12_1839,k_12_1840,k_12_1841,k_12_1842,k_12_1843,k_12_1844,k_12_1845,k_12_1846,k_12_1847,k_12_1848,k_12_1849,k_12_1850,k_12_1851,k_12_1852,k_12_1853,k_12_1854,k_12_1855,k_12_1856,k_12_1857,k_12_1858,k_12_1859,k_12_1860,k_12_1861,k_12_1862,k_12_1863,k_12_1864,k_12_1865,k_12_1866,k_12_1867,k_12_1868,k_12_1869,k_12_1870,k_12_1871,k_12_1872,k_12_1873,k_12_1874,k_12_1875,k_12_1876,k_12_1877,k_12_1878,k_12_1879,k_12_1880,k_12_1881,k_12_1882,k_12_1883,k_12_1884,k_12_1885,k_12_1886,k_12_1887,k_12_1888,k_12_1889,k_12_1890,k_12_1891,k_12_1892,k_12_1893,k_12_1894,k_12_1895,k_12_1896,k_12_1897,k_12_1898,k_12_1899,k_12_1900,k_12_1901,k_12_1902,k_12_1903,k_12_1904,k_12_1905,k_12_1906,k_12_1907,k_12_1908,k_12_1909,k_12_1910,k_12_1911,k_12_1912,k_12_1913,k_12_1914,k_12_1915,k_12_1916,k_12_1917,k_12_1918,k_12_1919,k_12_1920,k_12_1921,k_12_1922,k_12_1923,k_12_1924,k_12_1925,k_12_1926,k_12_1927,k_12_1928,k_12_1929,k_12_1930,k_12_1931,k_12_1932,k_12_1933,k_12_1934,k_12_1935,k_12_1936,k_12_1937,k_12_1938,k_12_1939,k_12_1940,k_12_1941,k_12_1942,k_12_1943,k_12_1944,k_12_1945,k_12_1946,k_12_1947,k_12_1948,k_12_1949,k_12_1950,k_12_1951,k_12_1952,k_12_1953,k_12_1954,k_12_1955,k_12_1956,k_12_1957,k_12_1958,k_12_1959,k_12_1960,k_12_1961,k_12_1962,k_12_1963,k_12_1964,k_12_1965,k_12_1966,k_12_1967,k_12_1968,k_12_1969,k_12_1970,k_12_1971,k_12_1972,k_12_1973,k_12_1974,k_12_1975,k_12_1976,k_12_1977,k_12_1978,k_12_1979,k_12_1980,k_12_1981,k_12_1982,k_12_1983,k_12_1984,k_12_1985,k_12_1986,k_12_1987,k_12_1988,k_12_1989,k_12_1990,k_12_1991,k_12_1992,k_12_1993,k_12_1994,k_12_1995,k_12_1996,k_12_1997,k_12_1998,k_12_1999,k_12_2000,k_12_2001,k_12_2002,k_12_2003,k_12_2004,k_12_2005,k_12_2006,k_12_2007,k_12_2008,k_12_2009,k_12_2010,k_12_2011,k_12_2012,k_12_2013,k_12_2014,k_12_2015,k_12_2016,k_12_2017,k_12_2018,k_12_2019,k_12_2020,k_12_2021,k_12_2022,k_12_2023,k_12_2024,k_12_2025,k_12_2026,k_12_2027,k_12_2028,k_12_2029,k_12_2030,k_12_2031,k_12_2032,k_12_2033,k_12_2034,k_12_2035,k_12_2036,k_12_2037,k_12_2038,k_12_2039,k_12_2040,k_12_2041,k_12_2042,k_12_2043,k_12_2044,k_12_2045,k_12_2046,k_12_2047,k_12_2048,k_12_2049,k_12_2050,k_12_2051,k_12_2052,k_12_2053,k_12_2054,k_12_2055,k_12_2056,k_12_2057,k_12_2058,k_12_2059,k_12_2060,k_12_2061,k_12_2062,k_12_2063,k_12_2064,k_12_2065,k_12_2066,k_12_2067,k_12_2068,k_12_2069,k_12_2070,k_12_2071,k_12_2072,k_12_2073,k_12_2074,k_12_2075,k_12_2076,k_12_2077,k_12_2078,k_12_2079,k_12_2080,k_12_2081,k_12_2082,k_12_2083,k_12_2084,k_12_2085,k_12_2086,k_12_2087,k_12_2088,k_12_2089,k_12_2090,k_12_2091,k_12_2092,k_12_2093,k_12_2094,k_12_2095,k_12_2096,k_12_2097,k_12_2098,k_12_2099,k_12_2100,k_12_2101,k_12_2102,k_12_2103,k_12_2104,k_12_2105,k_12_2106,k_12_2107,k_12_2108,k_12_2109,k_12_2110,k_12_2111,k_12_2112,k_12_2113,k_12_2114,k_12_2115,k_12_2116,k_12_2117,k_12_2118,k_12_2119,k_12_2120,k_12_2121,k_12_2122,k_12_2123,k_12_2124,k_12_2125,k_12_2126,k_12_2127,k_12_2128,k_12_2129,k_12_2130,k_12_2131,k_12_2132,k_12_2133,k_12_2134,k_12_2135,k_12_2136,k_12_2137,k_12_2138,k_12_2139,k_12_2140,k_12_2141,k_12_2142,k_12_2143,k_12_2144,k_12_2145,k_12_2146,k_12_2147,k_12_2148,k_12_2149,k_12_2150,k_12_2151,k_12_2152,k_12_2153,k_12_2154,k_12_2155,k_12_2156,k_12_2157,k_12_2158,k_12_2159,k_12_2160,k_12_2161,k_12_2162,k_12_2163,k_12_2164,k_12_2165,k_12_2166,k_12_2167,k_12_2168,k_12_2169,k_12_2170,k_12_2171,k_12_2172,k_12_2173,k_12_2174,k_12_2175,k_12_2176,k_12_2177,k_12_2178,k_12_2179,k_12_2180,k_12_2181,k_12_2182,k_12_2183,k_12_2184,k_12_2185,k_12_2186,k_12_2187,k_12_2188,k_12_2189,k_12_2190,k_12_2191,k_12_2192,k_12_2193,k_12_2194,k_12_2195,k_12_2196,k_12_2197,k_12_2198,k_12_2199,k_12_2200,k_12_2201,k_12_2202,k_12_2203,k_12_2204,k_12_2205,k_12_2206,k_12_2207,k_12_2208,k_12_2209,k_12_2210,k_12_2211,k_12_2212,k_12_2213,k_12_2214,k_12_2215,k_12_2216,k_12_2217,k_12_2218,k_12_2219,k_12_2220,k_12_2221,k_12_2222,k_12_2223,k_12_2224,k_12_2225,k_12_2226,k_12_2227,k_12_2228,k_12_2229,k_12_2230,k_12_2231,k_12_2232,k_12_2233,k_12_2234,k_12_2235,k_12_2236,k_12_2237,k_12_2238,k_12_2239,k_12_2240,k_12_2241,k_12_2242,k_12_2243,k_12_2244,k_12_2245,k_12_2246,k_12_2247,k_12_2248,k_12_2249,k_12_2250,k_12_2251,k_12_2252,k_12_2253,k_12_2254,k_12_2255,k_12_2256,k_12_2257,k_12_2258,k_12_2259,k_12_2260,k_12_2261,k_12_2262,k_12_2263,k_12_2264,k_12_2265,k_12_2266,k_12_2267,k_12_2268,k_12_2269,k_12_2270,k_12_2271,k_12_2272,k_12_2273,k_12_2274,k_12_2275,k_12_2276,k_12_2277,k_12_2278,k_12_2279,k_12_2280,k_12_2281,k_12_2282,k_12_2283,k_12_2284,k_12_2285,k_12_2286,k_12_2287,k_12_2288,k_12_2289,k_12_2290,k_12_2291,k_12_2292,k_12_2293,k_12_2294,k_12_2295,k_12_2296,k_12_2297,k_12_2298,k_12_2299,k_12_2300,k_12_2301,k_12_2302,k_12_2303,k_12_2304,k_12_2305,k_12_2306,k_12_2307,k_12_2308,k_12_2309,k_12_2310,k_12_2311,k_12_2312,k_12_2313,k_12_2314,k_12_2315,k_12_2316,k_12_2317,k_12_2318,k_12_2319,k_12_2320,k_12_2321,k_12_2322,k_12_2323,k_12_2324,k_12_2325,k_12_2326,k_12_2327,k_12_2328,k_12_2329,k_12_2330,k_12_2331,k_12_2332,k_12_2333,k_12_2334,k_12_2335,k_12_2336,k_12_2337,k_12_2338,k_12_2339,k_12_2340,k_12_2341,k_12_2342,k_12_2343,k_12_2344,k_12_2345,k_12_2346,k_12_2347,k_12_2348,k_12_2349,k_12_2350,k_12_2351,k_12_2352,k_12_2353,k_12_2354,k_12_2355,k_12_2356,k_12_2357,k_12_2358,k_12_2359,k_12_2360,k_12_2361,k_12_2362,k_12_2363,k_12_2364,k_12_2365,k_12_2366,k_12_2367,k_12_2368,k_12_2369,k_12_2370,k_12_2371,k_12_2372,k_12_2373,k_12_2374,k_12_2375,k_12_2376,k_12_2377,k_12_2378,k_12_2379,k_12_2380,k_12_2381,k_12_2382,k_12_2383,k_12_2384,k_12_2385,k_12_2386,k_12_2387,k_12_2388,k_12_2389,k_12_2390,k_12_2391,k_12_2392,k_12_2393,k_12_2394,k_12_2395,k_12_2396,k_12_2397,k_12_2398,k_12_2399,k_12_2400,k_12_2401,k_12_2402,k_12_2403,k_12_2404,k_12_2405,k_12_2406,k_12_2407,k_12_2408,k_12_2409,k_12_2410,k_12_2411,k_12_2412,k_12_2413,k_12_2414,k_12_2415,k_12_2416,k_12_2417,k_12_2418,k_12_2419,k_12_2420,k_12_2421,k_12_2422,k_12_2423,k_12_2424,k_12_2425,k_12_2426,k_12_2427,k_12_2428,k_12_2429,k_12_2430,k_12_2431,k_12_2432,k_12_2433,k_12_2434,k_12_2435,k_12_2436,k_12_2437,k_12_2438,k_12_2439,k_12_2440,k_12_2441,k_12_2442,k_12_2443,k_12_2444,k_12_2445,k_12_2446,k_12_2447,k_12_2448,k_12_2449,k_12_2450,k_12_2451,k_12_2452,k_12_2453,k_12_2454,k_12_2455,k_12_2456,k_12_2457,k_12_2458,k_12_2459,k_12_2460,k_12_2461,k_12_2462,k_12_2463,k_12_2464,k_12_2465,k_12_2466,k_12_2467,k_12_2468,k_12_2469,k_12_2470,k_12_2471,k_12_2472,k_12_2473,k_12_2474,k_12_2475,k_12_2476,k_12_2477,k_12_2478,k_12_2479,k_12_2480,k_12_2481,k_12_2482,k_12_2483,k_12_2484,k_12_2485,k_12_2486,k_12_2487,k_12_2488,k_12_2489,k_12_2490,k_12_2491,k_12_2492,k_12_2493,k_12_2494,k_12_2495,k_12_2496,k_12_2497,k_12_2498,k_12_2499,k_12_2500,k_12_2501,k_12_2502,k_12_2503,k_12_2504,k_12_2505,k_12_2506,k_12_2507,k_12_2508,k_12_2509,k_12_2510,k_12_2511,k_12_2512,k_12_2513,k_12_2514,k_12_2515,k_12_2516,k_12_2517,k_12_2518,k_12_2519,k_12_2520,k_12_2521,k_12_2522,k_12_2523,k_12_2524,k_12_2525,k_12_2526,k_12_2527,k_12_2528,k_12_2529,k_12_2530,k_12_2531,k_12_2532,k_12_2533,k_12_2534,k_12_2535,k_12_2536,k_12_2537,k_12_2538,k_12_2539,k_12_2540,k_12_2541,k_12_2542,k_12_2543,k_12_2544,k_12_2545,k_12_2546,k_12_2547,k_12_2548,k_12_2549,k_12_2550,k_12_2551,k_12_2552,k_12_2553,k_12_2554,k_12_2555,k_12_2556,k_12_2557,k_12_2558,k_12_2559,k_12_2560,k_12_2561,k_12_2562,k_12_2563,k_12_2564,k_12_2565,k_12_2566,k_12_2567,k_12_2568,k_12_2569,k_12_2570,k_12_2571,k_12_2572,k_12_2573,k_12_2574,k_12_2575,k_12_2576,k_12_2577,k_12_2578,k_12_2579,k_12_2580,k_12_2581,k_12_2582,k_12_2583,k_12_2584,k_12_2585,k_12_2586,k_12_2587,k_12_2588,k_12_2589,k_12_2590,k_12_2591,k_12_2592,k_12_2593,k_12_2594,k_12_2595,k_12_2596,k_12_2597,k_12_2598,k_12_2599,k_12_2600,k_12_2601,k_12_2602,k_12_2603,k_12_2604,k_12_2605,k_12_2606,k_12_2607,k_12_2608,k_12_2609,k_12_2610,k_12_2611,k_12_2612,k_12_2613,k_12_2614,k_12_2615,k_12_2616,k_12_2617,k_12_2618,k_12_2619,k_12_2620,k_12_2621,k_12_2622,k_12_2623,k_12_2624,k_12_2625,k_12_2626,k_12_2627,k_12_2628,k_12_2629,k_12_2630,k_12_2631,k_12_2632,k_12_2633,k_12_2634,k_12_2635,k_12_2636,k_12_2637,k_12_2638,k_12_2639,k_12_2640,k_12_2641,k_12_2642,k_12_2643,k_12_2644,k_12_2645,k_12_2646,k_12_2647,k_12_2648,k_12_2649,k_12_2650,k_12_2651,k_12_2652,k_12_2653,k_12_2654,k_12_2655,k_12_2656,k_12_2657,k_12_2658,k_12_2659,k_12_2660,k_12_2661,k_12_2662,k_12_2663,k_12_2664,k_12_2665,k_12_2666,k_12_2667,k_12_2668,k_12_2669,k_12_2670,k_12_2671,k_12_2672,k_12_2673,k_12_2674,k_12_2675,k_12_2676,k_12_2677,k_12_2678,k_12_2679,k_12_2680,k_12_2681,k_12_2682,k_12_2683,k_12_2684,k_12_2685,k_12_2686,k_12_2687,k_12_2688,k_12_2689,k_12_2690,k_12_2691,k_12_2692,k_12_2693,k_12_2694,k_12_2695,k_12_2696,k_12_2697,k_12_2698,k_12_2699,k_12_2700,k_12_2701,k_12_2702,k_12_2703,k_12_2704,k_12_2705,k_12_2706,k_12_2707,k_12_2708,k_12_2709,k_12_2710,k_12_2711,k_12_2712,k_12_2713,k_12_2714,k_12_2715,k_12_2716,k_12_2717,k_12_2718,k_12_2719,k_12_2720,k_12_2721,k_12_2722,k_12_2723,k_12_2724,k_12_2725,k_12_2726,k_12_2727,k_12_2728,k_12_2729,k_12_2730,k_12_2731,k_12_2732,k_12_2733,k_12_2734,k_12_2735,k_12_2736,k_12_2737,k_12_2738,k_12_2739,k_12_2740,k_12_2741,k_12_2742,k_12_2743,k_12_2744,k_12_2745,k_12_2746,k_12_2747,k_12_2748,k_12_2749,k_12_2750,k_12_2751,k_12_2752,k_12_2753,k_12_2754,k_12_2755,k_12_2756,k_12_2757,k_12_2758,k_12_2759,k_12_2760,k_12_2761,k_12_2762,k_12_2763,k_12_2764,k_12_2765,k_12_2766,k_12_2767,k_12_2768,k_12_2769,k_12_2770,k_12_2771,k_12_2772,k_12_2773,k_12_2774,k_12_2775,k_12_2776,k_12_2777,k_12_2778,k_12_2779,k_12_2780,k_12_2781,k_12_2782,k_12_2783,k_12_2784,k_12_2785,k_12_2786,k_12_2787,k_12_2788,k_12_2789,k_12_2790,k_12_2791,k_12_2792,k_12_2793,k_12_2794,k_12_2795,k_12_2796,k_12_2797,k_12_2798,k_12_2799,k_12_2800,k_12_2801,k_12_2802,k_12_2803,k_12_2804,k_12_2805,k_12_2806,k_12_2807,k_12_2808,k_12_2809,k_12_2810,k_12_2811,k_12_2812,k_12_2813,k_12_2814,k_12_2815,k_12_2816,k_12_2817,k_12_2818,k_12_2819,k_12_2820,k_12_2821,k_12_2822,k_12_2823,k_12_2824,k_12_2825,k_12_2826,k_12_2827,k_12_2828,k_12_2829,k_12_2830,k_12_2831,k_12_2832,k_12_2833,k_12_2834,k_12_2835,k_12_2836,k_12_2837,k_12_2838,k_12_2839,k_12_2840,k_12_2841,k_12_2842,k_12_2843,k_12_2844,k_12_2845,k_12_2846,k_12_2847,k_12_2848,k_12_2849,k_12_2850,k_12_2851,k_12_2852,k_12_2853,k_12_2854,k_12_2855,k_12_2856,k_12_2857,k_12_2858,k_12_2859,k_12_2860,k_12_2861,k_12_2862,k_12_2863,k_12_2864,k_12_2865,k_12_2866,k_12_2867,k_12_2868,k_12_2869,k_12_2870,k_12_2871,k_12_2872,k_12_2873,k_12_2874,k_12_2875,k_12_2876,k_12_2877,k_12_2878,k_12_2879,k_12_2880,k_12_2881,k_12_2882,k_12_2883,k_12_2884,k_12_2885,k_12_2886,k_12_2887,k_12_2888,k_12_2889,k_12_2890,k_12_2891,k_12_2892,k_12_2893,k_12_2894,k_12_2895,k_12_2896,k_12_2897,k_12_2898,k_12_2899,k_12_2900,k_12_2901,k_12_2902,k_12_2903,k_12_2904,k_12_2905,k_12_2906,k_12_2907,k_12_2908,k_12_2909,k_12_2910,k_12_2911,k_12_2912,k_12_2913,k_12_2914,k_12_2915,k_12_2916,k_12_2917,k_12_2918,k_12_2919,k_12_2920,k_12_2921,k_12_2922,k_12_2923,k_12_2924,k_12_2925,k_12_2926,k_12_2927,k_12_2928,k_12_2929,k_12_2930,k_12_2931,k_12_2932,k_12_2933,k_12_2934,k_12_2935,k_12_2936,k_12_2937,k_12_2938,k_12_2939,k_12_2940,k_12_2941,k_12_2942,k_12_2943,k_12_2944,k_12_2945,k_12_2946,k_12_2947,k_12_2948,k_12_2949,k_12_2950,k_12_2951,k_12_2952,k_12_2953,k_12_2954,k_12_2955,k_12_2956,k_12_2957,k_12_2958,k_12_2959,k_12_2960,k_12_2961,k_12_2962,k_12_2963,k_12_2964,k_12_2965,k_12_2966,k_12_2967,k_12_2968,k_12_2969,k_12_2970,k_12_2971,k_12_2972,k_12_2973,k_12_2974,k_12_2975,k_12_2976,k_12_2977,k_12_2978,k_12_2979,k_12_2980,k_12_2981,k_12_2982,k_12_2983,k_12_2984,k_12_2985,k_12_2986,k_12_2987,k_12_2988,k_12_2989,k_12_2990,k_12_2991,k_12_2992,k_12_2993,k_12_2994,k_12_2995,k_12_2996,k_12_2997,k_12_2998,k_12_2999,k_12_3000,k_12_3001,k_12_3002,k_12_3003,k_12_3004,k_12_3005,k_12_3006,k_12_3007,k_12_3008,k_12_3009,k_12_3010,k_12_3011,k_12_3012,k_12_3013,k_12_3014,k_12_3015,k_12_3016,k_12_3017,k_12_3018,k_12_3019,k_12_3020,k_12_3021,k_12_3022,k_12_3023,k_12_3024,k_12_3025,k_12_3026,k_12_3027,k_12_3028,k_12_3029,k_12_3030,k_12_3031,k_12_3032,k_12_3033,k_12_3034,k_12_3035,k_12_3036,k_12_3037,k_12_3038,k_12_3039,k_12_3040,k_12_3041,k_12_3042,k_12_3043,k_12_3044,k_12_3045,k_12_3046,k_12_3047,k_12_3048,k_12_3049,k_12_3050,k_12_3051,k_12_3052,k_12_3053,k_12_3054,k_12_3055,k_12_3056,k_12_3057,k_12_3058,k_12_3059,k_12_3060,k_12_3061,k_12_3062,k_12_3063,k_12_3064,k_12_3065,k_12_3066,k_12_3067,k_12_3068,k_12_3069,k_12_3070,k_12_3071,k_12_3072,k_12_3073,k_12_3074,k_12_3075,k_12_3076,k_12_3077,k_12_3078,k_12_3079,k_12_3080,k_12_3081,k_12_3082,k_12_3083,k_12_3084,k_12_3085,k_12_3086,k_12_3087,k_12_3088,k_12_3089,k_12_3090,k_12_3091,k_12_3092,k_12_3093,k_12_3094,k_12_3095,k_12_3096,k_12_3097,k_12_3098,k_12_3099,k_12_3100,k_12_3101,k_12_3102,k_12_3103,k_12_3104,k_12_3105,k_12_3106,k_12_3107,k_12_3108,k_12_3109,k_12_3110,k_12_3111,k_12_3112,k_12_3113,k_12_3114,k_12_3115,k_12_3116,k_12_3117,k_12_3118,k_12_3119,k_12_3120,k_12_3121,k_12_3122,k_12_3123,k_12_3124,k_12_3125,k_12_3126,k_12_3127,k_12_3128,k_12_3129,k_12_3130,k_12_3131,k_12_3132,k_12_3133,k_12_3134,k_12_3135,k_12_3136,k_12_3137,k_12_3138,k_12_3139,k_12_3140,k_12_3141,k_12_3142,k_12_3143,k_12_3144,k_12_3145,k_12_3146,k_12_3147,k_12_3148,k_12_3149,k_12_3150,k_12_3151,k_12_3152,k_12_3153,k_12_3154,k_12_3155,k_12_3156,k_12_3157,k_12_3158,k_12_3159,k_12_3160,k_12_3161,k_12_3162,k_12_3163,k_12_3164,k_12_3165,k_12_3166,k_12_3167,k_12_3168,k_12_3169,k_12_3170,k_12_3171,k_12_3172,k_12_3173,k_12_3174,k_12_3175,k_12_3176,k_12_3177,k_12_3178,k_12_3179,k_12_3180,k_12_3181,k_12_3182,k_12_3183,k_12_3184,k_12_3185,k_12_3186,k_12_3187,k_12_3188,k_12_3189,k_12_3190,k_12_3191,k_12_3192,k_12_3193,k_12_3194,k_12_3195,k_12_3196,k_12_3197,k_12_3198,k_12_3199,k_12_3200,k_12_3201,k_12_3202,k_12_3203,k_12_3204,k_12_3205,k_12_3206,k_12_3207,k_12_3208,k_12_3209,k_12_3210,k_12_3211,k_12_3212,k_12_3213,k_12_3214,k_12_3215,k_12_3216,k_12_3217,k_12_3218,k_12_3219,k_12_3220,k_12_3221,k_12_3222,k_12_3223,k_12_3224,k_12_3225,k_12_3226,k_12_3227,k_12_3228,k_12_3229,k_12_3230,k_12_3231,k_12_3232,k_12_3233,k_12_3234,k_12_3235,k_12_3236,k_12_3237,k_12_3238,k_12_3239,k_12_3240,k_12_3241,k_12_3242,k_12_3243,k_12_3244,k_12_3245,k_12_3246,k_12_3247,k_12_3248,k_12_3249,k_12_3250,k_12_3251,k_12_3252,k_12_3253,k_12_3254,k_12_3255,k_12_3256,k_12_3257,k_12_3258,k_12_3259,k_12_3260,k_12_3261,k_12_3262,k_12_3263,k_12_3264,k_12_3265,k_12_3266,k_12_3267,k_12_3268,k_12_3269,k_12_3270,k_12_3271,k_12_3272,k_12_3273,k_12_3274,k_12_3275,k_12_3276,k_12_3277,k_12_3278,k_12_3279,k_12_3280,k_12_3281,k_12_3282,k_12_3283,k_12_3284,k_12_3285,k_12_3286,k_12_3287,k_12_3288,k_12_3289,k_12_3290,k_12_3291,k_12_3292,k_12_3293,k_12_3294,k_12_3295,k_12_3296,k_12_3297,k_12_3298,k_12_3299,k_12_3300,k_12_3301,k_12_3302,k_12_3303,k_12_3304,k_12_3305,k_12_3306,k_12_3307,k_12_3308,k_12_3309,k_12_3310,k_12_3311,k_12_3312,k_12_3313,k_12_3314,k_12_3315,k_12_3316,k_12_3317,k_12_3318,k_12_3319,k_12_3320,k_12_3321,k_12_3322,k_12_3323,k_12_3324,k_12_3325,k_12_3326,k_12_3327,k_12_3328,k_12_3329,k_12_3330,k_12_3331,k_12_3332,k_12_3333,k_12_3334,k_12_3335,k_12_3336,k_12_3337,k_12_3338,k_12_3339,k_12_3340,k_12_3341,k_12_3342,k_12_3343,k_12_3344,k_12_3345,k_12_3346,k_12_3347,k_12_3348,k_12_3349,k_12_3350,k_12_3351,k_12_3352,k_12_3353,k_12_3354,k_12_3355,k_12_3356,k_12_3357,k_12_3358,k_12_3359,k_12_3360,k_12_3361,k_12_3362,k_12_3363,k_12_3364,k_12_3365,k_12_3366,k_12_3367,k_12_3368,k_12_3369,k_12_3370,k_12_3371,k_12_3372,k_12_3373,k_12_3374,k_12_3375,k_12_3376,k_12_3377,k_12_3378,k_12_3379,k_12_3380,k_12_3381,k_12_3382,k_12_3383,k_12_3384,k_12_3385,k_12_3386,k_12_3387,k_12_3388,k_12_3389,k_12_3390,k_12_3391,k_12_3392,k_12_3393,k_12_3394,k_12_3395,k_12_3396,k_12_3397,k_12_3398,k_12_3399,k_12_3400,k_12_3401,k_12_3402,k_12_3403,k_12_3404,k_12_3405,k_12_3406,k_12_3407,k_12_3408,k_12_3409,k_12_3410,k_12_3411,k_12_3412,k_12_3413,k_12_3414,k_12_3415,k_12_3416,k_12_3417,k_12_3418,k_12_3419,k_12_3420,k_12_3421,k_12_3422,k_12_3423,k_12_3424,k_12_3425,k_12_3426,k_12_3427,k_12_3428,k_12_3429,k_12_3430,k_12_3431,k_12_3432,k_12_3433,k_12_3434,k_12_3435,k_12_3436,k_12_3437,k_12_3438,k_12_3439,k_12_3440,k_12_3441,k_12_3442,k_12_3443,k_12_3444,k_12_3445,k_12_3446,k_12_3447,k_12_3448,k_12_3449,k_12_3450,k_12_3451,k_12_3452,k_12_3453,k_12_3454,k_12_3455,k_12_3456,k_12_3457,k_12_3458,k_12_3459,k_12_3460,k_12_3461,k_12_3462,k_12_3463,k_12_3464,k_12_3465,k_12_3466,k_12_3467,k_12_3468,k_12_3469,k_12_3470,k_12_3471,k_12_3472,k_12_3473,k_12_3474,k_12_3475,k_12_3476,k_12_3477,k_12_3478,k_12_3479,k_12_3480,k_12_3481,k_12_3482,k_12_3483,k_12_3484,k_12_3485,k_12_3486,k_12_3487,k_12_3488,k_12_3489,k_12_3490,k_12_3491,k_12_3492,k_12_3493,k_12_3494,k_12_3495,k_12_3496,k_12_3497,k_12_3498,k_12_3499,k_12_3500,k_12_3501,k_12_3502,k_12_3503,k_12_3504,k_12_3505,k_12_3506,k_12_3507,k_12_3508,k_12_3509,k_12_3510,k_12_3511,k_12_3512,k_12_3513,k_12_3514,k_12_3515,k_12_3516,k_12_3517,k_12_3518,k_12_3519,k_12_3520,k_12_3521,k_12_3522,k_12_3523,k_12_3524,k_12_3525,k_12_3526,k_12_3527,k_12_3528,k_12_3529,k_12_3530,k_12_3531,k_12_3532,k_12_3533,k_12_3534,k_12_3535,k_12_3536,k_12_3537,k_12_3538,k_12_3539,k_12_3540,k_12_3541,k_12_3542,k_12_3543,k_12_3544,k_12_3545,k_12_3546,k_12_3547,k_12_3548,k_12_3549,k_12_3550,k_12_3551,k_12_3552,k_12_3553,k_12_3554,k_12_3555,k_12_3556,k_12_3557,k_12_3558,k_12_3559,k_12_3560,k_12_3561,k_12_3562,k_12_3563,k_12_3564,k_12_3565,k_12_3566,k_12_3567,k_12_3568,k_12_3569,k_12_3570,k_12_3571,k_12_3572,k_12_3573,k_12_3574,k_12_3575,k_12_3576,k_12_3577,k_12_3578,k_12_3579,k_12_3580,k_12_3581,k_12_3582,k_12_3583,k_12_3584,k_12_3585,k_12_3586,k_12_3587,k_12_3588,k_12_3589,k_12_3590,k_12_3591,k_12_3592,k_12_3593,k_12_3594,k_12_3595,k_12_3596,k_12_3597,k_12_3598,k_12_3599,k_12_3600,k_12_3601,k_12_3602,k_12_3603,k_12_3604,k_12_3605,k_12_3606,k_12_3607,k_12_3608,k_12_3609,k_12_3610,k_12_3611,k_12_3612,k_12_3613,k_12_3614,k_12_3615,k_12_3616,k_12_3617,k_12_3618,k_12_3619,k_12_3620,k_12_3621,k_12_3622,k_12_3623,k_12_3624,k_12_3625,k_12_3626,k_12_3627,k_12_3628,k_12_3629,k_12_3630,k_12_3631,k_12_3632,k_12_3633,k_12_3634,k_12_3635,k_12_3636,k_12_3637,k_12_3638,k_12_3639,k_12_3640,k_12_3641,k_12_3642,k_12_3643,k_12_3644,k_12_3645,k_12_3646,k_12_3647,k_12_3648,k_12_3649,k_12_3650,k_12_3651,k_12_3652,k_12_3653,k_12_3654,k_12_3655,k_12_3656,k_12_3657,k_12_3658,k_12_3659,k_12_3660,k_12_3661,k_12_3662,k_12_3663,k_12_3664,k_12_3665,k_12_3666,k_12_3667,k_12_3668,k_12_3669,k_12_3670,k_12_3671,k_12_3672,k_12_3673,k_12_3674,k_12_3675,k_12_3676,k_12_3677,k_12_3678,k_12_3679,k_12_3680,k_12_3681,k_12_3682,k_12_3683,k_12_3684,k_12_3685,k_12_3686,k_12_3687,k_12_3688,k_12_3689,k_12_3690,k_12_3691,k_12_3692,k_12_3693,k_12_3694,k_12_3695,k_12_3696,k_12_3697,k_12_3698,k_12_3699,k_12_3700,k_12_3701,k_12_3702,k_12_3703,k_12_3704,k_12_3705,k_12_3706,k_12_3707,k_12_3708,k_12_3709,k_12_3710,k_12_3711,k_12_3712,k_12_3713,k_12_3714,k_12_3715,k_12_3716,k_12_3717,k_12_3718,k_12_3719,k_12_3720,k_12_3721,k_12_3722,k_12_3723,k_12_3724,k_12_3725,k_12_3726,k_12_3727,k_12_3728,k_12_3729,k_12_3730,k_12_3731,k_12_3732,k_12_3733,k_12_3734,k_12_3735,k_12_3736,k_12_3737,k_12_3738,k_12_3739,k_12_3740,k_12_3741,k_12_3742,k_12_3743,k_12_3744,k_12_3745,k_12_3746,k_12_3747,k_12_3748,k_12_3749,k_12_3750,k_12_3751,k_12_3752,k_12_3753,k_12_3754,k_12_3755,k_12_3756,k_12_3757,k_12_3758,k_12_3759,k_12_3760,k_12_3761,k_12_3762,k_12_3763,k_12_3764,k_12_3765,k_12_3766,k_12_3767,k_12_3768,k_12_3769,k_12_3770,k_12_3771,k_12_3772,k_12_3773,k_12_3774,k_12_3775,k_12_3776,k_12_3777,k_12_3778,k_12_3779,k_12_3780,k_12_3781,k_12_3782,k_12_3783,k_12_3784,k_12_3785,k_12_3786,k_12_3787,k_12_3788,k_12_3789,k_12_3790,k_12_3791,k_12_3792,k_12_3793,k_12_3794,k_12_3795,k_12_3796,k_12_3797,k_12_3798,k_12_3799,k_12_3800,k_12_3801,k_12_3802,k_12_3803,k_12_3804,k_12_3805,k_12_3806,k_12_3807,k_12_3808,k_12_3809,k_12_3810,k_12_3811,k_12_3812,k_12_3813,k_12_3814,k_12_3815,k_12_3816,k_12_3817,k_12_3818,k_12_3819,k_12_3820,k_12_3821,k_12_3822,k_12_3823,k_12_3824,k_12_3825,k_12_3826,k_12_3827,k_12_3828,k_12_3829,k_12_3830,k_12_3831,k_12_3832,k_12_3833,k_12_3834,k_12_3835,k_12_3836,k_12_3837,k_12_3838,k_12_3839,k_12_3840,k_12_3841,k_12_3842,k_12_3843,k_12_3844,k_12_3845,k_12_3846,k_12_3847,k_12_3848,k_12_3849,k_12_3850,k_12_3851,k_12_3852,k_12_3853,k_12_3854,k_12_3855,k_12_3856,k_12_3857,k_12_3858,k_12_3859,k_12_3860,k_12_3861,k_12_3862,k_12_3863,k_12_3864,k_12_3865,k_12_3866,k_12_3867,k_12_3868,k_12_3869,k_12_3870,k_12_3871,k_12_3872,k_12_3873,k_12_3874,k_12_3875,k_12_3876,k_12_3877,k_12_3878,k_12_3879,k_12_3880,k_12_3881,k_12_3882,k_12_3883,k_12_3884,k_12_3885,k_12_3886,k_12_3887,k_12_3888,k_12_3889,k_12_3890,k_12_3891,k_12_3892,k_12_3893,k_12_3894,k_12_3895,k_12_3896,k_12_3897,k_12_3898,k_12_3899,k_12_3900,k_12_3901,k_12_3902,k_12_3903,k_12_3904,k_12_3905,k_12_3906,k_12_3907,k_12_3908,k_12_3909,k_12_3910,k_12_3911,k_12_3912,k_12_3913,k_12_3914,k_12_3915,k_12_3916,k_12_3917,k_12_3918,k_12_3919,k_12_3920,k_12_3921,k_12_3922,k_12_3923,k_12_3924,k_12_3925,k_12_3926,k_12_3927,k_12_3928,k_12_3929,k_12_3930,k_12_3931,k_12_3932,k_12_3933,k_12_3934,k_12_3935,k_12_3936,k_12_3937,k_12_3938,k_12_3939,k_12_3940,k_12_3941,k_12_3942,k_12_3943,k_12_3944,k_12_3945,k_12_3946,k_12_3947,k_12_3948,k_12_3949,k_12_3950,k_12_3951,k_12_3952,k_12_3953,k_12_3954,k_12_3955,k_12_3956,k_12_3957,k_12_3958,k_12_3959,k_12_3960,k_12_3961,k_12_3962,k_12_3963,k_12_3964,k_12_3965,k_12_3966,k_12_3967,k_12_3968,k_12_3969,k_12_3970,k_12_3971,k_12_3972,k_12_3973,k_12_3974,k_12_3975,k_12_3976,k_12_3977,k_12_3978,k_12_3979,k_12_3980,k_12_3981,k_12_3982,k_12_3983,k_12_3984,k_12_3985,k_12_3986,k_12_3987,k_12_3988,k_12_3989,k_12_3990,k_12_3991,k_12_3992,k_12_3993,k_12_3994,k_12_3995,k_12_3996,k_12_3997,k_12_3998,k_12_3999,k_12_4000,k_12_4001,k_12_4002,k_12_4003,k_12_4004,k_12_4005,k_12_4006,k_12_4007,k_12_4008,k_12_4009,k_12_4010,k_12_4011,k_12_4012,k_12_4013,k_12_4014,k_12_4015,k_12_4016,k_12_4017,k_12_4018,k_12_4019,k_12_4020,k_12_4021,k_12_4022,k_12_4023,k_12_4024,k_12_4025,k_12_4026,k_12_4027,k_12_4028,k_12_4029,k_12_4030,k_12_4031,k_12_4032,k_12_4033,k_12_4034,k_12_4035,k_12_4036,k_12_4037,k_12_4038,k_12_4039,k_12_4040,k_12_4041,k_12_4042,k_12_4043,k_12_4044,k_12_4045,k_12_4046,k_12_4047,k_12_4048,k_12_4049,k_12_4050,k_12_4051,k_12_4052,k_12_4053,k_12_4054,k_12_4055,k_12_4056,k_12_4057,k_12_4058,k_12_4059,k_12_4060,k_12_4061,k_12_4062,k_12_4063,k_12_4064,k_12_4065,k_12_4066,k_12_4067,k_12_4068,k_12_4069,k_12_4070,k_12_4071,k_12_4072,k_12_4073,k_12_4074,k_12_4075,k_12_4076,k_12_4077,k_12_4078,k_12_4079,k_12_4080,k_12_4081,k_12_4082,k_12_4083,k_12_4084,k_12_4085,k_12_4086,k_12_4087,k_12_4088,k_12_4089,k_12_4090,k_12_4091,k_12_4092,k_12_4093,k_12_4094,k_12_4095,
input c_0_0, c_0_1,
input c_1_0, c_1_1,
input c_2_0, c_2_1,
input c_3_0, c_3_1,
input c_4_0, c_4_1,
input c_5_0, c_5_1,
input c_6_0, c_6_1,
input c_7_0, c_7_1,
input c_8_0, c_8_1,
input c_9_0, c_9_1,
input c_10_0, c_10_1,
input c_11_0, c_11_1,
input c_12_0, c_12_1
);
wire k_1_0,k_1_1;
wire k_2_0,k_2_1,k_2_2,k_2_3;
wire k_3_0,k_3_1,k_3_2,k_3_3,k_3_4,k_3_5,k_3_6,k_3_7;
wire k_4_0,k_4_1,k_4_2,k_4_3,k_4_4,k_4_5,k_4_6,k_4_7,k_4_8,k_4_9,k_4_10,k_4_11,k_4_12,k_4_13,k_4_14,k_4_15;
wire k_5_0,k_5_1,k_5_2,k_5_3,k_5_4,k_5_5,k_5_6,k_5_7,k_5_8,k_5_9,k_5_10,k_5_11,k_5_12,k_5_13,k_5_14,k_5_15,k_5_16,k_5_17,k_5_18,k_5_19,k_5_20,k_5_21,k_5_22,k_5_23,k_5_24,k_5_25,k_5_26,k_5_27,k_5_28,k_5_29,k_5_30,k_5_31;
wire k_6_0,k_6_1,k_6_2,k_6_3,k_6_4,k_6_5,k_6_6,k_6_7,k_6_8,k_6_9,k_6_10,k_6_11,k_6_12,k_6_13,k_6_14,k_6_15,k_6_16,k_6_17,k_6_18,k_6_19,k_6_20,k_6_21,k_6_22,k_6_23,k_6_24,k_6_25,k_6_26,k_6_27,k_6_28,k_6_29,k_6_30,k_6_31,k_6_32,k_6_33,k_6_34,k_6_35,k_6_36,k_6_37,k_6_38,k_6_39,k_6_40,k_6_41,k_6_42,k_6_43,k_6_44,k_6_45,k_6_46,k_6_47,k_6_48,k_6_49,k_6_50,k_6_51,k_6_52,k_6_53,k_6_54,k_6_55,k_6_56,k_6_57,k_6_58,k_6_59,k_6_60,k_6_61,k_6_62,k_6_63;
wire k_7_0,k_7_1,k_7_2,k_7_3,k_7_4,k_7_5,k_7_6,k_7_7,k_7_8,k_7_9,k_7_10,k_7_11,k_7_12,k_7_13,k_7_14,k_7_15,k_7_16,k_7_17,k_7_18,k_7_19,k_7_20,k_7_21,k_7_22,k_7_23,k_7_24,k_7_25,k_7_26,k_7_27,k_7_28,k_7_29,k_7_30,k_7_31,k_7_32,k_7_33,k_7_34,k_7_35,k_7_36,k_7_37,k_7_38,k_7_39,k_7_40,k_7_41,k_7_42,k_7_43,k_7_44,k_7_45,k_7_46,k_7_47,k_7_48,k_7_49,k_7_50,k_7_51,k_7_52,k_7_53,k_7_54,k_7_55,k_7_56,k_7_57,k_7_58,k_7_59,k_7_60,k_7_61,k_7_62,k_7_63,k_7_64,k_7_65,k_7_66,k_7_67,k_7_68,k_7_69,k_7_70,k_7_71,k_7_72,k_7_73,k_7_74,k_7_75,k_7_76,k_7_77,k_7_78,k_7_79,k_7_80,k_7_81,k_7_82,k_7_83,k_7_84,k_7_85,k_7_86,k_7_87,k_7_88,k_7_89,k_7_90,k_7_91,k_7_92,k_7_93,k_7_94,k_7_95,k_7_96,k_7_97,k_7_98,k_7_99,k_7_100,k_7_101,k_7_102,k_7_103,k_7_104,k_7_105,k_7_106,k_7_107,k_7_108,k_7_109,k_7_110,k_7_111,k_7_112,k_7_113,k_7_114,k_7_115,k_7_116,k_7_117,k_7_118,k_7_119,k_7_120,k_7_121,k_7_122,k_7_123,k_7_124,k_7_125,k_7_126,k_7_127;
wire k_8_0,k_8_1,k_8_2,k_8_3,k_8_4,k_8_5,k_8_6,k_8_7,k_8_8,k_8_9,k_8_10,k_8_11,k_8_12,k_8_13,k_8_14,k_8_15,k_8_16,k_8_17,k_8_18,k_8_19,k_8_20,k_8_21,k_8_22,k_8_23,k_8_24,k_8_25,k_8_26,k_8_27,k_8_28,k_8_29,k_8_30,k_8_31,k_8_32,k_8_33,k_8_34,k_8_35,k_8_36,k_8_37,k_8_38,k_8_39,k_8_40,k_8_41,k_8_42,k_8_43,k_8_44,k_8_45,k_8_46,k_8_47,k_8_48,k_8_49,k_8_50,k_8_51,k_8_52,k_8_53,k_8_54,k_8_55,k_8_56,k_8_57,k_8_58,k_8_59,k_8_60,k_8_61,k_8_62,k_8_63,k_8_64,k_8_65,k_8_66,k_8_67,k_8_68,k_8_69,k_8_70,k_8_71,k_8_72,k_8_73,k_8_74,k_8_75,k_8_76,k_8_77,k_8_78,k_8_79,k_8_80,k_8_81,k_8_82,k_8_83,k_8_84,k_8_85,k_8_86,k_8_87,k_8_88,k_8_89,k_8_90,k_8_91,k_8_92,k_8_93,k_8_94,k_8_95,k_8_96,k_8_97,k_8_98,k_8_99,k_8_100,k_8_101,k_8_102,k_8_103,k_8_104,k_8_105,k_8_106,k_8_107,k_8_108,k_8_109,k_8_110,k_8_111,k_8_112,k_8_113,k_8_114,k_8_115,k_8_116,k_8_117,k_8_118,k_8_119,k_8_120,k_8_121,k_8_122,k_8_123,k_8_124,k_8_125,k_8_126,k_8_127,k_8_128,k_8_129,k_8_130,k_8_131,k_8_132,k_8_133,k_8_134,k_8_135,k_8_136,k_8_137,k_8_138,k_8_139,k_8_140,k_8_141,k_8_142,k_8_143,k_8_144,k_8_145,k_8_146,k_8_147,k_8_148,k_8_149,k_8_150,k_8_151,k_8_152,k_8_153,k_8_154,k_8_155,k_8_156,k_8_157,k_8_158,k_8_159,k_8_160,k_8_161,k_8_162,k_8_163,k_8_164,k_8_165,k_8_166,k_8_167,k_8_168,k_8_169,k_8_170,k_8_171,k_8_172,k_8_173,k_8_174,k_8_175,k_8_176,k_8_177,k_8_178,k_8_179,k_8_180,k_8_181,k_8_182,k_8_183,k_8_184,k_8_185,k_8_186,k_8_187,k_8_188,k_8_189,k_8_190,k_8_191,k_8_192,k_8_193,k_8_194,k_8_195,k_8_196,k_8_197,k_8_198,k_8_199,k_8_200,k_8_201,k_8_202,k_8_203,k_8_204,k_8_205,k_8_206,k_8_207,k_8_208,k_8_209,k_8_210,k_8_211,k_8_212,k_8_213,k_8_214,k_8_215,k_8_216,k_8_217,k_8_218,k_8_219,k_8_220,k_8_221,k_8_222,k_8_223,k_8_224,k_8_225,k_8_226,k_8_227,k_8_228,k_8_229,k_8_230,k_8_231,k_8_232,k_8_233,k_8_234,k_8_235,k_8_236,k_8_237,k_8_238,k_8_239,k_8_240,k_8_241,k_8_242,k_8_243,k_8_244,k_8_245,k_8_246,k_8_247,k_8_248,k_8_249,k_8_250,k_8_251,k_8_252,k_8_253,k_8_254,k_8_255;
wire k_9_0,k_9_1,k_9_2,k_9_3,k_9_4,k_9_5,k_9_6,k_9_7,k_9_8,k_9_9,k_9_10,k_9_11,k_9_12,k_9_13,k_9_14,k_9_15,k_9_16,k_9_17,k_9_18,k_9_19,k_9_20,k_9_21,k_9_22,k_9_23,k_9_24,k_9_25,k_9_26,k_9_27,k_9_28,k_9_29,k_9_30,k_9_31,k_9_32,k_9_33,k_9_34,k_9_35,k_9_36,k_9_37,k_9_38,k_9_39,k_9_40,k_9_41,k_9_42,k_9_43,k_9_44,k_9_45,k_9_46,k_9_47,k_9_48,k_9_49,k_9_50,k_9_51,k_9_52,k_9_53,k_9_54,k_9_55,k_9_56,k_9_57,k_9_58,k_9_59,k_9_60,k_9_61,k_9_62,k_9_63,k_9_64,k_9_65,k_9_66,k_9_67,k_9_68,k_9_69,k_9_70,k_9_71,k_9_72,k_9_73,k_9_74,k_9_75,k_9_76,k_9_77,k_9_78,k_9_79,k_9_80,k_9_81,k_9_82,k_9_83,k_9_84,k_9_85,k_9_86,k_9_87,k_9_88,k_9_89,k_9_90,k_9_91,k_9_92,k_9_93,k_9_94,k_9_95,k_9_96,k_9_97,k_9_98,k_9_99,k_9_100,k_9_101,k_9_102,k_9_103,k_9_104,k_9_105,k_9_106,k_9_107,k_9_108,k_9_109,k_9_110,k_9_111,k_9_112,k_9_113,k_9_114,k_9_115,k_9_116,k_9_117,k_9_118,k_9_119,k_9_120,k_9_121,k_9_122,k_9_123,k_9_124,k_9_125,k_9_126,k_9_127,k_9_128,k_9_129,k_9_130,k_9_131,k_9_132,k_9_133,k_9_134,k_9_135,k_9_136,k_9_137,k_9_138,k_9_139,k_9_140,k_9_141,k_9_142,k_9_143,k_9_144,k_9_145,k_9_146,k_9_147,k_9_148,k_9_149,k_9_150,k_9_151,k_9_152,k_9_153,k_9_154,k_9_155,k_9_156,k_9_157,k_9_158,k_9_159,k_9_160,k_9_161,k_9_162,k_9_163,k_9_164,k_9_165,k_9_166,k_9_167,k_9_168,k_9_169,k_9_170,k_9_171,k_9_172,k_9_173,k_9_174,k_9_175,k_9_176,k_9_177,k_9_178,k_9_179,k_9_180,k_9_181,k_9_182,k_9_183,k_9_184,k_9_185,k_9_186,k_9_187,k_9_188,k_9_189,k_9_190,k_9_191,k_9_192,k_9_193,k_9_194,k_9_195,k_9_196,k_9_197,k_9_198,k_9_199,k_9_200,k_9_201,k_9_202,k_9_203,k_9_204,k_9_205,k_9_206,k_9_207,k_9_208,k_9_209,k_9_210,k_9_211,k_9_212,k_9_213,k_9_214,k_9_215,k_9_216,k_9_217,k_9_218,k_9_219,k_9_220,k_9_221,k_9_222,k_9_223,k_9_224,k_9_225,k_9_226,k_9_227,k_9_228,k_9_229,k_9_230,k_9_231,k_9_232,k_9_233,k_9_234,k_9_235,k_9_236,k_9_237,k_9_238,k_9_239,k_9_240,k_9_241,k_9_242,k_9_243,k_9_244,k_9_245,k_9_246,k_9_247,k_9_248,k_9_249,k_9_250,k_9_251,k_9_252,k_9_253,k_9_254,k_9_255,k_9_256,k_9_257,k_9_258,k_9_259,k_9_260,k_9_261,k_9_262,k_9_263,k_9_264,k_9_265,k_9_266,k_9_267,k_9_268,k_9_269,k_9_270,k_9_271,k_9_272,k_9_273,k_9_274,k_9_275,k_9_276,k_9_277,k_9_278,k_9_279,k_9_280,k_9_281,k_9_282,k_9_283,k_9_284,k_9_285,k_9_286,k_9_287,k_9_288,k_9_289,k_9_290,k_9_291,k_9_292,k_9_293,k_9_294,k_9_295,k_9_296,k_9_297,k_9_298,k_9_299,k_9_300,k_9_301,k_9_302,k_9_303,k_9_304,k_9_305,k_9_306,k_9_307,k_9_308,k_9_309,k_9_310,k_9_311,k_9_312,k_9_313,k_9_314,k_9_315,k_9_316,k_9_317,k_9_318,k_9_319,k_9_320,k_9_321,k_9_322,k_9_323,k_9_324,k_9_325,k_9_326,k_9_327,k_9_328,k_9_329,k_9_330,k_9_331,k_9_332,k_9_333,k_9_334,k_9_335,k_9_336,k_9_337,k_9_338,k_9_339,k_9_340,k_9_341,k_9_342,k_9_343,k_9_344,k_9_345,k_9_346,k_9_347,k_9_348,k_9_349,k_9_350,k_9_351,k_9_352,k_9_353,k_9_354,k_9_355,k_9_356,k_9_357,k_9_358,k_9_359,k_9_360,k_9_361,k_9_362,k_9_363,k_9_364,k_9_365,k_9_366,k_9_367,k_9_368,k_9_369,k_9_370,k_9_371,k_9_372,k_9_373,k_9_374,k_9_375,k_9_376,k_9_377,k_9_378,k_9_379,k_9_380,k_9_381,k_9_382,k_9_383,k_9_384,k_9_385,k_9_386,k_9_387,k_9_388,k_9_389,k_9_390,k_9_391,k_9_392,k_9_393,k_9_394,k_9_395,k_9_396,k_9_397,k_9_398,k_9_399,k_9_400,k_9_401,k_9_402,k_9_403,k_9_404,k_9_405,k_9_406,k_9_407,k_9_408,k_9_409,k_9_410,k_9_411,k_9_412,k_9_413,k_9_414,k_9_415,k_9_416,k_9_417,k_9_418,k_9_419,k_9_420,k_9_421,k_9_422,k_9_423,k_9_424,k_9_425,k_9_426,k_9_427,k_9_428,k_9_429,k_9_430,k_9_431,k_9_432,k_9_433,k_9_434,k_9_435,k_9_436,k_9_437,k_9_438,k_9_439,k_9_440,k_9_441,k_9_442,k_9_443,k_9_444,k_9_445,k_9_446,k_9_447,k_9_448,k_9_449,k_9_450,k_9_451,k_9_452,k_9_453,k_9_454,k_9_455,k_9_456,k_9_457,k_9_458,k_9_459,k_9_460,k_9_461,k_9_462,k_9_463,k_9_464,k_9_465,k_9_466,k_9_467,k_9_468,k_9_469,k_9_470,k_9_471,k_9_472,k_9_473,k_9_474,k_9_475,k_9_476,k_9_477,k_9_478,k_9_479,k_9_480,k_9_481,k_9_482,k_9_483,k_9_484,k_9_485,k_9_486,k_9_487,k_9_488,k_9_489,k_9_490,k_9_491,k_9_492,k_9_493,k_9_494,k_9_495,k_9_496,k_9_497,k_9_498,k_9_499,k_9_500,k_9_501,k_9_502,k_9_503,k_9_504,k_9_505,k_9_506,k_9_507,k_9_508,k_9_509,k_9_510,k_9_511;
wire k_10_0,k_10_1,k_10_2,k_10_3,k_10_4,k_10_5,k_10_6,k_10_7,k_10_8,k_10_9,k_10_10,k_10_11,k_10_12,k_10_13,k_10_14,k_10_15,k_10_16,k_10_17,k_10_18,k_10_19,k_10_20,k_10_21,k_10_22,k_10_23,k_10_24,k_10_25,k_10_26,k_10_27,k_10_28,k_10_29,k_10_30,k_10_31,k_10_32,k_10_33,k_10_34,k_10_35,k_10_36,k_10_37,k_10_38,k_10_39,k_10_40,k_10_41,k_10_42,k_10_43,k_10_44,k_10_45,k_10_46,k_10_47,k_10_48,k_10_49,k_10_50,k_10_51,k_10_52,k_10_53,k_10_54,k_10_55,k_10_56,k_10_57,k_10_58,k_10_59,k_10_60,k_10_61,k_10_62,k_10_63,k_10_64,k_10_65,k_10_66,k_10_67,k_10_68,k_10_69,k_10_70,k_10_71,k_10_72,k_10_73,k_10_74,k_10_75,k_10_76,k_10_77,k_10_78,k_10_79,k_10_80,k_10_81,k_10_82,k_10_83,k_10_84,k_10_85,k_10_86,k_10_87,k_10_88,k_10_89,k_10_90,k_10_91,k_10_92,k_10_93,k_10_94,k_10_95,k_10_96,k_10_97,k_10_98,k_10_99,k_10_100,k_10_101,k_10_102,k_10_103,k_10_104,k_10_105,k_10_106,k_10_107,k_10_108,k_10_109,k_10_110,k_10_111,k_10_112,k_10_113,k_10_114,k_10_115,k_10_116,k_10_117,k_10_118,k_10_119,k_10_120,k_10_121,k_10_122,k_10_123,k_10_124,k_10_125,k_10_126,k_10_127,k_10_128,k_10_129,k_10_130,k_10_131,k_10_132,k_10_133,k_10_134,k_10_135,k_10_136,k_10_137,k_10_138,k_10_139,k_10_140,k_10_141,k_10_142,k_10_143,k_10_144,k_10_145,k_10_146,k_10_147,k_10_148,k_10_149,k_10_150,k_10_151,k_10_152,k_10_153,k_10_154,k_10_155,k_10_156,k_10_157,k_10_158,k_10_159,k_10_160,k_10_161,k_10_162,k_10_163,k_10_164,k_10_165,k_10_166,k_10_167,k_10_168,k_10_169,k_10_170,k_10_171,k_10_172,k_10_173,k_10_174,k_10_175,k_10_176,k_10_177,k_10_178,k_10_179,k_10_180,k_10_181,k_10_182,k_10_183,k_10_184,k_10_185,k_10_186,k_10_187,k_10_188,k_10_189,k_10_190,k_10_191,k_10_192,k_10_193,k_10_194,k_10_195,k_10_196,k_10_197,k_10_198,k_10_199,k_10_200,k_10_201,k_10_202,k_10_203,k_10_204,k_10_205,k_10_206,k_10_207,k_10_208,k_10_209,k_10_210,k_10_211,k_10_212,k_10_213,k_10_214,k_10_215,k_10_216,k_10_217,k_10_218,k_10_219,k_10_220,k_10_221,k_10_222,k_10_223,k_10_224,k_10_225,k_10_226,k_10_227,k_10_228,k_10_229,k_10_230,k_10_231,k_10_232,k_10_233,k_10_234,k_10_235,k_10_236,k_10_237,k_10_238,k_10_239,k_10_240,k_10_241,k_10_242,k_10_243,k_10_244,k_10_245,k_10_246,k_10_247,k_10_248,k_10_249,k_10_250,k_10_251,k_10_252,k_10_253,k_10_254,k_10_255,k_10_256,k_10_257,k_10_258,k_10_259,k_10_260,k_10_261,k_10_262,k_10_263,k_10_264,k_10_265,k_10_266,k_10_267,k_10_268,k_10_269,k_10_270,k_10_271,k_10_272,k_10_273,k_10_274,k_10_275,k_10_276,k_10_277,k_10_278,k_10_279,k_10_280,k_10_281,k_10_282,k_10_283,k_10_284,k_10_285,k_10_286,k_10_287,k_10_288,k_10_289,k_10_290,k_10_291,k_10_292,k_10_293,k_10_294,k_10_295,k_10_296,k_10_297,k_10_298,k_10_299,k_10_300,k_10_301,k_10_302,k_10_303,k_10_304,k_10_305,k_10_306,k_10_307,k_10_308,k_10_309,k_10_310,k_10_311,k_10_312,k_10_313,k_10_314,k_10_315,k_10_316,k_10_317,k_10_318,k_10_319,k_10_320,k_10_321,k_10_322,k_10_323,k_10_324,k_10_325,k_10_326,k_10_327,k_10_328,k_10_329,k_10_330,k_10_331,k_10_332,k_10_333,k_10_334,k_10_335,k_10_336,k_10_337,k_10_338,k_10_339,k_10_340,k_10_341,k_10_342,k_10_343,k_10_344,k_10_345,k_10_346,k_10_347,k_10_348,k_10_349,k_10_350,k_10_351,k_10_352,k_10_353,k_10_354,k_10_355,k_10_356,k_10_357,k_10_358,k_10_359,k_10_360,k_10_361,k_10_362,k_10_363,k_10_364,k_10_365,k_10_366,k_10_367,k_10_368,k_10_369,k_10_370,k_10_371,k_10_372,k_10_373,k_10_374,k_10_375,k_10_376,k_10_377,k_10_378,k_10_379,k_10_380,k_10_381,k_10_382,k_10_383,k_10_384,k_10_385,k_10_386,k_10_387,k_10_388,k_10_389,k_10_390,k_10_391,k_10_392,k_10_393,k_10_394,k_10_395,k_10_396,k_10_397,k_10_398,k_10_399,k_10_400,k_10_401,k_10_402,k_10_403,k_10_404,k_10_405,k_10_406,k_10_407,k_10_408,k_10_409,k_10_410,k_10_411,k_10_412,k_10_413,k_10_414,k_10_415,k_10_416,k_10_417,k_10_418,k_10_419,k_10_420,k_10_421,k_10_422,k_10_423,k_10_424,k_10_425,k_10_426,k_10_427,k_10_428,k_10_429,k_10_430,k_10_431,k_10_432,k_10_433,k_10_434,k_10_435,k_10_436,k_10_437,k_10_438,k_10_439,k_10_440,k_10_441,k_10_442,k_10_443,k_10_444,k_10_445,k_10_446,k_10_447,k_10_448,k_10_449,k_10_450,k_10_451,k_10_452,k_10_453,k_10_454,k_10_455,k_10_456,k_10_457,k_10_458,k_10_459,k_10_460,k_10_461,k_10_462,k_10_463,k_10_464,k_10_465,k_10_466,k_10_467,k_10_468,k_10_469,k_10_470,k_10_471,k_10_472,k_10_473,k_10_474,k_10_475,k_10_476,k_10_477,k_10_478,k_10_479,k_10_480,k_10_481,k_10_482,k_10_483,k_10_484,k_10_485,k_10_486,k_10_487,k_10_488,k_10_489,k_10_490,k_10_491,k_10_492,k_10_493,k_10_494,k_10_495,k_10_496,k_10_497,k_10_498,k_10_499,k_10_500,k_10_501,k_10_502,k_10_503,k_10_504,k_10_505,k_10_506,k_10_507,k_10_508,k_10_509,k_10_510,k_10_511,k_10_512,k_10_513,k_10_514,k_10_515,k_10_516,k_10_517,k_10_518,k_10_519,k_10_520,k_10_521,k_10_522,k_10_523,k_10_524,k_10_525,k_10_526,k_10_527,k_10_528,k_10_529,k_10_530,k_10_531,k_10_532,k_10_533,k_10_534,k_10_535,k_10_536,k_10_537,k_10_538,k_10_539,k_10_540,k_10_541,k_10_542,k_10_543,k_10_544,k_10_545,k_10_546,k_10_547,k_10_548,k_10_549,k_10_550,k_10_551,k_10_552,k_10_553,k_10_554,k_10_555,k_10_556,k_10_557,k_10_558,k_10_559,k_10_560,k_10_561,k_10_562,k_10_563,k_10_564,k_10_565,k_10_566,k_10_567,k_10_568,k_10_569,k_10_570,k_10_571,k_10_572,k_10_573,k_10_574,k_10_575,k_10_576,k_10_577,k_10_578,k_10_579,k_10_580,k_10_581,k_10_582,k_10_583,k_10_584,k_10_585,k_10_586,k_10_587,k_10_588,k_10_589,k_10_590,k_10_591,k_10_592,k_10_593,k_10_594,k_10_595,k_10_596,k_10_597,k_10_598,k_10_599,k_10_600,k_10_601,k_10_602,k_10_603,k_10_604,k_10_605,k_10_606,k_10_607,k_10_608,k_10_609,k_10_610,k_10_611,k_10_612,k_10_613,k_10_614,k_10_615,k_10_616,k_10_617,k_10_618,k_10_619,k_10_620,k_10_621,k_10_622,k_10_623,k_10_624,k_10_625,k_10_626,k_10_627,k_10_628,k_10_629,k_10_630,k_10_631,k_10_632,k_10_633,k_10_634,k_10_635,k_10_636,k_10_637,k_10_638,k_10_639,k_10_640,k_10_641,k_10_642,k_10_643,k_10_644,k_10_645,k_10_646,k_10_647,k_10_648,k_10_649,k_10_650,k_10_651,k_10_652,k_10_653,k_10_654,k_10_655,k_10_656,k_10_657,k_10_658,k_10_659,k_10_660,k_10_661,k_10_662,k_10_663,k_10_664,k_10_665,k_10_666,k_10_667,k_10_668,k_10_669,k_10_670,k_10_671,k_10_672,k_10_673,k_10_674,k_10_675,k_10_676,k_10_677,k_10_678,k_10_679,k_10_680,k_10_681,k_10_682,k_10_683,k_10_684,k_10_685,k_10_686,k_10_687,k_10_688,k_10_689,k_10_690,k_10_691,k_10_692,k_10_693,k_10_694,k_10_695,k_10_696,k_10_697,k_10_698,k_10_699,k_10_700,k_10_701,k_10_702,k_10_703,k_10_704,k_10_705,k_10_706,k_10_707,k_10_708,k_10_709,k_10_710,k_10_711,k_10_712,k_10_713,k_10_714,k_10_715,k_10_716,k_10_717,k_10_718,k_10_719,k_10_720,k_10_721,k_10_722,k_10_723,k_10_724,k_10_725,k_10_726,k_10_727,k_10_728,k_10_729,k_10_730,k_10_731,k_10_732,k_10_733,k_10_734,k_10_735,k_10_736,k_10_737,k_10_738,k_10_739,k_10_740,k_10_741,k_10_742,k_10_743,k_10_744,k_10_745,k_10_746,k_10_747,k_10_748,k_10_749,k_10_750,k_10_751,k_10_752,k_10_753,k_10_754,k_10_755,k_10_756,k_10_757,k_10_758,k_10_759,k_10_760,k_10_761,k_10_762,k_10_763,k_10_764,k_10_765,k_10_766,k_10_767,k_10_768,k_10_769,k_10_770,k_10_771,k_10_772,k_10_773,k_10_774,k_10_775,k_10_776,k_10_777,k_10_778,k_10_779,k_10_780,k_10_781,k_10_782,k_10_783,k_10_784,k_10_785,k_10_786,k_10_787,k_10_788,k_10_789,k_10_790,k_10_791,k_10_792,k_10_793,k_10_794,k_10_795,k_10_796,k_10_797,k_10_798,k_10_799,k_10_800,k_10_801,k_10_802,k_10_803,k_10_804,k_10_805,k_10_806,k_10_807,k_10_808,k_10_809,k_10_810,k_10_811,k_10_812,k_10_813,k_10_814,k_10_815,k_10_816,k_10_817,k_10_818,k_10_819,k_10_820,k_10_821,k_10_822,k_10_823,k_10_824,k_10_825,k_10_826,k_10_827,k_10_828,k_10_829,k_10_830,k_10_831,k_10_832,k_10_833,k_10_834,k_10_835,k_10_836,k_10_837,k_10_838,k_10_839,k_10_840,k_10_841,k_10_842,k_10_843,k_10_844,k_10_845,k_10_846,k_10_847,k_10_848,k_10_849,k_10_850,k_10_851,k_10_852,k_10_853,k_10_854,k_10_855,k_10_856,k_10_857,k_10_858,k_10_859,k_10_860,k_10_861,k_10_862,k_10_863,k_10_864,k_10_865,k_10_866,k_10_867,k_10_868,k_10_869,k_10_870,k_10_871,k_10_872,k_10_873,k_10_874,k_10_875,k_10_876,k_10_877,k_10_878,k_10_879,k_10_880,k_10_881,k_10_882,k_10_883,k_10_884,k_10_885,k_10_886,k_10_887,k_10_888,k_10_889,k_10_890,k_10_891,k_10_892,k_10_893,k_10_894,k_10_895,k_10_896,k_10_897,k_10_898,k_10_899,k_10_900,k_10_901,k_10_902,k_10_903,k_10_904,k_10_905,k_10_906,k_10_907,k_10_908,k_10_909,k_10_910,k_10_911,k_10_912,k_10_913,k_10_914,k_10_915,k_10_916,k_10_917,k_10_918,k_10_919,k_10_920,k_10_921,k_10_922,k_10_923,k_10_924,k_10_925,k_10_926,k_10_927,k_10_928,k_10_929,k_10_930,k_10_931,k_10_932,k_10_933,k_10_934,k_10_935,k_10_936,k_10_937,k_10_938,k_10_939,k_10_940,k_10_941,k_10_942,k_10_943,k_10_944,k_10_945,k_10_946,k_10_947,k_10_948,k_10_949,k_10_950,k_10_951,k_10_952,k_10_953,k_10_954,k_10_955,k_10_956,k_10_957,k_10_958,k_10_959,k_10_960,k_10_961,k_10_962,k_10_963,k_10_964,k_10_965,k_10_966,k_10_967,k_10_968,k_10_969,k_10_970,k_10_971,k_10_972,k_10_973,k_10_974,k_10_975,k_10_976,k_10_977,k_10_978,k_10_979,k_10_980,k_10_981,k_10_982,k_10_983,k_10_984,k_10_985,k_10_986,k_10_987,k_10_988,k_10_989,k_10_990,k_10_991,k_10_992,k_10_993,k_10_994,k_10_995,k_10_996,k_10_997,k_10_998,k_10_999,k_10_1000,k_10_1001,k_10_1002,k_10_1003,k_10_1004,k_10_1005,k_10_1006,k_10_1007,k_10_1008,k_10_1009,k_10_1010,k_10_1011,k_10_1012,k_10_1013,k_10_1014,k_10_1015,k_10_1016,k_10_1017,k_10_1018,k_10_1019,k_10_1020,k_10_1021,k_10_1022,k_10_1023;
wire k_11_0,k_11_1,k_11_2,k_11_3,k_11_4,k_11_5,k_11_6,k_11_7,k_11_8,k_11_9,k_11_10,k_11_11,k_11_12,k_11_13,k_11_14,k_11_15,k_11_16,k_11_17,k_11_18,k_11_19,k_11_20,k_11_21,k_11_22,k_11_23,k_11_24,k_11_25,k_11_26,k_11_27,k_11_28,k_11_29,k_11_30,k_11_31,k_11_32,k_11_33,k_11_34,k_11_35,k_11_36,k_11_37,k_11_38,k_11_39,k_11_40,k_11_41,k_11_42,k_11_43,k_11_44,k_11_45,k_11_46,k_11_47,k_11_48,k_11_49,k_11_50,k_11_51,k_11_52,k_11_53,k_11_54,k_11_55,k_11_56,k_11_57,k_11_58,k_11_59,k_11_60,k_11_61,k_11_62,k_11_63,k_11_64,k_11_65,k_11_66,k_11_67,k_11_68,k_11_69,k_11_70,k_11_71,k_11_72,k_11_73,k_11_74,k_11_75,k_11_76,k_11_77,k_11_78,k_11_79,k_11_80,k_11_81,k_11_82,k_11_83,k_11_84,k_11_85,k_11_86,k_11_87,k_11_88,k_11_89,k_11_90,k_11_91,k_11_92,k_11_93,k_11_94,k_11_95,k_11_96,k_11_97,k_11_98,k_11_99,k_11_100,k_11_101,k_11_102,k_11_103,k_11_104,k_11_105,k_11_106,k_11_107,k_11_108,k_11_109,k_11_110,k_11_111,k_11_112,k_11_113,k_11_114,k_11_115,k_11_116,k_11_117,k_11_118,k_11_119,k_11_120,k_11_121,k_11_122,k_11_123,k_11_124,k_11_125,k_11_126,k_11_127,k_11_128,k_11_129,k_11_130,k_11_131,k_11_132,k_11_133,k_11_134,k_11_135,k_11_136,k_11_137,k_11_138,k_11_139,k_11_140,k_11_141,k_11_142,k_11_143,k_11_144,k_11_145,k_11_146,k_11_147,k_11_148,k_11_149,k_11_150,k_11_151,k_11_152,k_11_153,k_11_154,k_11_155,k_11_156,k_11_157,k_11_158,k_11_159,k_11_160,k_11_161,k_11_162,k_11_163,k_11_164,k_11_165,k_11_166,k_11_167,k_11_168,k_11_169,k_11_170,k_11_171,k_11_172,k_11_173,k_11_174,k_11_175,k_11_176,k_11_177,k_11_178,k_11_179,k_11_180,k_11_181,k_11_182,k_11_183,k_11_184,k_11_185,k_11_186,k_11_187,k_11_188,k_11_189,k_11_190,k_11_191,k_11_192,k_11_193,k_11_194,k_11_195,k_11_196,k_11_197,k_11_198,k_11_199,k_11_200,k_11_201,k_11_202,k_11_203,k_11_204,k_11_205,k_11_206,k_11_207,k_11_208,k_11_209,k_11_210,k_11_211,k_11_212,k_11_213,k_11_214,k_11_215,k_11_216,k_11_217,k_11_218,k_11_219,k_11_220,k_11_221,k_11_222,k_11_223,k_11_224,k_11_225,k_11_226,k_11_227,k_11_228,k_11_229,k_11_230,k_11_231,k_11_232,k_11_233,k_11_234,k_11_235,k_11_236,k_11_237,k_11_238,k_11_239,k_11_240,k_11_241,k_11_242,k_11_243,k_11_244,k_11_245,k_11_246,k_11_247,k_11_248,k_11_249,k_11_250,k_11_251,k_11_252,k_11_253,k_11_254,k_11_255,k_11_256,k_11_257,k_11_258,k_11_259,k_11_260,k_11_261,k_11_262,k_11_263,k_11_264,k_11_265,k_11_266,k_11_267,k_11_268,k_11_269,k_11_270,k_11_271,k_11_272,k_11_273,k_11_274,k_11_275,k_11_276,k_11_277,k_11_278,k_11_279,k_11_280,k_11_281,k_11_282,k_11_283,k_11_284,k_11_285,k_11_286,k_11_287,k_11_288,k_11_289,k_11_290,k_11_291,k_11_292,k_11_293,k_11_294,k_11_295,k_11_296,k_11_297,k_11_298,k_11_299,k_11_300,k_11_301,k_11_302,k_11_303,k_11_304,k_11_305,k_11_306,k_11_307,k_11_308,k_11_309,k_11_310,k_11_311,k_11_312,k_11_313,k_11_314,k_11_315,k_11_316,k_11_317,k_11_318,k_11_319,k_11_320,k_11_321,k_11_322,k_11_323,k_11_324,k_11_325,k_11_326,k_11_327,k_11_328,k_11_329,k_11_330,k_11_331,k_11_332,k_11_333,k_11_334,k_11_335,k_11_336,k_11_337,k_11_338,k_11_339,k_11_340,k_11_341,k_11_342,k_11_343,k_11_344,k_11_345,k_11_346,k_11_347,k_11_348,k_11_349,k_11_350,k_11_351,k_11_352,k_11_353,k_11_354,k_11_355,k_11_356,k_11_357,k_11_358,k_11_359,k_11_360,k_11_361,k_11_362,k_11_363,k_11_364,k_11_365,k_11_366,k_11_367,k_11_368,k_11_369,k_11_370,k_11_371,k_11_372,k_11_373,k_11_374,k_11_375,k_11_376,k_11_377,k_11_378,k_11_379,k_11_380,k_11_381,k_11_382,k_11_383,k_11_384,k_11_385,k_11_386,k_11_387,k_11_388,k_11_389,k_11_390,k_11_391,k_11_392,k_11_393,k_11_394,k_11_395,k_11_396,k_11_397,k_11_398,k_11_399,k_11_400,k_11_401,k_11_402,k_11_403,k_11_404,k_11_405,k_11_406,k_11_407,k_11_408,k_11_409,k_11_410,k_11_411,k_11_412,k_11_413,k_11_414,k_11_415,k_11_416,k_11_417,k_11_418,k_11_419,k_11_420,k_11_421,k_11_422,k_11_423,k_11_424,k_11_425,k_11_426,k_11_427,k_11_428,k_11_429,k_11_430,k_11_431,k_11_432,k_11_433,k_11_434,k_11_435,k_11_436,k_11_437,k_11_438,k_11_439,k_11_440,k_11_441,k_11_442,k_11_443,k_11_444,k_11_445,k_11_446,k_11_447,k_11_448,k_11_449,k_11_450,k_11_451,k_11_452,k_11_453,k_11_454,k_11_455,k_11_456,k_11_457,k_11_458,k_11_459,k_11_460,k_11_461,k_11_462,k_11_463,k_11_464,k_11_465,k_11_466,k_11_467,k_11_468,k_11_469,k_11_470,k_11_471,k_11_472,k_11_473,k_11_474,k_11_475,k_11_476,k_11_477,k_11_478,k_11_479,k_11_480,k_11_481,k_11_482,k_11_483,k_11_484,k_11_485,k_11_486,k_11_487,k_11_488,k_11_489,k_11_490,k_11_491,k_11_492,k_11_493,k_11_494,k_11_495,k_11_496,k_11_497,k_11_498,k_11_499,k_11_500,k_11_501,k_11_502,k_11_503,k_11_504,k_11_505,k_11_506,k_11_507,k_11_508,k_11_509,k_11_510,k_11_511,k_11_512,k_11_513,k_11_514,k_11_515,k_11_516,k_11_517,k_11_518,k_11_519,k_11_520,k_11_521,k_11_522,k_11_523,k_11_524,k_11_525,k_11_526,k_11_527,k_11_528,k_11_529,k_11_530,k_11_531,k_11_532,k_11_533,k_11_534,k_11_535,k_11_536,k_11_537,k_11_538,k_11_539,k_11_540,k_11_541,k_11_542,k_11_543,k_11_544,k_11_545,k_11_546,k_11_547,k_11_548,k_11_549,k_11_550,k_11_551,k_11_552,k_11_553,k_11_554,k_11_555,k_11_556,k_11_557,k_11_558,k_11_559,k_11_560,k_11_561,k_11_562,k_11_563,k_11_564,k_11_565,k_11_566,k_11_567,k_11_568,k_11_569,k_11_570,k_11_571,k_11_572,k_11_573,k_11_574,k_11_575,k_11_576,k_11_577,k_11_578,k_11_579,k_11_580,k_11_581,k_11_582,k_11_583,k_11_584,k_11_585,k_11_586,k_11_587,k_11_588,k_11_589,k_11_590,k_11_591,k_11_592,k_11_593,k_11_594,k_11_595,k_11_596,k_11_597,k_11_598,k_11_599,k_11_600,k_11_601,k_11_602,k_11_603,k_11_604,k_11_605,k_11_606,k_11_607,k_11_608,k_11_609,k_11_610,k_11_611,k_11_612,k_11_613,k_11_614,k_11_615,k_11_616,k_11_617,k_11_618,k_11_619,k_11_620,k_11_621,k_11_622,k_11_623,k_11_624,k_11_625,k_11_626,k_11_627,k_11_628,k_11_629,k_11_630,k_11_631,k_11_632,k_11_633,k_11_634,k_11_635,k_11_636,k_11_637,k_11_638,k_11_639,k_11_640,k_11_641,k_11_642,k_11_643,k_11_644,k_11_645,k_11_646,k_11_647,k_11_648,k_11_649,k_11_650,k_11_651,k_11_652,k_11_653,k_11_654,k_11_655,k_11_656,k_11_657,k_11_658,k_11_659,k_11_660,k_11_661,k_11_662,k_11_663,k_11_664,k_11_665,k_11_666,k_11_667,k_11_668,k_11_669,k_11_670,k_11_671,k_11_672,k_11_673,k_11_674,k_11_675,k_11_676,k_11_677,k_11_678,k_11_679,k_11_680,k_11_681,k_11_682,k_11_683,k_11_684,k_11_685,k_11_686,k_11_687,k_11_688,k_11_689,k_11_690,k_11_691,k_11_692,k_11_693,k_11_694,k_11_695,k_11_696,k_11_697,k_11_698,k_11_699,k_11_700,k_11_701,k_11_702,k_11_703,k_11_704,k_11_705,k_11_706,k_11_707,k_11_708,k_11_709,k_11_710,k_11_711,k_11_712,k_11_713,k_11_714,k_11_715,k_11_716,k_11_717,k_11_718,k_11_719,k_11_720,k_11_721,k_11_722,k_11_723,k_11_724,k_11_725,k_11_726,k_11_727,k_11_728,k_11_729,k_11_730,k_11_731,k_11_732,k_11_733,k_11_734,k_11_735,k_11_736,k_11_737,k_11_738,k_11_739,k_11_740,k_11_741,k_11_742,k_11_743,k_11_744,k_11_745,k_11_746,k_11_747,k_11_748,k_11_749,k_11_750,k_11_751,k_11_752,k_11_753,k_11_754,k_11_755,k_11_756,k_11_757,k_11_758,k_11_759,k_11_760,k_11_761,k_11_762,k_11_763,k_11_764,k_11_765,k_11_766,k_11_767,k_11_768,k_11_769,k_11_770,k_11_771,k_11_772,k_11_773,k_11_774,k_11_775,k_11_776,k_11_777,k_11_778,k_11_779,k_11_780,k_11_781,k_11_782,k_11_783,k_11_784,k_11_785,k_11_786,k_11_787,k_11_788,k_11_789,k_11_790,k_11_791,k_11_792,k_11_793,k_11_794,k_11_795,k_11_796,k_11_797,k_11_798,k_11_799,k_11_800,k_11_801,k_11_802,k_11_803,k_11_804,k_11_805,k_11_806,k_11_807,k_11_808,k_11_809,k_11_810,k_11_811,k_11_812,k_11_813,k_11_814,k_11_815,k_11_816,k_11_817,k_11_818,k_11_819,k_11_820,k_11_821,k_11_822,k_11_823,k_11_824,k_11_825,k_11_826,k_11_827,k_11_828,k_11_829,k_11_830,k_11_831,k_11_832,k_11_833,k_11_834,k_11_835,k_11_836,k_11_837,k_11_838,k_11_839,k_11_840,k_11_841,k_11_842,k_11_843,k_11_844,k_11_845,k_11_846,k_11_847,k_11_848,k_11_849,k_11_850,k_11_851,k_11_852,k_11_853,k_11_854,k_11_855,k_11_856,k_11_857,k_11_858,k_11_859,k_11_860,k_11_861,k_11_862,k_11_863,k_11_864,k_11_865,k_11_866,k_11_867,k_11_868,k_11_869,k_11_870,k_11_871,k_11_872,k_11_873,k_11_874,k_11_875,k_11_876,k_11_877,k_11_878,k_11_879,k_11_880,k_11_881,k_11_882,k_11_883,k_11_884,k_11_885,k_11_886,k_11_887,k_11_888,k_11_889,k_11_890,k_11_891,k_11_892,k_11_893,k_11_894,k_11_895,k_11_896,k_11_897,k_11_898,k_11_899,k_11_900,k_11_901,k_11_902,k_11_903,k_11_904,k_11_905,k_11_906,k_11_907,k_11_908,k_11_909,k_11_910,k_11_911,k_11_912,k_11_913,k_11_914,k_11_915,k_11_916,k_11_917,k_11_918,k_11_919,k_11_920,k_11_921,k_11_922,k_11_923,k_11_924,k_11_925,k_11_926,k_11_927,k_11_928,k_11_929,k_11_930,k_11_931,k_11_932,k_11_933,k_11_934,k_11_935,k_11_936,k_11_937,k_11_938,k_11_939,k_11_940,k_11_941,k_11_942,k_11_943,k_11_944,k_11_945,k_11_946,k_11_947,k_11_948,k_11_949,k_11_950,k_11_951,k_11_952,k_11_953,k_11_954,k_11_955,k_11_956,k_11_957,k_11_958,k_11_959,k_11_960,k_11_961,k_11_962,k_11_963,k_11_964,k_11_965,k_11_966,k_11_967,k_11_968,k_11_969,k_11_970,k_11_971,k_11_972,k_11_973,k_11_974,k_11_975,k_11_976,k_11_977,k_11_978,k_11_979,k_11_980,k_11_981,k_11_982,k_11_983,k_11_984,k_11_985,k_11_986,k_11_987,k_11_988,k_11_989,k_11_990,k_11_991,k_11_992,k_11_993,k_11_994,k_11_995,k_11_996,k_11_997,k_11_998,k_11_999,k_11_1000,k_11_1001,k_11_1002,k_11_1003,k_11_1004,k_11_1005,k_11_1006,k_11_1007,k_11_1008,k_11_1009,k_11_1010,k_11_1011,k_11_1012,k_11_1013,k_11_1014,k_11_1015,k_11_1016,k_11_1017,k_11_1018,k_11_1019,k_11_1020,k_11_1021,k_11_1022,k_11_1023,k_11_1024,k_11_1025,k_11_1026,k_11_1027,k_11_1028,k_11_1029,k_11_1030,k_11_1031,k_11_1032,k_11_1033,k_11_1034,k_11_1035,k_11_1036,k_11_1037,k_11_1038,k_11_1039,k_11_1040,k_11_1041,k_11_1042,k_11_1043,k_11_1044,k_11_1045,k_11_1046,k_11_1047,k_11_1048,k_11_1049,k_11_1050,k_11_1051,k_11_1052,k_11_1053,k_11_1054,k_11_1055,k_11_1056,k_11_1057,k_11_1058,k_11_1059,k_11_1060,k_11_1061,k_11_1062,k_11_1063,k_11_1064,k_11_1065,k_11_1066,k_11_1067,k_11_1068,k_11_1069,k_11_1070,k_11_1071,k_11_1072,k_11_1073,k_11_1074,k_11_1075,k_11_1076,k_11_1077,k_11_1078,k_11_1079,k_11_1080,k_11_1081,k_11_1082,k_11_1083,k_11_1084,k_11_1085,k_11_1086,k_11_1087,k_11_1088,k_11_1089,k_11_1090,k_11_1091,k_11_1092,k_11_1093,k_11_1094,k_11_1095,k_11_1096,k_11_1097,k_11_1098,k_11_1099,k_11_1100,k_11_1101,k_11_1102,k_11_1103,k_11_1104,k_11_1105,k_11_1106,k_11_1107,k_11_1108,k_11_1109,k_11_1110,k_11_1111,k_11_1112,k_11_1113,k_11_1114,k_11_1115,k_11_1116,k_11_1117,k_11_1118,k_11_1119,k_11_1120,k_11_1121,k_11_1122,k_11_1123,k_11_1124,k_11_1125,k_11_1126,k_11_1127,k_11_1128,k_11_1129,k_11_1130,k_11_1131,k_11_1132,k_11_1133,k_11_1134,k_11_1135,k_11_1136,k_11_1137,k_11_1138,k_11_1139,k_11_1140,k_11_1141,k_11_1142,k_11_1143,k_11_1144,k_11_1145,k_11_1146,k_11_1147,k_11_1148,k_11_1149,k_11_1150,k_11_1151,k_11_1152,k_11_1153,k_11_1154,k_11_1155,k_11_1156,k_11_1157,k_11_1158,k_11_1159,k_11_1160,k_11_1161,k_11_1162,k_11_1163,k_11_1164,k_11_1165,k_11_1166,k_11_1167,k_11_1168,k_11_1169,k_11_1170,k_11_1171,k_11_1172,k_11_1173,k_11_1174,k_11_1175,k_11_1176,k_11_1177,k_11_1178,k_11_1179,k_11_1180,k_11_1181,k_11_1182,k_11_1183,k_11_1184,k_11_1185,k_11_1186,k_11_1187,k_11_1188,k_11_1189,k_11_1190,k_11_1191,k_11_1192,k_11_1193,k_11_1194,k_11_1195,k_11_1196,k_11_1197,k_11_1198,k_11_1199,k_11_1200,k_11_1201,k_11_1202,k_11_1203,k_11_1204,k_11_1205,k_11_1206,k_11_1207,k_11_1208,k_11_1209,k_11_1210,k_11_1211,k_11_1212,k_11_1213,k_11_1214,k_11_1215,k_11_1216,k_11_1217,k_11_1218,k_11_1219,k_11_1220,k_11_1221,k_11_1222,k_11_1223,k_11_1224,k_11_1225,k_11_1226,k_11_1227,k_11_1228,k_11_1229,k_11_1230,k_11_1231,k_11_1232,k_11_1233,k_11_1234,k_11_1235,k_11_1236,k_11_1237,k_11_1238,k_11_1239,k_11_1240,k_11_1241,k_11_1242,k_11_1243,k_11_1244,k_11_1245,k_11_1246,k_11_1247,k_11_1248,k_11_1249,k_11_1250,k_11_1251,k_11_1252,k_11_1253,k_11_1254,k_11_1255,k_11_1256,k_11_1257,k_11_1258,k_11_1259,k_11_1260,k_11_1261,k_11_1262,k_11_1263,k_11_1264,k_11_1265,k_11_1266,k_11_1267,k_11_1268,k_11_1269,k_11_1270,k_11_1271,k_11_1272,k_11_1273,k_11_1274,k_11_1275,k_11_1276,k_11_1277,k_11_1278,k_11_1279,k_11_1280,k_11_1281,k_11_1282,k_11_1283,k_11_1284,k_11_1285,k_11_1286,k_11_1287,k_11_1288,k_11_1289,k_11_1290,k_11_1291,k_11_1292,k_11_1293,k_11_1294,k_11_1295,k_11_1296,k_11_1297,k_11_1298,k_11_1299,k_11_1300,k_11_1301,k_11_1302,k_11_1303,k_11_1304,k_11_1305,k_11_1306,k_11_1307,k_11_1308,k_11_1309,k_11_1310,k_11_1311,k_11_1312,k_11_1313,k_11_1314,k_11_1315,k_11_1316,k_11_1317,k_11_1318,k_11_1319,k_11_1320,k_11_1321,k_11_1322,k_11_1323,k_11_1324,k_11_1325,k_11_1326,k_11_1327,k_11_1328,k_11_1329,k_11_1330,k_11_1331,k_11_1332,k_11_1333,k_11_1334,k_11_1335,k_11_1336,k_11_1337,k_11_1338,k_11_1339,k_11_1340,k_11_1341,k_11_1342,k_11_1343,k_11_1344,k_11_1345,k_11_1346,k_11_1347,k_11_1348,k_11_1349,k_11_1350,k_11_1351,k_11_1352,k_11_1353,k_11_1354,k_11_1355,k_11_1356,k_11_1357,k_11_1358,k_11_1359,k_11_1360,k_11_1361,k_11_1362,k_11_1363,k_11_1364,k_11_1365,k_11_1366,k_11_1367,k_11_1368,k_11_1369,k_11_1370,k_11_1371,k_11_1372,k_11_1373,k_11_1374,k_11_1375,k_11_1376,k_11_1377,k_11_1378,k_11_1379,k_11_1380,k_11_1381,k_11_1382,k_11_1383,k_11_1384,k_11_1385,k_11_1386,k_11_1387,k_11_1388,k_11_1389,k_11_1390,k_11_1391,k_11_1392,k_11_1393,k_11_1394,k_11_1395,k_11_1396,k_11_1397,k_11_1398,k_11_1399,k_11_1400,k_11_1401,k_11_1402,k_11_1403,k_11_1404,k_11_1405,k_11_1406,k_11_1407,k_11_1408,k_11_1409,k_11_1410,k_11_1411,k_11_1412,k_11_1413,k_11_1414,k_11_1415,k_11_1416,k_11_1417,k_11_1418,k_11_1419,k_11_1420,k_11_1421,k_11_1422,k_11_1423,k_11_1424,k_11_1425,k_11_1426,k_11_1427,k_11_1428,k_11_1429,k_11_1430,k_11_1431,k_11_1432,k_11_1433,k_11_1434,k_11_1435,k_11_1436,k_11_1437,k_11_1438,k_11_1439,k_11_1440,k_11_1441,k_11_1442,k_11_1443,k_11_1444,k_11_1445,k_11_1446,k_11_1447,k_11_1448,k_11_1449,k_11_1450,k_11_1451,k_11_1452,k_11_1453,k_11_1454,k_11_1455,k_11_1456,k_11_1457,k_11_1458,k_11_1459,k_11_1460,k_11_1461,k_11_1462,k_11_1463,k_11_1464,k_11_1465,k_11_1466,k_11_1467,k_11_1468,k_11_1469,k_11_1470,k_11_1471,k_11_1472,k_11_1473,k_11_1474,k_11_1475,k_11_1476,k_11_1477,k_11_1478,k_11_1479,k_11_1480,k_11_1481,k_11_1482,k_11_1483,k_11_1484,k_11_1485,k_11_1486,k_11_1487,k_11_1488,k_11_1489,k_11_1490,k_11_1491,k_11_1492,k_11_1493,k_11_1494,k_11_1495,k_11_1496,k_11_1497,k_11_1498,k_11_1499,k_11_1500,k_11_1501,k_11_1502,k_11_1503,k_11_1504,k_11_1505,k_11_1506,k_11_1507,k_11_1508,k_11_1509,k_11_1510,k_11_1511,k_11_1512,k_11_1513,k_11_1514,k_11_1515,k_11_1516,k_11_1517,k_11_1518,k_11_1519,k_11_1520,k_11_1521,k_11_1522,k_11_1523,k_11_1524,k_11_1525,k_11_1526,k_11_1527,k_11_1528,k_11_1529,k_11_1530,k_11_1531,k_11_1532,k_11_1533,k_11_1534,k_11_1535,k_11_1536,k_11_1537,k_11_1538,k_11_1539,k_11_1540,k_11_1541,k_11_1542,k_11_1543,k_11_1544,k_11_1545,k_11_1546,k_11_1547,k_11_1548,k_11_1549,k_11_1550,k_11_1551,k_11_1552,k_11_1553,k_11_1554,k_11_1555,k_11_1556,k_11_1557,k_11_1558,k_11_1559,k_11_1560,k_11_1561,k_11_1562,k_11_1563,k_11_1564,k_11_1565,k_11_1566,k_11_1567,k_11_1568,k_11_1569,k_11_1570,k_11_1571,k_11_1572,k_11_1573,k_11_1574,k_11_1575,k_11_1576,k_11_1577,k_11_1578,k_11_1579,k_11_1580,k_11_1581,k_11_1582,k_11_1583,k_11_1584,k_11_1585,k_11_1586,k_11_1587,k_11_1588,k_11_1589,k_11_1590,k_11_1591,k_11_1592,k_11_1593,k_11_1594,k_11_1595,k_11_1596,k_11_1597,k_11_1598,k_11_1599,k_11_1600,k_11_1601,k_11_1602,k_11_1603,k_11_1604,k_11_1605,k_11_1606,k_11_1607,k_11_1608,k_11_1609,k_11_1610,k_11_1611,k_11_1612,k_11_1613,k_11_1614,k_11_1615,k_11_1616,k_11_1617,k_11_1618,k_11_1619,k_11_1620,k_11_1621,k_11_1622,k_11_1623,k_11_1624,k_11_1625,k_11_1626,k_11_1627,k_11_1628,k_11_1629,k_11_1630,k_11_1631,k_11_1632,k_11_1633,k_11_1634,k_11_1635,k_11_1636,k_11_1637,k_11_1638,k_11_1639,k_11_1640,k_11_1641,k_11_1642,k_11_1643,k_11_1644,k_11_1645,k_11_1646,k_11_1647,k_11_1648,k_11_1649,k_11_1650,k_11_1651,k_11_1652,k_11_1653,k_11_1654,k_11_1655,k_11_1656,k_11_1657,k_11_1658,k_11_1659,k_11_1660,k_11_1661,k_11_1662,k_11_1663,k_11_1664,k_11_1665,k_11_1666,k_11_1667,k_11_1668,k_11_1669,k_11_1670,k_11_1671,k_11_1672,k_11_1673,k_11_1674,k_11_1675,k_11_1676,k_11_1677,k_11_1678,k_11_1679,k_11_1680,k_11_1681,k_11_1682,k_11_1683,k_11_1684,k_11_1685,k_11_1686,k_11_1687,k_11_1688,k_11_1689,k_11_1690,k_11_1691,k_11_1692,k_11_1693,k_11_1694,k_11_1695,k_11_1696,k_11_1697,k_11_1698,k_11_1699,k_11_1700,k_11_1701,k_11_1702,k_11_1703,k_11_1704,k_11_1705,k_11_1706,k_11_1707,k_11_1708,k_11_1709,k_11_1710,k_11_1711,k_11_1712,k_11_1713,k_11_1714,k_11_1715,k_11_1716,k_11_1717,k_11_1718,k_11_1719,k_11_1720,k_11_1721,k_11_1722,k_11_1723,k_11_1724,k_11_1725,k_11_1726,k_11_1727,k_11_1728,k_11_1729,k_11_1730,k_11_1731,k_11_1732,k_11_1733,k_11_1734,k_11_1735,k_11_1736,k_11_1737,k_11_1738,k_11_1739,k_11_1740,k_11_1741,k_11_1742,k_11_1743,k_11_1744,k_11_1745,k_11_1746,k_11_1747,k_11_1748,k_11_1749,k_11_1750,k_11_1751,k_11_1752,k_11_1753,k_11_1754,k_11_1755,k_11_1756,k_11_1757,k_11_1758,k_11_1759,k_11_1760,k_11_1761,k_11_1762,k_11_1763,k_11_1764,k_11_1765,k_11_1766,k_11_1767,k_11_1768,k_11_1769,k_11_1770,k_11_1771,k_11_1772,k_11_1773,k_11_1774,k_11_1775,k_11_1776,k_11_1777,k_11_1778,k_11_1779,k_11_1780,k_11_1781,k_11_1782,k_11_1783,k_11_1784,k_11_1785,k_11_1786,k_11_1787,k_11_1788,k_11_1789,k_11_1790,k_11_1791,k_11_1792,k_11_1793,k_11_1794,k_11_1795,k_11_1796,k_11_1797,k_11_1798,k_11_1799,k_11_1800,k_11_1801,k_11_1802,k_11_1803,k_11_1804,k_11_1805,k_11_1806,k_11_1807,k_11_1808,k_11_1809,k_11_1810,k_11_1811,k_11_1812,k_11_1813,k_11_1814,k_11_1815,k_11_1816,k_11_1817,k_11_1818,k_11_1819,k_11_1820,k_11_1821,k_11_1822,k_11_1823,k_11_1824,k_11_1825,k_11_1826,k_11_1827,k_11_1828,k_11_1829,k_11_1830,k_11_1831,k_11_1832,k_11_1833,k_11_1834,k_11_1835,k_11_1836,k_11_1837,k_11_1838,k_11_1839,k_11_1840,k_11_1841,k_11_1842,k_11_1843,k_11_1844,k_11_1845,k_11_1846,k_11_1847,k_11_1848,k_11_1849,k_11_1850,k_11_1851,k_11_1852,k_11_1853,k_11_1854,k_11_1855,k_11_1856,k_11_1857,k_11_1858,k_11_1859,k_11_1860,k_11_1861,k_11_1862,k_11_1863,k_11_1864,k_11_1865,k_11_1866,k_11_1867,k_11_1868,k_11_1869,k_11_1870,k_11_1871,k_11_1872,k_11_1873,k_11_1874,k_11_1875,k_11_1876,k_11_1877,k_11_1878,k_11_1879,k_11_1880,k_11_1881,k_11_1882,k_11_1883,k_11_1884,k_11_1885,k_11_1886,k_11_1887,k_11_1888,k_11_1889,k_11_1890,k_11_1891,k_11_1892,k_11_1893,k_11_1894,k_11_1895,k_11_1896,k_11_1897,k_11_1898,k_11_1899,k_11_1900,k_11_1901,k_11_1902,k_11_1903,k_11_1904,k_11_1905,k_11_1906,k_11_1907,k_11_1908,k_11_1909,k_11_1910,k_11_1911,k_11_1912,k_11_1913,k_11_1914,k_11_1915,k_11_1916,k_11_1917,k_11_1918,k_11_1919,k_11_1920,k_11_1921,k_11_1922,k_11_1923,k_11_1924,k_11_1925,k_11_1926,k_11_1927,k_11_1928,k_11_1929,k_11_1930,k_11_1931,k_11_1932,k_11_1933,k_11_1934,k_11_1935,k_11_1936,k_11_1937,k_11_1938,k_11_1939,k_11_1940,k_11_1941,k_11_1942,k_11_1943,k_11_1944,k_11_1945,k_11_1946,k_11_1947,k_11_1948,k_11_1949,k_11_1950,k_11_1951,k_11_1952,k_11_1953,k_11_1954,k_11_1955,k_11_1956,k_11_1957,k_11_1958,k_11_1959,k_11_1960,k_11_1961,k_11_1962,k_11_1963,k_11_1964,k_11_1965,k_11_1966,k_11_1967,k_11_1968,k_11_1969,k_11_1970,k_11_1971,k_11_1972,k_11_1973,k_11_1974,k_11_1975,k_11_1976,k_11_1977,k_11_1978,k_11_1979,k_11_1980,k_11_1981,k_11_1982,k_11_1983,k_11_1984,k_11_1985,k_11_1986,k_11_1987,k_11_1988,k_11_1989,k_11_1990,k_11_1991,k_11_1992,k_11_1993,k_11_1994,k_11_1995,k_11_1996,k_11_1997,k_11_1998,k_11_1999,k_11_2000,k_11_2001,k_11_2002,k_11_2003,k_11_2004,k_11_2005,k_11_2006,k_11_2007,k_11_2008,k_11_2009,k_11_2010,k_11_2011,k_11_2012,k_11_2013,k_11_2014,k_11_2015,k_11_2016,k_11_2017,k_11_2018,k_11_2019,k_11_2020,k_11_2021,k_11_2022,k_11_2023,k_11_2024,k_11_2025,k_11_2026,k_11_2027,k_11_2028,k_11_2029,k_11_2030,k_11_2031,k_11_2032,k_11_2033,k_11_2034,k_11_2035,k_11_2036,k_11_2037,k_11_2038,k_11_2039,k_11_2040,k_11_2041,k_11_2042,k_11_2043,k_11_2044,k_11_2045,k_11_2046,k_11_2047;
valve v_1_0 (.fluid_in(k_1_0), .fluid_out(k_0_0), .air_in(c_1_0));
valve v_1_1 (.fluid_in(k_1_1), .fluid_out(k_0_0), .air_in(c_1_1));
valve v_2_0 (.fluid_in(k_2_0), .fluid_out(k_1_0), .air_in(c_2_0));
valve v_2_1 (.fluid_in(k_2_1), .fluid_out(k_1_0), .air_in(c_2_1));
valve v_2_2 (.fluid_in(k_2_2), .fluid_out(k_1_1), .air_in(c_2_0));
valve v_2_3 (.fluid_in(k_2_3), .fluid_out(k_1_1), .air_in(c_2_1));
valve v_3_0 (.fluid_in(k_3_0), .fluid_out(k_2_0), .air_in(c_3_0));
valve v_3_1 (.fluid_in(k_3_1), .fluid_out(k_2_0), .air_in(c_3_1));
valve v_3_2 (.fluid_in(k_3_2), .fluid_out(k_2_1), .air_in(c_3_0));
valve v_3_3 (.fluid_in(k_3_3), .fluid_out(k_2_1), .air_in(c_3_1));
valve v_3_4 (.fluid_in(k_3_4), .fluid_out(k_2_2), .air_in(c_3_0));
valve v_3_5 (.fluid_in(k_3_5), .fluid_out(k_2_2), .air_in(c_3_1));
valve v_3_6 (.fluid_in(k_3_6), .fluid_out(k_2_3), .air_in(c_3_0));
valve v_3_7 (.fluid_in(k_3_7), .fluid_out(k_2_3), .air_in(c_3_1));
valve v_4_0 (.fluid_in(k_4_0), .fluid_out(k_3_0), .air_in(c_4_0));
valve v_4_1 (.fluid_in(k_4_1), .fluid_out(k_3_0), .air_in(c_4_1));
valve v_4_2 (.fluid_in(k_4_2), .fluid_out(k_3_1), .air_in(c_4_0));
valve v_4_3 (.fluid_in(k_4_3), .fluid_out(k_3_1), .air_in(c_4_1));
valve v_4_4 (.fluid_in(k_4_4), .fluid_out(k_3_2), .air_in(c_4_0));
valve v_4_5 (.fluid_in(k_4_5), .fluid_out(k_3_2), .air_in(c_4_1));
valve v_4_6 (.fluid_in(k_4_6), .fluid_out(k_3_3), .air_in(c_4_0));
valve v_4_7 (.fluid_in(k_4_7), .fluid_out(k_3_3), .air_in(c_4_1));
valve v_4_8 (.fluid_in(k_4_8), .fluid_out(k_3_4), .air_in(c_4_0));
valve v_4_9 (.fluid_in(k_4_9), .fluid_out(k_3_4), .air_in(c_4_1));
valve v_4_10 (.fluid_in(k_4_10), .fluid_out(k_3_5), .air_in(c_4_0));
valve v_4_11 (.fluid_in(k_4_11), .fluid_out(k_3_5), .air_in(c_4_1));
valve v_4_12 (.fluid_in(k_4_12), .fluid_out(k_3_6), .air_in(c_4_0));
valve v_4_13 (.fluid_in(k_4_13), .fluid_out(k_3_6), .air_in(c_4_1));
valve v_4_14 (.fluid_in(k_4_14), .fluid_out(k_3_7), .air_in(c_4_0));
valve v_4_15 (.fluid_in(k_4_15), .fluid_out(k_3_7), .air_in(c_4_1));
valve v_5_0 (.fluid_in(k_5_0), .fluid_out(k_4_0), .air_in(c_5_0));
valve v_5_1 (.fluid_in(k_5_1), .fluid_out(k_4_0), .air_in(c_5_1));
valve v_5_2 (.fluid_in(k_5_2), .fluid_out(k_4_1), .air_in(c_5_0));
valve v_5_3 (.fluid_in(k_5_3), .fluid_out(k_4_1), .air_in(c_5_1));
valve v_5_4 (.fluid_in(k_5_4), .fluid_out(k_4_2), .air_in(c_5_0));
valve v_5_5 (.fluid_in(k_5_5), .fluid_out(k_4_2), .air_in(c_5_1));
valve v_5_6 (.fluid_in(k_5_6), .fluid_out(k_4_3), .air_in(c_5_0));
valve v_5_7 (.fluid_in(k_5_7), .fluid_out(k_4_3), .air_in(c_5_1));
valve v_5_8 (.fluid_in(k_5_8), .fluid_out(k_4_4), .air_in(c_5_0));
valve v_5_9 (.fluid_in(k_5_9), .fluid_out(k_4_4), .air_in(c_5_1));
valve v_5_10 (.fluid_in(k_5_10), .fluid_out(k_4_5), .air_in(c_5_0));
valve v_5_11 (.fluid_in(k_5_11), .fluid_out(k_4_5), .air_in(c_5_1));
valve v_5_12 (.fluid_in(k_5_12), .fluid_out(k_4_6), .air_in(c_5_0));
valve v_5_13 (.fluid_in(k_5_13), .fluid_out(k_4_6), .air_in(c_5_1));
valve v_5_14 (.fluid_in(k_5_14), .fluid_out(k_4_7), .air_in(c_5_0));
valve v_5_15 (.fluid_in(k_5_15), .fluid_out(k_4_7), .air_in(c_5_1));
valve v_5_16 (.fluid_in(k_5_16), .fluid_out(k_4_8), .air_in(c_5_0));
valve v_5_17 (.fluid_in(k_5_17), .fluid_out(k_4_8), .air_in(c_5_1));
valve v_5_18 (.fluid_in(k_5_18), .fluid_out(k_4_9), .air_in(c_5_0));
valve v_5_19 (.fluid_in(k_5_19), .fluid_out(k_4_9), .air_in(c_5_1));
valve v_5_20 (.fluid_in(k_5_20), .fluid_out(k_4_10), .air_in(c_5_0));
valve v_5_21 (.fluid_in(k_5_21), .fluid_out(k_4_10), .air_in(c_5_1));
valve v_5_22 (.fluid_in(k_5_22), .fluid_out(k_4_11), .air_in(c_5_0));
valve v_5_23 (.fluid_in(k_5_23), .fluid_out(k_4_11), .air_in(c_5_1));
valve v_5_24 (.fluid_in(k_5_24), .fluid_out(k_4_12), .air_in(c_5_0));
valve v_5_25 (.fluid_in(k_5_25), .fluid_out(k_4_12), .air_in(c_5_1));
valve v_5_26 (.fluid_in(k_5_26), .fluid_out(k_4_13), .air_in(c_5_0));
valve v_5_27 (.fluid_in(k_5_27), .fluid_out(k_4_13), .air_in(c_5_1));
valve v_5_28 (.fluid_in(k_5_28), .fluid_out(k_4_14), .air_in(c_5_0));
valve v_5_29 (.fluid_in(k_5_29), .fluid_out(k_4_14), .air_in(c_5_1));
valve v_5_30 (.fluid_in(k_5_30), .fluid_out(k_4_15), .air_in(c_5_0));
valve v_5_31 (.fluid_in(k_5_31), .fluid_out(k_4_15), .air_in(c_5_1));
valve v_6_0 (.fluid_in(k_6_0), .fluid_out(k_5_0), .air_in(c_6_0));
valve v_6_1 (.fluid_in(k_6_1), .fluid_out(k_5_0), .air_in(c_6_1));
valve v_6_2 (.fluid_in(k_6_2), .fluid_out(k_5_1), .air_in(c_6_0));
valve v_6_3 (.fluid_in(k_6_3), .fluid_out(k_5_1), .air_in(c_6_1));
valve v_6_4 (.fluid_in(k_6_4), .fluid_out(k_5_2), .air_in(c_6_0));
valve v_6_5 (.fluid_in(k_6_5), .fluid_out(k_5_2), .air_in(c_6_1));
valve v_6_6 (.fluid_in(k_6_6), .fluid_out(k_5_3), .air_in(c_6_0));
valve v_6_7 (.fluid_in(k_6_7), .fluid_out(k_5_3), .air_in(c_6_1));
valve v_6_8 (.fluid_in(k_6_8), .fluid_out(k_5_4), .air_in(c_6_0));
valve v_6_9 (.fluid_in(k_6_9), .fluid_out(k_5_4), .air_in(c_6_1));
valve v_6_10 (.fluid_in(k_6_10), .fluid_out(k_5_5), .air_in(c_6_0));
valve v_6_11 (.fluid_in(k_6_11), .fluid_out(k_5_5), .air_in(c_6_1));
valve v_6_12 (.fluid_in(k_6_12), .fluid_out(k_5_6), .air_in(c_6_0));
valve v_6_13 (.fluid_in(k_6_13), .fluid_out(k_5_6), .air_in(c_6_1));
valve v_6_14 (.fluid_in(k_6_14), .fluid_out(k_5_7), .air_in(c_6_0));
valve v_6_15 (.fluid_in(k_6_15), .fluid_out(k_5_7), .air_in(c_6_1));
valve v_6_16 (.fluid_in(k_6_16), .fluid_out(k_5_8), .air_in(c_6_0));
valve v_6_17 (.fluid_in(k_6_17), .fluid_out(k_5_8), .air_in(c_6_1));
valve v_6_18 (.fluid_in(k_6_18), .fluid_out(k_5_9), .air_in(c_6_0));
valve v_6_19 (.fluid_in(k_6_19), .fluid_out(k_5_9), .air_in(c_6_1));
valve v_6_20 (.fluid_in(k_6_20), .fluid_out(k_5_10), .air_in(c_6_0));
valve v_6_21 (.fluid_in(k_6_21), .fluid_out(k_5_10), .air_in(c_6_1));
valve v_6_22 (.fluid_in(k_6_22), .fluid_out(k_5_11), .air_in(c_6_0));
valve v_6_23 (.fluid_in(k_6_23), .fluid_out(k_5_11), .air_in(c_6_1));
valve v_6_24 (.fluid_in(k_6_24), .fluid_out(k_5_12), .air_in(c_6_0));
valve v_6_25 (.fluid_in(k_6_25), .fluid_out(k_5_12), .air_in(c_6_1));
valve v_6_26 (.fluid_in(k_6_26), .fluid_out(k_5_13), .air_in(c_6_0));
valve v_6_27 (.fluid_in(k_6_27), .fluid_out(k_5_13), .air_in(c_6_1));
valve v_6_28 (.fluid_in(k_6_28), .fluid_out(k_5_14), .air_in(c_6_0));
valve v_6_29 (.fluid_in(k_6_29), .fluid_out(k_5_14), .air_in(c_6_1));
valve v_6_30 (.fluid_in(k_6_30), .fluid_out(k_5_15), .air_in(c_6_0));
valve v_6_31 (.fluid_in(k_6_31), .fluid_out(k_5_15), .air_in(c_6_1));
valve v_6_32 (.fluid_in(k_6_32), .fluid_out(k_5_16), .air_in(c_6_0));
valve v_6_33 (.fluid_in(k_6_33), .fluid_out(k_5_16), .air_in(c_6_1));
valve v_6_34 (.fluid_in(k_6_34), .fluid_out(k_5_17), .air_in(c_6_0));
valve v_6_35 (.fluid_in(k_6_35), .fluid_out(k_5_17), .air_in(c_6_1));
valve v_6_36 (.fluid_in(k_6_36), .fluid_out(k_5_18), .air_in(c_6_0));
valve v_6_37 (.fluid_in(k_6_37), .fluid_out(k_5_18), .air_in(c_6_1));
valve v_6_38 (.fluid_in(k_6_38), .fluid_out(k_5_19), .air_in(c_6_0));
valve v_6_39 (.fluid_in(k_6_39), .fluid_out(k_5_19), .air_in(c_6_1));
valve v_6_40 (.fluid_in(k_6_40), .fluid_out(k_5_20), .air_in(c_6_0));
valve v_6_41 (.fluid_in(k_6_41), .fluid_out(k_5_20), .air_in(c_6_1));
valve v_6_42 (.fluid_in(k_6_42), .fluid_out(k_5_21), .air_in(c_6_0));
valve v_6_43 (.fluid_in(k_6_43), .fluid_out(k_5_21), .air_in(c_6_1));
valve v_6_44 (.fluid_in(k_6_44), .fluid_out(k_5_22), .air_in(c_6_0));
valve v_6_45 (.fluid_in(k_6_45), .fluid_out(k_5_22), .air_in(c_6_1));
valve v_6_46 (.fluid_in(k_6_46), .fluid_out(k_5_23), .air_in(c_6_0));
valve v_6_47 (.fluid_in(k_6_47), .fluid_out(k_5_23), .air_in(c_6_1));
valve v_6_48 (.fluid_in(k_6_48), .fluid_out(k_5_24), .air_in(c_6_0));
valve v_6_49 (.fluid_in(k_6_49), .fluid_out(k_5_24), .air_in(c_6_1));
valve v_6_50 (.fluid_in(k_6_50), .fluid_out(k_5_25), .air_in(c_6_0));
valve v_6_51 (.fluid_in(k_6_51), .fluid_out(k_5_25), .air_in(c_6_1));
valve v_6_52 (.fluid_in(k_6_52), .fluid_out(k_5_26), .air_in(c_6_0));
valve v_6_53 (.fluid_in(k_6_53), .fluid_out(k_5_26), .air_in(c_6_1));
valve v_6_54 (.fluid_in(k_6_54), .fluid_out(k_5_27), .air_in(c_6_0));
valve v_6_55 (.fluid_in(k_6_55), .fluid_out(k_5_27), .air_in(c_6_1));
valve v_6_56 (.fluid_in(k_6_56), .fluid_out(k_5_28), .air_in(c_6_0));
valve v_6_57 (.fluid_in(k_6_57), .fluid_out(k_5_28), .air_in(c_6_1));
valve v_6_58 (.fluid_in(k_6_58), .fluid_out(k_5_29), .air_in(c_6_0));
valve v_6_59 (.fluid_in(k_6_59), .fluid_out(k_5_29), .air_in(c_6_1));
valve v_6_60 (.fluid_in(k_6_60), .fluid_out(k_5_30), .air_in(c_6_0));
valve v_6_61 (.fluid_in(k_6_61), .fluid_out(k_5_30), .air_in(c_6_1));
valve v_6_62 (.fluid_in(k_6_62), .fluid_out(k_5_31), .air_in(c_6_0));
valve v_6_63 (.fluid_in(k_6_63), .fluid_out(k_5_31), .air_in(c_6_1));
valve v_7_0 (.fluid_in(k_7_0), .fluid_out(k_6_0), .air_in(c_7_0));
valve v_7_1 (.fluid_in(k_7_1), .fluid_out(k_6_0), .air_in(c_7_1));
valve v_7_2 (.fluid_in(k_7_2), .fluid_out(k_6_1), .air_in(c_7_0));
valve v_7_3 (.fluid_in(k_7_3), .fluid_out(k_6_1), .air_in(c_7_1));
valve v_7_4 (.fluid_in(k_7_4), .fluid_out(k_6_2), .air_in(c_7_0));
valve v_7_5 (.fluid_in(k_7_5), .fluid_out(k_6_2), .air_in(c_7_1));
valve v_7_6 (.fluid_in(k_7_6), .fluid_out(k_6_3), .air_in(c_7_0));
valve v_7_7 (.fluid_in(k_7_7), .fluid_out(k_6_3), .air_in(c_7_1));
valve v_7_8 (.fluid_in(k_7_8), .fluid_out(k_6_4), .air_in(c_7_0));
valve v_7_9 (.fluid_in(k_7_9), .fluid_out(k_6_4), .air_in(c_7_1));
valve v_7_10 (.fluid_in(k_7_10), .fluid_out(k_6_5), .air_in(c_7_0));
valve v_7_11 (.fluid_in(k_7_11), .fluid_out(k_6_5), .air_in(c_7_1));
valve v_7_12 (.fluid_in(k_7_12), .fluid_out(k_6_6), .air_in(c_7_0));
valve v_7_13 (.fluid_in(k_7_13), .fluid_out(k_6_6), .air_in(c_7_1));
valve v_7_14 (.fluid_in(k_7_14), .fluid_out(k_6_7), .air_in(c_7_0));
valve v_7_15 (.fluid_in(k_7_15), .fluid_out(k_6_7), .air_in(c_7_1));
valve v_7_16 (.fluid_in(k_7_16), .fluid_out(k_6_8), .air_in(c_7_0));
valve v_7_17 (.fluid_in(k_7_17), .fluid_out(k_6_8), .air_in(c_7_1));
valve v_7_18 (.fluid_in(k_7_18), .fluid_out(k_6_9), .air_in(c_7_0));
valve v_7_19 (.fluid_in(k_7_19), .fluid_out(k_6_9), .air_in(c_7_1));
valve v_7_20 (.fluid_in(k_7_20), .fluid_out(k_6_10), .air_in(c_7_0));
valve v_7_21 (.fluid_in(k_7_21), .fluid_out(k_6_10), .air_in(c_7_1));
valve v_7_22 (.fluid_in(k_7_22), .fluid_out(k_6_11), .air_in(c_7_0));
valve v_7_23 (.fluid_in(k_7_23), .fluid_out(k_6_11), .air_in(c_7_1));
valve v_7_24 (.fluid_in(k_7_24), .fluid_out(k_6_12), .air_in(c_7_0));
valve v_7_25 (.fluid_in(k_7_25), .fluid_out(k_6_12), .air_in(c_7_1));
valve v_7_26 (.fluid_in(k_7_26), .fluid_out(k_6_13), .air_in(c_7_0));
valve v_7_27 (.fluid_in(k_7_27), .fluid_out(k_6_13), .air_in(c_7_1));
valve v_7_28 (.fluid_in(k_7_28), .fluid_out(k_6_14), .air_in(c_7_0));
valve v_7_29 (.fluid_in(k_7_29), .fluid_out(k_6_14), .air_in(c_7_1));
valve v_7_30 (.fluid_in(k_7_30), .fluid_out(k_6_15), .air_in(c_7_0));
valve v_7_31 (.fluid_in(k_7_31), .fluid_out(k_6_15), .air_in(c_7_1));
valve v_7_32 (.fluid_in(k_7_32), .fluid_out(k_6_16), .air_in(c_7_0));
valve v_7_33 (.fluid_in(k_7_33), .fluid_out(k_6_16), .air_in(c_7_1));
valve v_7_34 (.fluid_in(k_7_34), .fluid_out(k_6_17), .air_in(c_7_0));
valve v_7_35 (.fluid_in(k_7_35), .fluid_out(k_6_17), .air_in(c_7_1));
valve v_7_36 (.fluid_in(k_7_36), .fluid_out(k_6_18), .air_in(c_7_0));
valve v_7_37 (.fluid_in(k_7_37), .fluid_out(k_6_18), .air_in(c_7_1));
valve v_7_38 (.fluid_in(k_7_38), .fluid_out(k_6_19), .air_in(c_7_0));
valve v_7_39 (.fluid_in(k_7_39), .fluid_out(k_6_19), .air_in(c_7_1));
valve v_7_40 (.fluid_in(k_7_40), .fluid_out(k_6_20), .air_in(c_7_0));
valve v_7_41 (.fluid_in(k_7_41), .fluid_out(k_6_20), .air_in(c_7_1));
valve v_7_42 (.fluid_in(k_7_42), .fluid_out(k_6_21), .air_in(c_7_0));
valve v_7_43 (.fluid_in(k_7_43), .fluid_out(k_6_21), .air_in(c_7_1));
valve v_7_44 (.fluid_in(k_7_44), .fluid_out(k_6_22), .air_in(c_7_0));
valve v_7_45 (.fluid_in(k_7_45), .fluid_out(k_6_22), .air_in(c_7_1));
valve v_7_46 (.fluid_in(k_7_46), .fluid_out(k_6_23), .air_in(c_7_0));
valve v_7_47 (.fluid_in(k_7_47), .fluid_out(k_6_23), .air_in(c_7_1));
valve v_7_48 (.fluid_in(k_7_48), .fluid_out(k_6_24), .air_in(c_7_0));
valve v_7_49 (.fluid_in(k_7_49), .fluid_out(k_6_24), .air_in(c_7_1));
valve v_7_50 (.fluid_in(k_7_50), .fluid_out(k_6_25), .air_in(c_7_0));
valve v_7_51 (.fluid_in(k_7_51), .fluid_out(k_6_25), .air_in(c_7_1));
valve v_7_52 (.fluid_in(k_7_52), .fluid_out(k_6_26), .air_in(c_7_0));
valve v_7_53 (.fluid_in(k_7_53), .fluid_out(k_6_26), .air_in(c_7_1));
valve v_7_54 (.fluid_in(k_7_54), .fluid_out(k_6_27), .air_in(c_7_0));
valve v_7_55 (.fluid_in(k_7_55), .fluid_out(k_6_27), .air_in(c_7_1));
valve v_7_56 (.fluid_in(k_7_56), .fluid_out(k_6_28), .air_in(c_7_0));
valve v_7_57 (.fluid_in(k_7_57), .fluid_out(k_6_28), .air_in(c_7_1));
valve v_7_58 (.fluid_in(k_7_58), .fluid_out(k_6_29), .air_in(c_7_0));
valve v_7_59 (.fluid_in(k_7_59), .fluid_out(k_6_29), .air_in(c_7_1));
valve v_7_60 (.fluid_in(k_7_60), .fluid_out(k_6_30), .air_in(c_7_0));
valve v_7_61 (.fluid_in(k_7_61), .fluid_out(k_6_30), .air_in(c_7_1));
valve v_7_62 (.fluid_in(k_7_62), .fluid_out(k_6_31), .air_in(c_7_0));
valve v_7_63 (.fluid_in(k_7_63), .fluid_out(k_6_31), .air_in(c_7_1));
valve v_7_64 (.fluid_in(k_7_64), .fluid_out(k_6_32), .air_in(c_7_0));
valve v_7_65 (.fluid_in(k_7_65), .fluid_out(k_6_32), .air_in(c_7_1));
valve v_7_66 (.fluid_in(k_7_66), .fluid_out(k_6_33), .air_in(c_7_0));
valve v_7_67 (.fluid_in(k_7_67), .fluid_out(k_6_33), .air_in(c_7_1));
valve v_7_68 (.fluid_in(k_7_68), .fluid_out(k_6_34), .air_in(c_7_0));
valve v_7_69 (.fluid_in(k_7_69), .fluid_out(k_6_34), .air_in(c_7_1));
valve v_7_70 (.fluid_in(k_7_70), .fluid_out(k_6_35), .air_in(c_7_0));
valve v_7_71 (.fluid_in(k_7_71), .fluid_out(k_6_35), .air_in(c_7_1));
valve v_7_72 (.fluid_in(k_7_72), .fluid_out(k_6_36), .air_in(c_7_0));
valve v_7_73 (.fluid_in(k_7_73), .fluid_out(k_6_36), .air_in(c_7_1));
valve v_7_74 (.fluid_in(k_7_74), .fluid_out(k_6_37), .air_in(c_7_0));
valve v_7_75 (.fluid_in(k_7_75), .fluid_out(k_6_37), .air_in(c_7_1));
valve v_7_76 (.fluid_in(k_7_76), .fluid_out(k_6_38), .air_in(c_7_0));
valve v_7_77 (.fluid_in(k_7_77), .fluid_out(k_6_38), .air_in(c_7_1));
valve v_7_78 (.fluid_in(k_7_78), .fluid_out(k_6_39), .air_in(c_7_0));
valve v_7_79 (.fluid_in(k_7_79), .fluid_out(k_6_39), .air_in(c_7_1));
valve v_7_80 (.fluid_in(k_7_80), .fluid_out(k_6_40), .air_in(c_7_0));
valve v_7_81 (.fluid_in(k_7_81), .fluid_out(k_6_40), .air_in(c_7_1));
valve v_7_82 (.fluid_in(k_7_82), .fluid_out(k_6_41), .air_in(c_7_0));
valve v_7_83 (.fluid_in(k_7_83), .fluid_out(k_6_41), .air_in(c_7_1));
valve v_7_84 (.fluid_in(k_7_84), .fluid_out(k_6_42), .air_in(c_7_0));
valve v_7_85 (.fluid_in(k_7_85), .fluid_out(k_6_42), .air_in(c_7_1));
valve v_7_86 (.fluid_in(k_7_86), .fluid_out(k_6_43), .air_in(c_7_0));
valve v_7_87 (.fluid_in(k_7_87), .fluid_out(k_6_43), .air_in(c_7_1));
valve v_7_88 (.fluid_in(k_7_88), .fluid_out(k_6_44), .air_in(c_7_0));
valve v_7_89 (.fluid_in(k_7_89), .fluid_out(k_6_44), .air_in(c_7_1));
valve v_7_90 (.fluid_in(k_7_90), .fluid_out(k_6_45), .air_in(c_7_0));
valve v_7_91 (.fluid_in(k_7_91), .fluid_out(k_6_45), .air_in(c_7_1));
valve v_7_92 (.fluid_in(k_7_92), .fluid_out(k_6_46), .air_in(c_7_0));
valve v_7_93 (.fluid_in(k_7_93), .fluid_out(k_6_46), .air_in(c_7_1));
valve v_7_94 (.fluid_in(k_7_94), .fluid_out(k_6_47), .air_in(c_7_0));
valve v_7_95 (.fluid_in(k_7_95), .fluid_out(k_6_47), .air_in(c_7_1));
valve v_7_96 (.fluid_in(k_7_96), .fluid_out(k_6_48), .air_in(c_7_0));
valve v_7_97 (.fluid_in(k_7_97), .fluid_out(k_6_48), .air_in(c_7_1));
valve v_7_98 (.fluid_in(k_7_98), .fluid_out(k_6_49), .air_in(c_7_0));
valve v_7_99 (.fluid_in(k_7_99), .fluid_out(k_6_49), .air_in(c_7_1));
valve v_7_100 (.fluid_in(k_7_100), .fluid_out(k_6_50), .air_in(c_7_0));
valve v_7_101 (.fluid_in(k_7_101), .fluid_out(k_6_50), .air_in(c_7_1));
valve v_7_102 (.fluid_in(k_7_102), .fluid_out(k_6_51), .air_in(c_7_0));
valve v_7_103 (.fluid_in(k_7_103), .fluid_out(k_6_51), .air_in(c_7_1));
valve v_7_104 (.fluid_in(k_7_104), .fluid_out(k_6_52), .air_in(c_7_0));
valve v_7_105 (.fluid_in(k_7_105), .fluid_out(k_6_52), .air_in(c_7_1));
valve v_7_106 (.fluid_in(k_7_106), .fluid_out(k_6_53), .air_in(c_7_0));
valve v_7_107 (.fluid_in(k_7_107), .fluid_out(k_6_53), .air_in(c_7_1));
valve v_7_108 (.fluid_in(k_7_108), .fluid_out(k_6_54), .air_in(c_7_0));
valve v_7_109 (.fluid_in(k_7_109), .fluid_out(k_6_54), .air_in(c_7_1));
valve v_7_110 (.fluid_in(k_7_110), .fluid_out(k_6_55), .air_in(c_7_0));
valve v_7_111 (.fluid_in(k_7_111), .fluid_out(k_6_55), .air_in(c_7_1));
valve v_7_112 (.fluid_in(k_7_112), .fluid_out(k_6_56), .air_in(c_7_0));
valve v_7_113 (.fluid_in(k_7_113), .fluid_out(k_6_56), .air_in(c_7_1));
valve v_7_114 (.fluid_in(k_7_114), .fluid_out(k_6_57), .air_in(c_7_0));
valve v_7_115 (.fluid_in(k_7_115), .fluid_out(k_6_57), .air_in(c_7_1));
valve v_7_116 (.fluid_in(k_7_116), .fluid_out(k_6_58), .air_in(c_7_0));
valve v_7_117 (.fluid_in(k_7_117), .fluid_out(k_6_58), .air_in(c_7_1));
valve v_7_118 (.fluid_in(k_7_118), .fluid_out(k_6_59), .air_in(c_7_0));
valve v_7_119 (.fluid_in(k_7_119), .fluid_out(k_6_59), .air_in(c_7_1));
valve v_7_120 (.fluid_in(k_7_120), .fluid_out(k_6_60), .air_in(c_7_0));
valve v_7_121 (.fluid_in(k_7_121), .fluid_out(k_6_60), .air_in(c_7_1));
valve v_7_122 (.fluid_in(k_7_122), .fluid_out(k_6_61), .air_in(c_7_0));
valve v_7_123 (.fluid_in(k_7_123), .fluid_out(k_6_61), .air_in(c_7_1));
valve v_7_124 (.fluid_in(k_7_124), .fluid_out(k_6_62), .air_in(c_7_0));
valve v_7_125 (.fluid_in(k_7_125), .fluid_out(k_6_62), .air_in(c_7_1));
valve v_7_126 (.fluid_in(k_7_126), .fluid_out(k_6_63), .air_in(c_7_0));
valve v_7_127 (.fluid_in(k_7_127), .fluid_out(k_6_63), .air_in(c_7_1));
valve v_8_0 (.fluid_in(k_8_0), .fluid_out(k_7_0), .air_in(c_8_0));
valve v_8_1 (.fluid_in(k_8_1), .fluid_out(k_7_0), .air_in(c_8_1));
valve v_8_2 (.fluid_in(k_8_2), .fluid_out(k_7_1), .air_in(c_8_0));
valve v_8_3 (.fluid_in(k_8_3), .fluid_out(k_7_1), .air_in(c_8_1));
valve v_8_4 (.fluid_in(k_8_4), .fluid_out(k_7_2), .air_in(c_8_0));
valve v_8_5 (.fluid_in(k_8_5), .fluid_out(k_7_2), .air_in(c_8_1));
valve v_8_6 (.fluid_in(k_8_6), .fluid_out(k_7_3), .air_in(c_8_0));
valve v_8_7 (.fluid_in(k_8_7), .fluid_out(k_7_3), .air_in(c_8_1));
valve v_8_8 (.fluid_in(k_8_8), .fluid_out(k_7_4), .air_in(c_8_0));
valve v_8_9 (.fluid_in(k_8_9), .fluid_out(k_7_4), .air_in(c_8_1));
valve v_8_10 (.fluid_in(k_8_10), .fluid_out(k_7_5), .air_in(c_8_0));
valve v_8_11 (.fluid_in(k_8_11), .fluid_out(k_7_5), .air_in(c_8_1));
valve v_8_12 (.fluid_in(k_8_12), .fluid_out(k_7_6), .air_in(c_8_0));
valve v_8_13 (.fluid_in(k_8_13), .fluid_out(k_7_6), .air_in(c_8_1));
valve v_8_14 (.fluid_in(k_8_14), .fluid_out(k_7_7), .air_in(c_8_0));
valve v_8_15 (.fluid_in(k_8_15), .fluid_out(k_7_7), .air_in(c_8_1));
valve v_8_16 (.fluid_in(k_8_16), .fluid_out(k_7_8), .air_in(c_8_0));
valve v_8_17 (.fluid_in(k_8_17), .fluid_out(k_7_8), .air_in(c_8_1));
valve v_8_18 (.fluid_in(k_8_18), .fluid_out(k_7_9), .air_in(c_8_0));
valve v_8_19 (.fluid_in(k_8_19), .fluid_out(k_7_9), .air_in(c_8_1));
valve v_8_20 (.fluid_in(k_8_20), .fluid_out(k_7_10), .air_in(c_8_0));
valve v_8_21 (.fluid_in(k_8_21), .fluid_out(k_7_10), .air_in(c_8_1));
valve v_8_22 (.fluid_in(k_8_22), .fluid_out(k_7_11), .air_in(c_8_0));
valve v_8_23 (.fluid_in(k_8_23), .fluid_out(k_7_11), .air_in(c_8_1));
valve v_8_24 (.fluid_in(k_8_24), .fluid_out(k_7_12), .air_in(c_8_0));
valve v_8_25 (.fluid_in(k_8_25), .fluid_out(k_7_12), .air_in(c_8_1));
valve v_8_26 (.fluid_in(k_8_26), .fluid_out(k_7_13), .air_in(c_8_0));
valve v_8_27 (.fluid_in(k_8_27), .fluid_out(k_7_13), .air_in(c_8_1));
valve v_8_28 (.fluid_in(k_8_28), .fluid_out(k_7_14), .air_in(c_8_0));
valve v_8_29 (.fluid_in(k_8_29), .fluid_out(k_7_14), .air_in(c_8_1));
valve v_8_30 (.fluid_in(k_8_30), .fluid_out(k_7_15), .air_in(c_8_0));
valve v_8_31 (.fluid_in(k_8_31), .fluid_out(k_7_15), .air_in(c_8_1));
valve v_8_32 (.fluid_in(k_8_32), .fluid_out(k_7_16), .air_in(c_8_0));
valve v_8_33 (.fluid_in(k_8_33), .fluid_out(k_7_16), .air_in(c_8_1));
valve v_8_34 (.fluid_in(k_8_34), .fluid_out(k_7_17), .air_in(c_8_0));
valve v_8_35 (.fluid_in(k_8_35), .fluid_out(k_7_17), .air_in(c_8_1));
valve v_8_36 (.fluid_in(k_8_36), .fluid_out(k_7_18), .air_in(c_8_0));
valve v_8_37 (.fluid_in(k_8_37), .fluid_out(k_7_18), .air_in(c_8_1));
valve v_8_38 (.fluid_in(k_8_38), .fluid_out(k_7_19), .air_in(c_8_0));
valve v_8_39 (.fluid_in(k_8_39), .fluid_out(k_7_19), .air_in(c_8_1));
valve v_8_40 (.fluid_in(k_8_40), .fluid_out(k_7_20), .air_in(c_8_0));
valve v_8_41 (.fluid_in(k_8_41), .fluid_out(k_7_20), .air_in(c_8_1));
valve v_8_42 (.fluid_in(k_8_42), .fluid_out(k_7_21), .air_in(c_8_0));
valve v_8_43 (.fluid_in(k_8_43), .fluid_out(k_7_21), .air_in(c_8_1));
valve v_8_44 (.fluid_in(k_8_44), .fluid_out(k_7_22), .air_in(c_8_0));
valve v_8_45 (.fluid_in(k_8_45), .fluid_out(k_7_22), .air_in(c_8_1));
valve v_8_46 (.fluid_in(k_8_46), .fluid_out(k_7_23), .air_in(c_8_0));
valve v_8_47 (.fluid_in(k_8_47), .fluid_out(k_7_23), .air_in(c_8_1));
valve v_8_48 (.fluid_in(k_8_48), .fluid_out(k_7_24), .air_in(c_8_0));
valve v_8_49 (.fluid_in(k_8_49), .fluid_out(k_7_24), .air_in(c_8_1));
valve v_8_50 (.fluid_in(k_8_50), .fluid_out(k_7_25), .air_in(c_8_0));
valve v_8_51 (.fluid_in(k_8_51), .fluid_out(k_7_25), .air_in(c_8_1));
valve v_8_52 (.fluid_in(k_8_52), .fluid_out(k_7_26), .air_in(c_8_0));
valve v_8_53 (.fluid_in(k_8_53), .fluid_out(k_7_26), .air_in(c_8_1));
valve v_8_54 (.fluid_in(k_8_54), .fluid_out(k_7_27), .air_in(c_8_0));
valve v_8_55 (.fluid_in(k_8_55), .fluid_out(k_7_27), .air_in(c_8_1));
valve v_8_56 (.fluid_in(k_8_56), .fluid_out(k_7_28), .air_in(c_8_0));
valve v_8_57 (.fluid_in(k_8_57), .fluid_out(k_7_28), .air_in(c_8_1));
valve v_8_58 (.fluid_in(k_8_58), .fluid_out(k_7_29), .air_in(c_8_0));
valve v_8_59 (.fluid_in(k_8_59), .fluid_out(k_7_29), .air_in(c_8_1));
valve v_8_60 (.fluid_in(k_8_60), .fluid_out(k_7_30), .air_in(c_8_0));
valve v_8_61 (.fluid_in(k_8_61), .fluid_out(k_7_30), .air_in(c_8_1));
valve v_8_62 (.fluid_in(k_8_62), .fluid_out(k_7_31), .air_in(c_8_0));
valve v_8_63 (.fluid_in(k_8_63), .fluid_out(k_7_31), .air_in(c_8_1));
valve v_8_64 (.fluid_in(k_8_64), .fluid_out(k_7_32), .air_in(c_8_0));
valve v_8_65 (.fluid_in(k_8_65), .fluid_out(k_7_32), .air_in(c_8_1));
valve v_8_66 (.fluid_in(k_8_66), .fluid_out(k_7_33), .air_in(c_8_0));
valve v_8_67 (.fluid_in(k_8_67), .fluid_out(k_7_33), .air_in(c_8_1));
valve v_8_68 (.fluid_in(k_8_68), .fluid_out(k_7_34), .air_in(c_8_0));
valve v_8_69 (.fluid_in(k_8_69), .fluid_out(k_7_34), .air_in(c_8_1));
valve v_8_70 (.fluid_in(k_8_70), .fluid_out(k_7_35), .air_in(c_8_0));
valve v_8_71 (.fluid_in(k_8_71), .fluid_out(k_7_35), .air_in(c_8_1));
valve v_8_72 (.fluid_in(k_8_72), .fluid_out(k_7_36), .air_in(c_8_0));
valve v_8_73 (.fluid_in(k_8_73), .fluid_out(k_7_36), .air_in(c_8_1));
valve v_8_74 (.fluid_in(k_8_74), .fluid_out(k_7_37), .air_in(c_8_0));
valve v_8_75 (.fluid_in(k_8_75), .fluid_out(k_7_37), .air_in(c_8_1));
valve v_8_76 (.fluid_in(k_8_76), .fluid_out(k_7_38), .air_in(c_8_0));
valve v_8_77 (.fluid_in(k_8_77), .fluid_out(k_7_38), .air_in(c_8_1));
valve v_8_78 (.fluid_in(k_8_78), .fluid_out(k_7_39), .air_in(c_8_0));
valve v_8_79 (.fluid_in(k_8_79), .fluid_out(k_7_39), .air_in(c_8_1));
valve v_8_80 (.fluid_in(k_8_80), .fluid_out(k_7_40), .air_in(c_8_0));
valve v_8_81 (.fluid_in(k_8_81), .fluid_out(k_7_40), .air_in(c_8_1));
valve v_8_82 (.fluid_in(k_8_82), .fluid_out(k_7_41), .air_in(c_8_0));
valve v_8_83 (.fluid_in(k_8_83), .fluid_out(k_7_41), .air_in(c_8_1));
valve v_8_84 (.fluid_in(k_8_84), .fluid_out(k_7_42), .air_in(c_8_0));
valve v_8_85 (.fluid_in(k_8_85), .fluid_out(k_7_42), .air_in(c_8_1));
valve v_8_86 (.fluid_in(k_8_86), .fluid_out(k_7_43), .air_in(c_8_0));
valve v_8_87 (.fluid_in(k_8_87), .fluid_out(k_7_43), .air_in(c_8_1));
valve v_8_88 (.fluid_in(k_8_88), .fluid_out(k_7_44), .air_in(c_8_0));
valve v_8_89 (.fluid_in(k_8_89), .fluid_out(k_7_44), .air_in(c_8_1));
valve v_8_90 (.fluid_in(k_8_90), .fluid_out(k_7_45), .air_in(c_8_0));
valve v_8_91 (.fluid_in(k_8_91), .fluid_out(k_7_45), .air_in(c_8_1));
valve v_8_92 (.fluid_in(k_8_92), .fluid_out(k_7_46), .air_in(c_8_0));
valve v_8_93 (.fluid_in(k_8_93), .fluid_out(k_7_46), .air_in(c_8_1));
valve v_8_94 (.fluid_in(k_8_94), .fluid_out(k_7_47), .air_in(c_8_0));
valve v_8_95 (.fluid_in(k_8_95), .fluid_out(k_7_47), .air_in(c_8_1));
valve v_8_96 (.fluid_in(k_8_96), .fluid_out(k_7_48), .air_in(c_8_0));
valve v_8_97 (.fluid_in(k_8_97), .fluid_out(k_7_48), .air_in(c_8_1));
valve v_8_98 (.fluid_in(k_8_98), .fluid_out(k_7_49), .air_in(c_8_0));
valve v_8_99 (.fluid_in(k_8_99), .fluid_out(k_7_49), .air_in(c_8_1));
valve v_8_100 (.fluid_in(k_8_100), .fluid_out(k_7_50), .air_in(c_8_0));
valve v_8_101 (.fluid_in(k_8_101), .fluid_out(k_7_50), .air_in(c_8_1));
valve v_8_102 (.fluid_in(k_8_102), .fluid_out(k_7_51), .air_in(c_8_0));
valve v_8_103 (.fluid_in(k_8_103), .fluid_out(k_7_51), .air_in(c_8_1));
valve v_8_104 (.fluid_in(k_8_104), .fluid_out(k_7_52), .air_in(c_8_0));
valve v_8_105 (.fluid_in(k_8_105), .fluid_out(k_7_52), .air_in(c_8_1));
valve v_8_106 (.fluid_in(k_8_106), .fluid_out(k_7_53), .air_in(c_8_0));
valve v_8_107 (.fluid_in(k_8_107), .fluid_out(k_7_53), .air_in(c_8_1));
valve v_8_108 (.fluid_in(k_8_108), .fluid_out(k_7_54), .air_in(c_8_0));
valve v_8_109 (.fluid_in(k_8_109), .fluid_out(k_7_54), .air_in(c_8_1));
valve v_8_110 (.fluid_in(k_8_110), .fluid_out(k_7_55), .air_in(c_8_0));
valve v_8_111 (.fluid_in(k_8_111), .fluid_out(k_7_55), .air_in(c_8_1));
valve v_8_112 (.fluid_in(k_8_112), .fluid_out(k_7_56), .air_in(c_8_0));
valve v_8_113 (.fluid_in(k_8_113), .fluid_out(k_7_56), .air_in(c_8_1));
valve v_8_114 (.fluid_in(k_8_114), .fluid_out(k_7_57), .air_in(c_8_0));
valve v_8_115 (.fluid_in(k_8_115), .fluid_out(k_7_57), .air_in(c_8_1));
valve v_8_116 (.fluid_in(k_8_116), .fluid_out(k_7_58), .air_in(c_8_0));
valve v_8_117 (.fluid_in(k_8_117), .fluid_out(k_7_58), .air_in(c_8_1));
valve v_8_118 (.fluid_in(k_8_118), .fluid_out(k_7_59), .air_in(c_8_0));
valve v_8_119 (.fluid_in(k_8_119), .fluid_out(k_7_59), .air_in(c_8_1));
valve v_8_120 (.fluid_in(k_8_120), .fluid_out(k_7_60), .air_in(c_8_0));
valve v_8_121 (.fluid_in(k_8_121), .fluid_out(k_7_60), .air_in(c_8_1));
valve v_8_122 (.fluid_in(k_8_122), .fluid_out(k_7_61), .air_in(c_8_0));
valve v_8_123 (.fluid_in(k_8_123), .fluid_out(k_7_61), .air_in(c_8_1));
valve v_8_124 (.fluid_in(k_8_124), .fluid_out(k_7_62), .air_in(c_8_0));
valve v_8_125 (.fluid_in(k_8_125), .fluid_out(k_7_62), .air_in(c_8_1));
valve v_8_126 (.fluid_in(k_8_126), .fluid_out(k_7_63), .air_in(c_8_0));
valve v_8_127 (.fluid_in(k_8_127), .fluid_out(k_7_63), .air_in(c_8_1));
valve v_8_128 (.fluid_in(k_8_128), .fluid_out(k_7_64), .air_in(c_8_0));
valve v_8_129 (.fluid_in(k_8_129), .fluid_out(k_7_64), .air_in(c_8_1));
valve v_8_130 (.fluid_in(k_8_130), .fluid_out(k_7_65), .air_in(c_8_0));
valve v_8_131 (.fluid_in(k_8_131), .fluid_out(k_7_65), .air_in(c_8_1));
valve v_8_132 (.fluid_in(k_8_132), .fluid_out(k_7_66), .air_in(c_8_0));
valve v_8_133 (.fluid_in(k_8_133), .fluid_out(k_7_66), .air_in(c_8_1));
valve v_8_134 (.fluid_in(k_8_134), .fluid_out(k_7_67), .air_in(c_8_0));
valve v_8_135 (.fluid_in(k_8_135), .fluid_out(k_7_67), .air_in(c_8_1));
valve v_8_136 (.fluid_in(k_8_136), .fluid_out(k_7_68), .air_in(c_8_0));
valve v_8_137 (.fluid_in(k_8_137), .fluid_out(k_7_68), .air_in(c_8_1));
valve v_8_138 (.fluid_in(k_8_138), .fluid_out(k_7_69), .air_in(c_8_0));
valve v_8_139 (.fluid_in(k_8_139), .fluid_out(k_7_69), .air_in(c_8_1));
valve v_8_140 (.fluid_in(k_8_140), .fluid_out(k_7_70), .air_in(c_8_0));
valve v_8_141 (.fluid_in(k_8_141), .fluid_out(k_7_70), .air_in(c_8_1));
valve v_8_142 (.fluid_in(k_8_142), .fluid_out(k_7_71), .air_in(c_8_0));
valve v_8_143 (.fluid_in(k_8_143), .fluid_out(k_7_71), .air_in(c_8_1));
valve v_8_144 (.fluid_in(k_8_144), .fluid_out(k_7_72), .air_in(c_8_0));
valve v_8_145 (.fluid_in(k_8_145), .fluid_out(k_7_72), .air_in(c_8_1));
valve v_8_146 (.fluid_in(k_8_146), .fluid_out(k_7_73), .air_in(c_8_0));
valve v_8_147 (.fluid_in(k_8_147), .fluid_out(k_7_73), .air_in(c_8_1));
valve v_8_148 (.fluid_in(k_8_148), .fluid_out(k_7_74), .air_in(c_8_0));
valve v_8_149 (.fluid_in(k_8_149), .fluid_out(k_7_74), .air_in(c_8_1));
valve v_8_150 (.fluid_in(k_8_150), .fluid_out(k_7_75), .air_in(c_8_0));
valve v_8_151 (.fluid_in(k_8_151), .fluid_out(k_7_75), .air_in(c_8_1));
valve v_8_152 (.fluid_in(k_8_152), .fluid_out(k_7_76), .air_in(c_8_0));
valve v_8_153 (.fluid_in(k_8_153), .fluid_out(k_7_76), .air_in(c_8_1));
valve v_8_154 (.fluid_in(k_8_154), .fluid_out(k_7_77), .air_in(c_8_0));
valve v_8_155 (.fluid_in(k_8_155), .fluid_out(k_7_77), .air_in(c_8_1));
valve v_8_156 (.fluid_in(k_8_156), .fluid_out(k_7_78), .air_in(c_8_0));
valve v_8_157 (.fluid_in(k_8_157), .fluid_out(k_7_78), .air_in(c_8_1));
valve v_8_158 (.fluid_in(k_8_158), .fluid_out(k_7_79), .air_in(c_8_0));
valve v_8_159 (.fluid_in(k_8_159), .fluid_out(k_7_79), .air_in(c_8_1));
valve v_8_160 (.fluid_in(k_8_160), .fluid_out(k_7_80), .air_in(c_8_0));
valve v_8_161 (.fluid_in(k_8_161), .fluid_out(k_7_80), .air_in(c_8_1));
valve v_8_162 (.fluid_in(k_8_162), .fluid_out(k_7_81), .air_in(c_8_0));
valve v_8_163 (.fluid_in(k_8_163), .fluid_out(k_7_81), .air_in(c_8_1));
valve v_8_164 (.fluid_in(k_8_164), .fluid_out(k_7_82), .air_in(c_8_0));
valve v_8_165 (.fluid_in(k_8_165), .fluid_out(k_7_82), .air_in(c_8_1));
valve v_8_166 (.fluid_in(k_8_166), .fluid_out(k_7_83), .air_in(c_8_0));
valve v_8_167 (.fluid_in(k_8_167), .fluid_out(k_7_83), .air_in(c_8_1));
valve v_8_168 (.fluid_in(k_8_168), .fluid_out(k_7_84), .air_in(c_8_0));
valve v_8_169 (.fluid_in(k_8_169), .fluid_out(k_7_84), .air_in(c_8_1));
valve v_8_170 (.fluid_in(k_8_170), .fluid_out(k_7_85), .air_in(c_8_0));
valve v_8_171 (.fluid_in(k_8_171), .fluid_out(k_7_85), .air_in(c_8_1));
valve v_8_172 (.fluid_in(k_8_172), .fluid_out(k_7_86), .air_in(c_8_0));
valve v_8_173 (.fluid_in(k_8_173), .fluid_out(k_7_86), .air_in(c_8_1));
valve v_8_174 (.fluid_in(k_8_174), .fluid_out(k_7_87), .air_in(c_8_0));
valve v_8_175 (.fluid_in(k_8_175), .fluid_out(k_7_87), .air_in(c_8_1));
valve v_8_176 (.fluid_in(k_8_176), .fluid_out(k_7_88), .air_in(c_8_0));
valve v_8_177 (.fluid_in(k_8_177), .fluid_out(k_7_88), .air_in(c_8_1));
valve v_8_178 (.fluid_in(k_8_178), .fluid_out(k_7_89), .air_in(c_8_0));
valve v_8_179 (.fluid_in(k_8_179), .fluid_out(k_7_89), .air_in(c_8_1));
valve v_8_180 (.fluid_in(k_8_180), .fluid_out(k_7_90), .air_in(c_8_0));
valve v_8_181 (.fluid_in(k_8_181), .fluid_out(k_7_90), .air_in(c_8_1));
valve v_8_182 (.fluid_in(k_8_182), .fluid_out(k_7_91), .air_in(c_8_0));
valve v_8_183 (.fluid_in(k_8_183), .fluid_out(k_7_91), .air_in(c_8_1));
valve v_8_184 (.fluid_in(k_8_184), .fluid_out(k_7_92), .air_in(c_8_0));
valve v_8_185 (.fluid_in(k_8_185), .fluid_out(k_7_92), .air_in(c_8_1));
valve v_8_186 (.fluid_in(k_8_186), .fluid_out(k_7_93), .air_in(c_8_0));
valve v_8_187 (.fluid_in(k_8_187), .fluid_out(k_7_93), .air_in(c_8_1));
valve v_8_188 (.fluid_in(k_8_188), .fluid_out(k_7_94), .air_in(c_8_0));
valve v_8_189 (.fluid_in(k_8_189), .fluid_out(k_7_94), .air_in(c_8_1));
valve v_8_190 (.fluid_in(k_8_190), .fluid_out(k_7_95), .air_in(c_8_0));
valve v_8_191 (.fluid_in(k_8_191), .fluid_out(k_7_95), .air_in(c_8_1));
valve v_8_192 (.fluid_in(k_8_192), .fluid_out(k_7_96), .air_in(c_8_0));
valve v_8_193 (.fluid_in(k_8_193), .fluid_out(k_7_96), .air_in(c_8_1));
valve v_8_194 (.fluid_in(k_8_194), .fluid_out(k_7_97), .air_in(c_8_0));
valve v_8_195 (.fluid_in(k_8_195), .fluid_out(k_7_97), .air_in(c_8_1));
valve v_8_196 (.fluid_in(k_8_196), .fluid_out(k_7_98), .air_in(c_8_0));
valve v_8_197 (.fluid_in(k_8_197), .fluid_out(k_7_98), .air_in(c_8_1));
valve v_8_198 (.fluid_in(k_8_198), .fluid_out(k_7_99), .air_in(c_8_0));
valve v_8_199 (.fluid_in(k_8_199), .fluid_out(k_7_99), .air_in(c_8_1));
valve v_8_200 (.fluid_in(k_8_200), .fluid_out(k_7_100), .air_in(c_8_0));
valve v_8_201 (.fluid_in(k_8_201), .fluid_out(k_7_100), .air_in(c_8_1));
valve v_8_202 (.fluid_in(k_8_202), .fluid_out(k_7_101), .air_in(c_8_0));
valve v_8_203 (.fluid_in(k_8_203), .fluid_out(k_7_101), .air_in(c_8_1));
valve v_8_204 (.fluid_in(k_8_204), .fluid_out(k_7_102), .air_in(c_8_0));
valve v_8_205 (.fluid_in(k_8_205), .fluid_out(k_7_102), .air_in(c_8_1));
valve v_8_206 (.fluid_in(k_8_206), .fluid_out(k_7_103), .air_in(c_8_0));
valve v_8_207 (.fluid_in(k_8_207), .fluid_out(k_7_103), .air_in(c_8_1));
valve v_8_208 (.fluid_in(k_8_208), .fluid_out(k_7_104), .air_in(c_8_0));
valve v_8_209 (.fluid_in(k_8_209), .fluid_out(k_7_104), .air_in(c_8_1));
valve v_8_210 (.fluid_in(k_8_210), .fluid_out(k_7_105), .air_in(c_8_0));
valve v_8_211 (.fluid_in(k_8_211), .fluid_out(k_7_105), .air_in(c_8_1));
valve v_8_212 (.fluid_in(k_8_212), .fluid_out(k_7_106), .air_in(c_8_0));
valve v_8_213 (.fluid_in(k_8_213), .fluid_out(k_7_106), .air_in(c_8_1));
valve v_8_214 (.fluid_in(k_8_214), .fluid_out(k_7_107), .air_in(c_8_0));
valve v_8_215 (.fluid_in(k_8_215), .fluid_out(k_7_107), .air_in(c_8_1));
valve v_8_216 (.fluid_in(k_8_216), .fluid_out(k_7_108), .air_in(c_8_0));
valve v_8_217 (.fluid_in(k_8_217), .fluid_out(k_7_108), .air_in(c_8_1));
valve v_8_218 (.fluid_in(k_8_218), .fluid_out(k_7_109), .air_in(c_8_0));
valve v_8_219 (.fluid_in(k_8_219), .fluid_out(k_7_109), .air_in(c_8_1));
valve v_8_220 (.fluid_in(k_8_220), .fluid_out(k_7_110), .air_in(c_8_0));
valve v_8_221 (.fluid_in(k_8_221), .fluid_out(k_7_110), .air_in(c_8_1));
valve v_8_222 (.fluid_in(k_8_222), .fluid_out(k_7_111), .air_in(c_8_0));
valve v_8_223 (.fluid_in(k_8_223), .fluid_out(k_7_111), .air_in(c_8_1));
valve v_8_224 (.fluid_in(k_8_224), .fluid_out(k_7_112), .air_in(c_8_0));
valve v_8_225 (.fluid_in(k_8_225), .fluid_out(k_7_112), .air_in(c_8_1));
valve v_8_226 (.fluid_in(k_8_226), .fluid_out(k_7_113), .air_in(c_8_0));
valve v_8_227 (.fluid_in(k_8_227), .fluid_out(k_7_113), .air_in(c_8_1));
valve v_8_228 (.fluid_in(k_8_228), .fluid_out(k_7_114), .air_in(c_8_0));
valve v_8_229 (.fluid_in(k_8_229), .fluid_out(k_7_114), .air_in(c_8_1));
valve v_8_230 (.fluid_in(k_8_230), .fluid_out(k_7_115), .air_in(c_8_0));
valve v_8_231 (.fluid_in(k_8_231), .fluid_out(k_7_115), .air_in(c_8_1));
valve v_8_232 (.fluid_in(k_8_232), .fluid_out(k_7_116), .air_in(c_8_0));
valve v_8_233 (.fluid_in(k_8_233), .fluid_out(k_7_116), .air_in(c_8_1));
valve v_8_234 (.fluid_in(k_8_234), .fluid_out(k_7_117), .air_in(c_8_0));
valve v_8_235 (.fluid_in(k_8_235), .fluid_out(k_7_117), .air_in(c_8_1));
valve v_8_236 (.fluid_in(k_8_236), .fluid_out(k_7_118), .air_in(c_8_0));
valve v_8_237 (.fluid_in(k_8_237), .fluid_out(k_7_118), .air_in(c_8_1));
valve v_8_238 (.fluid_in(k_8_238), .fluid_out(k_7_119), .air_in(c_8_0));
valve v_8_239 (.fluid_in(k_8_239), .fluid_out(k_7_119), .air_in(c_8_1));
valve v_8_240 (.fluid_in(k_8_240), .fluid_out(k_7_120), .air_in(c_8_0));
valve v_8_241 (.fluid_in(k_8_241), .fluid_out(k_7_120), .air_in(c_8_1));
valve v_8_242 (.fluid_in(k_8_242), .fluid_out(k_7_121), .air_in(c_8_0));
valve v_8_243 (.fluid_in(k_8_243), .fluid_out(k_7_121), .air_in(c_8_1));
valve v_8_244 (.fluid_in(k_8_244), .fluid_out(k_7_122), .air_in(c_8_0));
valve v_8_245 (.fluid_in(k_8_245), .fluid_out(k_7_122), .air_in(c_8_1));
valve v_8_246 (.fluid_in(k_8_246), .fluid_out(k_7_123), .air_in(c_8_0));
valve v_8_247 (.fluid_in(k_8_247), .fluid_out(k_7_123), .air_in(c_8_1));
valve v_8_248 (.fluid_in(k_8_248), .fluid_out(k_7_124), .air_in(c_8_0));
valve v_8_249 (.fluid_in(k_8_249), .fluid_out(k_7_124), .air_in(c_8_1));
valve v_8_250 (.fluid_in(k_8_250), .fluid_out(k_7_125), .air_in(c_8_0));
valve v_8_251 (.fluid_in(k_8_251), .fluid_out(k_7_125), .air_in(c_8_1));
valve v_8_252 (.fluid_in(k_8_252), .fluid_out(k_7_126), .air_in(c_8_0));
valve v_8_253 (.fluid_in(k_8_253), .fluid_out(k_7_126), .air_in(c_8_1));
valve v_8_254 (.fluid_in(k_8_254), .fluid_out(k_7_127), .air_in(c_8_0));
valve v_8_255 (.fluid_in(k_8_255), .fluid_out(k_7_127), .air_in(c_8_1));
valve v_9_0 (.fluid_in(k_9_0), .fluid_out(k_8_0), .air_in(c_9_0));
valve v_9_1 (.fluid_in(k_9_1), .fluid_out(k_8_0), .air_in(c_9_1));
valve v_9_2 (.fluid_in(k_9_2), .fluid_out(k_8_1), .air_in(c_9_0));
valve v_9_3 (.fluid_in(k_9_3), .fluid_out(k_8_1), .air_in(c_9_1));
valve v_9_4 (.fluid_in(k_9_4), .fluid_out(k_8_2), .air_in(c_9_0));
valve v_9_5 (.fluid_in(k_9_5), .fluid_out(k_8_2), .air_in(c_9_1));
valve v_9_6 (.fluid_in(k_9_6), .fluid_out(k_8_3), .air_in(c_9_0));
valve v_9_7 (.fluid_in(k_9_7), .fluid_out(k_8_3), .air_in(c_9_1));
valve v_9_8 (.fluid_in(k_9_8), .fluid_out(k_8_4), .air_in(c_9_0));
valve v_9_9 (.fluid_in(k_9_9), .fluid_out(k_8_4), .air_in(c_9_1));
valve v_9_10 (.fluid_in(k_9_10), .fluid_out(k_8_5), .air_in(c_9_0));
valve v_9_11 (.fluid_in(k_9_11), .fluid_out(k_8_5), .air_in(c_9_1));
valve v_9_12 (.fluid_in(k_9_12), .fluid_out(k_8_6), .air_in(c_9_0));
valve v_9_13 (.fluid_in(k_9_13), .fluid_out(k_8_6), .air_in(c_9_1));
valve v_9_14 (.fluid_in(k_9_14), .fluid_out(k_8_7), .air_in(c_9_0));
valve v_9_15 (.fluid_in(k_9_15), .fluid_out(k_8_7), .air_in(c_9_1));
valve v_9_16 (.fluid_in(k_9_16), .fluid_out(k_8_8), .air_in(c_9_0));
valve v_9_17 (.fluid_in(k_9_17), .fluid_out(k_8_8), .air_in(c_9_1));
valve v_9_18 (.fluid_in(k_9_18), .fluid_out(k_8_9), .air_in(c_9_0));
valve v_9_19 (.fluid_in(k_9_19), .fluid_out(k_8_9), .air_in(c_9_1));
valve v_9_20 (.fluid_in(k_9_20), .fluid_out(k_8_10), .air_in(c_9_0));
valve v_9_21 (.fluid_in(k_9_21), .fluid_out(k_8_10), .air_in(c_9_1));
valve v_9_22 (.fluid_in(k_9_22), .fluid_out(k_8_11), .air_in(c_9_0));
valve v_9_23 (.fluid_in(k_9_23), .fluid_out(k_8_11), .air_in(c_9_1));
valve v_9_24 (.fluid_in(k_9_24), .fluid_out(k_8_12), .air_in(c_9_0));
valve v_9_25 (.fluid_in(k_9_25), .fluid_out(k_8_12), .air_in(c_9_1));
valve v_9_26 (.fluid_in(k_9_26), .fluid_out(k_8_13), .air_in(c_9_0));
valve v_9_27 (.fluid_in(k_9_27), .fluid_out(k_8_13), .air_in(c_9_1));
valve v_9_28 (.fluid_in(k_9_28), .fluid_out(k_8_14), .air_in(c_9_0));
valve v_9_29 (.fluid_in(k_9_29), .fluid_out(k_8_14), .air_in(c_9_1));
valve v_9_30 (.fluid_in(k_9_30), .fluid_out(k_8_15), .air_in(c_9_0));
valve v_9_31 (.fluid_in(k_9_31), .fluid_out(k_8_15), .air_in(c_9_1));
valve v_9_32 (.fluid_in(k_9_32), .fluid_out(k_8_16), .air_in(c_9_0));
valve v_9_33 (.fluid_in(k_9_33), .fluid_out(k_8_16), .air_in(c_9_1));
valve v_9_34 (.fluid_in(k_9_34), .fluid_out(k_8_17), .air_in(c_9_0));
valve v_9_35 (.fluid_in(k_9_35), .fluid_out(k_8_17), .air_in(c_9_1));
valve v_9_36 (.fluid_in(k_9_36), .fluid_out(k_8_18), .air_in(c_9_0));
valve v_9_37 (.fluid_in(k_9_37), .fluid_out(k_8_18), .air_in(c_9_1));
valve v_9_38 (.fluid_in(k_9_38), .fluid_out(k_8_19), .air_in(c_9_0));
valve v_9_39 (.fluid_in(k_9_39), .fluid_out(k_8_19), .air_in(c_9_1));
valve v_9_40 (.fluid_in(k_9_40), .fluid_out(k_8_20), .air_in(c_9_0));
valve v_9_41 (.fluid_in(k_9_41), .fluid_out(k_8_20), .air_in(c_9_1));
valve v_9_42 (.fluid_in(k_9_42), .fluid_out(k_8_21), .air_in(c_9_0));
valve v_9_43 (.fluid_in(k_9_43), .fluid_out(k_8_21), .air_in(c_9_1));
valve v_9_44 (.fluid_in(k_9_44), .fluid_out(k_8_22), .air_in(c_9_0));
valve v_9_45 (.fluid_in(k_9_45), .fluid_out(k_8_22), .air_in(c_9_1));
valve v_9_46 (.fluid_in(k_9_46), .fluid_out(k_8_23), .air_in(c_9_0));
valve v_9_47 (.fluid_in(k_9_47), .fluid_out(k_8_23), .air_in(c_9_1));
valve v_9_48 (.fluid_in(k_9_48), .fluid_out(k_8_24), .air_in(c_9_0));
valve v_9_49 (.fluid_in(k_9_49), .fluid_out(k_8_24), .air_in(c_9_1));
valve v_9_50 (.fluid_in(k_9_50), .fluid_out(k_8_25), .air_in(c_9_0));
valve v_9_51 (.fluid_in(k_9_51), .fluid_out(k_8_25), .air_in(c_9_1));
valve v_9_52 (.fluid_in(k_9_52), .fluid_out(k_8_26), .air_in(c_9_0));
valve v_9_53 (.fluid_in(k_9_53), .fluid_out(k_8_26), .air_in(c_9_1));
valve v_9_54 (.fluid_in(k_9_54), .fluid_out(k_8_27), .air_in(c_9_0));
valve v_9_55 (.fluid_in(k_9_55), .fluid_out(k_8_27), .air_in(c_9_1));
valve v_9_56 (.fluid_in(k_9_56), .fluid_out(k_8_28), .air_in(c_9_0));
valve v_9_57 (.fluid_in(k_9_57), .fluid_out(k_8_28), .air_in(c_9_1));
valve v_9_58 (.fluid_in(k_9_58), .fluid_out(k_8_29), .air_in(c_9_0));
valve v_9_59 (.fluid_in(k_9_59), .fluid_out(k_8_29), .air_in(c_9_1));
valve v_9_60 (.fluid_in(k_9_60), .fluid_out(k_8_30), .air_in(c_9_0));
valve v_9_61 (.fluid_in(k_9_61), .fluid_out(k_8_30), .air_in(c_9_1));
valve v_9_62 (.fluid_in(k_9_62), .fluid_out(k_8_31), .air_in(c_9_0));
valve v_9_63 (.fluid_in(k_9_63), .fluid_out(k_8_31), .air_in(c_9_1));
valve v_9_64 (.fluid_in(k_9_64), .fluid_out(k_8_32), .air_in(c_9_0));
valve v_9_65 (.fluid_in(k_9_65), .fluid_out(k_8_32), .air_in(c_9_1));
valve v_9_66 (.fluid_in(k_9_66), .fluid_out(k_8_33), .air_in(c_9_0));
valve v_9_67 (.fluid_in(k_9_67), .fluid_out(k_8_33), .air_in(c_9_1));
valve v_9_68 (.fluid_in(k_9_68), .fluid_out(k_8_34), .air_in(c_9_0));
valve v_9_69 (.fluid_in(k_9_69), .fluid_out(k_8_34), .air_in(c_9_1));
valve v_9_70 (.fluid_in(k_9_70), .fluid_out(k_8_35), .air_in(c_9_0));
valve v_9_71 (.fluid_in(k_9_71), .fluid_out(k_8_35), .air_in(c_9_1));
valve v_9_72 (.fluid_in(k_9_72), .fluid_out(k_8_36), .air_in(c_9_0));
valve v_9_73 (.fluid_in(k_9_73), .fluid_out(k_8_36), .air_in(c_9_1));
valve v_9_74 (.fluid_in(k_9_74), .fluid_out(k_8_37), .air_in(c_9_0));
valve v_9_75 (.fluid_in(k_9_75), .fluid_out(k_8_37), .air_in(c_9_1));
valve v_9_76 (.fluid_in(k_9_76), .fluid_out(k_8_38), .air_in(c_9_0));
valve v_9_77 (.fluid_in(k_9_77), .fluid_out(k_8_38), .air_in(c_9_1));
valve v_9_78 (.fluid_in(k_9_78), .fluid_out(k_8_39), .air_in(c_9_0));
valve v_9_79 (.fluid_in(k_9_79), .fluid_out(k_8_39), .air_in(c_9_1));
valve v_9_80 (.fluid_in(k_9_80), .fluid_out(k_8_40), .air_in(c_9_0));
valve v_9_81 (.fluid_in(k_9_81), .fluid_out(k_8_40), .air_in(c_9_1));
valve v_9_82 (.fluid_in(k_9_82), .fluid_out(k_8_41), .air_in(c_9_0));
valve v_9_83 (.fluid_in(k_9_83), .fluid_out(k_8_41), .air_in(c_9_1));
valve v_9_84 (.fluid_in(k_9_84), .fluid_out(k_8_42), .air_in(c_9_0));
valve v_9_85 (.fluid_in(k_9_85), .fluid_out(k_8_42), .air_in(c_9_1));
valve v_9_86 (.fluid_in(k_9_86), .fluid_out(k_8_43), .air_in(c_9_0));
valve v_9_87 (.fluid_in(k_9_87), .fluid_out(k_8_43), .air_in(c_9_1));
valve v_9_88 (.fluid_in(k_9_88), .fluid_out(k_8_44), .air_in(c_9_0));
valve v_9_89 (.fluid_in(k_9_89), .fluid_out(k_8_44), .air_in(c_9_1));
valve v_9_90 (.fluid_in(k_9_90), .fluid_out(k_8_45), .air_in(c_9_0));
valve v_9_91 (.fluid_in(k_9_91), .fluid_out(k_8_45), .air_in(c_9_1));
valve v_9_92 (.fluid_in(k_9_92), .fluid_out(k_8_46), .air_in(c_9_0));
valve v_9_93 (.fluid_in(k_9_93), .fluid_out(k_8_46), .air_in(c_9_1));
valve v_9_94 (.fluid_in(k_9_94), .fluid_out(k_8_47), .air_in(c_9_0));
valve v_9_95 (.fluid_in(k_9_95), .fluid_out(k_8_47), .air_in(c_9_1));
valve v_9_96 (.fluid_in(k_9_96), .fluid_out(k_8_48), .air_in(c_9_0));
valve v_9_97 (.fluid_in(k_9_97), .fluid_out(k_8_48), .air_in(c_9_1));
valve v_9_98 (.fluid_in(k_9_98), .fluid_out(k_8_49), .air_in(c_9_0));
valve v_9_99 (.fluid_in(k_9_99), .fluid_out(k_8_49), .air_in(c_9_1));
valve v_9_100 (.fluid_in(k_9_100), .fluid_out(k_8_50), .air_in(c_9_0));
valve v_9_101 (.fluid_in(k_9_101), .fluid_out(k_8_50), .air_in(c_9_1));
valve v_9_102 (.fluid_in(k_9_102), .fluid_out(k_8_51), .air_in(c_9_0));
valve v_9_103 (.fluid_in(k_9_103), .fluid_out(k_8_51), .air_in(c_9_1));
valve v_9_104 (.fluid_in(k_9_104), .fluid_out(k_8_52), .air_in(c_9_0));
valve v_9_105 (.fluid_in(k_9_105), .fluid_out(k_8_52), .air_in(c_9_1));
valve v_9_106 (.fluid_in(k_9_106), .fluid_out(k_8_53), .air_in(c_9_0));
valve v_9_107 (.fluid_in(k_9_107), .fluid_out(k_8_53), .air_in(c_9_1));
valve v_9_108 (.fluid_in(k_9_108), .fluid_out(k_8_54), .air_in(c_9_0));
valve v_9_109 (.fluid_in(k_9_109), .fluid_out(k_8_54), .air_in(c_9_1));
valve v_9_110 (.fluid_in(k_9_110), .fluid_out(k_8_55), .air_in(c_9_0));
valve v_9_111 (.fluid_in(k_9_111), .fluid_out(k_8_55), .air_in(c_9_1));
valve v_9_112 (.fluid_in(k_9_112), .fluid_out(k_8_56), .air_in(c_9_0));
valve v_9_113 (.fluid_in(k_9_113), .fluid_out(k_8_56), .air_in(c_9_1));
valve v_9_114 (.fluid_in(k_9_114), .fluid_out(k_8_57), .air_in(c_9_0));
valve v_9_115 (.fluid_in(k_9_115), .fluid_out(k_8_57), .air_in(c_9_1));
valve v_9_116 (.fluid_in(k_9_116), .fluid_out(k_8_58), .air_in(c_9_0));
valve v_9_117 (.fluid_in(k_9_117), .fluid_out(k_8_58), .air_in(c_9_1));
valve v_9_118 (.fluid_in(k_9_118), .fluid_out(k_8_59), .air_in(c_9_0));
valve v_9_119 (.fluid_in(k_9_119), .fluid_out(k_8_59), .air_in(c_9_1));
valve v_9_120 (.fluid_in(k_9_120), .fluid_out(k_8_60), .air_in(c_9_0));
valve v_9_121 (.fluid_in(k_9_121), .fluid_out(k_8_60), .air_in(c_9_1));
valve v_9_122 (.fluid_in(k_9_122), .fluid_out(k_8_61), .air_in(c_9_0));
valve v_9_123 (.fluid_in(k_9_123), .fluid_out(k_8_61), .air_in(c_9_1));
valve v_9_124 (.fluid_in(k_9_124), .fluid_out(k_8_62), .air_in(c_9_0));
valve v_9_125 (.fluid_in(k_9_125), .fluid_out(k_8_62), .air_in(c_9_1));
valve v_9_126 (.fluid_in(k_9_126), .fluid_out(k_8_63), .air_in(c_9_0));
valve v_9_127 (.fluid_in(k_9_127), .fluid_out(k_8_63), .air_in(c_9_1));
valve v_9_128 (.fluid_in(k_9_128), .fluid_out(k_8_64), .air_in(c_9_0));
valve v_9_129 (.fluid_in(k_9_129), .fluid_out(k_8_64), .air_in(c_9_1));
valve v_9_130 (.fluid_in(k_9_130), .fluid_out(k_8_65), .air_in(c_9_0));
valve v_9_131 (.fluid_in(k_9_131), .fluid_out(k_8_65), .air_in(c_9_1));
valve v_9_132 (.fluid_in(k_9_132), .fluid_out(k_8_66), .air_in(c_9_0));
valve v_9_133 (.fluid_in(k_9_133), .fluid_out(k_8_66), .air_in(c_9_1));
valve v_9_134 (.fluid_in(k_9_134), .fluid_out(k_8_67), .air_in(c_9_0));
valve v_9_135 (.fluid_in(k_9_135), .fluid_out(k_8_67), .air_in(c_9_1));
valve v_9_136 (.fluid_in(k_9_136), .fluid_out(k_8_68), .air_in(c_9_0));
valve v_9_137 (.fluid_in(k_9_137), .fluid_out(k_8_68), .air_in(c_9_1));
valve v_9_138 (.fluid_in(k_9_138), .fluid_out(k_8_69), .air_in(c_9_0));
valve v_9_139 (.fluid_in(k_9_139), .fluid_out(k_8_69), .air_in(c_9_1));
valve v_9_140 (.fluid_in(k_9_140), .fluid_out(k_8_70), .air_in(c_9_0));
valve v_9_141 (.fluid_in(k_9_141), .fluid_out(k_8_70), .air_in(c_9_1));
valve v_9_142 (.fluid_in(k_9_142), .fluid_out(k_8_71), .air_in(c_9_0));
valve v_9_143 (.fluid_in(k_9_143), .fluid_out(k_8_71), .air_in(c_9_1));
valve v_9_144 (.fluid_in(k_9_144), .fluid_out(k_8_72), .air_in(c_9_0));
valve v_9_145 (.fluid_in(k_9_145), .fluid_out(k_8_72), .air_in(c_9_1));
valve v_9_146 (.fluid_in(k_9_146), .fluid_out(k_8_73), .air_in(c_9_0));
valve v_9_147 (.fluid_in(k_9_147), .fluid_out(k_8_73), .air_in(c_9_1));
valve v_9_148 (.fluid_in(k_9_148), .fluid_out(k_8_74), .air_in(c_9_0));
valve v_9_149 (.fluid_in(k_9_149), .fluid_out(k_8_74), .air_in(c_9_1));
valve v_9_150 (.fluid_in(k_9_150), .fluid_out(k_8_75), .air_in(c_9_0));
valve v_9_151 (.fluid_in(k_9_151), .fluid_out(k_8_75), .air_in(c_9_1));
valve v_9_152 (.fluid_in(k_9_152), .fluid_out(k_8_76), .air_in(c_9_0));
valve v_9_153 (.fluid_in(k_9_153), .fluid_out(k_8_76), .air_in(c_9_1));
valve v_9_154 (.fluid_in(k_9_154), .fluid_out(k_8_77), .air_in(c_9_0));
valve v_9_155 (.fluid_in(k_9_155), .fluid_out(k_8_77), .air_in(c_9_1));
valve v_9_156 (.fluid_in(k_9_156), .fluid_out(k_8_78), .air_in(c_9_0));
valve v_9_157 (.fluid_in(k_9_157), .fluid_out(k_8_78), .air_in(c_9_1));
valve v_9_158 (.fluid_in(k_9_158), .fluid_out(k_8_79), .air_in(c_9_0));
valve v_9_159 (.fluid_in(k_9_159), .fluid_out(k_8_79), .air_in(c_9_1));
valve v_9_160 (.fluid_in(k_9_160), .fluid_out(k_8_80), .air_in(c_9_0));
valve v_9_161 (.fluid_in(k_9_161), .fluid_out(k_8_80), .air_in(c_9_1));
valve v_9_162 (.fluid_in(k_9_162), .fluid_out(k_8_81), .air_in(c_9_0));
valve v_9_163 (.fluid_in(k_9_163), .fluid_out(k_8_81), .air_in(c_9_1));
valve v_9_164 (.fluid_in(k_9_164), .fluid_out(k_8_82), .air_in(c_9_0));
valve v_9_165 (.fluid_in(k_9_165), .fluid_out(k_8_82), .air_in(c_9_1));
valve v_9_166 (.fluid_in(k_9_166), .fluid_out(k_8_83), .air_in(c_9_0));
valve v_9_167 (.fluid_in(k_9_167), .fluid_out(k_8_83), .air_in(c_9_1));
valve v_9_168 (.fluid_in(k_9_168), .fluid_out(k_8_84), .air_in(c_9_0));
valve v_9_169 (.fluid_in(k_9_169), .fluid_out(k_8_84), .air_in(c_9_1));
valve v_9_170 (.fluid_in(k_9_170), .fluid_out(k_8_85), .air_in(c_9_0));
valve v_9_171 (.fluid_in(k_9_171), .fluid_out(k_8_85), .air_in(c_9_1));
valve v_9_172 (.fluid_in(k_9_172), .fluid_out(k_8_86), .air_in(c_9_0));
valve v_9_173 (.fluid_in(k_9_173), .fluid_out(k_8_86), .air_in(c_9_1));
valve v_9_174 (.fluid_in(k_9_174), .fluid_out(k_8_87), .air_in(c_9_0));
valve v_9_175 (.fluid_in(k_9_175), .fluid_out(k_8_87), .air_in(c_9_1));
valve v_9_176 (.fluid_in(k_9_176), .fluid_out(k_8_88), .air_in(c_9_0));
valve v_9_177 (.fluid_in(k_9_177), .fluid_out(k_8_88), .air_in(c_9_1));
valve v_9_178 (.fluid_in(k_9_178), .fluid_out(k_8_89), .air_in(c_9_0));
valve v_9_179 (.fluid_in(k_9_179), .fluid_out(k_8_89), .air_in(c_9_1));
valve v_9_180 (.fluid_in(k_9_180), .fluid_out(k_8_90), .air_in(c_9_0));
valve v_9_181 (.fluid_in(k_9_181), .fluid_out(k_8_90), .air_in(c_9_1));
valve v_9_182 (.fluid_in(k_9_182), .fluid_out(k_8_91), .air_in(c_9_0));
valve v_9_183 (.fluid_in(k_9_183), .fluid_out(k_8_91), .air_in(c_9_1));
valve v_9_184 (.fluid_in(k_9_184), .fluid_out(k_8_92), .air_in(c_9_0));
valve v_9_185 (.fluid_in(k_9_185), .fluid_out(k_8_92), .air_in(c_9_1));
valve v_9_186 (.fluid_in(k_9_186), .fluid_out(k_8_93), .air_in(c_9_0));
valve v_9_187 (.fluid_in(k_9_187), .fluid_out(k_8_93), .air_in(c_9_1));
valve v_9_188 (.fluid_in(k_9_188), .fluid_out(k_8_94), .air_in(c_9_0));
valve v_9_189 (.fluid_in(k_9_189), .fluid_out(k_8_94), .air_in(c_9_1));
valve v_9_190 (.fluid_in(k_9_190), .fluid_out(k_8_95), .air_in(c_9_0));
valve v_9_191 (.fluid_in(k_9_191), .fluid_out(k_8_95), .air_in(c_9_1));
valve v_9_192 (.fluid_in(k_9_192), .fluid_out(k_8_96), .air_in(c_9_0));
valve v_9_193 (.fluid_in(k_9_193), .fluid_out(k_8_96), .air_in(c_9_1));
valve v_9_194 (.fluid_in(k_9_194), .fluid_out(k_8_97), .air_in(c_9_0));
valve v_9_195 (.fluid_in(k_9_195), .fluid_out(k_8_97), .air_in(c_9_1));
valve v_9_196 (.fluid_in(k_9_196), .fluid_out(k_8_98), .air_in(c_9_0));
valve v_9_197 (.fluid_in(k_9_197), .fluid_out(k_8_98), .air_in(c_9_1));
valve v_9_198 (.fluid_in(k_9_198), .fluid_out(k_8_99), .air_in(c_9_0));
valve v_9_199 (.fluid_in(k_9_199), .fluid_out(k_8_99), .air_in(c_9_1));
valve v_9_200 (.fluid_in(k_9_200), .fluid_out(k_8_100), .air_in(c_9_0));
valve v_9_201 (.fluid_in(k_9_201), .fluid_out(k_8_100), .air_in(c_9_1));
valve v_9_202 (.fluid_in(k_9_202), .fluid_out(k_8_101), .air_in(c_9_0));
valve v_9_203 (.fluid_in(k_9_203), .fluid_out(k_8_101), .air_in(c_9_1));
valve v_9_204 (.fluid_in(k_9_204), .fluid_out(k_8_102), .air_in(c_9_0));
valve v_9_205 (.fluid_in(k_9_205), .fluid_out(k_8_102), .air_in(c_9_1));
valve v_9_206 (.fluid_in(k_9_206), .fluid_out(k_8_103), .air_in(c_9_0));
valve v_9_207 (.fluid_in(k_9_207), .fluid_out(k_8_103), .air_in(c_9_1));
valve v_9_208 (.fluid_in(k_9_208), .fluid_out(k_8_104), .air_in(c_9_0));
valve v_9_209 (.fluid_in(k_9_209), .fluid_out(k_8_104), .air_in(c_9_1));
valve v_9_210 (.fluid_in(k_9_210), .fluid_out(k_8_105), .air_in(c_9_0));
valve v_9_211 (.fluid_in(k_9_211), .fluid_out(k_8_105), .air_in(c_9_1));
valve v_9_212 (.fluid_in(k_9_212), .fluid_out(k_8_106), .air_in(c_9_0));
valve v_9_213 (.fluid_in(k_9_213), .fluid_out(k_8_106), .air_in(c_9_1));
valve v_9_214 (.fluid_in(k_9_214), .fluid_out(k_8_107), .air_in(c_9_0));
valve v_9_215 (.fluid_in(k_9_215), .fluid_out(k_8_107), .air_in(c_9_1));
valve v_9_216 (.fluid_in(k_9_216), .fluid_out(k_8_108), .air_in(c_9_0));
valve v_9_217 (.fluid_in(k_9_217), .fluid_out(k_8_108), .air_in(c_9_1));
valve v_9_218 (.fluid_in(k_9_218), .fluid_out(k_8_109), .air_in(c_9_0));
valve v_9_219 (.fluid_in(k_9_219), .fluid_out(k_8_109), .air_in(c_9_1));
valve v_9_220 (.fluid_in(k_9_220), .fluid_out(k_8_110), .air_in(c_9_0));
valve v_9_221 (.fluid_in(k_9_221), .fluid_out(k_8_110), .air_in(c_9_1));
valve v_9_222 (.fluid_in(k_9_222), .fluid_out(k_8_111), .air_in(c_9_0));
valve v_9_223 (.fluid_in(k_9_223), .fluid_out(k_8_111), .air_in(c_9_1));
valve v_9_224 (.fluid_in(k_9_224), .fluid_out(k_8_112), .air_in(c_9_0));
valve v_9_225 (.fluid_in(k_9_225), .fluid_out(k_8_112), .air_in(c_9_1));
valve v_9_226 (.fluid_in(k_9_226), .fluid_out(k_8_113), .air_in(c_9_0));
valve v_9_227 (.fluid_in(k_9_227), .fluid_out(k_8_113), .air_in(c_9_1));
valve v_9_228 (.fluid_in(k_9_228), .fluid_out(k_8_114), .air_in(c_9_0));
valve v_9_229 (.fluid_in(k_9_229), .fluid_out(k_8_114), .air_in(c_9_1));
valve v_9_230 (.fluid_in(k_9_230), .fluid_out(k_8_115), .air_in(c_9_0));
valve v_9_231 (.fluid_in(k_9_231), .fluid_out(k_8_115), .air_in(c_9_1));
valve v_9_232 (.fluid_in(k_9_232), .fluid_out(k_8_116), .air_in(c_9_0));
valve v_9_233 (.fluid_in(k_9_233), .fluid_out(k_8_116), .air_in(c_9_1));
valve v_9_234 (.fluid_in(k_9_234), .fluid_out(k_8_117), .air_in(c_9_0));
valve v_9_235 (.fluid_in(k_9_235), .fluid_out(k_8_117), .air_in(c_9_1));
valve v_9_236 (.fluid_in(k_9_236), .fluid_out(k_8_118), .air_in(c_9_0));
valve v_9_237 (.fluid_in(k_9_237), .fluid_out(k_8_118), .air_in(c_9_1));
valve v_9_238 (.fluid_in(k_9_238), .fluid_out(k_8_119), .air_in(c_9_0));
valve v_9_239 (.fluid_in(k_9_239), .fluid_out(k_8_119), .air_in(c_9_1));
valve v_9_240 (.fluid_in(k_9_240), .fluid_out(k_8_120), .air_in(c_9_0));
valve v_9_241 (.fluid_in(k_9_241), .fluid_out(k_8_120), .air_in(c_9_1));
valve v_9_242 (.fluid_in(k_9_242), .fluid_out(k_8_121), .air_in(c_9_0));
valve v_9_243 (.fluid_in(k_9_243), .fluid_out(k_8_121), .air_in(c_9_1));
valve v_9_244 (.fluid_in(k_9_244), .fluid_out(k_8_122), .air_in(c_9_0));
valve v_9_245 (.fluid_in(k_9_245), .fluid_out(k_8_122), .air_in(c_9_1));
valve v_9_246 (.fluid_in(k_9_246), .fluid_out(k_8_123), .air_in(c_9_0));
valve v_9_247 (.fluid_in(k_9_247), .fluid_out(k_8_123), .air_in(c_9_1));
valve v_9_248 (.fluid_in(k_9_248), .fluid_out(k_8_124), .air_in(c_9_0));
valve v_9_249 (.fluid_in(k_9_249), .fluid_out(k_8_124), .air_in(c_9_1));
valve v_9_250 (.fluid_in(k_9_250), .fluid_out(k_8_125), .air_in(c_9_0));
valve v_9_251 (.fluid_in(k_9_251), .fluid_out(k_8_125), .air_in(c_9_1));
valve v_9_252 (.fluid_in(k_9_252), .fluid_out(k_8_126), .air_in(c_9_0));
valve v_9_253 (.fluid_in(k_9_253), .fluid_out(k_8_126), .air_in(c_9_1));
valve v_9_254 (.fluid_in(k_9_254), .fluid_out(k_8_127), .air_in(c_9_0));
valve v_9_255 (.fluid_in(k_9_255), .fluid_out(k_8_127), .air_in(c_9_1));
valve v_9_256 (.fluid_in(k_9_256), .fluid_out(k_8_128), .air_in(c_9_0));
valve v_9_257 (.fluid_in(k_9_257), .fluid_out(k_8_128), .air_in(c_9_1));
valve v_9_258 (.fluid_in(k_9_258), .fluid_out(k_8_129), .air_in(c_9_0));
valve v_9_259 (.fluid_in(k_9_259), .fluid_out(k_8_129), .air_in(c_9_1));
valve v_9_260 (.fluid_in(k_9_260), .fluid_out(k_8_130), .air_in(c_9_0));
valve v_9_261 (.fluid_in(k_9_261), .fluid_out(k_8_130), .air_in(c_9_1));
valve v_9_262 (.fluid_in(k_9_262), .fluid_out(k_8_131), .air_in(c_9_0));
valve v_9_263 (.fluid_in(k_9_263), .fluid_out(k_8_131), .air_in(c_9_1));
valve v_9_264 (.fluid_in(k_9_264), .fluid_out(k_8_132), .air_in(c_9_0));
valve v_9_265 (.fluid_in(k_9_265), .fluid_out(k_8_132), .air_in(c_9_1));
valve v_9_266 (.fluid_in(k_9_266), .fluid_out(k_8_133), .air_in(c_9_0));
valve v_9_267 (.fluid_in(k_9_267), .fluid_out(k_8_133), .air_in(c_9_1));
valve v_9_268 (.fluid_in(k_9_268), .fluid_out(k_8_134), .air_in(c_9_0));
valve v_9_269 (.fluid_in(k_9_269), .fluid_out(k_8_134), .air_in(c_9_1));
valve v_9_270 (.fluid_in(k_9_270), .fluid_out(k_8_135), .air_in(c_9_0));
valve v_9_271 (.fluid_in(k_9_271), .fluid_out(k_8_135), .air_in(c_9_1));
valve v_9_272 (.fluid_in(k_9_272), .fluid_out(k_8_136), .air_in(c_9_0));
valve v_9_273 (.fluid_in(k_9_273), .fluid_out(k_8_136), .air_in(c_9_1));
valve v_9_274 (.fluid_in(k_9_274), .fluid_out(k_8_137), .air_in(c_9_0));
valve v_9_275 (.fluid_in(k_9_275), .fluid_out(k_8_137), .air_in(c_9_1));
valve v_9_276 (.fluid_in(k_9_276), .fluid_out(k_8_138), .air_in(c_9_0));
valve v_9_277 (.fluid_in(k_9_277), .fluid_out(k_8_138), .air_in(c_9_1));
valve v_9_278 (.fluid_in(k_9_278), .fluid_out(k_8_139), .air_in(c_9_0));
valve v_9_279 (.fluid_in(k_9_279), .fluid_out(k_8_139), .air_in(c_9_1));
valve v_9_280 (.fluid_in(k_9_280), .fluid_out(k_8_140), .air_in(c_9_0));
valve v_9_281 (.fluid_in(k_9_281), .fluid_out(k_8_140), .air_in(c_9_1));
valve v_9_282 (.fluid_in(k_9_282), .fluid_out(k_8_141), .air_in(c_9_0));
valve v_9_283 (.fluid_in(k_9_283), .fluid_out(k_8_141), .air_in(c_9_1));
valve v_9_284 (.fluid_in(k_9_284), .fluid_out(k_8_142), .air_in(c_9_0));
valve v_9_285 (.fluid_in(k_9_285), .fluid_out(k_8_142), .air_in(c_9_1));
valve v_9_286 (.fluid_in(k_9_286), .fluid_out(k_8_143), .air_in(c_9_0));
valve v_9_287 (.fluid_in(k_9_287), .fluid_out(k_8_143), .air_in(c_9_1));
valve v_9_288 (.fluid_in(k_9_288), .fluid_out(k_8_144), .air_in(c_9_0));
valve v_9_289 (.fluid_in(k_9_289), .fluid_out(k_8_144), .air_in(c_9_1));
valve v_9_290 (.fluid_in(k_9_290), .fluid_out(k_8_145), .air_in(c_9_0));
valve v_9_291 (.fluid_in(k_9_291), .fluid_out(k_8_145), .air_in(c_9_1));
valve v_9_292 (.fluid_in(k_9_292), .fluid_out(k_8_146), .air_in(c_9_0));
valve v_9_293 (.fluid_in(k_9_293), .fluid_out(k_8_146), .air_in(c_9_1));
valve v_9_294 (.fluid_in(k_9_294), .fluid_out(k_8_147), .air_in(c_9_0));
valve v_9_295 (.fluid_in(k_9_295), .fluid_out(k_8_147), .air_in(c_9_1));
valve v_9_296 (.fluid_in(k_9_296), .fluid_out(k_8_148), .air_in(c_9_0));
valve v_9_297 (.fluid_in(k_9_297), .fluid_out(k_8_148), .air_in(c_9_1));
valve v_9_298 (.fluid_in(k_9_298), .fluid_out(k_8_149), .air_in(c_9_0));
valve v_9_299 (.fluid_in(k_9_299), .fluid_out(k_8_149), .air_in(c_9_1));
valve v_9_300 (.fluid_in(k_9_300), .fluid_out(k_8_150), .air_in(c_9_0));
valve v_9_301 (.fluid_in(k_9_301), .fluid_out(k_8_150), .air_in(c_9_1));
valve v_9_302 (.fluid_in(k_9_302), .fluid_out(k_8_151), .air_in(c_9_0));
valve v_9_303 (.fluid_in(k_9_303), .fluid_out(k_8_151), .air_in(c_9_1));
valve v_9_304 (.fluid_in(k_9_304), .fluid_out(k_8_152), .air_in(c_9_0));
valve v_9_305 (.fluid_in(k_9_305), .fluid_out(k_8_152), .air_in(c_9_1));
valve v_9_306 (.fluid_in(k_9_306), .fluid_out(k_8_153), .air_in(c_9_0));
valve v_9_307 (.fluid_in(k_9_307), .fluid_out(k_8_153), .air_in(c_9_1));
valve v_9_308 (.fluid_in(k_9_308), .fluid_out(k_8_154), .air_in(c_9_0));
valve v_9_309 (.fluid_in(k_9_309), .fluid_out(k_8_154), .air_in(c_9_1));
valve v_9_310 (.fluid_in(k_9_310), .fluid_out(k_8_155), .air_in(c_9_0));
valve v_9_311 (.fluid_in(k_9_311), .fluid_out(k_8_155), .air_in(c_9_1));
valve v_9_312 (.fluid_in(k_9_312), .fluid_out(k_8_156), .air_in(c_9_0));
valve v_9_313 (.fluid_in(k_9_313), .fluid_out(k_8_156), .air_in(c_9_1));
valve v_9_314 (.fluid_in(k_9_314), .fluid_out(k_8_157), .air_in(c_9_0));
valve v_9_315 (.fluid_in(k_9_315), .fluid_out(k_8_157), .air_in(c_9_1));
valve v_9_316 (.fluid_in(k_9_316), .fluid_out(k_8_158), .air_in(c_9_0));
valve v_9_317 (.fluid_in(k_9_317), .fluid_out(k_8_158), .air_in(c_9_1));
valve v_9_318 (.fluid_in(k_9_318), .fluid_out(k_8_159), .air_in(c_9_0));
valve v_9_319 (.fluid_in(k_9_319), .fluid_out(k_8_159), .air_in(c_9_1));
valve v_9_320 (.fluid_in(k_9_320), .fluid_out(k_8_160), .air_in(c_9_0));
valve v_9_321 (.fluid_in(k_9_321), .fluid_out(k_8_160), .air_in(c_9_1));
valve v_9_322 (.fluid_in(k_9_322), .fluid_out(k_8_161), .air_in(c_9_0));
valve v_9_323 (.fluid_in(k_9_323), .fluid_out(k_8_161), .air_in(c_9_1));
valve v_9_324 (.fluid_in(k_9_324), .fluid_out(k_8_162), .air_in(c_9_0));
valve v_9_325 (.fluid_in(k_9_325), .fluid_out(k_8_162), .air_in(c_9_1));
valve v_9_326 (.fluid_in(k_9_326), .fluid_out(k_8_163), .air_in(c_9_0));
valve v_9_327 (.fluid_in(k_9_327), .fluid_out(k_8_163), .air_in(c_9_1));
valve v_9_328 (.fluid_in(k_9_328), .fluid_out(k_8_164), .air_in(c_9_0));
valve v_9_329 (.fluid_in(k_9_329), .fluid_out(k_8_164), .air_in(c_9_1));
valve v_9_330 (.fluid_in(k_9_330), .fluid_out(k_8_165), .air_in(c_9_0));
valve v_9_331 (.fluid_in(k_9_331), .fluid_out(k_8_165), .air_in(c_9_1));
valve v_9_332 (.fluid_in(k_9_332), .fluid_out(k_8_166), .air_in(c_9_0));
valve v_9_333 (.fluid_in(k_9_333), .fluid_out(k_8_166), .air_in(c_9_1));
valve v_9_334 (.fluid_in(k_9_334), .fluid_out(k_8_167), .air_in(c_9_0));
valve v_9_335 (.fluid_in(k_9_335), .fluid_out(k_8_167), .air_in(c_9_1));
valve v_9_336 (.fluid_in(k_9_336), .fluid_out(k_8_168), .air_in(c_9_0));
valve v_9_337 (.fluid_in(k_9_337), .fluid_out(k_8_168), .air_in(c_9_1));
valve v_9_338 (.fluid_in(k_9_338), .fluid_out(k_8_169), .air_in(c_9_0));
valve v_9_339 (.fluid_in(k_9_339), .fluid_out(k_8_169), .air_in(c_9_1));
valve v_9_340 (.fluid_in(k_9_340), .fluid_out(k_8_170), .air_in(c_9_0));
valve v_9_341 (.fluid_in(k_9_341), .fluid_out(k_8_170), .air_in(c_9_1));
valve v_9_342 (.fluid_in(k_9_342), .fluid_out(k_8_171), .air_in(c_9_0));
valve v_9_343 (.fluid_in(k_9_343), .fluid_out(k_8_171), .air_in(c_9_1));
valve v_9_344 (.fluid_in(k_9_344), .fluid_out(k_8_172), .air_in(c_9_0));
valve v_9_345 (.fluid_in(k_9_345), .fluid_out(k_8_172), .air_in(c_9_1));
valve v_9_346 (.fluid_in(k_9_346), .fluid_out(k_8_173), .air_in(c_9_0));
valve v_9_347 (.fluid_in(k_9_347), .fluid_out(k_8_173), .air_in(c_9_1));
valve v_9_348 (.fluid_in(k_9_348), .fluid_out(k_8_174), .air_in(c_9_0));
valve v_9_349 (.fluid_in(k_9_349), .fluid_out(k_8_174), .air_in(c_9_1));
valve v_9_350 (.fluid_in(k_9_350), .fluid_out(k_8_175), .air_in(c_9_0));
valve v_9_351 (.fluid_in(k_9_351), .fluid_out(k_8_175), .air_in(c_9_1));
valve v_9_352 (.fluid_in(k_9_352), .fluid_out(k_8_176), .air_in(c_9_0));
valve v_9_353 (.fluid_in(k_9_353), .fluid_out(k_8_176), .air_in(c_9_1));
valve v_9_354 (.fluid_in(k_9_354), .fluid_out(k_8_177), .air_in(c_9_0));
valve v_9_355 (.fluid_in(k_9_355), .fluid_out(k_8_177), .air_in(c_9_1));
valve v_9_356 (.fluid_in(k_9_356), .fluid_out(k_8_178), .air_in(c_9_0));
valve v_9_357 (.fluid_in(k_9_357), .fluid_out(k_8_178), .air_in(c_9_1));
valve v_9_358 (.fluid_in(k_9_358), .fluid_out(k_8_179), .air_in(c_9_0));
valve v_9_359 (.fluid_in(k_9_359), .fluid_out(k_8_179), .air_in(c_9_1));
valve v_9_360 (.fluid_in(k_9_360), .fluid_out(k_8_180), .air_in(c_9_0));
valve v_9_361 (.fluid_in(k_9_361), .fluid_out(k_8_180), .air_in(c_9_1));
valve v_9_362 (.fluid_in(k_9_362), .fluid_out(k_8_181), .air_in(c_9_0));
valve v_9_363 (.fluid_in(k_9_363), .fluid_out(k_8_181), .air_in(c_9_1));
valve v_9_364 (.fluid_in(k_9_364), .fluid_out(k_8_182), .air_in(c_9_0));
valve v_9_365 (.fluid_in(k_9_365), .fluid_out(k_8_182), .air_in(c_9_1));
valve v_9_366 (.fluid_in(k_9_366), .fluid_out(k_8_183), .air_in(c_9_0));
valve v_9_367 (.fluid_in(k_9_367), .fluid_out(k_8_183), .air_in(c_9_1));
valve v_9_368 (.fluid_in(k_9_368), .fluid_out(k_8_184), .air_in(c_9_0));
valve v_9_369 (.fluid_in(k_9_369), .fluid_out(k_8_184), .air_in(c_9_1));
valve v_9_370 (.fluid_in(k_9_370), .fluid_out(k_8_185), .air_in(c_9_0));
valve v_9_371 (.fluid_in(k_9_371), .fluid_out(k_8_185), .air_in(c_9_1));
valve v_9_372 (.fluid_in(k_9_372), .fluid_out(k_8_186), .air_in(c_9_0));
valve v_9_373 (.fluid_in(k_9_373), .fluid_out(k_8_186), .air_in(c_9_1));
valve v_9_374 (.fluid_in(k_9_374), .fluid_out(k_8_187), .air_in(c_9_0));
valve v_9_375 (.fluid_in(k_9_375), .fluid_out(k_8_187), .air_in(c_9_1));
valve v_9_376 (.fluid_in(k_9_376), .fluid_out(k_8_188), .air_in(c_9_0));
valve v_9_377 (.fluid_in(k_9_377), .fluid_out(k_8_188), .air_in(c_9_1));
valve v_9_378 (.fluid_in(k_9_378), .fluid_out(k_8_189), .air_in(c_9_0));
valve v_9_379 (.fluid_in(k_9_379), .fluid_out(k_8_189), .air_in(c_9_1));
valve v_9_380 (.fluid_in(k_9_380), .fluid_out(k_8_190), .air_in(c_9_0));
valve v_9_381 (.fluid_in(k_9_381), .fluid_out(k_8_190), .air_in(c_9_1));
valve v_9_382 (.fluid_in(k_9_382), .fluid_out(k_8_191), .air_in(c_9_0));
valve v_9_383 (.fluid_in(k_9_383), .fluid_out(k_8_191), .air_in(c_9_1));
valve v_9_384 (.fluid_in(k_9_384), .fluid_out(k_8_192), .air_in(c_9_0));
valve v_9_385 (.fluid_in(k_9_385), .fluid_out(k_8_192), .air_in(c_9_1));
valve v_9_386 (.fluid_in(k_9_386), .fluid_out(k_8_193), .air_in(c_9_0));
valve v_9_387 (.fluid_in(k_9_387), .fluid_out(k_8_193), .air_in(c_9_1));
valve v_9_388 (.fluid_in(k_9_388), .fluid_out(k_8_194), .air_in(c_9_0));
valve v_9_389 (.fluid_in(k_9_389), .fluid_out(k_8_194), .air_in(c_9_1));
valve v_9_390 (.fluid_in(k_9_390), .fluid_out(k_8_195), .air_in(c_9_0));
valve v_9_391 (.fluid_in(k_9_391), .fluid_out(k_8_195), .air_in(c_9_1));
valve v_9_392 (.fluid_in(k_9_392), .fluid_out(k_8_196), .air_in(c_9_0));
valve v_9_393 (.fluid_in(k_9_393), .fluid_out(k_8_196), .air_in(c_9_1));
valve v_9_394 (.fluid_in(k_9_394), .fluid_out(k_8_197), .air_in(c_9_0));
valve v_9_395 (.fluid_in(k_9_395), .fluid_out(k_8_197), .air_in(c_9_1));
valve v_9_396 (.fluid_in(k_9_396), .fluid_out(k_8_198), .air_in(c_9_0));
valve v_9_397 (.fluid_in(k_9_397), .fluid_out(k_8_198), .air_in(c_9_1));
valve v_9_398 (.fluid_in(k_9_398), .fluid_out(k_8_199), .air_in(c_9_0));
valve v_9_399 (.fluid_in(k_9_399), .fluid_out(k_8_199), .air_in(c_9_1));
valve v_9_400 (.fluid_in(k_9_400), .fluid_out(k_8_200), .air_in(c_9_0));
valve v_9_401 (.fluid_in(k_9_401), .fluid_out(k_8_200), .air_in(c_9_1));
valve v_9_402 (.fluid_in(k_9_402), .fluid_out(k_8_201), .air_in(c_9_0));
valve v_9_403 (.fluid_in(k_9_403), .fluid_out(k_8_201), .air_in(c_9_1));
valve v_9_404 (.fluid_in(k_9_404), .fluid_out(k_8_202), .air_in(c_9_0));
valve v_9_405 (.fluid_in(k_9_405), .fluid_out(k_8_202), .air_in(c_9_1));
valve v_9_406 (.fluid_in(k_9_406), .fluid_out(k_8_203), .air_in(c_9_0));
valve v_9_407 (.fluid_in(k_9_407), .fluid_out(k_8_203), .air_in(c_9_1));
valve v_9_408 (.fluid_in(k_9_408), .fluid_out(k_8_204), .air_in(c_9_0));
valve v_9_409 (.fluid_in(k_9_409), .fluid_out(k_8_204), .air_in(c_9_1));
valve v_9_410 (.fluid_in(k_9_410), .fluid_out(k_8_205), .air_in(c_9_0));
valve v_9_411 (.fluid_in(k_9_411), .fluid_out(k_8_205), .air_in(c_9_1));
valve v_9_412 (.fluid_in(k_9_412), .fluid_out(k_8_206), .air_in(c_9_0));
valve v_9_413 (.fluid_in(k_9_413), .fluid_out(k_8_206), .air_in(c_9_1));
valve v_9_414 (.fluid_in(k_9_414), .fluid_out(k_8_207), .air_in(c_9_0));
valve v_9_415 (.fluid_in(k_9_415), .fluid_out(k_8_207), .air_in(c_9_1));
valve v_9_416 (.fluid_in(k_9_416), .fluid_out(k_8_208), .air_in(c_9_0));
valve v_9_417 (.fluid_in(k_9_417), .fluid_out(k_8_208), .air_in(c_9_1));
valve v_9_418 (.fluid_in(k_9_418), .fluid_out(k_8_209), .air_in(c_9_0));
valve v_9_419 (.fluid_in(k_9_419), .fluid_out(k_8_209), .air_in(c_9_1));
valve v_9_420 (.fluid_in(k_9_420), .fluid_out(k_8_210), .air_in(c_9_0));
valve v_9_421 (.fluid_in(k_9_421), .fluid_out(k_8_210), .air_in(c_9_1));
valve v_9_422 (.fluid_in(k_9_422), .fluid_out(k_8_211), .air_in(c_9_0));
valve v_9_423 (.fluid_in(k_9_423), .fluid_out(k_8_211), .air_in(c_9_1));
valve v_9_424 (.fluid_in(k_9_424), .fluid_out(k_8_212), .air_in(c_9_0));
valve v_9_425 (.fluid_in(k_9_425), .fluid_out(k_8_212), .air_in(c_9_1));
valve v_9_426 (.fluid_in(k_9_426), .fluid_out(k_8_213), .air_in(c_9_0));
valve v_9_427 (.fluid_in(k_9_427), .fluid_out(k_8_213), .air_in(c_9_1));
valve v_9_428 (.fluid_in(k_9_428), .fluid_out(k_8_214), .air_in(c_9_0));
valve v_9_429 (.fluid_in(k_9_429), .fluid_out(k_8_214), .air_in(c_9_1));
valve v_9_430 (.fluid_in(k_9_430), .fluid_out(k_8_215), .air_in(c_9_0));
valve v_9_431 (.fluid_in(k_9_431), .fluid_out(k_8_215), .air_in(c_9_1));
valve v_9_432 (.fluid_in(k_9_432), .fluid_out(k_8_216), .air_in(c_9_0));
valve v_9_433 (.fluid_in(k_9_433), .fluid_out(k_8_216), .air_in(c_9_1));
valve v_9_434 (.fluid_in(k_9_434), .fluid_out(k_8_217), .air_in(c_9_0));
valve v_9_435 (.fluid_in(k_9_435), .fluid_out(k_8_217), .air_in(c_9_1));
valve v_9_436 (.fluid_in(k_9_436), .fluid_out(k_8_218), .air_in(c_9_0));
valve v_9_437 (.fluid_in(k_9_437), .fluid_out(k_8_218), .air_in(c_9_1));
valve v_9_438 (.fluid_in(k_9_438), .fluid_out(k_8_219), .air_in(c_9_0));
valve v_9_439 (.fluid_in(k_9_439), .fluid_out(k_8_219), .air_in(c_9_1));
valve v_9_440 (.fluid_in(k_9_440), .fluid_out(k_8_220), .air_in(c_9_0));
valve v_9_441 (.fluid_in(k_9_441), .fluid_out(k_8_220), .air_in(c_9_1));
valve v_9_442 (.fluid_in(k_9_442), .fluid_out(k_8_221), .air_in(c_9_0));
valve v_9_443 (.fluid_in(k_9_443), .fluid_out(k_8_221), .air_in(c_9_1));
valve v_9_444 (.fluid_in(k_9_444), .fluid_out(k_8_222), .air_in(c_9_0));
valve v_9_445 (.fluid_in(k_9_445), .fluid_out(k_8_222), .air_in(c_9_1));
valve v_9_446 (.fluid_in(k_9_446), .fluid_out(k_8_223), .air_in(c_9_0));
valve v_9_447 (.fluid_in(k_9_447), .fluid_out(k_8_223), .air_in(c_9_1));
valve v_9_448 (.fluid_in(k_9_448), .fluid_out(k_8_224), .air_in(c_9_0));
valve v_9_449 (.fluid_in(k_9_449), .fluid_out(k_8_224), .air_in(c_9_1));
valve v_9_450 (.fluid_in(k_9_450), .fluid_out(k_8_225), .air_in(c_9_0));
valve v_9_451 (.fluid_in(k_9_451), .fluid_out(k_8_225), .air_in(c_9_1));
valve v_9_452 (.fluid_in(k_9_452), .fluid_out(k_8_226), .air_in(c_9_0));
valve v_9_453 (.fluid_in(k_9_453), .fluid_out(k_8_226), .air_in(c_9_1));
valve v_9_454 (.fluid_in(k_9_454), .fluid_out(k_8_227), .air_in(c_9_0));
valve v_9_455 (.fluid_in(k_9_455), .fluid_out(k_8_227), .air_in(c_9_1));
valve v_9_456 (.fluid_in(k_9_456), .fluid_out(k_8_228), .air_in(c_9_0));
valve v_9_457 (.fluid_in(k_9_457), .fluid_out(k_8_228), .air_in(c_9_1));
valve v_9_458 (.fluid_in(k_9_458), .fluid_out(k_8_229), .air_in(c_9_0));
valve v_9_459 (.fluid_in(k_9_459), .fluid_out(k_8_229), .air_in(c_9_1));
valve v_9_460 (.fluid_in(k_9_460), .fluid_out(k_8_230), .air_in(c_9_0));
valve v_9_461 (.fluid_in(k_9_461), .fluid_out(k_8_230), .air_in(c_9_1));
valve v_9_462 (.fluid_in(k_9_462), .fluid_out(k_8_231), .air_in(c_9_0));
valve v_9_463 (.fluid_in(k_9_463), .fluid_out(k_8_231), .air_in(c_9_1));
valve v_9_464 (.fluid_in(k_9_464), .fluid_out(k_8_232), .air_in(c_9_0));
valve v_9_465 (.fluid_in(k_9_465), .fluid_out(k_8_232), .air_in(c_9_1));
valve v_9_466 (.fluid_in(k_9_466), .fluid_out(k_8_233), .air_in(c_9_0));
valve v_9_467 (.fluid_in(k_9_467), .fluid_out(k_8_233), .air_in(c_9_1));
valve v_9_468 (.fluid_in(k_9_468), .fluid_out(k_8_234), .air_in(c_9_0));
valve v_9_469 (.fluid_in(k_9_469), .fluid_out(k_8_234), .air_in(c_9_1));
valve v_9_470 (.fluid_in(k_9_470), .fluid_out(k_8_235), .air_in(c_9_0));
valve v_9_471 (.fluid_in(k_9_471), .fluid_out(k_8_235), .air_in(c_9_1));
valve v_9_472 (.fluid_in(k_9_472), .fluid_out(k_8_236), .air_in(c_9_0));
valve v_9_473 (.fluid_in(k_9_473), .fluid_out(k_8_236), .air_in(c_9_1));
valve v_9_474 (.fluid_in(k_9_474), .fluid_out(k_8_237), .air_in(c_9_0));
valve v_9_475 (.fluid_in(k_9_475), .fluid_out(k_8_237), .air_in(c_9_1));
valve v_9_476 (.fluid_in(k_9_476), .fluid_out(k_8_238), .air_in(c_9_0));
valve v_9_477 (.fluid_in(k_9_477), .fluid_out(k_8_238), .air_in(c_9_1));
valve v_9_478 (.fluid_in(k_9_478), .fluid_out(k_8_239), .air_in(c_9_0));
valve v_9_479 (.fluid_in(k_9_479), .fluid_out(k_8_239), .air_in(c_9_1));
valve v_9_480 (.fluid_in(k_9_480), .fluid_out(k_8_240), .air_in(c_9_0));
valve v_9_481 (.fluid_in(k_9_481), .fluid_out(k_8_240), .air_in(c_9_1));
valve v_9_482 (.fluid_in(k_9_482), .fluid_out(k_8_241), .air_in(c_9_0));
valve v_9_483 (.fluid_in(k_9_483), .fluid_out(k_8_241), .air_in(c_9_1));
valve v_9_484 (.fluid_in(k_9_484), .fluid_out(k_8_242), .air_in(c_9_0));
valve v_9_485 (.fluid_in(k_9_485), .fluid_out(k_8_242), .air_in(c_9_1));
valve v_9_486 (.fluid_in(k_9_486), .fluid_out(k_8_243), .air_in(c_9_0));
valve v_9_487 (.fluid_in(k_9_487), .fluid_out(k_8_243), .air_in(c_9_1));
valve v_9_488 (.fluid_in(k_9_488), .fluid_out(k_8_244), .air_in(c_9_0));
valve v_9_489 (.fluid_in(k_9_489), .fluid_out(k_8_244), .air_in(c_9_1));
valve v_9_490 (.fluid_in(k_9_490), .fluid_out(k_8_245), .air_in(c_9_0));
valve v_9_491 (.fluid_in(k_9_491), .fluid_out(k_8_245), .air_in(c_9_1));
valve v_9_492 (.fluid_in(k_9_492), .fluid_out(k_8_246), .air_in(c_9_0));
valve v_9_493 (.fluid_in(k_9_493), .fluid_out(k_8_246), .air_in(c_9_1));
valve v_9_494 (.fluid_in(k_9_494), .fluid_out(k_8_247), .air_in(c_9_0));
valve v_9_495 (.fluid_in(k_9_495), .fluid_out(k_8_247), .air_in(c_9_1));
valve v_9_496 (.fluid_in(k_9_496), .fluid_out(k_8_248), .air_in(c_9_0));
valve v_9_497 (.fluid_in(k_9_497), .fluid_out(k_8_248), .air_in(c_9_1));
valve v_9_498 (.fluid_in(k_9_498), .fluid_out(k_8_249), .air_in(c_9_0));
valve v_9_499 (.fluid_in(k_9_499), .fluid_out(k_8_249), .air_in(c_9_1));
valve v_9_500 (.fluid_in(k_9_500), .fluid_out(k_8_250), .air_in(c_9_0));
valve v_9_501 (.fluid_in(k_9_501), .fluid_out(k_8_250), .air_in(c_9_1));
valve v_9_502 (.fluid_in(k_9_502), .fluid_out(k_8_251), .air_in(c_9_0));
valve v_9_503 (.fluid_in(k_9_503), .fluid_out(k_8_251), .air_in(c_9_1));
valve v_9_504 (.fluid_in(k_9_504), .fluid_out(k_8_252), .air_in(c_9_0));
valve v_9_505 (.fluid_in(k_9_505), .fluid_out(k_8_252), .air_in(c_9_1));
valve v_9_506 (.fluid_in(k_9_506), .fluid_out(k_8_253), .air_in(c_9_0));
valve v_9_507 (.fluid_in(k_9_507), .fluid_out(k_8_253), .air_in(c_9_1));
valve v_9_508 (.fluid_in(k_9_508), .fluid_out(k_8_254), .air_in(c_9_0));
valve v_9_509 (.fluid_in(k_9_509), .fluid_out(k_8_254), .air_in(c_9_1));
valve v_9_510 (.fluid_in(k_9_510), .fluid_out(k_8_255), .air_in(c_9_0));
valve v_9_511 (.fluid_in(k_9_511), .fluid_out(k_8_255), .air_in(c_9_1));
valve v_10_0 (.fluid_in(k_10_0), .fluid_out(k_9_0), .air_in(c_10_0));
valve v_10_1 (.fluid_in(k_10_1), .fluid_out(k_9_0), .air_in(c_10_1));
valve v_10_2 (.fluid_in(k_10_2), .fluid_out(k_9_1), .air_in(c_10_0));
valve v_10_3 (.fluid_in(k_10_3), .fluid_out(k_9_1), .air_in(c_10_1));
valve v_10_4 (.fluid_in(k_10_4), .fluid_out(k_9_2), .air_in(c_10_0));
valve v_10_5 (.fluid_in(k_10_5), .fluid_out(k_9_2), .air_in(c_10_1));
valve v_10_6 (.fluid_in(k_10_6), .fluid_out(k_9_3), .air_in(c_10_0));
valve v_10_7 (.fluid_in(k_10_7), .fluid_out(k_9_3), .air_in(c_10_1));
valve v_10_8 (.fluid_in(k_10_8), .fluid_out(k_9_4), .air_in(c_10_0));
valve v_10_9 (.fluid_in(k_10_9), .fluid_out(k_9_4), .air_in(c_10_1));
valve v_10_10 (.fluid_in(k_10_10), .fluid_out(k_9_5), .air_in(c_10_0));
valve v_10_11 (.fluid_in(k_10_11), .fluid_out(k_9_5), .air_in(c_10_1));
valve v_10_12 (.fluid_in(k_10_12), .fluid_out(k_9_6), .air_in(c_10_0));
valve v_10_13 (.fluid_in(k_10_13), .fluid_out(k_9_6), .air_in(c_10_1));
valve v_10_14 (.fluid_in(k_10_14), .fluid_out(k_9_7), .air_in(c_10_0));
valve v_10_15 (.fluid_in(k_10_15), .fluid_out(k_9_7), .air_in(c_10_1));
valve v_10_16 (.fluid_in(k_10_16), .fluid_out(k_9_8), .air_in(c_10_0));
valve v_10_17 (.fluid_in(k_10_17), .fluid_out(k_9_8), .air_in(c_10_1));
valve v_10_18 (.fluid_in(k_10_18), .fluid_out(k_9_9), .air_in(c_10_0));
valve v_10_19 (.fluid_in(k_10_19), .fluid_out(k_9_9), .air_in(c_10_1));
valve v_10_20 (.fluid_in(k_10_20), .fluid_out(k_9_10), .air_in(c_10_0));
valve v_10_21 (.fluid_in(k_10_21), .fluid_out(k_9_10), .air_in(c_10_1));
valve v_10_22 (.fluid_in(k_10_22), .fluid_out(k_9_11), .air_in(c_10_0));
valve v_10_23 (.fluid_in(k_10_23), .fluid_out(k_9_11), .air_in(c_10_1));
valve v_10_24 (.fluid_in(k_10_24), .fluid_out(k_9_12), .air_in(c_10_0));
valve v_10_25 (.fluid_in(k_10_25), .fluid_out(k_9_12), .air_in(c_10_1));
valve v_10_26 (.fluid_in(k_10_26), .fluid_out(k_9_13), .air_in(c_10_0));
valve v_10_27 (.fluid_in(k_10_27), .fluid_out(k_9_13), .air_in(c_10_1));
valve v_10_28 (.fluid_in(k_10_28), .fluid_out(k_9_14), .air_in(c_10_0));
valve v_10_29 (.fluid_in(k_10_29), .fluid_out(k_9_14), .air_in(c_10_1));
valve v_10_30 (.fluid_in(k_10_30), .fluid_out(k_9_15), .air_in(c_10_0));
valve v_10_31 (.fluid_in(k_10_31), .fluid_out(k_9_15), .air_in(c_10_1));
valve v_10_32 (.fluid_in(k_10_32), .fluid_out(k_9_16), .air_in(c_10_0));
valve v_10_33 (.fluid_in(k_10_33), .fluid_out(k_9_16), .air_in(c_10_1));
valve v_10_34 (.fluid_in(k_10_34), .fluid_out(k_9_17), .air_in(c_10_0));
valve v_10_35 (.fluid_in(k_10_35), .fluid_out(k_9_17), .air_in(c_10_1));
valve v_10_36 (.fluid_in(k_10_36), .fluid_out(k_9_18), .air_in(c_10_0));
valve v_10_37 (.fluid_in(k_10_37), .fluid_out(k_9_18), .air_in(c_10_1));
valve v_10_38 (.fluid_in(k_10_38), .fluid_out(k_9_19), .air_in(c_10_0));
valve v_10_39 (.fluid_in(k_10_39), .fluid_out(k_9_19), .air_in(c_10_1));
valve v_10_40 (.fluid_in(k_10_40), .fluid_out(k_9_20), .air_in(c_10_0));
valve v_10_41 (.fluid_in(k_10_41), .fluid_out(k_9_20), .air_in(c_10_1));
valve v_10_42 (.fluid_in(k_10_42), .fluid_out(k_9_21), .air_in(c_10_0));
valve v_10_43 (.fluid_in(k_10_43), .fluid_out(k_9_21), .air_in(c_10_1));
valve v_10_44 (.fluid_in(k_10_44), .fluid_out(k_9_22), .air_in(c_10_0));
valve v_10_45 (.fluid_in(k_10_45), .fluid_out(k_9_22), .air_in(c_10_1));
valve v_10_46 (.fluid_in(k_10_46), .fluid_out(k_9_23), .air_in(c_10_0));
valve v_10_47 (.fluid_in(k_10_47), .fluid_out(k_9_23), .air_in(c_10_1));
valve v_10_48 (.fluid_in(k_10_48), .fluid_out(k_9_24), .air_in(c_10_0));
valve v_10_49 (.fluid_in(k_10_49), .fluid_out(k_9_24), .air_in(c_10_1));
valve v_10_50 (.fluid_in(k_10_50), .fluid_out(k_9_25), .air_in(c_10_0));
valve v_10_51 (.fluid_in(k_10_51), .fluid_out(k_9_25), .air_in(c_10_1));
valve v_10_52 (.fluid_in(k_10_52), .fluid_out(k_9_26), .air_in(c_10_0));
valve v_10_53 (.fluid_in(k_10_53), .fluid_out(k_9_26), .air_in(c_10_1));
valve v_10_54 (.fluid_in(k_10_54), .fluid_out(k_9_27), .air_in(c_10_0));
valve v_10_55 (.fluid_in(k_10_55), .fluid_out(k_9_27), .air_in(c_10_1));
valve v_10_56 (.fluid_in(k_10_56), .fluid_out(k_9_28), .air_in(c_10_0));
valve v_10_57 (.fluid_in(k_10_57), .fluid_out(k_9_28), .air_in(c_10_1));
valve v_10_58 (.fluid_in(k_10_58), .fluid_out(k_9_29), .air_in(c_10_0));
valve v_10_59 (.fluid_in(k_10_59), .fluid_out(k_9_29), .air_in(c_10_1));
valve v_10_60 (.fluid_in(k_10_60), .fluid_out(k_9_30), .air_in(c_10_0));
valve v_10_61 (.fluid_in(k_10_61), .fluid_out(k_9_30), .air_in(c_10_1));
valve v_10_62 (.fluid_in(k_10_62), .fluid_out(k_9_31), .air_in(c_10_0));
valve v_10_63 (.fluid_in(k_10_63), .fluid_out(k_9_31), .air_in(c_10_1));
valve v_10_64 (.fluid_in(k_10_64), .fluid_out(k_9_32), .air_in(c_10_0));
valve v_10_65 (.fluid_in(k_10_65), .fluid_out(k_9_32), .air_in(c_10_1));
valve v_10_66 (.fluid_in(k_10_66), .fluid_out(k_9_33), .air_in(c_10_0));
valve v_10_67 (.fluid_in(k_10_67), .fluid_out(k_9_33), .air_in(c_10_1));
valve v_10_68 (.fluid_in(k_10_68), .fluid_out(k_9_34), .air_in(c_10_0));
valve v_10_69 (.fluid_in(k_10_69), .fluid_out(k_9_34), .air_in(c_10_1));
valve v_10_70 (.fluid_in(k_10_70), .fluid_out(k_9_35), .air_in(c_10_0));
valve v_10_71 (.fluid_in(k_10_71), .fluid_out(k_9_35), .air_in(c_10_1));
valve v_10_72 (.fluid_in(k_10_72), .fluid_out(k_9_36), .air_in(c_10_0));
valve v_10_73 (.fluid_in(k_10_73), .fluid_out(k_9_36), .air_in(c_10_1));
valve v_10_74 (.fluid_in(k_10_74), .fluid_out(k_9_37), .air_in(c_10_0));
valve v_10_75 (.fluid_in(k_10_75), .fluid_out(k_9_37), .air_in(c_10_1));
valve v_10_76 (.fluid_in(k_10_76), .fluid_out(k_9_38), .air_in(c_10_0));
valve v_10_77 (.fluid_in(k_10_77), .fluid_out(k_9_38), .air_in(c_10_1));
valve v_10_78 (.fluid_in(k_10_78), .fluid_out(k_9_39), .air_in(c_10_0));
valve v_10_79 (.fluid_in(k_10_79), .fluid_out(k_9_39), .air_in(c_10_1));
valve v_10_80 (.fluid_in(k_10_80), .fluid_out(k_9_40), .air_in(c_10_0));
valve v_10_81 (.fluid_in(k_10_81), .fluid_out(k_9_40), .air_in(c_10_1));
valve v_10_82 (.fluid_in(k_10_82), .fluid_out(k_9_41), .air_in(c_10_0));
valve v_10_83 (.fluid_in(k_10_83), .fluid_out(k_9_41), .air_in(c_10_1));
valve v_10_84 (.fluid_in(k_10_84), .fluid_out(k_9_42), .air_in(c_10_0));
valve v_10_85 (.fluid_in(k_10_85), .fluid_out(k_9_42), .air_in(c_10_1));
valve v_10_86 (.fluid_in(k_10_86), .fluid_out(k_9_43), .air_in(c_10_0));
valve v_10_87 (.fluid_in(k_10_87), .fluid_out(k_9_43), .air_in(c_10_1));
valve v_10_88 (.fluid_in(k_10_88), .fluid_out(k_9_44), .air_in(c_10_0));
valve v_10_89 (.fluid_in(k_10_89), .fluid_out(k_9_44), .air_in(c_10_1));
valve v_10_90 (.fluid_in(k_10_90), .fluid_out(k_9_45), .air_in(c_10_0));
valve v_10_91 (.fluid_in(k_10_91), .fluid_out(k_9_45), .air_in(c_10_1));
valve v_10_92 (.fluid_in(k_10_92), .fluid_out(k_9_46), .air_in(c_10_0));
valve v_10_93 (.fluid_in(k_10_93), .fluid_out(k_9_46), .air_in(c_10_1));
valve v_10_94 (.fluid_in(k_10_94), .fluid_out(k_9_47), .air_in(c_10_0));
valve v_10_95 (.fluid_in(k_10_95), .fluid_out(k_9_47), .air_in(c_10_1));
valve v_10_96 (.fluid_in(k_10_96), .fluid_out(k_9_48), .air_in(c_10_0));
valve v_10_97 (.fluid_in(k_10_97), .fluid_out(k_9_48), .air_in(c_10_1));
valve v_10_98 (.fluid_in(k_10_98), .fluid_out(k_9_49), .air_in(c_10_0));
valve v_10_99 (.fluid_in(k_10_99), .fluid_out(k_9_49), .air_in(c_10_1));
valve v_10_100 (.fluid_in(k_10_100), .fluid_out(k_9_50), .air_in(c_10_0));
valve v_10_101 (.fluid_in(k_10_101), .fluid_out(k_9_50), .air_in(c_10_1));
valve v_10_102 (.fluid_in(k_10_102), .fluid_out(k_9_51), .air_in(c_10_0));
valve v_10_103 (.fluid_in(k_10_103), .fluid_out(k_9_51), .air_in(c_10_1));
valve v_10_104 (.fluid_in(k_10_104), .fluid_out(k_9_52), .air_in(c_10_0));
valve v_10_105 (.fluid_in(k_10_105), .fluid_out(k_9_52), .air_in(c_10_1));
valve v_10_106 (.fluid_in(k_10_106), .fluid_out(k_9_53), .air_in(c_10_0));
valve v_10_107 (.fluid_in(k_10_107), .fluid_out(k_9_53), .air_in(c_10_1));
valve v_10_108 (.fluid_in(k_10_108), .fluid_out(k_9_54), .air_in(c_10_0));
valve v_10_109 (.fluid_in(k_10_109), .fluid_out(k_9_54), .air_in(c_10_1));
valve v_10_110 (.fluid_in(k_10_110), .fluid_out(k_9_55), .air_in(c_10_0));
valve v_10_111 (.fluid_in(k_10_111), .fluid_out(k_9_55), .air_in(c_10_1));
valve v_10_112 (.fluid_in(k_10_112), .fluid_out(k_9_56), .air_in(c_10_0));
valve v_10_113 (.fluid_in(k_10_113), .fluid_out(k_9_56), .air_in(c_10_1));
valve v_10_114 (.fluid_in(k_10_114), .fluid_out(k_9_57), .air_in(c_10_0));
valve v_10_115 (.fluid_in(k_10_115), .fluid_out(k_9_57), .air_in(c_10_1));
valve v_10_116 (.fluid_in(k_10_116), .fluid_out(k_9_58), .air_in(c_10_0));
valve v_10_117 (.fluid_in(k_10_117), .fluid_out(k_9_58), .air_in(c_10_1));
valve v_10_118 (.fluid_in(k_10_118), .fluid_out(k_9_59), .air_in(c_10_0));
valve v_10_119 (.fluid_in(k_10_119), .fluid_out(k_9_59), .air_in(c_10_1));
valve v_10_120 (.fluid_in(k_10_120), .fluid_out(k_9_60), .air_in(c_10_0));
valve v_10_121 (.fluid_in(k_10_121), .fluid_out(k_9_60), .air_in(c_10_1));
valve v_10_122 (.fluid_in(k_10_122), .fluid_out(k_9_61), .air_in(c_10_0));
valve v_10_123 (.fluid_in(k_10_123), .fluid_out(k_9_61), .air_in(c_10_1));
valve v_10_124 (.fluid_in(k_10_124), .fluid_out(k_9_62), .air_in(c_10_0));
valve v_10_125 (.fluid_in(k_10_125), .fluid_out(k_9_62), .air_in(c_10_1));
valve v_10_126 (.fluid_in(k_10_126), .fluid_out(k_9_63), .air_in(c_10_0));
valve v_10_127 (.fluid_in(k_10_127), .fluid_out(k_9_63), .air_in(c_10_1));
valve v_10_128 (.fluid_in(k_10_128), .fluid_out(k_9_64), .air_in(c_10_0));
valve v_10_129 (.fluid_in(k_10_129), .fluid_out(k_9_64), .air_in(c_10_1));
valve v_10_130 (.fluid_in(k_10_130), .fluid_out(k_9_65), .air_in(c_10_0));
valve v_10_131 (.fluid_in(k_10_131), .fluid_out(k_9_65), .air_in(c_10_1));
valve v_10_132 (.fluid_in(k_10_132), .fluid_out(k_9_66), .air_in(c_10_0));
valve v_10_133 (.fluid_in(k_10_133), .fluid_out(k_9_66), .air_in(c_10_1));
valve v_10_134 (.fluid_in(k_10_134), .fluid_out(k_9_67), .air_in(c_10_0));
valve v_10_135 (.fluid_in(k_10_135), .fluid_out(k_9_67), .air_in(c_10_1));
valve v_10_136 (.fluid_in(k_10_136), .fluid_out(k_9_68), .air_in(c_10_0));
valve v_10_137 (.fluid_in(k_10_137), .fluid_out(k_9_68), .air_in(c_10_1));
valve v_10_138 (.fluid_in(k_10_138), .fluid_out(k_9_69), .air_in(c_10_0));
valve v_10_139 (.fluid_in(k_10_139), .fluid_out(k_9_69), .air_in(c_10_1));
valve v_10_140 (.fluid_in(k_10_140), .fluid_out(k_9_70), .air_in(c_10_0));
valve v_10_141 (.fluid_in(k_10_141), .fluid_out(k_9_70), .air_in(c_10_1));
valve v_10_142 (.fluid_in(k_10_142), .fluid_out(k_9_71), .air_in(c_10_0));
valve v_10_143 (.fluid_in(k_10_143), .fluid_out(k_9_71), .air_in(c_10_1));
valve v_10_144 (.fluid_in(k_10_144), .fluid_out(k_9_72), .air_in(c_10_0));
valve v_10_145 (.fluid_in(k_10_145), .fluid_out(k_9_72), .air_in(c_10_1));
valve v_10_146 (.fluid_in(k_10_146), .fluid_out(k_9_73), .air_in(c_10_0));
valve v_10_147 (.fluid_in(k_10_147), .fluid_out(k_9_73), .air_in(c_10_1));
valve v_10_148 (.fluid_in(k_10_148), .fluid_out(k_9_74), .air_in(c_10_0));
valve v_10_149 (.fluid_in(k_10_149), .fluid_out(k_9_74), .air_in(c_10_1));
valve v_10_150 (.fluid_in(k_10_150), .fluid_out(k_9_75), .air_in(c_10_0));
valve v_10_151 (.fluid_in(k_10_151), .fluid_out(k_9_75), .air_in(c_10_1));
valve v_10_152 (.fluid_in(k_10_152), .fluid_out(k_9_76), .air_in(c_10_0));
valve v_10_153 (.fluid_in(k_10_153), .fluid_out(k_9_76), .air_in(c_10_1));
valve v_10_154 (.fluid_in(k_10_154), .fluid_out(k_9_77), .air_in(c_10_0));
valve v_10_155 (.fluid_in(k_10_155), .fluid_out(k_9_77), .air_in(c_10_1));
valve v_10_156 (.fluid_in(k_10_156), .fluid_out(k_9_78), .air_in(c_10_0));
valve v_10_157 (.fluid_in(k_10_157), .fluid_out(k_9_78), .air_in(c_10_1));
valve v_10_158 (.fluid_in(k_10_158), .fluid_out(k_9_79), .air_in(c_10_0));
valve v_10_159 (.fluid_in(k_10_159), .fluid_out(k_9_79), .air_in(c_10_1));
valve v_10_160 (.fluid_in(k_10_160), .fluid_out(k_9_80), .air_in(c_10_0));
valve v_10_161 (.fluid_in(k_10_161), .fluid_out(k_9_80), .air_in(c_10_1));
valve v_10_162 (.fluid_in(k_10_162), .fluid_out(k_9_81), .air_in(c_10_0));
valve v_10_163 (.fluid_in(k_10_163), .fluid_out(k_9_81), .air_in(c_10_1));
valve v_10_164 (.fluid_in(k_10_164), .fluid_out(k_9_82), .air_in(c_10_0));
valve v_10_165 (.fluid_in(k_10_165), .fluid_out(k_9_82), .air_in(c_10_1));
valve v_10_166 (.fluid_in(k_10_166), .fluid_out(k_9_83), .air_in(c_10_0));
valve v_10_167 (.fluid_in(k_10_167), .fluid_out(k_9_83), .air_in(c_10_1));
valve v_10_168 (.fluid_in(k_10_168), .fluid_out(k_9_84), .air_in(c_10_0));
valve v_10_169 (.fluid_in(k_10_169), .fluid_out(k_9_84), .air_in(c_10_1));
valve v_10_170 (.fluid_in(k_10_170), .fluid_out(k_9_85), .air_in(c_10_0));
valve v_10_171 (.fluid_in(k_10_171), .fluid_out(k_9_85), .air_in(c_10_1));
valve v_10_172 (.fluid_in(k_10_172), .fluid_out(k_9_86), .air_in(c_10_0));
valve v_10_173 (.fluid_in(k_10_173), .fluid_out(k_9_86), .air_in(c_10_1));
valve v_10_174 (.fluid_in(k_10_174), .fluid_out(k_9_87), .air_in(c_10_0));
valve v_10_175 (.fluid_in(k_10_175), .fluid_out(k_9_87), .air_in(c_10_1));
valve v_10_176 (.fluid_in(k_10_176), .fluid_out(k_9_88), .air_in(c_10_0));
valve v_10_177 (.fluid_in(k_10_177), .fluid_out(k_9_88), .air_in(c_10_1));
valve v_10_178 (.fluid_in(k_10_178), .fluid_out(k_9_89), .air_in(c_10_0));
valve v_10_179 (.fluid_in(k_10_179), .fluid_out(k_9_89), .air_in(c_10_1));
valve v_10_180 (.fluid_in(k_10_180), .fluid_out(k_9_90), .air_in(c_10_0));
valve v_10_181 (.fluid_in(k_10_181), .fluid_out(k_9_90), .air_in(c_10_1));
valve v_10_182 (.fluid_in(k_10_182), .fluid_out(k_9_91), .air_in(c_10_0));
valve v_10_183 (.fluid_in(k_10_183), .fluid_out(k_9_91), .air_in(c_10_1));
valve v_10_184 (.fluid_in(k_10_184), .fluid_out(k_9_92), .air_in(c_10_0));
valve v_10_185 (.fluid_in(k_10_185), .fluid_out(k_9_92), .air_in(c_10_1));
valve v_10_186 (.fluid_in(k_10_186), .fluid_out(k_9_93), .air_in(c_10_0));
valve v_10_187 (.fluid_in(k_10_187), .fluid_out(k_9_93), .air_in(c_10_1));
valve v_10_188 (.fluid_in(k_10_188), .fluid_out(k_9_94), .air_in(c_10_0));
valve v_10_189 (.fluid_in(k_10_189), .fluid_out(k_9_94), .air_in(c_10_1));
valve v_10_190 (.fluid_in(k_10_190), .fluid_out(k_9_95), .air_in(c_10_0));
valve v_10_191 (.fluid_in(k_10_191), .fluid_out(k_9_95), .air_in(c_10_1));
valve v_10_192 (.fluid_in(k_10_192), .fluid_out(k_9_96), .air_in(c_10_0));
valve v_10_193 (.fluid_in(k_10_193), .fluid_out(k_9_96), .air_in(c_10_1));
valve v_10_194 (.fluid_in(k_10_194), .fluid_out(k_9_97), .air_in(c_10_0));
valve v_10_195 (.fluid_in(k_10_195), .fluid_out(k_9_97), .air_in(c_10_1));
valve v_10_196 (.fluid_in(k_10_196), .fluid_out(k_9_98), .air_in(c_10_0));
valve v_10_197 (.fluid_in(k_10_197), .fluid_out(k_9_98), .air_in(c_10_1));
valve v_10_198 (.fluid_in(k_10_198), .fluid_out(k_9_99), .air_in(c_10_0));
valve v_10_199 (.fluid_in(k_10_199), .fluid_out(k_9_99), .air_in(c_10_1));
valve v_10_200 (.fluid_in(k_10_200), .fluid_out(k_9_100), .air_in(c_10_0));
valve v_10_201 (.fluid_in(k_10_201), .fluid_out(k_9_100), .air_in(c_10_1));
valve v_10_202 (.fluid_in(k_10_202), .fluid_out(k_9_101), .air_in(c_10_0));
valve v_10_203 (.fluid_in(k_10_203), .fluid_out(k_9_101), .air_in(c_10_1));
valve v_10_204 (.fluid_in(k_10_204), .fluid_out(k_9_102), .air_in(c_10_0));
valve v_10_205 (.fluid_in(k_10_205), .fluid_out(k_9_102), .air_in(c_10_1));
valve v_10_206 (.fluid_in(k_10_206), .fluid_out(k_9_103), .air_in(c_10_0));
valve v_10_207 (.fluid_in(k_10_207), .fluid_out(k_9_103), .air_in(c_10_1));
valve v_10_208 (.fluid_in(k_10_208), .fluid_out(k_9_104), .air_in(c_10_0));
valve v_10_209 (.fluid_in(k_10_209), .fluid_out(k_9_104), .air_in(c_10_1));
valve v_10_210 (.fluid_in(k_10_210), .fluid_out(k_9_105), .air_in(c_10_0));
valve v_10_211 (.fluid_in(k_10_211), .fluid_out(k_9_105), .air_in(c_10_1));
valve v_10_212 (.fluid_in(k_10_212), .fluid_out(k_9_106), .air_in(c_10_0));
valve v_10_213 (.fluid_in(k_10_213), .fluid_out(k_9_106), .air_in(c_10_1));
valve v_10_214 (.fluid_in(k_10_214), .fluid_out(k_9_107), .air_in(c_10_0));
valve v_10_215 (.fluid_in(k_10_215), .fluid_out(k_9_107), .air_in(c_10_1));
valve v_10_216 (.fluid_in(k_10_216), .fluid_out(k_9_108), .air_in(c_10_0));
valve v_10_217 (.fluid_in(k_10_217), .fluid_out(k_9_108), .air_in(c_10_1));
valve v_10_218 (.fluid_in(k_10_218), .fluid_out(k_9_109), .air_in(c_10_0));
valve v_10_219 (.fluid_in(k_10_219), .fluid_out(k_9_109), .air_in(c_10_1));
valve v_10_220 (.fluid_in(k_10_220), .fluid_out(k_9_110), .air_in(c_10_0));
valve v_10_221 (.fluid_in(k_10_221), .fluid_out(k_9_110), .air_in(c_10_1));
valve v_10_222 (.fluid_in(k_10_222), .fluid_out(k_9_111), .air_in(c_10_0));
valve v_10_223 (.fluid_in(k_10_223), .fluid_out(k_9_111), .air_in(c_10_1));
valve v_10_224 (.fluid_in(k_10_224), .fluid_out(k_9_112), .air_in(c_10_0));
valve v_10_225 (.fluid_in(k_10_225), .fluid_out(k_9_112), .air_in(c_10_1));
valve v_10_226 (.fluid_in(k_10_226), .fluid_out(k_9_113), .air_in(c_10_0));
valve v_10_227 (.fluid_in(k_10_227), .fluid_out(k_9_113), .air_in(c_10_1));
valve v_10_228 (.fluid_in(k_10_228), .fluid_out(k_9_114), .air_in(c_10_0));
valve v_10_229 (.fluid_in(k_10_229), .fluid_out(k_9_114), .air_in(c_10_1));
valve v_10_230 (.fluid_in(k_10_230), .fluid_out(k_9_115), .air_in(c_10_0));
valve v_10_231 (.fluid_in(k_10_231), .fluid_out(k_9_115), .air_in(c_10_1));
valve v_10_232 (.fluid_in(k_10_232), .fluid_out(k_9_116), .air_in(c_10_0));
valve v_10_233 (.fluid_in(k_10_233), .fluid_out(k_9_116), .air_in(c_10_1));
valve v_10_234 (.fluid_in(k_10_234), .fluid_out(k_9_117), .air_in(c_10_0));
valve v_10_235 (.fluid_in(k_10_235), .fluid_out(k_9_117), .air_in(c_10_1));
valve v_10_236 (.fluid_in(k_10_236), .fluid_out(k_9_118), .air_in(c_10_0));
valve v_10_237 (.fluid_in(k_10_237), .fluid_out(k_9_118), .air_in(c_10_1));
valve v_10_238 (.fluid_in(k_10_238), .fluid_out(k_9_119), .air_in(c_10_0));
valve v_10_239 (.fluid_in(k_10_239), .fluid_out(k_9_119), .air_in(c_10_1));
valve v_10_240 (.fluid_in(k_10_240), .fluid_out(k_9_120), .air_in(c_10_0));
valve v_10_241 (.fluid_in(k_10_241), .fluid_out(k_9_120), .air_in(c_10_1));
valve v_10_242 (.fluid_in(k_10_242), .fluid_out(k_9_121), .air_in(c_10_0));
valve v_10_243 (.fluid_in(k_10_243), .fluid_out(k_9_121), .air_in(c_10_1));
valve v_10_244 (.fluid_in(k_10_244), .fluid_out(k_9_122), .air_in(c_10_0));
valve v_10_245 (.fluid_in(k_10_245), .fluid_out(k_9_122), .air_in(c_10_1));
valve v_10_246 (.fluid_in(k_10_246), .fluid_out(k_9_123), .air_in(c_10_0));
valve v_10_247 (.fluid_in(k_10_247), .fluid_out(k_9_123), .air_in(c_10_1));
valve v_10_248 (.fluid_in(k_10_248), .fluid_out(k_9_124), .air_in(c_10_0));
valve v_10_249 (.fluid_in(k_10_249), .fluid_out(k_9_124), .air_in(c_10_1));
valve v_10_250 (.fluid_in(k_10_250), .fluid_out(k_9_125), .air_in(c_10_0));
valve v_10_251 (.fluid_in(k_10_251), .fluid_out(k_9_125), .air_in(c_10_1));
valve v_10_252 (.fluid_in(k_10_252), .fluid_out(k_9_126), .air_in(c_10_0));
valve v_10_253 (.fluid_in(k_10_253), .fluid_out(k_9_126), .air_in(c_10_1));
valve v_10_254 (.fluid_in(k_10_254), .fluid_out(k_9_127), .air_in(c_10_0));
valve v_10_255 (.fluid_in(k_10_255), .fluid_out(k_9_127), .air_in(c_10_1));
valve v_10_256 (.fluid_in(k_10_256), .fluid_out(k_9_128), .air_in(c_10_0));
valve v_10_257 (.fluid_in(k_10_257), .fluid_out(k_9_128), .air_in(c_10_1));
valve v_10_258 (.fluid_in(k_10_258), .fluid_out(k_9_129), .air_in(c_10_0));
valve v_10_259 (.fluid_in(k_10_259), .fluid_out(k_9_129), .air_in(c_10_1));
valve v_10_260 (.fluid_in(k_10_260), .fluid_out(k_9_130), .air_in(c_10_0));
valve v_10_261 (.fluid_in(k_10_261), .fluid_out(k_9_130), .air_in(c_10_1));
valve v_10_262 (.fluid_in(k_10_262), .fluid_out(k_9_131), .air_in(c_10_0));
valve v_10_263 (.fluid_in(k_10_263), .fluid_out(k_9_131), .air_in(c_10_1));
valve v_10_264 (.fluid_in(k_10_264), .fluid_out(k_9_132), .air_in(c_10_0));
valve v_10_265 (.fluid_in(k_10_265), .fluid_out(k_9_132), .air_in(c_10_1));
valve v_10_266 (.fluid_in(k_10_266), .fluid_out(k_9_133), .air_in(c_10_0));
valve v_10_267 (.fluid_in(k_10_267), .fluid_out(k_9_133), .air_in(c_10_1));
valve v_10_268 (.fluid_in(k_10_268), .fluid_out(k_9_134), .air_in(c_10_0));
valve v_10_269 (.fluid_in(k_10_269), .fluid_out(k_9_134), .air_in(c_10_1));
valve v_10_270 (.fluid_in(k_10_270), .fluid_out(k_9_135), .air_in(c_10_0));
valve v_10_271 (.fluid_in(k_10_271), .fluid_out(k_9_135), .air_in(c_10_1));
valve v_10_272 (.fluid_in(k_10_272), .fluid_out(k_9_136), .air_in(c_10_0));
valve v_10_273 (.fluid_in(k_10_273), .fluid_out(k_9_136), .air_in(c_10_1));
valve v_10_274 (.fluid_in(k_10_274), .fluid_out(k_9_137), .air_in(c_10_0));
valve v_10_275 (.fluid_in(k_10_275), .fluid_out(k_9_137), .air_in(c_10_1));
valve v_10_276 (.fluid_in(k_10_276), .fluid_out(k_9_138), .air_in(c_10_0));
valve v_10_277 (.fluid_in(k_10_277), .fluid_out(k_9_138), .air_in(c_10_1));
valve v_10_278 (.fluid_in(k_10_278), .fluid_out(k_9_139), .air_in(c_10_0));
valve v_10_279 (.fluid_in(k_10_279), .fluid_out(k_9_139), .air_in(c_10_1));
valve v_10_280 (.fluid_in(k_10_280), .fluid_out(k_9_140), .air_in(c_10_0));
valve v_10_281 (.fluid_in(k_10_281), .fluid_out(k_9_140), .air_in(c_10_1));
valve v_10_282 (.fluid_in(k_10_282), .fluid_out(k_9_141), .air_in(c_10_0));
valve v_10_283 (.fluid_in(k_10_283), .fluid_out(k_9_141), .air_in(c_10_1));
valve v_10_284 (.fluid_in(k_10_284), .fluid_out(k_9_142), .air_in(c_10_0));
valve v_10_285 (.fluid_in(k_10_285), .fluid_out(k_9_142), .air_in(c_10_1));
valve v_10_286 (.fluid_in(k_10_286), .fluid_out(k_9_143), .air_in(c_10_0));
valve v_10_287 (.fluid_in(k_10_287), .fluid_out(k_9_143), .air_in(c_10_1));
valve v_10_288 (.fluid_in(k_10_288), .fluid_out(k_9_144), .air_in(c_10_0));
valve v_10_289 (.fluid_in(k_10_289), .fluid_out(k_9_144), .air_in(c_10_1));
valve v_10_290 (.fluid_in(k_10_290), .fluid_out(k_9_145), .air_in(c_10_0));
valve v_10_291 (.fluid_in(k_10_291), .fluid_out(k_9_145), .air_in(c_10_1));
valve v_10_292 (.fluid_in(k_10_292), .fluid_out(k_9_146), .air_in(c_10_0));
valve v_10_293 (.fluid_in(k_10_293), .fluid_out(k_9_146), .air_in(c_10_1));
valve v_10_294 (.fluid_in(k_10_294), .fluid_out(k_9_147), .air_in(c_10_0));
valve v_10_295 (.fluid_in(k_10_295), .fluid_out(k_9_147), .air_in(c_10_1));
valve v_10_296 (.fluid_in(k_10_296), .fluid_out(k_9_148), .air_in(c_10_0));
valve v_10_297 (.fluid_in(k_10_297), .fluid_out(k_9_148), .air_in(c_10_1));
valve v_10_298 (.fluid_in(k_10_298), .fluid_out(k_9_149), .air_in(c_10_0));
valve v_10_299 (.fluid_in(k_10_299), .fluid_out(k_9_149), .air_in(c_10_1));
valve v_10_300 (.fluid_in(k_10_300), .fluid_out(k_9_150), .air_in(c_10_0));
valve v_10_301 (.fluid_in(k_10_301), .fluid_out(k_9_150), .air_in(c_10_1));
valve v_10_302 (.fluid_in(k_10_302), .fluid_out(k_9_151), .air_in(c_10_0));
valve v_10_303 (.fluid_in(k_10_303), .fluid_out(k_9_151), .air_in(c_10_1));
valve v_10_304 (.fluid_in(k_10_304), .fluid_out(k_9_152), .air_in(c_10_0));
valve v_10_305 (.fluid_in(k_10_305), .fluid_out(k_9_152), .air_in(c_10_1));
valve v_10_306 (.fluid_in(k_10_306), .fluid_out(k_9_153), .air_in(c_10_0));
valve v_10_307 (.fluid_in(k_10_307), .fluid_out(k_9_153), .air_in(c_10_1));
valve v_10_308 (.fluid_in(k_10_308), .fluid_out(k_9_154), .air_in(c_10_0));
valve v_10_309 (.fluid_in(k_10_309), .fluid_out(k_9_154), .air_in(c_10_1));
valve v_10_310 (.fluid_in(k_10_310), .fluid_out(k_9_155), .air_in(c_10_0));
valve v_10_311 (.fluid_in(k_10_311), .fluid_out(k_9_155), .air_in(c_10_1));
valve v_10_312 (.fluid_in(k_10_312), .fluid_out(k_9_156), .air_in(c_10_0));
valve v_10_313 (.fluid_in(k_10_313), .fluid_out(k_9_156), .air_in(c_10_1));
valve v_10_314 (.fluid_in(k_10_314), .fluid_out(k_9_157), .air_in(c_10_0));
valve v_10_315 (.fluid_in(k_10_315), .fluid_out(k_9_157), .air_in(c_10_1));
valve v_10_316 (.fluid_in(k_10_316), .fluid_out(k_9_158), .air_in(c_10_0));
valve v_10_317 (.fluid_in(k_10_317), .fluid_out(k_9_158), .air_in(c_10_1));
valve v_10_318 (.fluid_in(k_10_318), .fluid_out(k_9_159), .air_in(c_10_0));
valve v_10_319 (.fluid_in(k_10_319), .fluid_out(k_9_159), .air_in(c_10_1));
valve v_10_320 (.fluid_in(k_10_320), .fluid_out(k_9_160), .air_in(c_10_0));
valve v_10_321 (.fluid_in(k_10_321), .fluid_out(k_9_160), .air_in(c_10_1));
valve v_10_322 (.fluid_in(k_10_322), .fluid_out(k_9_161), .air_in(c_10_0));
valve v_10_323 (.fluid_in(k_10_323), .fluid_out(k_9_161), .air_in(c_10_1));
valve v_10_324 (.fluid_in(k_10_324), .fluid_out(k_9_162), .air_in(c_10_0));
valve v_10_325 (.fluid_in(k_10_325), .fluid_out(k_9_162), .air_in(c_10_1));
valve v_10_326 (.fluid_in(k_10_326), .fluid_out(k_9_163), .air_in(c_10_0));
valve v_10_327 (.fluid_in(k_10_327), .fluid_out(k_9_163), .air_in(c_10_1));
valve v_10_328 (.fluid_in(k_10_328), .fluid_out(k_9_164), .air_in(c_10_0));
valve v_10_329 (.fluid_in(k_10_329), .fluid_out(k_9_164), .air_in(c_10_1));
valve v_10_330 (.fluid_in(k_10_330), .fluid_out(k_9_165), .air_in(c_10_0));
valve v_10_331 (.fluid_in(k_10_331), .fluid_out(k_9_165), .air_in(c_10_1));
valve v_10_332 (.fluid_in(k_10_332), .fluid_out(k_9_166), .air_in(c_10_0));
valve v_10_333 (.fluid_in(k_10_333), .fluid_out(k_9_166), .air_in(c_10_1));
valve v_10_334 (.fluid_in(k_10_334), .fluid_out(k_9_167), .air_in(c_10_0));
valve v_10_335 (.fluid_in(k_10_335), .fluid_out(k_9_167), .air_in(c_10_1));
valve v_10_336 (.fluid_in(k_10_336), .fluid_out(k_9_168), .air_in(c_10_0));
valve v_10_337 (.fluid_in(k_10_337), .fluid_out(k_9_168), .air_in(c_10_1));
valve v_10_338 (.fluid_in(k_10_338), .fluid_out(k_9_169), .air_in(c_10_0));
valve v_10_339 (.fluid_in(k_10_339), .fluid_out(k_9_169), .air_in(c_10_1));
valve v_10_340 (.fluid_in(k_10_340), .fluid_out(k_9_170), .air_in(c_10_0));
valve v_10_341 (.fluid_in(k_10_341), .fluid_out(k_9_170), .air_in(c_10_1));
valve v_10_342 (.fluid_in(k_10_342), .fluid_out(k_9_171), .air_in(c_10_0));
valve v_10_343 (.fluid_in(k_10_343), .fluid_out(k_9_171), .air_in(c_10_1));
valve v_10_344 (.fluid_in(k_10_344), .fluid_out(k_9_172), .air_in(c_10_0));
valve v_10_345 (.fluid_in(k_10_345), .fluid_out(k_9_172), .air_in(c_10_1));
valve v_10_346 (.fluid_in(k_10_346), .fluid_out(k_9_173), .air_in(c_10_0));
valve v_10_347 (.fluid_in(k_10_347), .fluid_out(k_9_173), .air_in(c_10_1));
valve v_10_348 (.fluid_in(k_10_348), .fluid_out(k_9_174), .air_in(c_10_0));
valve v_10_349 (.fluid_in(k_10_349), .fluid_out(k_9_174), .air_in(c_10_1));
valve v_10_350 (.fluid_in(k_10_350), .fluid_out(k_9_175), .air_in(c_10_0));
valve v_10_351 (.fluid_in(k_10_351), .fluid_out(k_9_175), .air_in(c_10_1));
valve v_10_352 (.fluid_in(k_10_352), .fluid_out(k_9_176), .air_in(c_10_0));
valve v_10_353 (.fluid_in(k_10_353), .fluid_out(k_9_176), .air_in(c_10_1));
valve v_10_354 (.fluid_in(k_10_354), .fluid_out(k_9_177), .air_in(c_10_0));
valve v_10_355 (.fluid_in(k_10_355), .fluid_out(k_9_177), .air_in(c_10_1));
valve v_10_356 (.fluid_in(k_10_356), .fluid_out(k_9_178), .air_in(c_10_0));
valve v_10_357 (.fluid_in(k_10_357), .fluid_out(k_9_178), .air_in(c_10_1));
valve v_10_358 (.fluid_in(k_10_358), .fluid_out(k_9_179), .air_in(c_10_0));
valve v_10_359 (.fluid_in(k_10_359), .fluid_out(k_9_179), .air_in(c_10_1));
valve v_10_360 (.fluid_in(k_10_360), .fluid_out(k_9_180), .air_in(c_10_0));
valve v_10_361 (.fluid_in(k_10_361), .fluid_out(k_9_180), .air_in(c_10_1));
valve v_10_362 (.fluid_in(k_10_362), .fluid_out(k_9_181), .air_in(c_10_0));
valve v_10_363 (.fluid_in(k_10_363), .fluid_out(k_9_181), .air_in(c_10_1));
valve v_10_364 (.fluid_in(k_10_364), .fluid_out(k_9_182), .air_in(c_10_0));
valve v_10_365 (.fluid_in(k_10_365), .fluid_out(k_9_182), .air_in(c_10_1));
valve v_10_366 (.fluid_in(k_10_366), .fluid_out(k_9_183), .air_in(c_10_0));
valve v_10_367 (.fluid_in(k_10_367), .fluid_out(k_9_183), .air_in(c_10_1));
valve v_10_368 (.fluid_in(k_10_368), .fluid_out(k_9_184), .air_in(c_10_0));
valve v_10_369 (.fluid_in(k_10_369), .fluid_out(k_9_184), .air_in(c_10_1));
valve v_10_370 (.fluid_in(k_10_370), .fluid_out(k_9_185), .air_in(c_10_0));
valve v_10_371 (.fluid_in(k_10_371), .fluid_out(k_9_185), .air_in(c_10_1));
valve v_10_372 (.fluid_in(k_10_372), .fluid_out(k_9_186), .air_in(c_10_0));
valve v_10_373 (.fluid_in(k_10_373), .fluid_out(k_9_186), .air_in(c_10_1));
valve v_10_374 (.fluid_in(k_10_374), .fluid_out(k_9_187), .air_in(c_10_0));
valve v_10_375 (.fluid_in(k_10_375), .fluid_out(k_9_187), .air_in(c_10_1));
valve v_10_376 (.fluid_in(k_10_376), .fluid_out(k_9_188), .air_in(c_10_0));
valve v_10_377 (.fluid_in(k_10_377), .fluid_out(k_9_188), .air_in(c_10_1));
valve v_10_378 (.fluid_in(k_10_378), .fluid_out(k_9_189), .air_in(c_10_0));
valve v_10_379 (.fluid_in(k_10_379), .fluid_out(k_9_189), .air_in(c_10_1));
valve v_10_380 (.fluid_in(k_10_380), .fluid_out(k_9_190), .air_in(c_10_0));
valve v_10_381 (.fluid_in(k_10_381), .fluid_out(k_9_190), .air_in(c_10_1));
valve v_10_382 (.fluid_in(k_10_382), .fluid_out(k_9_191), .air_in(c_10_0));
valve v_10_383 (.fluid_in(k_10_383), .fluid_out(k_9_191), .air_in(c_10_1));
valve v_10_384 (.fluid_in(k_10_384), .fluid_out(k_9_192), .air_in(c_10_0));
valve v_10_385 (.fluid_in(k_10_385), .fluid_out(k_9_192), .air_in(c_10_1));
valve v_10_386 (.fluid_in(k_10_386), .fluid_out(k_9_193), .air_in(c_10_0));
valve v_10_387 (.fluid_in(k_10_387), .fluid_out(k_9_193), .air_in(c_10_1));
valve v_10_388 (.fluid_in(k_10_388), .fluid_out(k_9_194), .air_in(c_10_0));
valve v_10_389 (.fluid_in(k_10_389), .fluid_out(k_9_194), .air_in(c_10_1));
valve v_10_390 (.fluid_in(k_10_390), .fluid_out(k_9_195), .air_in(c_10_0));
valve v_10_391 (.fluid_in(k_10_391), .fluid_out(k_9_195), .air_in(c_10_1));
valve v_10_392 (.fluid_in(k_10_392), .fluid_out(k_9_196), .air_in(c_10_0));
valve v_10_393 (.fluid_in(k_10_393), .fluid_out(k_9_196), .air_in(c_10_1));
valve v_10_394 (.fluid_in(k_10_394), .fluid_out(k_9_197), .air_in(c_10_0));
valve v_10_395 (.fluid_in(k_10_395), .fluid_out(k_9_197), .air_in(c_10_1));
valve v_10_396 (.fluid_in(k_10_396), .fluid_out(k_9_198), .air_in(c_10_0));
valve v_10_397 (.fluid_in(k_10_397), .fluid_out(k_9_198), .air_in(c_10_1));
valve v_10_398 (.fluid_in(k_10_398), .fluid_out(k_9_199), .air_in(c_10_0));
valve v_10_399 (.fluid_in(k_10_399), .fluid_out(k_9_199), .air_in(c_10_1));
valve v_10_400 (.fluid_in(k_10_400), .fluid_out(k_9_200), .air_in(c_10_0));
valve v_10_401 (.fluid_in(k_10_401), .fluid_out(k_9_200), .air_in(c_10_1));
valve v_10_402 (.fluid_in(k_10_402), .fluid_out(k_9_201), .air_in(c_10_0));
valve v_10_403 (.fluid_in(k_10_403), .fluid_out(k_9_201), .air_in(c_10_1));
valve v_10_404 (.fluid_in(k_10_404), .fluid_out(k_9_202), .air_in(c_10_0));
valve v_10_405 (.fluid_in(k_10_405), .fluid_out(k_9_202), .air_in(c_10_1));
valve v_10_406 (.fluid_in(k_10_406), .fluid_out(k_9_203), .air_in(c_10_0));
valve v_10_407 (.fluid_in(k_10_407), .fluid_out(k_9_203), .air_in(c_10_1));
valve v_10_408 (.fluid_in(k_10_408), .fluid_out(k_9_204), .air_in(c_10_0));
valve v_10_409 (.fluid_in(k_10_409), .fluid_out(k_9_204), .air_in(c_10_1));
valve v_10_410 (.fluid_in(k_10_410), .fluid_out(k_9_205), .air_in(c_10_0));
valve v_10_411 (.fluid_in(k_10_411), .fluid_out(k_9_205), .air_in(c_10_1));
valve v_10_412 (.fluid_in(k_10_412), .fluid_out(k_9_206), .air_in(c_10_0));
valve v_10_413 (.fluid_in(k_10_413), .fluid_out(k_9_206), .air_in(c_10_1));
valve v_10_414 (.fluid_in(k_10_414), .fluid_out(k_9_207), .air_in(c_10_0));
valve v_10_415 (.fluid_in(k_10_415), .fluid_out(k_9_207), .air_in(c_10_1));
valve v_10_416 (.fluid_in(k_10_416), .fluid_out(k_9_208), .air_in(c_10_0));
valve v_10_417 (.fluid_in(k_10_417), .fluid_out(k_9_208), .air_in(c_10_1));
valve v_10_418 (.fluid_in(k_10_418), .fluid_out(k_9_209), .air_in(c_10_0));
valve v_10_419 (.fluid_in(k_10_419), .fluid_out(k_9_209), .air_in(c_10_1));
valve v_10_420 (.fluid_in(k_10_420), .fluid_out(k_9_210), .air_in(c_10_0));
valve v_10_421 (.fluid_in(k_10_421), .fluid_out(k_9_210), .air_in(c_10_1));
valve v_10_422 (.fluid_in(k_10_422), .fluid_out(k_9_211), .air_in(c_10_0));
valve v_10_423 (.fluid_in(k_10_423), .fluid_out(k_9_211), .air_in(c_10_1));
valve v_10_424 (.fluid_in(k_10_424), .fluid_out(k_9_212), .air_in(c_10_0));
valve v_10_425 (.fluid_in(k_10_425), .fluid_out(k_9_212), .air_in(c_10_1));
valve v_10_426 (.fluid_in(k_10_426), .fluid_out(k_9_213), .air_in(c_10_0));
valve v_10_427 (.fluid_in(k_10_427), .fluid_out(k_9_213), .air_in(c_10_1));
valve v_10_428 (.fluid_in(k_10_428), .fluid_out(k_9_214), .air_in(c_10_0));
valve v_10_429 (.fluid_in(k_10_429), .fluid_out(k_9_214), .air_in(c_10_1));
valve v_10_430 (.fluid_in(k_10_430), .fluid_out(k_9_215), .air_in(c_10_0));
valve v_10_431 (.fluid_in(k_10_431), .fluid_out(k_9_215), .air_in(c_10_1));
valve v_10_432 (.fluid_in(k_10_432), .fluid_out(k_9_216), .air_in(c_10_0));
valve v_10_433 (.fluid_in(k_10_433), .fluid_out(k_9_216), .air_in(c_10_1));
valve v_10_434 (.fluid_in(k_10_434), .fluid_out(k_9_217), .air_in(c_10_0));
valve v_10_435 (.fluid_in(k_10_435), .fluid_out(k_9_217), .air_in(c_10_1));
valve v_10_436 (.fluid_in(k_10_436), .fluid_out(k_9_218), .air_in(c_10_0));
valve v_10_437 (.fluid_in(k_10_437), .fluid_out(k_9_218), .air_in(c_10_1));
valve v_10_438 (.fluid_in(k_10_438), .fluid_out(k_9_219), .air_in(c_10_0));
valve v_10_439 (.fluid_in(k_10_439), .fluid_out(k_9_219), .air_in(c_10_1));
valve v_10_440 (.fluid_in(k_10_440), .fluid_out(k_9_220), .air_in(c_10_0));
valve v_10_441 (.fluid_in(k_10_441), .fluid_out(k_9_220), .air_in(c_10_1));
valve v_10_442 (.fluid_in(k_10_442), .fluid_out(k_9_221), .air_in(c_10_0));
valve v_10_443 (.fluid_in(k_10_443), .fluid_out(k_9_221), .air_in(c_10_1));
valve v_10_444 (.fluid_in(k_10_444), .fluid_out(k_9_222), .air_in(c_10_0));
valve v_10_445 (.fluid_in(k_10_445), .fluid_out(k_9_222), .air_in(c_10_1));
valve v_10_446 (.fluid_in(k_10_446), .fluid_out(k_9_223), .air_in(c_10_0));
valve v_10_447 (.fluid_in(k_10_447), .fluid_out(k_9_223), .air_in(c_10_1));
valve v_10_448 (.fluid_in(k_10_448), .fluid_out(k_9_224), .air_in(c_10_0));
valve v_10_449 (.fluid_in(k_10_449), .fluid_out(k_9_224), .air_in(c_10_1));
valve v_10_450 (.fluid_in(k_10_450), .fluid_out(k_9_225), .air_in(c_10_0));
valve v_10_451 (.fluid_in(k_10_451), .fluid_out(k_9_225), .air_in(c_10_1));
valve v_10_452 (.fluid_in(k_10_452), .fluid_out(k_9_226), .air_in(c_10_0));
valve v_10_453 (.fluid_in(k_10_453), .fluid_out(k_9_226), .air_in(c_10_1));
valve v_10_454 (.fluid_in(k_10_454), .fluid_out(k_9_227), .air_in(c_10_0));
valve v_10_455 (.fluid_in(k_10_455), .fluid_out(k_9_227), .air_in(c_10_1));
valve v_10_456 (.fluid_in(k_10_456), .fluid_out(k_9_228), .air_in(c_10_0));
valve v_10_457 (.fluid_in(k_10_457), .fluid_out(k_9_228), .air_in(c_10_1));
valve v_10_458 (.fluid_in(k_10_458), .fluid_out(k_9_229), .air_in(c_10_0));
valve v_10_459 (.fluid_in(k_10_459), .fluid_out(k_9_229), .air_in(c_10_1));
valve v_10_460 (.fluid_in(k_10_460), .fluid_out(k_9_230), .air_in(c_10_0));
valve v_10_461 (.fluid_in(k_10_461), .fluid_out(k_9_230), .air_in(c_10_1));
valve v_10_462 (.fluid_in(k_10_462), .fluid_out(k_9_231), .air_in(c_10_0));
valve v_10_463 (.fluid_in(k_10_463), .fluid_out(k_9_231), .air_in(c_10_1));
valve v_10_464 (.fluid_in(k_10_464), .fluid_out(k_9_232), .air_in(c_10_0));
valve v_10_465 (.fluid_in(k_10_465), .fluid_out(k_9_232), .air_in(c_10_1));
valve v_10_466 (.fluid_in(k_10_466), .fluid_out(k_9_233), .air_in(c_10_0));
valve v_10_467 (.fluid_in(k_10_467), .fluid_out(k_9_233), .air_in(c_10_1));
valve v_10_468 (.fluid_in(k_10_468), .fluid_out(k_9_234), .air_in(c_10_0));
valve v_10_469 (.fluid_in(k_10_469), .fluid_out(k_9_234), .air_in(c_10_1));
valve v_10_470 (.fluid_in(k_10_470), .fluid_out(k_9_235), .air_in(c_10_0));
valve v_10_471 (.fluid_in(k_10_471), .fluid_out(k_9_235), .air_in(c_10_1));
valve v_10_472 (.fluid_in(k_10_472), .fluid_out(k_9_236), .air_in(c_10_0));
valve v_10_473 (.fluid_in(k_10_473), .fluid_out(k_9_236), .air_in(c_10_1));
valve v_10_474 (.fluid_in(k_10_474), .fluid_out(k_9_237), .air_in(c_10_0));
valve v_10_475 (.fluid_in(k_10_475), .fluid_out(k_9_237), .air_in(c_10_1));
valve v_10_476 (.fluid_in(k_10_476), .fluid_out(k_9_238), .air_in(c_10_0));
valve v_10_477 (.fluid_in(k_10_477), .fluid_out(k_9_238), .air_in(c_10_1));
valve v_10_478 (.fluid_in(k_10_478), .fluid_out(k_9_239), .air_in(c_10_0));
valve v_10_479 (.fluid_in(k_10_479), .fluid_out(k_9_239), .air_in(c_10_1));
valve v_10_480 (.fluid_in(k_10_480), .fluid_out(k_9_240), .air_in(c_10_0));
valve v_10_481 (.fluid_in(k_10_481), .fluid_out(k_9_240), .air_in(c_10_1));
valve v_10_482 (.fluid_in(k_10_482), .fluid_out(k_9_241), .air_in(c_10_0));
valve v_10_483 (.fluid_in(k_10_483), .fluid_out(k_9_241), .air_in(c_10_1));
valve v_10_484 (.fluid_in(k_10_484), .fluid_out(k_9_242), .air_in(c_10_0));
valve v_10_485 (.fluid_in(k_10_485), .fluid_out(k_9_242), .air_in(c_10_1));
valve v_10_486 (.fluid_in(k_10_486), .fluid_out(k_9_243), .air_in(c_10_0));
valve v_10_487 (.fluid_in(k_10_487), .fluid_out(k_9_243), .air_in(c_10_1));
valve v_10_488 (.fluid_in(k_10_488), .fluid_out(k_9_244), .air_in(c_10_0));
valve v_10_489 (.fluid_in(k_10_489), .fluid_out(k_9_244), .air_in(c_10_1));
valve v_10_490 (.fluid_in(k_10_490), .fluid_out(k_9_245), .air_in(c_10_0));
valve v_10_491 (.fluid_in(k_10_491), .fluid_out(k_9_245), .air_in(c_10_1));
valve v_10_492 (.fluid_in(k_10_492), .fluid_out(k_9_246), .air_in(c_10_0));
valve v_10_493 (.fluid_in(k_10_493), .fluid_out(k_9_246), .air_in(c_10_1));
valve v_10_494 (.fluid_in(k_10_494), .fluid_out(k_9_247), .air_in(c_10_0));
valve v_10_495 (.fluid_in(k_10_495), .fluid_out(k_9_247), .air_in(c_10_1));
valve v_10_496 (.fluid_in(k_10_496), .fluid_out(k_9_248), .air_in(c_10_0));
valve v_10_497 (.fluid_in(k_10_497), .fluid_out(k_9_248), .air_in(c_10_1));
valve v_10_498 (.fluid_in(k_10_498), .fluid_out(k_9_249), .air_in(c_10_0));
valve v_10_499 (.fluid_in(k_10_499), .fluid_out(k_9_249), .air_in(c_10_1));
valve v_10_500 (.fluid_in(k_10_500), .fluid_out(k_9_250), .air_in(c_10_0));
valve v_10_501 (.fluid_in(k_10_501), .fluid_out(k_9_250), .air_in(c_10_1));
valve v_10_502 (.fluid_in(k_10_502), .fluid_out(k_9_251), .air_in(c_10_0));
valve v_10_503 (.fluid_in(k_10_503), .fluid_out(k_9_251), .air_in(c_10_1));
valve v_10_504 (.fluid_in(k_10_504), .fluid_out(k_9_252), .air_in(c_10_0));
valve v_10_505 (.fluid_in(k_10_505), .fluid_out(k_9_252), .air_in(c_10_1));
valve v_10_506 (.fluid_in(k_10_506), .fluid_out(k_9_253), .air_in(c_10_0));
valve v_10_507 (.fluid_in(k_10_507), .fluid_out(k_9_253), .air_in(c_10_1));
valve v_10_508 (.fluid_in(k_10_508), .fluid_out(k_9_254), .air_in(c_10_0));
valve v_10_509 (.fluid_in(k_10_509), .fluid_out(k_9_254), .air_in(c_10_1));
valve v_10_510 (.fluid_in(k_10_510), .fluid_out(k_9_255), .air_in(c_10_0));
valve v_10_511 (.fluid_in(k_10_511), .fluid_out(k_9_255), .air_in(c_10_1));
valve v_10_512 (.fluid_in(k_10_512), .fluid_out(k_9_256), .air_in(c_10_0));
valve v_10_513 (.fluid_in(k_10_513), .fluid_out(k_9_256), .air_in(c_10_1));
valve v_10_514 (.fluid_in(k_10_514), .fluid_out(k_9_257), .air_in(c_10_0));
valve v_10_515 (.fluid_in(k_10_515), .fluid_out(k_9_257), .air_in(c_10_1));
valve v_10_516 (.fluid_in(k_10_516), .fluid_out(k_9_258), .air_in(c_10_0));
valve v_10_517 (.fluid_in(k_10_517), .fluid_out(k_9_258), .air_in(c_10_1));
valve v_10_518 (.fluid_in(k_10_518), .fluid_out(k_9_259), .air_in(c_10_0));
valve v_10_519 (.fluid_in(k_10_519), .fluid_out(k_9_259), .air_in(c_10_1));
valve v_10_520 (.fluid_in(k_10_520), .fluid_out(k_9_260), .air_in(c_10_0));
valve v_10_521 (.fluid_in(k_10_521), .fluid_out(k_9_260), .air_in(c_10_1));
valve v_10_522 (.fluid_in(k_10_522), .fluid_out(k_9_261), .air_in(c_10_0));
valve v_10_523 (.fluid_in(k_10_523), .fluid_out(k_9_261), .air_in(c_10_1));
valve v_10_524 (.fluid_in(k_10_524), .fluid_out(k_9_262), .air_in(c_10_0));
valve v_10_525 (.fluid_in(k_10_525), .fluid_out(k_9_262), .air_in(c_10_1));
valve v_10_526 (.fluid_in(k_10_526), .fluid_out(k_9_263), .air_in(c_10_0));
valve v_10_527 (.fluid_in(k_10_527), .fluid_out(k_9_263), .air_in(c_10_1));
valve v_10_528 (.fluid_in(k_10_528), .fluid_out(k_9_264), .air_in(c_10_0));
valve v_10_529 (.fluid_in(k_10_529), .fluid_out(k_9_264), .air_in(c_10_1));
valve v_10_530 (.fluid_in(k_10_530), .fluid_out(k_9_265), .air_in(c_10_0));
valve v_10_531 (.fluid_in(k_10_531), .fluid_out(k_9_265), .air_in(c_10_1));
valve v_10_532 (.fluid_in(k_10_532), .fluid_out(k_9_266), .air_in(c_10_0));
valve v_10_533 (.fluid_in(k_10_533), .fluid_out(k_9_266), .air_in(c_10_1));
valve v_10_534 (.fluid_in(k_10_534), .fluid_out(k_9_267), .air_in(c_10_0));
valve v_10_535 (.fluid_in(k_10_535), .fluid_out(k_9_267), .air_in(c_10_1));
valve v_10_536 (.fluid_in(k_10_536), .fluid_out(k_9_268), .air_in(c_10_0));
valve v_10_537 (.fluid_in(k_10_537), .fluid_out(k_9_268), .air_in(c_10_1));
valve v_10_538 (.fluid_in(k_10_538), .fluid_out(k_9_269), .air_in(c_10_0));
valve v_10_539 (.fluid_in(k_10_539), .fluid_out(k_9_269), .air_in(c_10_1));
valve v_10_540 (.fluid_in(k_10_540), .fluid_out(k_9_270), .air_in(c_10_0));
valve v_10_541 (.fluid_in(k_10_541), .fluid_out(k_9_270), .air_in(c_10_1));
valve v_10_542 (.fluid_in(k_10_542), .fluid_out(k_9_271), .air_in(c_10_0));
valve v_10_543 (.fluid_in(k_10_543), .fluid_out(k_9_271), .air_in(c_10_1));
valve v_10_544 (.fluid_in(k_10_544), .fluid_out(k_9_272), .air_in(c_10_0));
valve v_10_545 (.fluid_in(k_10_545), .fluid_out(k_9_272), .air_in(c_10_1));
valve v_10_546 (.fluid_in(k_10_546), .fluid_out(k_9_273), .air_in(c_10_0));
valve v_10_547 (.fluid_in(k_10_547), .fluid_out(k_9_273), .air_in(c_10_1));
valve v_10_548 (.fluid_in(k_10_548), .fluid_out(k_9_274), .air_in(c_10_0));
valve v_10_549 (.fluid_in(k_10_549), .fluid_out(k_9_274), .air_in(c_10_1));
valve v_10_550 (.fluid_in(k_10_550), .fluid_out(k_9_275), .air_in(c_10_0));
valve v_10_551 (.fluid_in(k_10_551), .fluid_out(k_9_275), .air_in(c_10_1));
valve v_10_552 (.fluid_in(k_10_552), .fluid_out(k_9_276), .air_in(c_10_0));
valve v_10_553 (.fluid_in(k_10_553), .fluid_out(k_9_276), .air_in(c_10_1));
valve v_10_554 (.fluid_in(k_10_554), .fluid_out(k_9_277), .air_in(c_10_0));
valve v_10_555 (.fluid_in(k_10_555), .fluid_out(k_9_277), .air_in(c_10_1));
valve v_10_556 (.fluid_in(k_10_556), .fluid_out(k_9_278), .air_in(c_10_0));
valve v_10_557 (.fluid_in(k_10_557), .fluid_out(k_9_278), .air_in(c_10_1));
valve v_10_558 (.fluid_in(k_10_558), .fluid_out(k_9_279), .air_in(c_10_0));
valve v_10_559 (.fluid_in(k_10_559), .fluid_out(k_9_279), .air_in(c_10_1));
valve v_10_560 (.fluid_in(k_10_560), .fluid_out(k_9_280), .air_in(c_10_0));
valve v_10_561 (.fluid_in(k_10_561), .fluid_out(k_9_280), .air_in(c_10_1));
valve v_10_562 (.fluid_in(k_10_562), .fluid_out(k_9_281), .air_in(c_10_0));
valve v_10_563 (.fluid_in(k_10_563), .fluid_out(k_9_281), .air_in(c_10_1));
valve v_10_564 (.fluid_in(k_10_564), .fluid_out(k_9_282), .air_in(c_10_0));
valve v_10_565 (.fluid_in(k_10_565), .fluid_out(k_9_282), .air_in(c_10_1));
valve v_10_566 (.fluid_in(k_10_566), .fluid_out(k_9_283), .air_in(c_10_0));
valve v_10_567 (.fluid_in(k_10_567), .fluid_out(k_9_283), .air_in(c_10_1));
valve v_10_568 (.fluid_in(k_10_568), .fluid_out(k_9_284), .air_in(c_10_0));
valve v_10_569 (.fluid_in(k_10_569), .fluid_out(k_9_284), .air_in(c_10_1));
valve v_10_570 (.fluid_in(k_10_570), .fluid_out(k_9_285), .air_in(c_10_0));
valve v_10_571 (.fluid_in(k_10_571), .fluid_out(k_9_285), .air_in(c_10_1));
valve v_10_572 (.fluid_in(k_10_572), .fluid_out(k_9_286), .air_in(c_10_0));
valve v_10_573 (.fluid_in(k_10_573), .fluid_out(k_9_286), .air_in(c_10_1));
valve v_10_574 (.fluid_in(k_10_574), .fluid_out(k_9_287), .air_in(c_10_0));
valve v_10_575 (.fluid_in(k_10_575), .fluid_out(k_9_287), .air_in(c_10_1));
valve v_10_576 (.fluid_in(k_10_576), .fluid_out(k_9_288), .air_in(c_10_0));
valve v_10_577 (.fluid_in(k_10_577), .fluid_out(k_9_288), .air_in(c_10_1));
valve v_10_578 (.fluid_in(k_10_578), .fluid_out(k_9_289), .air_in(c_10_0));
valve v_10_579 (.fluid_in(k_10_579), .fluid_out(k_9_289), .air_in(c_10_1));
valve v_10_580 (.fluid_in(k_10_580), .fluid_out(k_9_290), .air_in(c_10_0));
valve v_10_581 (.fluid_in(k_10_581), .fluid_out(k_9_290), .air_in(c_10_1));
valve v_10_582 (.fluid_in(k_10_582), .fluid_out(k_9_291), .air_in(c_10_0));
valve v_10_583 (.fluid_in(k_10_583), .fluid_out(k_9_291), .air_in(c_10_1));
valve v_10_584 (.fluid_in(k_10_584), .fluid_out(k_9_292), .air_in(c_10_0));
valve v_10_585 (.fluid_in(k_10_585), .fluid_out(k_9_292), .air_in(c_10_1));
valve v_10_586 (.fluid_in(k_10_586), .fluid_out(k_9_293), .air_in(c_10_0));
valve v_10_587 (.fluid_in(k_10_587), .fluid_out(k_9_293), .air_in(c_10_1));
valve v_10_588 (.fluid_in(k_10_588), .fluid_out(k_9_294), .air_in(c_10_0));
valve v_10_589 (.fluid_in(k_10_589), .fluid_out(k_9_294), .air_in(c_10_1));
valve v_10_590 (.fluid_in(k_10_590), .fluid_out(k_9_295), .air_in(c_10_0));
valve v_10_591 (.fluid_in(k_10_591), .fluid_out(k_9_295), .air_in(c_10_1));
valve v_10_592 (.fluid_in(k_10_592), .fluid_out(k_9_296), .air_in(c_10_0));
valve v_10_593 (.fluid_in(k_10_593), .fluid_out(k_9_296), .air_in(c_10_1));
valve v_10_594 (.fluid_in(k_10_594), .fluid_out(k_9_297), .air_in(c_10_0));
valve v_10_595 (.fluid_in(k_10_595), .fluid_out(k_9_297), .air_in(c_10_1));
valve v_10_596 (.fluid_in(k_10_596), .fluid_out(k_9_298), .air_in(c_10_0));
valve v_10_597 (.fluid_in(k_10_597), .fluid_out(k_9_298), .air_in(c_10_1));
valve v_10_598 (.fluid_in(k_10_598), .fluid_out(k_9_299), .air_in(c_10_0));
valve v_10_599 (.fluid_in(k_10_599), .fluid_out(k_9_299), .air_in(c_10_1));
valve v_10_600 (.fluid_in(k_10_600), .fluid_out(k_9_300), .air_in(c_10_0));
valve v_10_601 (.fluid_in(k_10_601), .fluid_out(k_9_300), .air_in(c_10_1));
valve v_10_602 (.fluid_in(k_10_602), .fluid_out(k_9_301), .air_in(c_10_0));
valve v_10_603 (.fluid_in(k_10_603), .fluid_out(k_9_301), .air_in(c_10_1));
valve v_10_604 (.fluid_in(k_10_604), .fluid_out(k_9_302), .air_in(c_10_0));
valve v_10_605 (.fluid_in(k_10_605), .fluid_out(k_9_302), .air_in(c_10_1));
valve v_10_606 (.fluid_in(k_10_606), .fluid_out(k_9_303), .air_in(c_10_0));
valve v_10_607 (.fluid_in(k_10_607), .fluid_out(k_9_303), .air_in(c_10_1));
valve v_10_608 (.fluid_in(k_10_608), .fluid_out(k_9_304), .air_in(c_10_0));
valve v_10_609 (.fluid_in(k_10_609), .fluid_out(k_9_304), .air_in(c_10_1));
valve v_10_610 (.fluid_in(k_10_610), .fluid_out(k_9_305), .air_in(c_10_0));
valve v_10_611 (.fluid_in(k_10_611), .fluid_out(k_9_305), .air_in(c_10_1));
valve v_10_612 (.fluid_in(k_10_612), .fluid_out(k_9_306), .air_in(c_10_0));
valve v_10_613 (.fluid_in(k_10_613), .fluid_out(k_9_306), .air_in(c_10_1));
valve v_10_614 (.fluid_in(k_10_614), .fluid_out(k_9_307), .air_in(c_10_0));
valve v_10_615 (.fluid_in(k_10_615), .fluid_out(k_9_307), .air_in(c_10_1));
valve v_10_616 (.fluid_in(k_10_616), .fluid_out(k_9_308), .air_in(c_10_0));
valve v_10_617 (.fluid_in(k_10_617), .fluid_out(k_9_308), .air_in(c_10_1));
valve v_10_618 (.fluid_in(k_10_618), .fluid_out(k_9_309), .air_in(c_10_0));
valve v_10_619 (.fluid_in(k_10_619), .fluid_out(k_9_309), .air_in(c_10_1));
valve v_10_620 (.fluid_in(k_10_620), .fluid_out(k_9_310), .air_in(c_10_0));
valve v_10_621 (.fluid_in(k_10_621), .fluid_out(k_9_310), .air_in(c_10_1));
valve v_10_622 (.fluid_in(k_10_622), .fluid_out(k_9_311), .air_in(c_10_0));
valve v_10_623 (.fluid_in(k_10_623), .fluid_out(k_9_311), .air_in(c_10_1));
valve v_10_624 (.fluid_in(k_10_624), .fluid_out(k_9_312), .air_in(c_10_0));
valve v_10_625 (.fluid_in(k_10_625), .fluid_out(k_9_312), .air_in(c_10_1));
valve v_10_626 (.fluid_in(k_10_626), .fluid_out(k_9_313), .air_in(c_10_0));
valve v_10_627 (.fluid_in(k_10_627), .fluid_out(k_9_313), .air_in(c_10_1));
valve v_10_628 (.fluid_in(k_10_628), .fluid_out(k_9_314), .air_in(c_10_0));
valve v_10_629 (.fluid_in(k_10_629), .fluid_out(k_9_314), .air_in(c_10_1));
valve v_10_630 (.fluid_in(k_10_630), .fluid_out(k_9_315), .air_in(c_10_0));
valve v_10_631 (.fluid_in(k_10_631), .fluid_out(k_9_315), .air_in(c_10_1));
valve v_10_632 (.fluid_in(k_10_632), .fluid_out(k_9_316), .air_in(c_10_0));
valve v_10_633 (.fluid_in(k_10_633), .fluid_out(k_9_316), .air_in(c_10_1));
valve v_10_634 (.fluid_in(k_10_634), .fluid_out(k_9_317), .air_in(c_10_0));
valve v_10_635 (.fluid_in(k_10_635), .fluid_out(k_9_317), .air_in(c_10_1));
valve v_10_636 (.fluid_in(k_10_636), .fluid_out(k_9_318), .air_in(c_10_0));
valve v_10_637 (.fluid_in(k_10_637), .fluid_out(k_9_318), .air_in(c_10_1));
valve v_10_638 (.fluid_in(k_10_638), .fluid_out(k_9_319), .air_in(c_10_0));
valve v_10_639 (.fluid_in(k_10_639), .fluid_out(k_9_319), .air_in(c_10_1));
valve v_10_640 (.fluid_in(k_10_640), .fluid_out(k_9_320), .air_in(c_10_0));
valve v_10_641 (.fluid_in(k_10_641), .fluid_out(k_9_320), .air_in(c_10_1));
valve v_10_642 (.fluid_in(k_10_642), .fluid_out(k_9_321), .air_in(c_10_0));
valve v_10_643 (.fluid_in(k_10_643), .fluid_out(k_9_321), .air_in(c_10_1));
valve v_10_644 (.fluid_in(k_10_644), .fluid_out(k_9_322), .air_in(c_10_0));
valve v_10_645 (.fluid_in(k_10_645), .fluid_out(k_9_322), .air_in(c_10_1));
valve v_10_646 (.fluid_in(k_10_646), .fluid_out(k_9_323), .air_in(c_10_0));
valve v_10_647 (.fluid_in(k_10_647), .fluid_out(k_9_323), .air_in(c_10_1));
valve v_10_648 (.fluid_in(k_10_648), .fluid_out(k_9_324), .air_in(c_10_0));
valve v_10_649 (.fluid_in(k_10_649), .fluid_out(k_9_324), .air_in(c_10_1));
valve v_10_650 (.fluid_in(k_10_650), .fluid_out(k_9_325), .air_in(c_10_0));
valve v_10_651 (.fluid_in(k_10_651), .fluid_out(k_9_325), .air_in(c_10_1));
valve v_10_652 (.fluid_in(k_10_652), .fluid_out(k_9_326), .air_in(c_10_0));
valve v_10_653 (.fluid_in(k_10_653), .fluid_out(k_9_326), .air_in(c_10_1));
valve v_10_654 (.fluid_in(k_10_654), .fluid_out(k_9_327), .air_in(c_10_0));
valve v_10_655 (.fluid_in(k_10_655), .fluid_out(k_9_327), .air_in(c_10_1));
valve v_10_656 (.fluid_in(k_10_656), .fluid_out(k_9_328), .air_in(c_10_0));
valve v_10_657 (.fluid_in(k_10_657), .fluid_out(k_9_328), .air_in(c_10_1));
valve v_10_658 (.fluid_in(k_10_658), .fluid_out(k_9_329), .air_in(c_10_0));
valve v_10_659 (.fluid_in(k_10_659), .fluid_out(k_9_329), .air_in(c_10_1));
valve v_10_660 (.fluid_in(k_10_660), .fluid_out(k_9_330), .air_in(c_10_0));
valve v_10_661 (.fluid_in(k_10_661), .fluid_out(k_9_330), .air_in(c_10_1));
valve v_10_662 (.fluid_in(k_10_662), .fluid_out(k_9_331), .air_in(c_10_0));
valve v_10_663 (.fluid_in(k_10_663), .fluid_out(k_9_331), .air_in(c_10_1));
valve v_10_664 (.fluid_in(k_10_664), .fluid_out(k_9_332), .air_in(c_10_0));
valve v_10_665 (.fluid_in(k_10_665), .fluid_out(k_9_332), .air_in(c_10_1));
valve v_10_666 (.fluid_in(k_10_666), .fluid_out(k_9_333), .air_in(c_10_0));
valve v_10_667 (.fluid_in(k_10_667), .fluid_out(k_9_333), .air_in(c_10_1));
valve v_10_668 (.fluid_in(k_10_668), .fluid_out(k_9_334), .air_in(c_10_0));
valve v_10_669 (.fluid_in(k_10_669), .fluid_out(k_9_334), .air_in(c_10_1));
valve v_10_670 (.fluid_in(k_10_670), .fluid_out(k_9_335), .air_in(c_10_0));
valve v_10_671 (.fluid_in(k_10_671), .fluid_out(k_9_335), .air_in(c_10_1));
valve v_10_672 (.fluid_in(k_10_672), .fluid_out(k_9_336), .air_in(c_10_0));
valve v_10_673 (.fluid_in(k_10_673), .fluid_out(k_9_336), .air_in(c_10_1));
valve v_10_674 (.fluid_in(k_10_674), .fluid_out(k_9_337), .air_in(c_10_0));
valve v_10_675 (.fluid_in(k_10_675), .fluid_out(k_9_337), .air_in(c_10_1));
valve v_10_676 (.fluid_in(k_10_676), .fluid_out(k_9_338), .air_in(c_10_0));
valve v_10_677 (.fluid_in(k_10_677), .fluid_out(k_9_338), .air_in(c_10_1));
valve v_10_678 (.fluid_in(k_10_678), .fluid_out(k_9_339), .air_in(c_10_0));
valve v_10_679 (.fluid_in(k_10_679), .fluid_out(k_9_339), .air_in(c_10_1));
valve v_10_680 (.fluid_in(k_10_680), .fluid_out(k_9_340), .air_in(c_10_0));
valve v_10_681 (.fluid_in(k_10_681), .fluid_out(k_9_340), .air_in(c_10_1));
valve v_10_682 (.fluid_in(k_10_682), .fluid_out(k_9_341), .air_in(c_10_0));
valve v_10_683 (.fluid_in(k_10_683), .fluid_out(k_9_341), .air_in(c_10_1));
valve v_10_684 (.fluid_in(k_10_684), .fluid_out(k_9_342), .air_in(c_10_0));
valve v_10_685 (.fluid_in(k_10_685), .fluid_out(k_9_342), .air_in(c_10_1));
valve v_10_686 (.fluid_in(k_10_686), .fluid_out(k_9_343), .air_in(c_10_0));
valve v_10_687 (.fluid_in(k_10_687), .fluid_out(k_9_343), .air_in(c_10_1));
valve v_10_688 (.fluid_in(k_10_688), .fluid_out(k_9_344), .air_in(c_10_0));
valve v_10_689 (.fluid_in(k_10_689), .fluid_out(k_9_344), .air_in(c_10_1));
valve v_10_690 (.fluid_in(k_10_690), .fluid_out(k_9_345), .air_in(c_10_0));
valve v_10_691 (.fluid_in(k_10_691), .fluid_out(k_9_345), .air_in(c_10_1));
valve v_10_692 (.fluid_in(k_10_692), .fluid_out(k_9_346), .air_in(c_10_0));
valve v_10_693 (.fluid_in(k_10_693), .fluid_out(k_9_346), .air_in(c_10_1));
valve v_10_694 (.fluid_in(k_10_694), .fluid_out(k_9_347), .air_in(c_10_0));
valve v_10_695 (.fluid_in(k_10_695), .fluid_out(k_9_347), .air_in(c_10_1));
valve v_10_696 (.fluid_in(k_10_696), .fluid_out(k_9_348), .air_in(c_10_0));
valve v_10_697 (.fluid_in(k_10_697), .fluid_out(k_9_348), .air_in(c_10_1));
valve v_10_698 (.fluid_in(k_10_698), .fluid_out(k_9_349), .air_in(c_10_0));
valve v_10_699 (.fluid_in(k_10_699), .fluid_out(k_9_349), .air_in(c_10_1));
valve v_10_700 (.fluid_in(k_10_700), .fluid_out(k_9_350), .air_in(c_10_0));
valve v_10_701 (.fluid_in(k_10_701), .fluid_out(k_9_350), .air_in(c_10_1));
valve v_10_702 (.fluid_in(k_10_702), .fluid_out(k_9_351), .air_in(c_10_0));
valve v_10_703 (.fluid_in(k_10_703), .fluid_out(k_9_351), .air_in(c_10_1));
valve v_10_704 (.fluid_in(k_10_704), .fluid_out(k_9_352), .air_in(c_10_0));
valve v_10_705 (.fluid_in(k_10_705), .fluid_out(k_9_352), .air_in(c_10_1));
valve v_10_706 (.fluid_in(k_10_706), .fluid_out(k_9_353), .air_in(c_10_0));
valve v_10_707 (.fluid_in(k_10_707), .fluid_out(k_9_353), .air_in(c_10_1));
valve v_10_708 (.fluid_in(k_10_708), .fluid_out(k_9_354), .air_in(c_10_0));
valve v_10_709 (.fluid_in(k_10_709), .fluid_out(k_9_354), .air_in(c_10_1));
valve v_10_710 (.fluid_in(k_10_710), .fluid_out(k_9_355), .air_in(c_10_0));
valve v_10_711 (.fluid_in(k_10_711), .fluid_out(k_9_355), .air_in(c_10_1));
valve v_10_712 (.fluid_in(k_10_712), .fluid_out(k_9_356), .air_in(c_10_0));
valve v_10_713 (.fluid_in(k_10_713), .fluid_out(k_9_356), .air_in(c_10_1));
valve v_10_714 (.fluid_in(k_10_714), .fluid_out(k_9_357), .air_in(c_10_0));
valve v_10_715 (.fluid_in(k_10_715), .fluid_out(k_9_357), .air_in(c_10_1));
valve v_10_716 (.fluid_in(k_10_716), .fluid_out(k_9_358), .air_in(c_10_0));
valve v_10_717 (.fluid_in(k_10_717), .fluid_out(k_9_358), .air_in(c_10_1));
valve v_10_718 (.fluid_in(k_10_718), .fluid_out(k_9_359), .air_in(c_10_0));
valve v_10_719 (.fluid_in(k_10_719), .fluid_out(k_9_359), .air_in(c_10_1));
valve v_10_720 (.fluid_in(k_10_720), .fluid_out(k_9_360), .air_in(c_10_0));
valve v_10_721 (.fluid_in(k_10_721), .fluid_out(k_9_360), .air_in(c_10_1));
valve v_10_722 (.fluid_in(k_10_722), .fluid_out(k_9_361), .air_in(c_10_0));
valve v_10_723 (.fluid_in(k_10_723), .fluid_out(k_9_361), .air_in(c_10_1));
valve v_10_724 (.fluid_in(k_10_724), .fluid_out(k_9_362), .air_in(c_10_0));
valve v_10_725 (.fluid_in(k_10_725), .fluid_out(k_9_362), .air_in(c_10_1));
valve v_10_726 (.fluid_in(k_10_726), .fluid_out(k_9_363), .air_in(c_10_0));
valve v_10_727 (.fluid_in(k_10_727), .fluid_out(k_9_363), .air_in(c_10_1));
valve v_10_728 (.fluid_in(k_10_728), .fluid_out(k_9_364), .air_in(c_10_0));
valve v_10_729 (.fluid_in(k_10_729), .fluid_out(k_9_364), .air_in(c_10_1));
valve v_10_730 (.fluid_in(k_10_730), .fluid_out(k_9_365), .air_in(c_10_0));
valve v_10_731 (.fluid_in(k_10_731), .fluid_out(k_9_365), .air_in(c_10_1));
valve v_10_732 (.fluid_in(k_10_732), .fluid_out(k_9_366), .air_in(c_10_0));
valve v_10_733 (.fluid_in(k_10_733), .fluid_out(k_9_366), .air_in(c_10_1));
valve v_10_734 (.fluid_in(k_10_734), .fluid_out(k_9_367), .air_in(c_10_0));
valve v_10_735 (.fluid_in(k_10_735), .fluid_out(k_9_367), .air_in(c_10_1));
valve v_10_736 (.fluid_in(k_10_736), .fluid_out(k_9_368), .air_in(c_10_0));
valve v_10_737 (.fluid_in(k_10_737), .fluid_out(k_9_368), .air_in(c_10_1));
valve v_10_738 (.fluid_in(k_10_738), .fluid_out(k_9_369), .air_in(c_10_0));
valve v_10_739 (.fluid_in(k_10_739), .fluid_out(k_9_369), .air_in(c_10_1));
valve v_10_740 (.fluid_in(k_10_740), .fluid_out(k_9_370), .air_in(c_10_0));
valve v_10_741 (.fluid_in(k_10_741), .fluid_out(k_9_370), .air_in(c_10_1));
valve v_10_742 (.fluid_in(k_10_742), .fluid_out(k_9_371), .air_in(c_10_0));
valve v_10_743 (.fluid_in(k_10_743), .fluid_out(k_9_371), .air_in(c_10_1));
valve v_10_744 (.fluid_in(k_10_744), .fluid_out(k_9_372), .air_in(c_10_0));
valve v_10_745 (.fluid_in(k_10_745), .fluid_out(k_9_372), .air_in(c_10_1));
valve v_10_746 (.fluid_in(k_10_746), .fluid_out(k_9_373), .air_in(c_10_0));
valve v_10_747 (.fluid_in(k_10_747), .fluid_out(k_9_373), .air_in(c_10_1));
valve v_10_748 (.fluid_in(k_10_748), .fluid_out(k_9_374), .air_in(c_10_0));
valve v_10_749 (.fluid_in(k_10_749), .fluid_out(k_9_374), .air_in(c_10_1));
valve v_10_750 (.fluid_in(k_10_750), .fluid_out(k_9_375), .air_in(c_10_0));
valve v_10_751 (.fluid_in(k_10_751), .fluid_out(k_9_375), .air_in(c_10_1));
valve v_10_752 (.fluid_in(k_10_752), .fluid_out(k_9_376), .air_in(c_10_0));
valve v_10_753 (.fluid_in(k_10_753), .fluid_out(k_9_376), .air_in(c_10_1));
valve v_10_754 (.fluid_in(k_10_754), .fluid_out(k_9_377), .air_in(c_10_0));
valve v_10_755 (.fluid_in(k_10_755), .fluid_out(k_9_377), .air_in(c_10_1));
valve v_10_756 (.fluid_in(k_10_756), .fluid_out(k_9_378), .air_in(c_10_0));
valve v_10_757 (.fluid_in(k_10_757), .fluid_out(k_9_378), .air_in(c_10_1));
valve v_10_758 (.fluid_in(k_10_758), .fluid_out(k_9_379), .air_in(c_10_0));
valve v_10_759 (.fluid_in(k_10_759), .fluid_out(k_9_379), .air_in(c_10_1));
valve v_10_760 (.fluid_in(k_10_760), .fluid_out(k_9_380), .air_in(c_10_0));
valve v_10_761 (.fluid_in(k_10_761), .fluid_out(k_9_380), .air_in(c_10_1));
valve v_10_762 (.fluid_in(k_10_762), .fluid_out(k_9_381), .air_in(c_10_0));
valve v_10_763 (.fluid_in(k_10_763), .fluid_out(k_9_381), .air_in(c_10_1));
valve v_10_764 (.fluid_in(k_10_764), .fluid_out(k_9_382), .air_in(c_10_0));
valve v_10_765 (.fluid_in(k_10_765), .fluid_out(k_9_382), .air_in(c_10_1));
valve v_10_766 (.fluid_in(k_10_766), .fluid_out(k_9_383), .air_in(c_10_0));
valve v_10_767 (.fluid_in(k_10_767), .fluid_out(k_9_383), .air_in(c_10_1));
valve v_10_768 (.fluid_in(k_10_768), .fluid_out(k_9_384), .air_in(c_10_0));
valve v_10_769 (.fluid_in(k_10_769), .fluid_out(k_9_384), .air_in(c_10_1));
valve v_10_770 (.fluid_in(k_10_770), .fluid_out(k_9_385), .air_in(c_10_0));
valve v_10_771 (.fluid_in(k_10_771), .fluid_out(k_9_385), .air_in(c_10_1));
valve v_10_772 (.fluid_in(k_10_772), .fluid_out(k_9_386), .air_in(c_10_0));
valve v_10_773 (.fluid_in(k_10_773), .fluid_out(k_9_386), .air_in(c_10_1));
valve v_10_774 (.fluid_in(k_10_774), .fluid_out(k_9_387), .air_in(c_10_0));
valve v_10_775 (.fluid_in(k_10_775), .fluid_out(k_9_387), .air_in(c_10_1));
valve v_10_776 (.fluid_in(k_10_776), .fluid_out(k_9_388), .air_in(c_10_0));
valve v_10_777 (.fluid_in(k_10_777), .fluid_out(k_9_388), .air_in(c_10_1));
valve v_10_778 (.fluid_in(k_10_778), .fluid_out(k_9_389), .air_in(c_10_0));
valve v_10_779 (.fluid_in(k_10_779), .fluid_out(k_9_389), .air_in(c_10_1));
valve v_10_780 (.fluid_in(k_10_780), .fluid_out(k_9_390), .air_in(c_10_0));
valve v_10_781 (.fluid_in(k_10_781), .fluid_out(k_9_390), .air_in(c_10_1));
valve v_10_782 (.fluid_in(k_10_782), .fluid_out(k_9_391), .air_in(c_10_0));
valve v_10_783 (.fluid_in(k_10_783), .fluid_out(k_9_391), .air_in(c_10_1));
valve v_10_784 (.fluid_in(k_10_784), .fluid_out(k_9_392), .air_in(c_10_0));
valve v_10_785 (.fluid_in(k_10_785), .fluid_out(k_9_392), .air_in(c_10_1));
valve v_10_786 (.fluid_in(k_10_786), .fluid_out(k_9_393), .air_in(c_10_0));
valve v_10_787 (.fluid_in(k_10_787), .fluid_out(k_9_393), .air_in(c_10_1));
valve v_10_788 (.fluid_in(k_10_788), .fluid_out(k_9_394), .air_in(c_10_0));
valve v_10_789 (.fluid_in(k_10_789), .fluid_out(k_9_394), .air_in(c_10_1));
valve v_10_790 (.fluid_in(k_10_790), .fluid_out(k_9_395), .air_in(c_10_0));
valve v_10_791 (.fluid_in(k_10_791), .fluid_out(k_9_395), .air_in(c_10_1));
valve v_10_792 (.fluid_in(k_10_792), .fluid_out(k_9_396), .air_in(c_10_0));
valve v_10_793 (.fluid_in(k_10_793), .fluid_out(k_9_396), .air_in(c_10_1));
valve v_10_794 (.fluid_in(k_10_794), .fluid_out(k_9_397), .air_in(c_10_0));
valve v_10_795 (.fluid_in(k_10_795), .fluid_out(k_9_397), .air_in(c_10_1));
valve v_10_796 (.fluid_in(k_10_796), .fluid_out(k_9_398), .air_in(c_10_0));
valve v_10_797 (.fluid_in(k_10_797), .fluid_out(k_9_398), .air_in(c_10_1));
valve v_10_798 (.fluid_in(k_10_798), .fluid_out(k_9_399), .air_in(c_10_0));
valve v_10_799 (.fluid_in(k_10_799), .fluid_out(k_9_399), .air_in(c_10_1));
valve v_10_800 (.fluid_in(k_10_800), .fluid_out(k_9_400), .air_in(c_10_0));
valve v_10_801 (.fluid_in(k_10_801), .fluid_out(k_9_400), .air_in(c_10_1));
valve v_10_802 (.fluid_in(k_10_802), .fluid_out(k_9_401), .air_in(c_10_0));
valve v_10_803 (.fluid_in(k_10_803), .fluid_out(k_9_401), .air_in(c_10_1));
valve v_10_804 (.fluid_in(k_10_804), .fluid_out(k_9_402), .air_in(c_10_0));
valve v_10_805 (.fluid_in(k_10_805), .fluid_out(k_9_402), .air_in(c_10_1));
valve v_10_806 (.fluid_in(k_10_806), .fluid_out(k_9_403), .air_in(c_10_0));
valve v_10_807 (.fluid_in(k_10_807), .fluid_out(k_9_403), .air_in(c_10_1));
valve v_10_808 (.fluid_in(k_10_808), .fluid_out(k_9_404), .air_in(c_10_0));
valve v_10_809 (.fluid_in(k_10_809), .fluid_out(k_9_404), .air_in(c_10_1));
valve v_10_810 (.fluid_in(k_10_810), .fluid_out(k_9_405), .air_in(c_10_0));
valve v_10_811 (.fluid_in(k_10_811), .fluid_out(k_9_405), .air_in(c_10_1));
valve v_10_812 (.fluid_in(k_10_812), .fluid_out(k_9_406), .air_in(c_10_0));
valve v_10_813 (.fluid_in(k_10_813), .fluid_out(k_9_406), .air_in(c_10_1));
valve v_10_814 (.fluid_in(k_10_814), .fluid_out(k_9_407), .air_in(c_10_0));
valve v_10_815 (.fluid_in(k_10_815), .fluid_out(k_9_407), .air_in(c_10_1));
valve v_10_816 (.fluid_in(k_10_816), .fluid_out(k_9_408), .air_in(c_10_0));
valve v_10_817 (.fluid_in(k_10_817), .fluid_out(k_9_408), .air_in(c_10_1));
valve v_10_818 (.fluid_in(k_10_818), .fluid_out(k_9_409), .air_in(c_10_0));
valve v_10_819 (.fluid_in(k_10_819), .fluid_out(k_9_409), .air_in(c_10_1));
valve v_10_820 (.fluid_in(k_10_820), .fluid_out(k_9_410), .air_in(c_10_0));
valve v_10_821 (.fluid_in(k_10_821), .fluid_out(k_9_410), .air_in(c_10_1));
valve v_10_822 (.fluid_in(k_10_822), .fluid_out(k_9_411), .air_in(c_10_0));
valve v_10_823 (.fluid_in(k_10_823), .fluid_out(k_9_411), .air_in(c_10_1));
valve v_10_824 (.fluid_in(k_10_824), .fluid_out(k_9_412), .air_in(c_10_0));
valve v_10_825 (.fluid_in(k_10_825), .fluid_out(k_9_412), .air_in(c_10_1));
valve v_10_826 (.fluid_in(k_10_826), .fluid_out(k_9_413), .air_in(c_10_0));
valve v_10_827 (.fluid_in(k_10_827), .fluid_out(k_9_413), .air_in(c_10_1));
valve v_10_828 (.fluid_in(k_10_828), .fluid_out(k_9_414), .air_in(c_10_0));
valve v_10_829 (.fluid_in(k_10_829), .fluid_out(k_9_414), .air_in(c_10_1));
valve v_10_830 (.fluid_in(k_10_830), .fluid_out(k_9_415), .air_in(c_10_0));
valve v_10_831 (.fluid_in(k_10_831), .fluid_out(k_9_415), .air_in(c_10_1));
valve v_10_832 (.fluid_in(k_10_832), .fluid_out(k_9_416), .air_in(c_10_0));
valve v_10_833 (.fluid_in(k_10_833), .fluid_out(k_9_416), .air_in(c_10_1));
valve v_10_834 (.fluid_in(k_10_834), .fluid_out(k_9_417), .air_in(c_10_0));
valve v_10_835 (.fluid_in(k_10_835), .fluid_out(k_9_417), .air_in(c_10_1));
valve v_10_836 (.fluid_in(k_10_836), .fluid_out(k_9_418), .air_in(c_10_0));
valve v_10_837 (.fluid_in(k_10_837), .fluid_out(k_9_418), .air_in(c_10_1));
valve v_10_838 (.fluid_in(k_10_838), .fluid_out(k_9_419), .air_in(c_10_0));
valve v_10_839 (.fluid_in(k_10_839), .fluid_out(k_9_419), .air_in(c_10_1));
valve v_10_840 (.fluid_in(k_10_840), .fluid_out(k_9_420), .air_in(c_10_0));
valve v_10_841 (.fluid_in(k_10_841), .fluid_out(k_9_420), .air_in(c_10_1));
valve v_10_842 (.fluid_in(k_10_842), .fluid_out(k_9_421), .air_in(c_10_0));
valve v_10_843 (.fluid_in(k_10_843), .fluid_out(k_9_421), .air_in(c_10_1));
valve v_10_844 (.fluid_in(k_10_844), .fluid_out(k_9_422), .air_in(c_10_0));
valve v_10_845 (.fluid_in(k_10_845), .fluid_out(k_9_422), .air_in(c_10_1));
valve v_10_846 (.fluid_in(k_10_846), .fluid_out(k_9_423), .air_in(c_10_0));
valve v_10_847 (.fluid_in(k_10_847), .fluid_out(k_9_423), .air_in(c_10_1));
valve v_10_848 (.fluid_in(k_10_848), .fluid_out(k_9_424), .air_in(c_10_0));
valve v_10_849 (.fluid_in(k_10_849), .fluid_out(k_9_424), .air_in(c_10_1));
valve v_10_850 (.fluid_in(k_10_850), .fluid_out(k_9_425), .air_in(c_10_0));
valve v_10_851 (.fluid_in(k_10_851), .fluid_out(k_9_425), .air_in(c_10_1));
valve v_10_852 (.fluid_in(k_10_852), .fluid_out(k_9_426), .air_in(c_10_0));
valve v_10_853 (.fluid_in(k_10_853), .fluid_out(k_9_426), .air_in(c_10_1));
valve v_10_854 (.fluid_in(k_10_854), .fluid_out(k_9_427), .air_in(c_10_0));
valve v_10_855 (.fluid_in(k_10_855), .fluid_out(k_9_427), .air_in(c_10_1));
valve v_10_856 (.fluid_in(k_10_856), .fluid_out(k_9_428), .air_in(c_10_0));
valve v_10_857 (.fluid_in(k_10_857), .fluid_out(k_9_428), .air_in(c_10_1));
valve v_10_858 (.fluid_in(k_10_858), .fluid_out(k_9_429), .air_in(c_10_0));
valve v_10_859 (.fluid_in(k_10_859), .fluid_out(k_9_429), .air_in(c_10_1));
valve v_10_860 (.fluid_in(k_10_860), .fluid_out(k_9_430), .air_in(c_10_0));
valve v_10_861 (.fluid_in(k_10_861), .fluid_out(k_9_430), .air_in(c_10_1));
valve v_10_862 (.fluid_in(k_10_862), .fluid_out(k_9_431), .air_in(c_10_0));
valve v_10_863 (.fluid_in(k_10_863), .fluid_out(k_9_431), .air_in(c_10_1));
valve v_10_864 (.fluid_in(k_10_864), .fluid_out(k_9_432), .air_in(c_10_0));
valve v_10_865 (.fluid_in(k_10_865), .fluid_out(k_9_432), .air_in(c_10_1));
valve v_10_866 (.fluid_in(k_10_866), .fluid_out(k_9_433), .air_in(c_10_0));
valve v_10_867 (.fluid_in(k_10_867), .fluid_out(k_9_433), .air_in(c_10_1));
valve v_10_868 (.fluid_in(k_10_868), .fluid_out(k_9_434), .air_in(c_10_0));
valve v_10_869 (.fluid_in(k_10_869), .fluid_out(k_9_434), .air_in(c_10_1));
valve v_10_870 (.fluid_in(k_10_870), .fluid_out(k_9_435), .air_in(c_10_0));
valve v_10_871 (.fluid_in(k_10_871), .fluid_out(k_9_435), .air_in(c_10_1));
valve v_10_872 (.fluid_in(k_10_872), .fluid_out(k_9_436), .air_in(c_10_0));
valve v_10_873 (.fluid_in(k_10_873), .fluid_out(k_9_436), .air_in(c_10_1));
valve v_10_874 (.fluid_in(k_10_874), .fluid_out(k_9_437), .air_in(c_10_0));
valve v_10_875 (.fluid_in(k_10_875), .fluid_out(k_9_437), .air_in(c_10_1));
valve v_10_876 (.fluid_in(k_10_876), .fluid_out(k_9_438), .air_in(c_10_0));
valve v_10_877 (.fluid_in(k_10_877), .fluid_out(k_9_438), .air_in(c_10_1));
valve v_10_878 (.fluid_in(k_10_878), .fluid_out(k_9_439), .air_in(c_10_0));
valve v_10_879 (.fluid_in(k_10_879), .fluid_out(k_9_439), .air_in(c_10_1));
valve v_10_880 (.fluid_in(k_10_880), .fluid_out(k_9_440), .air_in(c_10_0));
valve v_10_881 (.fluid_in(k_10_881), .fluid_out(k_9_440), .air_in(c_10_1));
valve v_10_882 (.fluid_in(k_10_882), .fluid_out(k_9_441), .air_in(c_10_0));
valve v_10_883 (.fluid_in(k_10_883), .fluid_out(k_9_441), .air_in(c_10_1));
valve v_10_884 (.fluid_in(k_10_884), .fluid_out(k_9_442), .air_in(c_10_0));
valve v_10_885 (.fluid_in(k_10_885), .fluid_out(k_9_442), .air_in(c_10_1));
valve v_10_886 (.fluid_in(k_10_886), .fluid_out(k_9_443), .air_in(c_10_0));
valve v_10_887 (.fluid_in(k_10_887), .fluid_out(k_9_443), .air_in(c_10_1));
valve v_10_888 (.fluid_in(k_10_888), .fluid_out(k_9_444), .air_in(c_10_0));
valve v_10_889 (.fluid_in(k_10_889), .fluid_out(k_9_444), .air_in(c_10_1));
valve v_10_890 (.fluid_in(k_10_890), .fluid_out(k_9_445), .air_in(c_10_0));
valve v_10_891 (.fluid_in(k_10_891), .fluid_out(k_9_445), .air_in(c_10_1));
valve v_10_892 (.fluid_in(k_10_892), .fluid_out(k_9_446), .air_in(c_10_0));
valve v_10_893 (.fluid_in(k_10_893), .fluid_out(k_9_446), .air_in(c_10_1));
valve v_10_894 (.fluid_in(k_10_894), .fluid_out(k_9_447), .air_in(c_10_0));
valve v_10_895 (.fluid_in(k_10_895), .fluid_out(k_9_447), .air_in(c_10_1));
valve v_10_896 (.fluid_in(k_10_896), .fluid_out(k_9_448), .air_in(c_10_0));
valve v_10_897 (.fluid_in(k_10_897), .fluid_out(k_9_448), .air_in(c_10_1));
valve v_10_898 (.fluid_in(k_10_898), .fluid_out(k_9_449), .air_in(c_10_0));
valve v_10_899 (.fluid_in(k_10_899), .fluid_out(k_9_449), .air_in(c_10_1));
valve v_10_900 (.fluid_in(k_10_900), .fluid_out(k_9_450), .air_in(c_10_0));
valve v_10_901 (.fluid_in(k_10_901), .fluid_out(k_9_450), .air_in(c_10_1));
valve v_10_902 (.fluid_in(k_10_902), .fluid_out(k_9_451), .air_in(c_10_0));
valve v_10_903 (.fluid_in(k_10_903), .fluid_out(k_9_451), .air_in(c_10_1));
valve v_10_904 (.fluid_in(k_10_904), .fluid_out(k_9_452), .air_in(c_10_0));
valve v_10_905 (.fluid_in(k_10_905), .fluid_out(k_9_452), .air_in(c_10_1));
valve v_10_906 (.fluid_in(k_10_906), .fluid_out(k_9_453), .air_in(c_10_0));
valve v_10_907 (.fluid_in(k_10_907), .fluid_out(k_9_453), .air_in(c_10_1));
valve v_10_908 (.fluid_in(k_10_908), .fluid_out(k_9_454), .air_in(c_10_0));
valve v_10_909 (.fluid_in(k_10_909), .fluid_out(k_9_454), .air_in(c_10_1));
valve v_10_910 (.fluid_in(k_10_910), .fluid_out(k_9_455), .air_in(c_10_0));
valve v_10_911 (.fluid_in(k_10_911), .fluid_out(k_9_455), .air_in(c_10_1));
valve v_10_912 (.fluid_in(k_10_912), .fluid_out(k_9_456), .air_in(c_10_0));
valve v_10_913 (.fluid_in(k_10_913), .fluid_out(k_9_456), .air_in(c_10_1));
valve v_10_914 (.fluid_in(k_10_914), .fluid_out(k_9_457), .air_in(c_10_0));
valve v_10_915 (.fluid_in(k_10_915), .fluid_out(k_9_457), .air_in(c_10_1));
valve v_10_916 (.fluid_in(k_10_916), .fluid_out(k_9_458), .air_in(c_10_0));
valve v_10_917 (.fluid_in(k_10_917), .fluid_out(k_9_458), .air_in(c_10_1));
valve v_10_918 (.fluid_in(k_10_918), .fluid_out(k_9_459), .air_in(c_10_0));
valve v_10_919 (.fluid_in(k_10_919), .fluid_out(k_9_459), .air_in(c_10_1));
valve v_10_920 (.fluid_in(k_10_920), .fluid_out(k_9_460), .air_in(c_10_0));
valve v_10_921 (.fluid_in(k_10_921), .fluid_out(k_9_460), .air_in(c_10_1));
valve v_10_922 (.fluid_in(k_10_922), .fluid_out(k_9_461), .air_in(c_10_0));
valve v_10_923 (.fluid_in(k_10_923), .fluid_out(k_9_461), .air_in(c_10_1));
valve v_10_924 (.fluid_in(k_10_924), .fluid_out(k_9_462), .air_in(c_10_0));
valve v_10_925 (.fluid_in(k_10_925), .fluid_out(k_9_462), .air_in(c_10_1));
valve v_10_926 (.fluid_in(k_10_926), .fluid_out(k_9_463), .air_in(c_10_0));
valve v_10_927 (.fluid_in(k_10_927), .fluid_out(k_9_463), .air_in(c_10_1));
valve v_10_928 (.fluid_in(k_10_928), .fluid_out(k_9_464), .air_in(c_10_0));
valve v_10_929 (.fluid_in(k_10_929), .fluid_out(k_9_464), .air_in(c_10_1));
valve v_10_930 (.fluid_in(k_10_930), .fluid_out(k_9_465), .air_in(c_10_0));
valve v_10_931 (.fluid_in(k_10_931), .fluid_out(k_9_465), .air_in(c_10_1));
valve v_10_932 (.fluid_in(k_10_932), .fluid_out(k_9_466), .air_in(c_10_0));
valve v_10_933 (.fluid_in(k_10_933), .fluid_out(k_9_466), .air_in(c_10_1));
valve v_10_934 (.fluid_in(k_10_934), .fluid_out(k_9_467), .air_in(c_10_0));
valve v_10_935 (.fluid_in(k_10_935), .fluid_out(k_9_467), .air_in(c_10_1));
valve v_10_936 (.fluid_in(k_10_936), .fluid_out(k_9_468), .air_in(c_10_0));
valve v_10_937 (.fluid_in(k_10_937), .fluid_out(k_9_468), .air_in(c_10_1));
valve v_10_938 (.fluid_in(k_10_938), .fluid_out(k_9_469), .air_in(c_10_0));
valve v_10_939 (.fluid_in(k_10_939), .fluid_out(k_9_469), .air_in(c_10_1));
valve v_10_940 (.fluid_in(k_10_940), .fluid_out(k_9_470), .air_in(c_10_0));
valve v_10_941 (.fluid_in(k_10_941), .fluid_out(k_9_470), .air_in(c_10_1));
valve v_10_942 (.fluid_in(k_10_942), .fluid_out(k_9_471), .air_in(c_10_0));
valve v_10_943 (.fluid_in(k_10_943), .fluid_out(k_9_471), .air_in(c_10_1));
valve v_10_944 (.fluid_in(k_10_944), .fluid_out(k_9_472), .air_in(c_10_0));
valve v_10_945 (.fluid_in(k_10_945), .fluid_out(k_9_472), .air_in(c_10_1));
valve v_10_946 (.fluid_in(k_10_946), .fluid_out(k_9_473), .air_in(c_10_0));
valve v_10_947 (.fluid_in(k_10_947), .fluid_out(k_9_473), .air_in(c_10_1));
valve v_10_948 (.fluid_in(k_10_948), .fluid_out(k_9_474), .air_in(c_10_0));
valve v_10_949 (.fluid_in(k_10_949), .fluid_out(k_9_474), .air_in(c_10_1));
valve v_10_950 (.fluid_in(k_10_950), .fluid_out(k_9_475), .air_in(c_10_0));
valve v_10_951 (.fluid_in(k_10_951), .fluid_out(k_9_475), .air_in(c_10_1));
valve v_10_952 (.fluid_in(k_10_952), .fluid_out(k_9_476), .air_in(c_10_0));
valve v_10_953 (.fluid_in(k_10_953), .fluid_out(k_9_476), .air_in(c_10_1));
valve v_10_954 (.fluid_in(k_10_954), .fluid_out(k_9_477), .air_in(c_10_0));
valve v_10_955 (.fluid_in(k_10_955), .fluid_out(k_9_477), .air_in(c_10_1));
valve v_10_956 (.fluid_in(k_10_956), .fluid_out(k_9_478), .air_in(c_10_0));
valve v_10_957 (.fluid_in(k_10_957), .fluid_out(k_9_478), .air_in(c_10_1));
valve v_10_958 (.fluid_in(k_10_958), .fluid_out(k_9_479), .air_in(c_10_0));
valve v_10_959 (.fluid_in(k_10_959), .fluid_out(k_9_479), .air_in(c_10_1));
valve v_10_960 (.fluid_in(k_10_960), .fluid_out(k_9_480), .air_in(c_10_0));
valve v_10_961 (.fluid_in(k_10_961), .fluid_out(k_9_480), .air_in(c_10_1));
valve v_10_962 (.fluid_in(k_10_962), .fluid_out(k_9_481), .air_in(c_10_0));
valve v_10_963 (.fluid_in(k_10_963), .fluid_out(k_9_481), .air_in(c_10_1));
valve v_10_964 (.fluid_in(k_10_964), .fluid_out(k_9_482), .air_in(c_10_0));
valve v_10_965 (.fluid_in(k_10_965), .fluid_out(k_9_482), .air_in(c_10_1));
valve v_10_966 (.fluid_in(k_10_966), .fluid_out(k_9_483), .air_in(c_10_0));
valve v_10_967 (.fluid_in(k_10_967), .fluid_out(k_9_483), .air_in(c_10_1));
valve v_10_968 (.fluid_in(k_10_968), .fluid_out(k_9_484), .air_in(c_10_0));
valve v_10_969 (.fluid_in(k_10_969), .fluid_out(k_9_484), .air_in(c_10_1));
valve v_10_970 (.fluid_in(k_10_970), .fluid_out(k_9_485), .air_in(c_10_0));
valve v_10_971 (.fluid_in(k_10_971), .fluid_out(k_9_485), .air_in(c_10_1));
valve v_10_972 (.fluid_in(k_10_972), .fluid_out(k_9_486), .air_in(c_10_0));
valve v_10_973 (.fluid_in(k_10_973), .fluid_out(k_9_486), .air_in(c_10_1));
valve v_10_974 (.fluid_in(k_10_974), .fluid_out(k_9_487), .air_in(c_10_0));
valve v_10_975 (.fluid_in(k_10_975), .fluid_out(k_9_487), .air_in(c_10_1));
valve v_10_976 (.fluid_in(k_10_976), .fluid_out(k_9_488), .air_in(c_10_0));
valve v_10_977 (.fluid_in(k_10_977), .fluid_out(k_9_488), .air_in(c_10_1));
valve v_10_978 (.fluid_in(k_10_978), .fluid_out(k_9_489), .air_in(c_10_0));
valve v_10_979 (.fluid_in(k_10_979), .fluid_out(k_9_489), .air_in(c_10_1));
valve v_10_980 (.fluid_in(k_10_980), .fluid_out(k_9_490), .air_in(c_10_0));
valve v_10_981 (.fluid_in(k_10_981), .fluid_out(k_9_490), .air_in(c_10_1));
valve v_10_982 (.fluid_in(k_10_982), .fluid_out(k_9_491), .air_in(c_10_0));
valve v_10_983 (.fluid_in(k_10_983), .fluid_out(k_9_491), .air_in(c_10_1));
valve v_10_984 (.fluid_in(k_10_984), .fluid_out(k_9_492), .air_in(c_10_0));
valve v_10_985 (.fluid_in(k_10_985), .fluid_out(k_9_492), .air_in(c_10_1));
valve v_10_986 (.fluid_in(k_10_986), .fluid_out(k_9_493), .air_in(c_10_0));
valve v_10_987 (.fluid_in(k_10_987), .fluid_out(k_9_493), .air_in(c_10_1));
valve v_10_988 (.fluid_in(k_10_988), .fluid_out(k_9_494), .air_in(c_10_0));
valve v_10_989 (.fluid_in(k_10_989), .fluid_out(k_9_494), .air_in(c_10_1));
valve v_10_990 (.fluid_in(k_10_990), .fluid_out(k_9_495), .air_in(c_10_0));
valve v_10_991 (.fluid_in(k_10_991), .fluid_out(k_9_495), .air_in(c_10_1));
valve v_10_992 (.fluid_in(k_10_992), .fluid_out(k_9_496), .air_in(c_10_0));
valve v_10_993 (.fluid_in(k_10_993), .fluid_out(k_9_496), .air_in(c_10_1));
valve v_10_994 (.fluid_in(k_10_994), .fluid_out(k_9_497), .air_in(c_10_0));
valve v_10_995 (.fluid_in(k_10_995), .fluid_out(k_9_497), .air_in(c_10_1));
valve v_10_996 (.fluid_in(k_10_996), .fluid_out(k_9_498), .air_in(c_10_0));
valve v_10_997 (.fluid_in(k_10_997), .fluid_out(k_9_498), .air_in(c_10_1));
valve v_10_998 (.fluid_in(k_10_998), .fluid_out(k_9_499), .air_in(c_10_0));
valve v_10_999 (.fluid_in(k_10_999), .fluid_out(k_9_499), .air_in(c_10_1));
valve v_10_1000 (.fluid_in(k_10_1000), .fluid_out(k_9_500), .air_in(c_10_0));
valve v_10_1001 (.fluid_in(k_10_1001), .fluid_out(k_9_500), .air_in(c_10_1));
valve v_10_1002 (.fluid_in(k_10_1002), .fluid_out(k_9_501), .air_in(c_10_0));
valve v_10_1003 (.fluid_in(k_10_1003), .fluid_out(k_9_501), .air_in(c_10_1));
valve v_10_1004 (.fluid_in(k_10_1004), .fluid_out(k_9_502), .air_in(c_10_0));
valve v_10_1005 (.fluid_in(k_10_1005), .fluid_out(k_9_502), .air_in(c_10_1));
valve v_10_1006 (.fluid_in(k_10_1006), .fluid_out(k_9_503), .air_in(c_10_0));
valve v_10_1007 (.fluid_in(k_10_1007), .fluid_out(k_9_503), .air_in(c_10_1));
valve v_10_1008 (.fluid_in(k_10_1008), .fluid_out(k_9_504), .air_in(c_10_0));
valve v_10_1009 (.fluid_in(k_10_1009), .fluid_out(k_9_504), .air_in(c_10_1));
valve v_10_1010 (.fluid_in(k_10_1010), .fluid_out(k_9_505), .air_in(c_10_0));
valve v_10_1011 (.fluid_in(k_10_1011), .fluid_out(k_9_505), .air_in(c_10_1));
valve v_10_1012 (.fluid_in(k_10_1012), .fluid_out(k_9_506), .air_in(c_10_0));
valve v_10_1013 (.fluid_in(k_10_1013), .fluid_out(k_9_506), .air_in(c_10_1));
valve v_10_1014 (.fluid_in(k_10_1014), .fluid_out(k_9_507), .air_in(c_10_0));
valve v_10_1015 (.fluid_in(k_10_1015), .fluid_out(k_9_507), .air_in(c_10_1));
valve v_10_1016 (.fluid_in(k_10_1016), .fluid_out(k_9_508), .air_in(c_10_0));
valve v_10_1017 (.fluid_in(k_10_1017), .fluid_out(k_9_508), .air_in(c_10_1));
valve v_10_1018 (.fluid_in(k_10_1018), .fluid_out(k_9_509), .air_in(c_10_0));
valve v_10_1019 (.fluid_in(k_10_1019), .fluid_out(k_9_509), .air_in(c_10_1));
valve v_10_1020 (.fluid_in(k_10_1020), .fluid_out(k_9_510), .air_in(c_10_0));
valve v_10_1021 (.fluid_in(k_10_1021), .fluid_out(k_9_510), .air_in(c_10_1));
valve v_10_1022 (.fluid_in(k_10_1022), .fluid_out(k_9_511), .air_in(c_10_0));
valve v_10_1023 (.fluid_in(k_10_1023), .fluid_out(k_9_511), .air_in(c_10_1));
valve v_11_0 (.fluid_in(k_11_0), .fluid_out(k_10_0), .air_in(c_11_0));
valve v_11_1 (.fluid_in(k_11_1), .fluid_out(k_10_0), .air_in(c_11_1));
valve v_11_2 (.fluid_in(k_11_2), .fluid_out(k_10_1), .air_in(c_11_0));
valve v_11_3 (.fluid_in(k_11_3), .fluid_out(k_10_1), .air_in(c_11_1));
valve v_11_4 (.fluid_in(k_11_4), .fluid_out(k_10_2), .air_in(c_11_0));
valve v_11_5 (.fluid_in(k_11_5), .fluid_out(k_10_2), .air_in(c_11_1));
valve v_11_6 (.fluid_in(k_11_6), .fluid_out(k_10_3), .air_in(c_11_0));
valve v_11_7 (.fluid_in(k_11_7), .fluid_out(k_10_3), .air_in(c_11_1));
valve v_11_8 (.fluid_in(k_11_8), .fluid_out(k_10_4), .air_in(c_11_0));
valve v_11_9 (.fluid_in(k_11_9), .fluid_out(k_10_4), .air_in(c_11_1));
valve v_11_10 (.fluid_in(k_11_10), .fluid_out(k_10_5), .air_in(c_11_0));
valve v_11_11 (.fluid_in(k_11_11), .fluid_out(k_10_5), .air_in(c_11_1));
valve v_11_12 (.fluid_in(k_11_12), .fluid_out(k_10_6), .air_in(c_11_0));
valve v_11_13 (.fluid_in(k_11_13), .fluid_out(k_10_6), .air_in(c_11_1));
valve v_11_14 (.fluid_in(k_11_14), .fluid_out(k_10_7), .air_in(c_11_0));
valve v_11_15 (.fluid_in(k_11_15), .fluid_out(k_10_7), .air_in(c_11_1));
valve v_11_16 (.fluid_in(k_11_16), .fluid_out(k_10_8), .air_in(c_11_0));
valve v_11_17 (.fluid_in(k_11_17), .fluid_out(k_10_8), .air_in(c_11_1));
valve v_11_18 (.fluid_in(k_11_18), .fluid_out(k_10_9), .air_in(c_11_0));
valve v_11_19 (.fluid_in(k_11_19), .fluid_out(k_10_9), .air_in(c_11_1));
valve v_11_20 (.fluid_in(k_11_20), .fluid_out(k_10_10), .air_in(c_11_0));
valve v_11_21 (.fluid_in(k_11_21), .fluid_out(k_10_10), .air_in(c_11_1));
valve v_11_22 (.fluid_in(k_11_22), .fluid_out(k_10_11), .air_in(c_11_0));
valve v_11_23 (.fluid_in(k_11_23), .fluid_out(k_10_11), .air_in(c_11_1));
valve v_11_24 (.fluid_in(k_11_24), .fluid_out(k_10_12), .air_in(c_11_0));
valve v_11_25 (.fluid_in(k_11_25), .fluid_out(k_10_12), .air_in(c_11_1));
valve v_11_26 (.fluid_in(k_11_26), .fluid_out(k_10_13), .air_in(c_11_0));
valve v_11_27 (.fluid_in(k_11_27), .fluid_out(k_10_13), .air_in(c_11_1));
valve v_11_28 (.fluid_in(k_11_28), .fluid_out(k_10_14), .air_in(c_11_0));
valve v_11_29 (.fluid_in(k_11_29), .fluid_out(k_10_14), .air_in(c_11_1));
valve v_11_30 (.fluid_in(k_11_30), .fluid_out(k_10_15), .air_in(c_11_0));
valve v_11_31 (.fluid_in(k_11_31), .fluid_out(k_10_15), .air_in(c_11_1));
valve v_11_32 (.fluid_in(k_11_32), .fluid_out(k_10_16), .air_in(c_11_0));
valve v_11_33 (.fluid_in(k_11_33), .fluid_out(k_10_16), .air_in(c_11_1));
valve v_11_34 (.fluid_in(k_11_34), .fluid_out(k_10_17), .air_in(c_11_0));
valve v_11_35 (.fluid_in(k_11_35), .fluid_out(k_10_17), .air_in(c_11_1));
valve v_11_36 (.fluid_in(k_11_36), .fluid_out(k_10_18), .air_in(c_11_0));
valve v_11_37 (.fluid_in(k_11_37), .fluid_out(k_10_18), .air_in(c_11_1));
valve v_11_38 (.fluid_in(k_11_38), .fluid_out(k_10_19), .air_in(c_11_0));
valve v_11_39 (.fluid_in(k_11_39), .fluid_out(k_10_19), .air_in(c_11_1));
valve v_11_40 (.fluid_in(k_11_40), .fluid_out(k_10_20), .air_in(c_11_0));
valve v_11_41 (.fluid_in(k_11_41), .fluid_out(k_10_20), .air_in(c_11_1));
valve v_11_42 (.fluid_in(k_11_42), .fluid_out(k_10_21), .air_in(c_11_0));
valve v_11_43 (.fluid_in(k_11_43), .fluid_out(k_10_21), .air_in(c_11_1));
valve v_11_44 (.fluid_in(k_11_44), .fluid_out(k_10_22), .air_in(c_11_0));
valve v_11_45 (.fluid_in(k_11_45), .fluid_out(k_10_22), .air_in(c_11_1));
valve v_11_46 (.fluid_in(k_11_46), .fluid_out(k_10_23), .air_in(c_11_0));
valve v_11_47 (.fluid_in(k_11_47), .fluid_out(k_10_23), .air_in(c_11_1));
valve v_11_48 (.fluid_in(k_11_48), .fluid_out(k_10_24), .air_in(c_11_0));
valve v_11_49 (.fluid_in(k_11_49), .fluid_out(k_10_24), .air_in(c_11_1));
valve v_11_50 (.fluid_in(k_11_50), .fluid_out(k_10_25), .air_in(c_11_0));
valve v_11_51 (.fluid_in(k_11_51), .fluid_out(k_10_25), .air_in(c_11_1));
valve v_11_52 (.fluid_in(k_11_52), .fluid_out(k_10_26), .air_in(c_11_0));
valve v_11_53 (.fluid_in(k_11_53), .fluid_out(k_10_26), .air_in(c_11_1));
valve v_11_54 (.fluid_in(k_11_54), .fluid_out(k_10_27), .air_in(c_11_0));
valve v_11_55 (.fluid_in(k_11_55), .fluid_out(k_10_27), .air_in(c_11_1));
valve v_11_56 (.fluid_in(k_11_56), .fluid_out(k_10_28), .air_in(c_11_0));
valve v_11_57 (.fluid_in(k_11_57), .fluid_out(k_10_28), .air_in(c_11_1));
valve v_11_58 (.fluid_in(k_11_58), .fluid_out(k_10_29), .air_in(c_11_0));
valve v_11_59 (.fluid_in(k_11_59), .fluid_out(k_10_29), .air_in(c_11_1));
valve v_11_60 (.fluid_in(k_11_60), .fluid_out(k_10_30), .air_in(c_11_0));
valve v_11_61 (.fluid_in(k_11_61), .fluid_out(k_10_30), .air_in(c_11_1));
valve v_11_62 (.fluid_in(k_11_62), .fluid_out(k_10_31), .air_in(c_11_0));
valve v_11_63 (.fluid_in(k_11_63), .fluid_out(k_10_31), .air_in(c_11_1));
valve v_11_64 (.fluid_in(k_11_64), .fluid_out(k_10_32), .air_in(c_11_0));
valve v_11_65 (.fluid_in(k_11_65), .fluid_out(k_10_32), .air_in(c_11_1));
valve v_11_66 (.fluid_in(k_11_66), .fluid_out(k_10_33), .air_in(c_11_0));
valve v_11_67 (.fluid_in(k_11_67), .fluid_out(k_10_33), .air_in(c_11_1));
valve v_11_68 (.fluid_in(k_11_68), .fluid_out(k_10_34), .air_in(c_11_0));
valve v_11_69 (.fluid_in(k_11_69), .fluid_out(k_10_34), .air_in(c_11_1));
valve v_11_70 (.fluid_in(k_11_70), .fluid_out(k_10_35), .air_in(c_11_0));
valve v_11_71 (.fluid_in(k_11_71), .fluid_out(k_10_35), .air_in(c_11_1));
valve v_11_72 (.fluid_in(k_11_72), .fluid_out(k_10_36), .air_in(c_11_0));
valve v_11_73 (.fluid_in(k_11_73), .fluid_out(k_10_36), .air_in(c_11_1));
valve v_11_74 (.fluid_in(k_11_74), .fluid_out(k_10_37), .air_in(c_11_0));
valve v_11_75 (.fluid_in(k_11_75), .fluid_out(k_10_37), .air_in(c_11_1));
valve v_11_76 (.fluid_in(k_11_76), .fluid_out(k_10_38), .air_in(c_11_0));
valve v_11_77 (.fluid_in(k_11_77), .fluid_out(k_10_38), .air_in(c_11_1));
valve v_11_78 (.fluid_in(k_11_78), .fluid_out(k_10_39), .air_in(c_11_0));
valve v_11_79 (.fluid_in(k_11_79), .fluid_out(k_10_39), .air_in(c_11_1));
valve v_11_80 (.fluid_in(k_11_80), .fluid_out(k_10_40), .air_in(c_11_0));
valve v_11_81 (.fluid_in(k_11_81), .fluid_out(k_10_40), .air_in(c_11_1));
valve v_11_82 (.fluid_in(k_11_82), .fluid_out(k_10_41), .air_in(c_11_0));
valve v_11_83 (.fluid_in(k_11_83), .fluid_out(k_10_41), .air_in(c_11_1));
valve v_11_84 (.fluid_in(k_11_84), .fluid_out(k_10_42), .air_in(c_11_0));
valve v_11_85 (.fluid_in(k_11_85), .fluid_out(k_10_42), .air_in(c_11_1));
valve v_11_86 (.fluid_in(k_11_86), .fluid_out(k_10_43), .air_in(c_11_0));
valve v_11_87 (.fluid_in(k_11_87), .fluid_out(k_10_43), .air_in(c_11_1));
valve v_11_88 (.fluid_in(k_11_88), .fluid_out(k_10_44), .air_in(c_11_0));
valve v_11_89 (.fluid_in(k_11_89), .fluid_out(k_10_44), .air_in(c_11_1));
valve v_11_90 (.fluid_in(k_11_90), .fluid_out(k_10_45), .air_in(c_11_0));
valve v_11_91 (.fluid_in(k_11_91), .fluid_out(k_10_45), .air_in(c_11_1));
valve v_11_92 (.fluid_in(k_11_92), .fluid_out(k_10_46), .air_in(c_11_0));
valve v_11_93 (.fluid_in(k_11_93), .fluid_out(k_10_46), .air_in(c_11_1));
valve v_11_94 (.fluid_in(k_11_94), .fluid_out(k_10_47), .air_in(c_11_0));
valve v_11_95 (.fluid_in(k_11_95), .fluid_out(k_10_47), .air_in(c_11_1));
valve v_11_96 (.fluid_in(k_11_96), .fluid_out(k_10_48), .air_in(c_11_0));
valve v_11_97 (.fluid_in(k_11_97), .fluid_out(k_10_48), .air_in(c_11_1));
valve v_11_98 (.fluid_in(k_11_98), .fluid_out(k_10_49), .air_in(c_11_0));
valve v_11_99 (.fluid_in(k_11_99), .fluid_out(k_10_49), .air_in(c_11_1));
valve v_11_100 (.fluid_in(k_11_100), .fluid_out(k_10_50), .air_in(c_11_0));
valve v_11_101 (.fluid_in(k_11_101), .fluid_out(k_10_50), .air_in(c_11_1));
valve v_11_102 (.fluid_in(k_11_102), .fluid_out(k_10_51), .air_in(c_11_0));
valve v_11_103 (.fluid_in(k_11_103), .fluid_out(k_10_51), .air_in(c_11_1));
valve v_11_104 (.fluid_in(k_11_104), .fluid_out(k_10_52), .air_in(c_11_0));
valve v_11_105 (.fluid_in(k_11_105), .fluid_out(k_10_52), .air_in(c_11_1));
valve v_11_106 (.fluid_in(k_11_106), .fluid_out(k_10_53), .air_in(c_11_0));
valve v_11_107 (.fluid_in(k_11_107), .fluid_out(k_10_53), .air_in(c_11_1));
valve v_11_108 (.fluid_in(k_11_108), .fluid_out(k_10_54), .air_in(c_11_0));
valve v_11_109 (.fluid_in(k_11_109), .fluid_out(k_10_54), .air_in(c_11_1));
valve v_11_110 (.fluid_in(k_11_110), .fluid_out(k_10_55), .air_in(c_11_0));
valve v_11_111 (.fluid_in(k_11_111), .fluid_out(k_10_55), .air_in(c_11_1));
valve v_11_112 (.fluid_in(k_11_112), .fluid_out(k_10_56), .air_in(c_11_0));
valve v_11_113 (.fluid_in(k_11_113), .fluid_out(k_10_56), .air_in(c_11_1));
valve v_11_114 (.fluid_in(k_11_114), .fluid_out(k_10_57), .air_in(c_11_0));
valve v_11_115 (.fluid_in(k_11_115), .fluid_out(k_10_57), .air_in(c_11_1));
valve v_11_116 (.fluid_in(k_11_116), .fluid_out(k_10_58), .air_in(c_11_0));
valve v_11_117 (.fluid_in(k_11_117), .fluid_out(k_10_58), .air_in(c_11_1));
valve v_11_118 (.fluid_in(k_11_118), .fluid_out(k_10_59), .air_in(c_11_0));
valve v_11_119 (.fluid_in(k_11_119), .fluid_out(k_10_59), .air_in(c_11_1));
valve v_11_120 (.fluid_in(k_11_120), .fluid_out(k_10_60), .air_in(c_11_0));
valve v_11_121 (.fluid_in(k_11_121), .fluid_out(k_10_60), .air_in(c_11_1));
valve v_11_122 (.fluid_in(k_11_122), .fluid_out(k_10_61), .air_in(c_11_0));
valve v_11_123 (.fluid_in(k_11_123), .fluid_out(k_10_61), .air_in(c_11_1));
valve v_11_124 (.fluid_in(k_11_124), .fluid_out(k_10_62), .air_in(c_11_0));
valve v_11_125 (.fluid_in(k_11_125), .fluid_out(k_10_62), .air_in(c_11_1));
valve v_11_126 (.fluid_in(k_11_126), .fluid_out(k_10_63), .air_in(c_11_0));
valve v_11_127 (.fluid_in(k_11_127), .fluid_out(k_10_63), .air_in(c_11_1));
valve v_11_128 (.fluid_in(k_11_128), .fluid_out(k_10_64), .air_in(c_11_0));
valve v_11_129 (.fluid_in(k_11_129), .fluid_out(k_10_64), .air_in(c_11_1));
valve v_11_130 (.fluid_in(k_11_130), .fluid_out(k_10_65), .air_in(c_11_0));
valve v_11_131 (.fluid_in(k_11_131), .fluid_out(k_10_65), .air_in(c_11_1));
valve v_11_132 (.fluid_in(k_11_132), .fluid_out(k_10_66), .air_in(c_11_0));
valve v_11_133 (.fluid_in(k_11_133), .fluid_out(k_10_66), .air_in(c_11_1));
valve v_11_134 (.fluid_in(k_11_134), .fluid_out(k_10_67), .air_in(c_11_0));
valve v_11_135 (.fluid_in(k_11_135), .fluid_out(k_10_67), .air_in(c_11_1));
valve v_11_136 (.fluid_in(k_11_136), .fluid_out(k_10_68), .air_in(c_11_0));
valve v_11_137 (.fluid_in(k_11_137), .fluid_out(k_10_68), .air_in(c_11_1));
valve v_11_138 (.fluid_in(k_11_138), .fluid_out(k_10_69), .air_in(c_11_0));
valve v_11_139 (.fluid_in(k_11_139), .fluid_out(k_10_69), .air_in(c_11_1));
valve v_11_140 (.fluid_in(k_11_140), .fluid_out(k_10_70), .air_in(c_11_0));
valve v_11_141 (.fluid_in(k_11_141), .fluid_out(k_10_70), .air_in(c_11_1));
valve v_11_142 (.fluid_in(k_11_142), .fluid_out(k_10_71), .air_in(c_11_0));
valve v_11_143 (.fluid_in(k_11_143), .fluid_out(k_10_71), .air_in(c_11_1));
valve v_11_144 (.fluid_in(k_11_144), .fluid_out(k_10_72), .air_in(c_11_0));
valve v_11_145 (.fluid_in(k_11_145), .fluid_out(k_10_72), .air_in(c_11_1));
valve v_11_146 (.fluid_in(k_11_146), .fluid_out(k_10_73), .air_in(c_11_0));
valve v_11_147 (.fluid_in(k_11_147), .fluid_out(k_10_73), .air_in(c_11_1));
valve v_11_148 (.fluid_in(k_11_148), .fluid_out(k_10_74), .air_in(c_11_0));
valve v_11_149 (.fluid_in(k_11_149), .fluid_out(k_10_74), .air_in(c_11_1));
valve v_11_150 (.fluid_in(k_11_150), .fluid_out(k_10_75), .air_in(c_11_0));
valve v_11_151 (.fluid_in(k_11_151), .fluid_out(k_10_75), .air_in(c_11_1));
valve v_11_152 (.fluid_in(k_11_152), .fluid_out(k_10_76), .air_in(c_11_0));
valve v_11_153 (.fluid_in(k_11_153), .fluid_out(k_10_76), .air_in(c_11_1));
valve v_11_154 (.fluid_in(k_11_154), .fluid_out(k_10_77), .air_in(c_11_0));
valve v_11_155 (.fluid_in(k_11_155), .fluid_out(k_10_77), .air_in(c_11_1));
valve v_11_156 (.fluid_in(k_11_156), .fluid_out(k_10_78), .air_in(c_11_0));
valve v_11_157 (.fluid_in(k_11_157), .fluid_out(k_10_78), .air_in(c_11_1));
valve v_11_158 (.fluid_in(k_11_158), .fluid_out(k_10_79), .air_in(c_11_0));
valve v_11_159 (.fluid_in(k_11_159), .fluid_out(k_10_79), .air_in(c_11_1));
valve v_11_160 (.fluid_in(k_11_160), .fluid_out(k_10_80), .air_in(c_11_0));
valve v_11_161 (.fluid_in(k_11_161), .fluid_out(k_10_80), .air_in(c_11_1));
valve v_11_162 (.fluid_in(k_11_162), .fluid_out(k_10_81), .air_in(c_11_0));
valve v_11_163 (.fluid_in(k_11_163), .fluid_out(k_10_81), .air_in(c_11_1));
valve v_11_164 (.fluid_in(k_11_164), .fluid_out(k_10_82), .air_in(c_11_0));
valve v_11_165 (.fluid_in(k_11_165), .fluid_out(k_10_82), .air_in(c_11_1));
valve v_11_166 (.fluid_in(k_11_166), .fluid_out(k_10_83), .air_in(c_11_0));
valve v_11_167 (.fluid_in(k_11_167), .fluid_out(k_10_83), .air_in(c_11_1));
valve v_11_168 (.fluid_in(k_11_168), .fluid_out(k_10_84), .air_in(c_11_0));
valve v_11_169 (.fluid_in(k_11_169), .fluid_out(k_10_84), .air_in(c_11_1));
valve v_11_170 (.fluid_in(k_11_170), .fluid_out(k_10_85), .air_in(c_11_0));
valve v_11_171 (.fluid_in(k_11_171), .fluid_out(k_10_85), .air_in(c_11_1));
valve v_11_172 (.fluid_in(k_11_172), .fluid_out(k_10_86), .air_in(c_11_0));
valve v_11_173 (.fluid_in(k_11_173), .fluid_out(k_10_86), .air_in(c_11_1));
valve v_11_174 (.fluid_in(k_11_174), .fluid_out(k_10_87), .air_in(c_11_0));
valve v_11_175 (.fluid_in(k_11_175), .fluid_out(k_10_87), .air_in(c_11_1));
valve v_11_176 (.fluid_in(k_11_176), .fluid_out(k_10_88), .air_in(c_11_0));
valve v_11_177 (.fluid_in(k_11_177), .fluid_out(k_10_88), .air_in(c_11_1));
valve v_11_178 (.fluid_in(k_11_178), .fluid_out(k_10_89), .air_in(c_11_0));
valve v_11_179 (.fluid_in(k_11_179), .fluid_out(k_10_89), .air_in(c_11_1));
valve v_11_180 (.fluid_in(k_11_180), .fluid_out(k_10_90), .air_in(c_11_0));
valve v_11_181 (.fluid_in(k_11_181), .fluid_out(k_10_90), .air_in(c_11_1));
valve v_11_182 (.fluid_in(k_11_182), .fluid_out(k_10_91), .air_in(c_11_0));
valve v_11_183 (.fluid_in(k_11_183), .fluid_out(k_10_91), .air_in(c_11_1));
valve v_11_184 (.fluid_in(k_11_184), .fluid_out(k_10_92), .air_in(c_11_0));
valve v_11_185 (.fluid_in(k_11_185), .fluid_out(k_10_92), .air_in(c_11_1));
valve v_11_186 (.fluid_in(k_11_186), .fluid_out(k_10_93), .air_in(c_11_0));
valve v_11_187 (.fluid_in(k_11_187), .fluid_out(k_10_93), .air_in(c_11_1));
valve v_11_188 (.fluid_in(k_11_188), .fluid_out(k_10_94), .air_in(c_11_0));
valve v_11_189 (.fluid_in(k_11_189), .fluid_out(k_10_94), .air_in(c_11_1));
valve v_11_190 (.fluid_in(k_11_190), .fluid_out(k_10_95), .air_in(c_11_0));
valve v_11_191 (.fluid_in(k_11_191), .fluid_out(k_10_95), .air_in(c_11_1));
valve v_11_192 (.fluid_in(k_11_192), .fluid_out(k_10_96), .air_in(c_11_0));
valve v_11_193 (.fluid_in(k_11_193), .fluid_out(k_10_96), .air_in(c_11_1));
valve v_11_194 (.fluid_in(k_11_194), .fluid_out(k_10_97), .air_in(c_11_0));
valve v_11_195 (.fluid_in(k_11_195), .fluid_out(k_10_97), .air_in(c_11_1));
valve v_11_196 (.fluid_in(k_11_196), .fluid_out(k_10_98), .air_in(c_11_0));
valve v_11_197 (.fluid_in(k_11_197), .fluid_out(k_10_98), .air_in(c_11_1));
valve v_11_198 (.fluid_in(k_11_198), .fluid_out(k_10_99), .air_in(c_11_0));
valve v_11_199 (.fluid_in(k_11_199), .fluid_out(k_10_99), .air_in(c_11_1));
valve v_11_200 (.fluid_in(k_11_200), .fluid_out(k_10_100), .air_in(c_11_0));
valve v_11_201 (.fluid_in(k_11_201), .fluid_out(k_10_100), .air_in(c_11_1));
valve v_11_202 (.fluid_in(k_11_202), .fluid_out(k_10_101), .air_in(c_11_0));
valve v_11_203 (.fluid_in(k_11_203), .fluid_out(k_10_101), .air_in(c_11_1));
valve v_11_204 (.fluid_in(k_11_204), .fluid_out(k_10_102), .air_in(c_11_0));
valve v_11_205 (.fluid_in(k_11_205), .fluid_out(k_10_102), .air_in(c_11_1));
valve v_11_206 (.fluid_in(k_11_206), .fluid_out(k_10_103), .air_in(c_11_0));
valve v_11_207 (.fluid_in(k_11_207), .fluid_out(k_10_103), .air_in(c_11_1));
valve v_11_208 (.fluid_in(k_11_208), .fluid_out(k_10_104), .air_in(c_11_0));
valve v_11_209 (.fluid_in(k_11_209), .fluid_out(k_10_104), .air_in(c_11_1));
valve v_11_210 (.fluid_in(k_11_210), .fluid_out(k_10_105), .air_in(c_11_0));
valve v_11_211 (.fluid_in(k_11_211), .fluid_out(k_10_105), .air_in(c_11_1));
valve v_11_212 (.fluid_in(k_11_212), .fluid_out(k_10_106), .air_in(c_11_0));
valve v_11_213 (.fluid_in(k_11_213), .fluid_out(k_10_106), .air_in(c_11_1));
valve v_11_214 (.fluid_in(k_11_214), .fluid_out(k_10_107), .air_in(c_11_0));
valve v_11_215 (.fluid_in(k_11_215), .fluid_out(k_10_107), .air_in(c_11_1));
valve v_11_216 (.fluid_in(k_11_216), .fluid_out(k_10_108), .air_in(c_11_0));
valve v_11_217 (.fluid_in(k_11_217), .fluid_out(k_10_108), .air_in(c_11_1));
valve v_11_218 (.fluid_in(k_11_218), .fluid_out(k_10_109), .air_in(c_11_0));
valve v_11_219 (.fluid_in(k_11_219), .fluid_out(k_10_109), .air_in(c_11_1));
valve v_11_220 (.fluid_in(k_11_220), .fluid_out(k_10_110), .air_in(c_11_0));
valve v_11_221 (.fluid_in(k_11_221), .fluid_out(k_10_110), .air_in(c_11_1));
valve v_11_222 (.fluid_in(k_11_222), .fluid_out(k_10_111), .air_in(c_11_0));
valve v_11_223 (.fluid_in(k_11_223), .fluid_out(k_10_111), .air_in(c_11_1));
valve v_11_224 (.fluid_in(k_11_224), .fluid_out(k_10_112), .air_in(c_11_0));
valve v_11_225 (.fluid_in(k_11_225), .fluid_out(k_10_112), .air_in(c_11_1));
valve v_11_226 (.fluid_in(k_11_226), .fluid_out(k_10_113), .air_in(c_11_0));
valve v_11_227 (.fluid_in(k_11_227), .fluid_out(k_10_113), .air_in(c_11_1));
valve v_11_228 (.fluid_in(k_11_228), .fluid_out(k_10_114), .air_in(c_11_0));
valve v_11_229 (.fluid_in(k_11_229), .fluid_out(k_10_114), .air_in(c_11_1));
valve v_11_230 (.fluid_in(k_11_230), .fluid_out(k_10_115), .air_in(c_11_0));
valve v_11_231 (.fluid_in(k_11_231), .fluid_out(k_10_115), .air_in(c_11_1));
valve v_11_232 (.fluid_in(k_11_232), .fluid_out(k_10_116), .air_in(c_11_0));
valve v_11_233 (.fluid_in(k_11_233), .fluid_out(k_10_116), .air_in(c_11_1));
valve v_11_234 (.fluid_in(k_11_234), .fluid_out(k_10_117), .air_in(c_11_0));
valve v_11_235 (.fluid_in(k_11_235), .fluid_out(k_10_117), .air_in(c_11_1));
valve v_11_236 (.fluid_in(k_11_236), .fluid_out(k_10_118), .air_in(c_11_0));
valve v_11_237 (.fluid_in(k_11_237), .fluid_out(k_10_118), .air_in(c_11_1));
valve v_11_238 (.fluid_in(k_11_238), .fluid_out(k_10_119), .air_in(c_11_0));
valve v_11_239 (.fluid_in(k_11_239), .fluid_out(k_10_119), .air_in(c_11_1));
valve v_11_240 (.fluid_in(k_11_240), .fluid_out(k_10_120), .air_in(c_11_0));
valve v_11_241 (.fluid_in(k_11_241), .fluid_out(k_10_120), .air_in(c_11_1));
valve v_11_242 (.fluid_in(k_11_242), .fluid_out(k_10_121), .air_in(c_11_0));
valve v_11_243 (.fluid_in(k_11_243), .fluid_out(k_10_121), .air_in(c_11_1));
valve v_11_244 (.fluid_in(k_11_244), .fluid_out(k_10_122), .air_in(c_11_0));
valve v_11_245 (.fluid_in(k_11_245), .fluid_out(k_10_122), .air_in(c_11_1));
valve v_11_246 (.fluid_in(k_11_246), .fluid_out(k_10_123), .air_in(c_11_0));
valve v_11_247 (.fluid_in(k_11_247), .fluid_out(k_10_123), .air_in(c_11_1));
valve v_11_248 (.fluid_in(k_11_248), .fluid_out(k_10_124), .air_in(c_11_0));
valve v_11_249 (.fluid_in(k_11_249), .fluid_out(k_10_124), .air_in(c_11_1));
valve v_11_250 (.fluid_in(k_11_250), .fluid_out(k_10_125), .air_in(c_11_0));
valve v_11_251 (.fluid_in(k_11_251), .fluid_out(k_10_125), .air_in(c_11_1));
valve v_11_252 (.fluid_in(k_11_252), .fluid_out(k_10_126), .air_in(c_11_0));
valve v_11_253 (.fluid_in(k_11_253), .fluid_out(k_10_126), .air_in(c_11_1));
valve v_11_254 (.fluid_in(k_11_254), .fluid_out(k_10_127), .air_in(c_11_0));
valve v_11_255 (.fluid_in(k_11_255), .fluid_out(k_10_127), .air_in(c_11_1));
valve v_11_256 (.fluid_in(k_11_256), .fluid_out(k_10_128), .air_in(c_11_0));
valve v_11_257 (.fluid_in(k_11_257), .fluid_out(k_10_128), .air_in(c_11_1));
valve v_11_258 (.fluid_in(k_11_258), .fluid_out(k_10_129), .air_in(c_11_0));
valve v_11_259 (.fluid_in(k_11_259), .fluid_out(k_10_129), .air_in(c_11_1));
valve v_11_260 (.fluid_in(k_11_260), .fluid_out(k_10_130), .air_in(c_11_0));
valve v_11_261 (.fluid_in(k_11_261), .fluid_out(k_10_130), .air_in(c_11_1));
valve v_11_262 (.fluid_in(k_11_262), .fluid_out(k_10_131), .air_in(c_11_0));
valve v_11_263 (.fluid_in(k_11_263), .fluid_out(k_10_131), .air_in(c_11_1));
valve v_11_264 (.fluid_in(k_11_264), .fluid_out(k_10_132), .air_in(c_11_0));
valve v_11_265 (.fluid_in(k_11_265), .fluid_out(k_10_132), .air_in(c_11_1));
valve v_11_266 (.fluid_in(k_11_266), .fluid_out(k_10_133), .air_in(c_11_0));
valve v_11_267 (.fluid_in(k_11_267), .fluid_out(k_10_133), .air_in(c_11_1));
valve v_11_268 (.fluid_in(k_11_268), .fluid_out(k_10_134), .air_in(c_11_0));
valve v_11_269 (.fluid_in(k_11_269), .fluid_out(k_10_134), .air_in(c_11_1));
valve v_11_270 (.fluid_in(k_11_270), .fluid_out(k_10_135), .air_in(c_11_0));
valve v_11_271 (.fluid_in(k_11_271), .fluid_out(k_10_135), .air_in(c_11_1));
valve v_11_272 (.fluid_in(k_11_272), .fluid_out(k_10_136), .air_in(c_11_0));
valve v_11_273 (.fluid_in(k_11_273), .fluid_out(k_10_136), .air_in(c_11_1));
valve v_11_274 (.fluid_in(k_11_274), .fluid_out(k_10_137), .air_in(c_11_0));
valve v_11_275 (.fluid_in(k_11_275), .fluid_out(k_10_137), .air_in(c_11_1));
valve v_11_276 (.fluid_in(k_11_276), .fluid_out(k_10_138), .air_in(c_11_0));
valve v_11_277 (.fluid_in(k_11_277), .fluid_out(k_10_138), .air_in(c_11_1));
valve v_11_278 (.fluid_in(k_11_278), .fluid_out(k_10_139), .air_in(c_11_0));
valve v_11_279 (.fluid_in(k_11_279), .fluid_out(k_10_139), .air_in(c_11_1));
valve v_11_280 (.fluid_in(k_11_280), .fluid_out(k_10_140), .air_in(c_11_0));
valve v_11_281 (.fluid_in(k_11_281), .fluid_out(k_10_140), .air_in(c_11_1));
valve v_11_282 (.fluid_in(k_11_282), .fluid_out(k_10_141), .air_in(c_11_0));
valve v_11_283 (.fluid_in(k_11_283), .fluid_out(k_10_141), .air_in(c_11_1));
valve v_11_284 (.fluid_in(k_11_284), .fluid_out(k_10_142), .air_in(c_11_0));
valve v_11_285 (.fluid_in(k_11_285), .fluid_out(k_10_142), .air_in(c_11_1));
valve v_11_286 (.fluid_in(k_11_286), .fluid_out(k_10_143), .air_in(c_11_0));
valve v_11_287 (.fluid_in(k_11_287), .fluid_out(k_10_143), .air_in(c_11_1));
valve v_11_288 (.fluid_in(k_11_288), .fluid_out(k_10_144), .air_in(c_11_0));
valve v_11_289 (.fluid_in(k_11_289), .fluid_out(k_10_144), .air_in(c_11_1));
valve v_11_290 (.fluid_in(k_11_290), .fluid_out(k_10_145), .air_in(c_11_0));
valve v_11_291 (.fluid_in(k_11_291), .fluid_out(k_10_145), .air_in(c_11_1));
valve v_11_292 (.fluid_in(k_11_292), .fluid_out(k_10_146), .air_in(c_11_0));
valve v_11_293 (.fluid_in(k_11_293), .fluid_out(k_10_146), .air_in(c_11_1));
valve v_11_294 (.fluid_in(k_11_294), .fluid_out(k_10_147), .air_in(c_11_0));
valve v_11_295 (.fluid_in(k_11_295), .fluid_out(k_10_147), .air_in(c_11_1));
valve v_11_296 (.fluid_in(k_11_296), .fluid_out(k_10_148), .air_in(c_11_0));
valve v_11_297 (.fluid_in(k_11_297), .fluid_out(k_10_148), .air_in(c_11_1));
valve v_11_298 (.fluid_in(k_11_298), .fluid_out(k_10_149), .air_in(c_11_0));
valve v_11_299 (.fluid_in(k_11_299), .fluid_out(k_10_149), .air_in(c_11_1));
valve v_11_300 (.fluid_in(k_11_300), .fluid_out(k_10_150), .air_in(c_11_0));
valve v_11_301 (.fluid_in(k_11_301), .fluid_out(k_10_150), .air_in(c_11_1));
valve v_11_302 (.fluid_in(k_11_302), .fluid_out(k_10_151), .air_in(c_11_0));
valve v_11_303 (.fluid_in(k_11_303), .fluid_out(k_10_151), .air_in(c_11_1));
valve v_11_304 (.fluid_in(k_11_304), .fluid_out(k_10_152), .air_in(c_11_0));
valve v_11_305 (.fluid_in(k_11_305), .fluid_out(k_10_152), .air_in(c_11_1));
valve v_11_306 (.fluid_in(k_11_306), .fluid_out(k_10_153), .air_in(c_11_0));
valve v_11_307 (.fluid_in(k_11_307), .fluid_out(k_10_153), .air_in(c_11_1));
valve v_11_308 (.fluid_in(k_11_308), .fluid_out(k_10_154), .air_in(c_11_0));
valve v_11_309 (.fluid_in(k_11_309), .fluid_out(k_10_154), .air_in(c_11_1));
valve v_11_310 (.fluid_in(k_11_310), .fluid_out(k_10_155), .air_in(c_11_0));
valve v_11_311 (.fluid_in(k_11_311), .fluid_out(k_10_155), .air_in(c_11_1));
valve v_11_312 (.fluid_in(k_11_312), .fluid_out(k_10_156), .air_in(c_11_0));
valve v_11_313 (.fluid_in(k_11_313), .fluid_out(k_10_156), .air_in(c_11_1));
valve v_11_314 (.fluid_in(k_11_314), .fluid_out(k_10_157), .air_in(c_11_0));
valve v_11_315 (.fluid_in(k_11_315), .fluid_out(k_10_157), .air_in(c_11_1));
valve v_11_316 (.fluid_in(k_11_316), .fluid_out(k_10_158), .air_in(c_11_0));
valve v_11_317 (.fluid_in(k_11_317), .fluid_out(k_10_158), .air_in(c_11_1));
valve v_11_318 (.fluid_in(k_11_318), .fluid_out(k_10_159), .air_in(c_11_0));
valve v_11_319 (.fluid_in(k_11_319), .fluid_out(k_10_159), .air_in(c_11_1));
valve v_11_320 (.fluid_in(k_11_320), .fluid_out(k_10_160), .air_in(c_11_0));
valve v_11_321 (.fluid_in(k_11_321), .fluid_out(k_10_160), .air_in(c_11_1));
valve v_11_322 (.fluid_in(k_11_322), .fluid_out(k_10_161), .air_in(c_11_0));
valve v_11_323 (.fluid_in(k_11_323), .fluid_out(k_10_161), .air_in(c_11_1));
valve v_11_324 (.fluid_in(k_11_324), .fluid_out(k_10_162), .air_in(c_11_0));
valve v_11_325 (.fluid_in(k_11_325), .fluid_out(k_10_162), .air_in(c_11_1));
valve v_11_326 (.fluid_in(k_11_326), .fluid_out(k_10_163), .air_in(c_11_0));
valve v_11_327 (.fluid_in(k_11_327), .fluid_out(k_10_163), .air_in(c_11_1));
valve v_11_328 (.fluid_in(k_11_328), .fluid_out(k_10_164), .air_in(c_11_0));
valve v_11_329 (.fluid_in(k_11_329), .fluid_out(k_10_164), .air_in(c_11_1));
valve v_11_330 (.fluid_in(k_11_330), .fluid_out(k_10_165), .air_in(c_11_0));
valve v_11_331 (.fluid_in(k_11_331), .fluid_out(k_10_165), .air_in(c_11_1));
valve v_11_332 (.fluid_in(k_11_332), .fluid_out(k_10_166), .air_in(c_11_0));
valve v_11_333 (.fluid_in(k_11_333), .fluid_out(k_10_166), .air_in(c_11_1));
valve v_11_334 (.fluid_in(k_11_334), .fluid_out(k_10_167), .air_in(c_11_0));
valve v_11_335 (.fluid_in(k_11_335), .fluid_out(k_10_167), .air_in(c_11_1));
valve v_11_336 (.fluid_in(k_11_336), .fluid_out(k_10_168), .air_in(c_11_0));
valve v_11_337 (.fluid_in(k_11_337), .fluid_out(k_10_168), .air_in(c_11_1));
valve v_11_338 (.fluid_in(k_11_338), .fluid_out(k_10_169), .air_in(c_11_0));
valve v_11_339 (.fluid_in(k_11_339), .fluid_out(k_10_169), .air_in(c_11_1));
valve v_11_340 (.fluid_in(k_11_340), .fluid_out(k_10_170), .air_in(c_11_0));
valve v_11_341 (.fluid_in(k_11_341), .fluid_out(k_10_170), .air_in(c_11_1));
valve v_11_342 (.fluid_in(k_11_342), .fluid_out(k_10_171), .air_in(c_11_0));
valve v_11_343 (.fluid_in(k_11_343), .fluid_out(k_10_171), .air_in(c_11_1));
valve v_11_344 (.fluid_in(k_11_344), .fluid_out(k_10_172), .air_in(c_11_0));
valve v_11_345 (.fluid_in(k_11_345), .fluid_out(k_10_172), .air_in(c_11_1));
valve v_11_346 (.fluid_in(k_11_346), .fluid_out(k_10_173), .air_in(c_11_0));
valve v_11_347 (.fluid_in(k_11_347), .fluid_out(k_10_173), .air_in(c_11_1));
valve v_11_348 (.fluid_in(k_11_348), .fluid_out(k_10_174), .air_in(c_11_0));
valve v_11_349 (.fluid_in(k_11_349), .fluid_out(k_10_174), .air_in(c_11_1));
valve v_11_350 (.fluid_in(k_11_350), .fluid_out(k_10_175), .air_in(c_11_0));
valve v_11_351 (.fluid_in(k_11_351), .fluid_out(k_10_175), .air_in(c_11_1));
valve v_11_352 (.fluid_in(k_11_352), .fluid_out(k_10_176), .air_in(c_11_0));
valve v_11_353 (.fluid_in(k_11_353), .fluid_out(k_10_176), .air_in(c_11_1));
valve v_11_354 (.fluid_in(k_11_354), .fluid_out(k_10_177), .air_in(c_11_0));
valve v_11_355 (.fluid_in(k_11_355), .fluid_out(k_10_177), .air_in(c_11_1));
valve v_11_356 (.fluid_in(k_11_356), .fluid_out(k_10_178), .air_in(c_11_0));
valve v_11_357 (.fluid_in(k_11_357), .fluid_out(k_10_178), .air_in(c_11_1));
valve v_11_358 (.fluid_in(k_11_358), .fluid_out(k_10_179), .air_in(c_11_0));
valve v_11_359 (.fluid_in(k_11_359), .fluid_out(k_10_179), .air_in(c_11_1));
valve v_11_360 (.fluid_in(k_11_360), .fluid_out(k_10_180), .air_in(c_11_0));
valve v_11_361 (.fluid_in(k_11_361), .fluid_out(k_10_180), .air_in(c_11_1));
valve v_11_362 (.fluid_in(k_11_362), .fluid_out(k_10_181), .air_in(c_11_0));
valve v_11_363 (.fluid_in(k_11_363), .fluid_out(k_10_181), .air_in(c_11_1));
valve v_11_364 (.fluid_in(k_11_364), .fluid_out(k_10_182), .air_in(c_11_0));
valve v_11_365 (.fluid_in(k_11_365), .fluid_out(k_10_182), .air_in(c_11_1));
valve v_11_366 (.fluid_in(k_11_366), .fluid_out(k_10_183), .air_in(c_11_0));
valve v_11_367 (.fluid_in(k_11_367), .fluid_out(k_10_183), .air_in(c_11_1));
valve v_11_368 (.fluid_in(k_11_368), .fluid_out(k_10_184), .air_in(c_11_0));
valve v_11_369 (.fluid_in(k_11_369), .fluid_out(k_10_184), .air_in(c_11_1));
valve v_11_370 (.fluid_in(k_11_370), .fluid_out(k_10_185), .air_in(c_11_0));
valve v_11_371 (.fluid_in(k_11_371), .fluid_out(k_10_185), .air_in(c_11_1));
valve v_11_372 (.fluid_in(k_11_372), .fluid_out(k_10_186), .air_in(c_11_0));
valve v_11_373 (.fluid_in(k_11_373), .fluid_out(k_10_186), .air_in(c_11_1));
valve v_11_374 (.fluid_in(k_11_374), .fluid_out(k_10_187), .air_in(c_11_0));
valve v_11_375 (.fluid_in(k_11_375), .fluid_out(k_10_187), .air_in(c_11_1));
valve v_11_376 (.fluid_in(k_11_376), .fluid_out(k_10_188), .air_in(c_11_0));
valve v_11_377 (.fluid_in(k_11_377), .fluid_out(k_10_188), .air_in(c_11_1));
valve v_11_378 (.fluid_in(k_11_378), .fluid_out(k_10_189), .air_in(c_11_0));
valve v_11_379 (.fluid_in(k_11_379), .fluid_out(k_10_189), .air_in(c_11_1));
valve v_11_380 (.fluid_in(k_11_380), .fluid_out(k_10_190), .air_in(c_11_0));
valve v_11_381 (.fluid_in(k_11_381), .fluid_out(k_10_190), .air_in(c_11_1));
valve v_11_382 (.fluid_in(k_11_382), .fluid_out(k_10_191), .air_in(c_11_0));
valve v_11_383 (.fluid_in(k_11_383), .fluid_out(k_10_191), .air_in(c_11_1));
valve v_11_384 (.fluid_in(k_11_384), .fluid_out(k_10_192), .air_in(c_11_0));
valve v_11_385 (.fluid_in(k_11_385), .fluid_out(k_10_192), .air_in(c_11_1));
valve v_11_386 (.fluid_in(k_11_386), .fluid_out(k_10_193), .air_in(c_11_0));
valve v_11_387 (.fluid_in(k_11_387), .fluid_out(k_10_193), .air_in(c_11_1));
valve v_11_388 (.fluid_in(k_11_388), .fluid_out(k_10_194), .air_in(c_11_0));
valve v_11_389 (.fluid_in(k_11_389), .fluid_out(k_10_194), .air_in(c_11_1));
valve v_11_390 (.fluid_in(k_11_390), .fluid_out(k_10_195), .air_in(c_11_0));
valve v_11_391 (.fluid_in(k_11_391), .fluid_out(k_10_195), .air_in(c_11_1));
valve v_11_392 (.fluid_in(k_11_392), .fluid_out(k_10_196), .air_in(c_11_0));
valve v_11_393 (.fluid_in(k_11_393), .fluid_out(k_10_196), .air_in(c_11_1));
valve v_11_394 (.fluid_in(k_11_394), .fluid_out(k_10_197), .air_in(c_11_0));
valve v_11_395 (.fluid_in(k_11_395), .fluid_out(k_10_197), .air_in(c_11_1));
valve v_11_396 (.fluid_in(k_11_396), .fluid_out(k_10_198), .air_in(c_11_0));
valve v_11_397 (.fluid_in(k_11_397), .fluid_out(k_10_198), .air_in(c_11_1));
valve v_11_398 (.fluid_in(k_11_398), .fluid_out(k_10_199), .air_in(c_11_0));
valve v_11_399 (.fluid_in(k_11_399), .fluid_out(k_10_199), .air_in(c_11_1));
valve v_11_400 (.fluid_in(k_11_400), .fluid_out(k_10_200), .air_in(c_11_0));
valve v_11_401 (.fluid_in(k_11_401), .fluid_out(k_10_200), .air_in(c_11_1));
valve v_11_402 (.fluid_in(k_11_402), .fluid_out(k_10_201), .air_in(c_11_0));
valve v_11_403 (.fluid_in(k_11_403), .fluid_out(k_10_201), .air_in(c_11_1));
valve v_11_404 (.fluid_in(k_11_404), .fluid_out(k_10_202), .air_in(c_11_0));
valve v_11_405 (.fluid_in(k_11_405), .fluid_out(k_10_202), .air_in(c_11_1));
valve v_11_406 (.fluid_in(k_11_406), .fluid_out(k_10_203), .air_in(c_11_0));
valve v_11_407 (.fluid_in(k_11_407), .fluid_out(k_10_203), .air_in(c_11_1));
valve v_11_408 (.fluid_in(k_11_408), .fluid_out(k_10_204), .air_in(c_11_0));
valve v_11_409 (.fluid_in(k_11_409), .fluid_out(k_10_204), .air_in(c_11_1));
valve v_11_410 (.fluid_in(k_11_410), .fluid_out(k_10_205), .air_in(c_11_0));
valve v_11_411 (.fluid_in(k_11_411), .fluid_out(k_10_205), .air_in(c_11_1));
valve v_11_412 (.fluid_in(k_11_412), .fluid_out(k_10_206), .air_in(c_11_0));
valve v_11_413 (.fluid_in(k_11_413), .fluid_out(k_10_206), .air_in(c_11_1));
valve v_11_414 (.fluid_in(k_11_414), .fluid_out(k_10_207), .air_in(c_11_0));
valve v_11_415 (.fluid_in(k_11_415), .fluid_out(k_10_207), .air_in(c_11_1));
valve v_11_416 (.fluid_in(k_11_416), .fluid_out(k_10_208), .air_in(c_11_0));
valve v_11_417 (.fluid_in(k_11_417), .fluid_out(k_10_208), .air_in(c_11_1));
valve v_11_418 (.fluid_in(k_11_418), .fluid_out(k_10_209), .air_in(c_11_0));
valve v_11_419 (.fluid_in(k_11_419), .fluid_out(k_10_209), .air_in(c_11_1));
valve v_11_420 (.fluid_in(k_11_420), .fluid_out(k_10_210), .air_in(c_11_0));
valve v_11_421 (.fluid_in(k_11_421), .fluid_out(k_10_210), .air_in(c_11_1));
valve v_11_422 (.fluid_in(k_11_422), .fluid_out(k_10_211), .air_in(c_11_0));
valve v_11_423 (.fluid_in(k_11_423), .fluid_out(k_10_211), .air_in(c_11_1));
valve v_11_424 (.fluid_in(k_11_424), .fluid_out(k_10_212), .air_in(c_11_0));
valve v_11_425 (.fluid_in(k_11_425), .fluid_out(k_10_212), .air_in(c_11_1));
valve v_11_426 (.fluid_in(k_11_426), .fluid_out(k_10_213), .air_in(c_11_0));
valve v_11_427 (.fluid_in(k_11_427), .fluid_out(k_10_213), .air_in(c_11_1));
valve v_11_428 (.fluid_in(k_11_428), .fluid_out(k_10_214), .air_in(c_11_0));
valve v_11_429 (.fluid_in(k_11_429), .fluid_out(k_10_214), .air_in(c_11_1));
valve v_11_430 (.fluid_in(k_11_430), .fluid_out(k_10_215), .air_in(c_11_0));
valve v_11_431 (.fluid_in(k_11_431), .fluid_out(k_10_215), .air_in(c_11_1));
valve v_11_432 (.fluid_in(k_11_432), .fluid_out(k_10_216), .air_in(c_11_0));
valve v_11_433 (.fluid_in(k_11_433), .fluid_out(k_10_216), .air_in(c_11_1));
valve v_11_434 (.fluid_in(k_11_434), .fluid_out(k_10_217), .air_in(c_11_0));
valve v_11_435 (.fluid_in(k_11_435), .fluid_out(k_10_217), .air_in(c_11_1));
valve v_11_436 (.fluid_in(k_11_436), .fluid_out(k_10_218), .air_in(c_11_0));
valve v_11_437 (.fluid_in(k_11_437), .fluid_out(k_10_218), .air_in(c_11_1));
valve v_11_438 (.fluid_in(k_11_438), .fluid_out(k_10_219), .air_in(c_11_0));
valve v_11_439 (.fluid_in(k_11_439), .fluid_out(k_10_219), .air_in(c_11_1));
valve v_11_440 (.fluid_in(k_11_440), .fluid_out(k_10_220), .air_in(c_11_0));
valve v_11_441 (.fluid_in(k_11_441), .fluid_out(k_10_220), .air_in(c_11_1));
valve v_11_442 (.fluid_in(k_11_442), .fluid_out(k_10_221), .air_in(c_11_0));
valve v_11_443 (.fluid_in(k_11_443), .fluid_out(k_10_221), .air_in(c_11_1));
valve v_11_444 (.fluid_in(k_11_444), .fluid_out(k_10_222), .air_in(c_11_0));
valve v_11_445 (.fluid_in(k_11_445), .fluid_out(k_10_222), .air_in(c_11_1));
valve v_11_446 (.fluid_in(k_11_446), .fluid_out(k_10_223), .air_in(c_11_0));
valve v_11_447 (.fluid_in(k_11_447), .fluid_out(k_10_223), .air_in(c_11_1));
valve v_11_448 (.fluid_in(k_11_448), .fluid_out(k_10_224), .air_in(c_11_0));
valve v_11_449 (.fluid_in(k_11_449), .fluid_out(k_10_224), .air_in(c_11_1));
valve v_11_450 (.fluid_in(k_11_450), .fluid_out(k_10_225), .air_in(c_11_0));
valve v_11_451 (.fluid_in(k_11_451), .fluid_out(k_10_225), .air_in(c_11_1));
valve v_11_452 (.fluid_in(k_11_452), .fluid_out(k_10_226), .air_in(c_11_0));
valve v_11_453 (.fluid_in(k_11_453), .fluid_out(k_10_226), .air_in(c_11_1));
valve v_11_454 (.fluid_in(k_11_454), .fluid_out(k_10_227), .air_in(c_11_0));
valve v_11_455 (.fluid_in(k_11_455), .fluid_out(k_10_227), .air_in(c_11_1));
valve v_11_456 (.fluid_in(k_11_456), .fluid_out(k_10_228), .air_in(c_11_0));
valve v_11_457 (.fluid_in(k_11_457), .fluid_out(k_10_228), .air_in(c_11_1));
valve v_11_458 (.fluid_in(k_11_458), .fluid_out(k_10_229), .air_in(c_11_0));
valve v_11_459 (.fluid_in(k_11_459), .fluid_out(k_10_229), .air_in(c_11_1));
valve v_11_460 (.fluid_in(k_11_460), .fluid_out(k_10_230), .air_in(c_11_0));
valve v_11_461 (.fluid_in(k_11_461), .fluid_out(k_10_230), .air_in(c_11_1));
valve v_11_462 (.fluid_in(k_11_462), .fluid_out(k_10_231), .air_in(c_11_0));
valve v_11_463 (.fluid_in(k_11_463), .fluid_out(k_10_231), .air_in(c_11_1));
valve v_11_464 (.fluid_in(k_11_464), .fluid_out(k_10_232), .air_in(c_11_0));
valve v_11_465 (.fluid_in(k_11_465), .fluid_out(k_10_232), .air_in(c_11_1));
valve v_11_466 (.fluid_in(k_11_466), .fluid_out(k_10_233), .air_in(c_11_0));
valve v_11_467 (.fluid_in(k_11_467), .fluid_out(k_10_233), .air_in(c_11_1));
valve v_11_468 (.fluid_in(k_11_468), .fluid_out(k_10_234), .air_in(c_11_0));
valve v_11_469 (.fluid_in(k_11_469), .fluid_out(k_10_234), .air_in(c_11_1));
valve v_11_470 (.fluid_in(k_11_470), .fluid_out(k_10_235), .air_in(c_11_0));
valve v_11_471 (.fluid_in(k_11_471), .fluid_out(k_10_235), .air_in(c_11_1));
valve v_11_472 (.fluid_in(k_11_472), .fluid_out(k_10_236), .air_in(c_11_0));
valve v_11_473 (.fluid_in(k_11_473), .fluid_out(k_10_236), .air_in(c_11_1));
valve v_11_474 (.fluid_in(k_11_474), .fluid_out(k_10_237), .air_in(c_11_0));
valve v_11_475 (.fluid_in(k_11_475), .fluid_out(k_10_237), .air_in(c_11_1));
valve v_11_476 (.fluid_in(k_11_476), .fluid_out(k_10_238), .air_in(c_11_0));
valve v_11_477 (.fluid_in(k_11_477), .fluid_out(k_10_238), .air_in(c_11_1));
valve v_11_478 (.fluid_in(k_11_478), .fluid_out(k_10_239), .air_in(c_11_0));
valve v_11_479 (.fluid_in(k_11_479), .fluid_out(k_10_239), .air_in(c_11_1));
valve v_11_480 (.fluid_in(k_11_480), .fluid_out(k_10_240), .air_in(c_11_0));
valve v_11_481 (.fluid_in(k_11_481), .fluid_out(k_10_240), .air_in(c_11_1));
valve v_11_482 (.fluid_in(k_11_482), .fluid_out(k_10_241), .air_in(c_11_0));
valve v_11_483 (.fluid_in(k_11_483), .fluid_out(k_10_241), .air_in(c_11_1));
valve v_11_484 (.fluid_in(k_11_484), .fluid_out(k_10_242), .air_in(c_11_0));
valve v_11_485 (.fluid_in(k_11_485), .fluid_out(k_10_242), .air_in(c_11_1));
valve v_11_486 (.fluid_in(k_11_486), .fluid_out(k_10_243), .air_in(c_11_0));
valve v_11_487 (.fluid_in(k_11_487), .fluid_out(k_10_243), .air_in(c_11_1));
valve v_11_488 (.fluid_in(k_11_488), .fluid_out(k_10_244), .air_in(c_11_0));
valve v_11_489 (.fluid_in(k_11_489), .fluid_out(k_10_244), .air_in(c_11_1));
valve v_11_490 (.fluid_in(k_11_490), .fluid_out(k_10_245), .air_in(c_11_0));
valve v_11_491 (.fluid_in(k_11_491), .fluid_out(k_10_245), .air_in(c_11_1));
valve v_11_492 (.fluid_in(k_11_492), .fluid_out(k_10_246), .air_in(c_11_0));
valve v_11_493 (.fluid_in(k_11_493), .fluid_out(k_10_246), .air_in(c_11_1));
valve v_11_494 (.fluid_in(k_11_494), .fluid_out(k_10_247), .air_in(c_11_0));
valve v_11_495 (.fluid_in(k_11_495), .fluid_out(k_10_247), .air_in(c_11_1));
valve v_11_496 (.fluid_in(k_11_496), .fluid_out(k_10_248), .air_in(c_11_0));
valve v_11_497 (.fluid_in(k_11_497), .fluid_out(k_10_248), .air_in(c_11_1));
valve v_11_498 (.fluid_in(k_11_498), .fluid_out(k_10_249), .air_in(c_11_0));
valve v_11_499 (.fluid_in(k_11_499), .fluid_out(k_10_249), .air_in(c_11_1));
valve v_11_500 (.fluid_in(k_11_500), .fluid_out(k_10_250), .air_in(c_11_0));
valve v_11_501 (.fluid_in(k_11_501), .fluid_out(k_10_250), .air_in(c_11_1));
valve v_11_502 (.fluid_in(k_11_502), .fluid_out(k_10_251), .air_in(c_11_0));
valve v_11_503 (.fluid_in(k_11_503), .fluid_out(k_10_251), .air_in(c_11_1));
valve v_11_504 (.fluid_in(k_11_504), .fluid_out(k_10_252), .air_in(c_11_0));
valve v_11_505 (.fluid_in(k_11_505), .fluid_out(k_10_252), .air_in(c_11_1));
valve v_11_506 (.fluid_in(k_11_506), .fluid_out(k_10_253), .air_in(c_11_0));
valve v_11_507 (.fluid_in(k_11_507), .fluid_out(k_10_253), .air_in(c_11_1));
valve v_11_508 (.fluid_in(k_11_508), .fluid_out(k_10_254), .air_in(c_11_0));
valve v_11_509 (.fluid_in(k_11_509), .fluid_out(k_10_254), .air_in(c_11_1));
valve v_11_510 (.fluid_in(k_11_510), .fluid_out(k_10_255), .air_in(c_11_0));
valve v_11_511 (.fluid_in(k_11_511), .fluid_out(k_10_255), .air_in(c_11_1));
valve v_11_512 (.fluid_in(k_11_512), .fluid_out(k_10_256), .air_in(c_11_0));
valve v_11_513 (.fluid_in(k_11_513), .fluid_out(k_10_256), .air_in(c_11_1));
valve v_11_514 (.fluid_in(k_11_514), .fluid_out(k_10_257), .air_in(c_11_0));
valve v_11_515 (.fluid_in(k_11_515), .fluid_out(k_10_257), .air_in(c_11_1));
valve v_11_516 (.fluid_in(k_11_516), .fluid_out(k_10_258), .air_in(c_11_0));
valve v_11_517 (.fluid_in(k_11_517), .fluid_out(k_10_258), .air_in(c_11_1));
valve v_11_518 (.fluid_in(k_11_518), .fluid_out(k_10_259), .air_in(c_11_0));
valve v_11_519 (.fluid_in(k_11_519), .fluid_out(k_10_259), .air_in(c_11_1));
valve v_11_520 (.fluid_in(k_11_520), .fluid_out(k_10_260), .air_in(c_11_0));
valve v_11_521 (.fluid_in(k_11_521), .fluid_out(k_10_260), .air_in(c_11_1));
valve v_11_522 (.fluid_in(k_11_522), .fluid_out(k_10_261), .air_in(c_11_0));
valve v_11_523 (.fluid_in(k_11_523), .fluid_out(k_10_261), .air_in(c_11_1));
valve v_11_524 (.fluid_in(k_11_524), .fluid_out(k_10_262), .air_in(c_11_0));
valve v_11_525 (.fluid_in(k_11_525), .fluid_out(k_10_262), .air_in(c_11_1));
valve v_11_526 (.fluid_in(k_11_526), .fluid_out(k_10_263), .air_in(c_11_0));
valve v_11_527 (.fluid_in(k_11_527), .fluid_out(k_10_263), .air_in(c_11_1));
valve v_11_528 (.fluid_in(k_11_528), .fluid_out(k_10_264), .air_in(c_11_0));
valve v_11_529 (.fluid_in(k_11_529), .fluid_out(k_10_264), .air_in(c_11_1));
valve v_11_530 (.fluid_in(k_11_530), .fluid_out(k_10_265), .air_in(c_11_0));
valve v_11_531 (.fluid_in(k_11_531), .fluid_out(k_10_265), .air_in(c_11_1));
valve v_11_532 (.fluid_in(k_11_532), .fluid_out(k_10_266), .air_in(c_11_0));
valve v_11_533 (.fluid_in(k_11_533), .fluid_out(k_10_266), .air_in(c_11_1));
valve v_11_534 (.fluid_in(k_11_534), .fluid_out(k_10_267), .air_in(c_11_0));
valve v_11_535 (.fluid_in(k_11_535), .fluid_out(k_10_267), .air_in(c_11_1));
valve v_11_536 (.fluid_in(k_11_536), .fluid_out(k_10_268), .air_in(c_11_0));
valve v_11_537 (.fluid_in(k_11_537), .fluid_out(k_10_268), .air_in(c_11_1));
valve v_11_538 (.fluid_in(k_11_538), .fluid_out(k_10_269), .air_in(c_11_0));
valve v_11_539 (.fluid_in(k_11_539), .fluid_out(k_10_269), .air_in(c_11_1));
valve v_11_540 (.fluid_in(k_11_540), .fluid_out(k_10_270), .air_in(c_11_0));
valve v_11_541 (.fluid_in(k_11_541), .fluid_out(k_10_270), .air_in(c_11_1));
valve v_11_542 (.fluid_in(k_11_542), .fluid_out(k_10_271), .air_in(c_11_0));
valve v_11_543 (.fluid_in(k_11_543), .fluid_out(k_10_271), .air_in(c_11_1));
valve v_11_544 (.fluid_in(k_11_544), .fluid_out(k_10_272), .air_in(c_11_0));
valve v_11_545 (.fluid_in(k_11_545), .fluid_out(k_10_272), .air_in(c_11_1));
valve v_11_546 (.fluid_in(k_11_546), .fluid_out(k_10_273), .air_in(c_11_0));
valve v_11_547 (.fluid_in(k_11_547), .fluid_out(k_10_273), .air_in(c_11_1));
valve v_11_548 (.fluid_in(k_11_548), .fluid_out(k_10_274), .air_in(c_11_0));
valve v_11_549 (.fluid_in(k_11_549), .fluid_out(k_10_274), .air_in(c_11_1));
valve v_11_550 (.fluid_in(k_11_550), .fluid_out(k_10_275), .air_in(c_11_0));
valve v_11_551 (.fluid_in(k_11_551), .fluid_out(k_10_275), .air_in(c_11_1));
valve v_11_552 (.fluid_in(k_11_552), .fluid_out(k_10_276), .air_in(c_11_0));
valve v_11_553 (.fluid_in(k_11_553), .fluid_out(k_10_276), .air_in(c_11_1));
valve v_11_554 (.fluid_in(k_11_554), .fluid_out(k_10_277), .air_in(c_11_0));
valve v_11_555 (.fluid_in(k_11_555), .fluid_out(k_10_277), .air_in(c_11_1));
valve v_11_556 (.fluid_in(k_11_556), .fluid_out(k_10_278), .air_in(c_11_0));
valve v_11_557 (.fluid_in(k_11_557), .fluid_out(k_10_278), .air_in(c_11_1));
valve v_11_558 (.fluid_in(k_11_558), .fluid_out(k_10_279), .air_in(c_11_0));
valve v_11_559 (.fluid_in(k_11_559), .fluid_out(k_10_279), .air_in(c_11_1));
valve v_11_560 (.fluid_in(k_11_560), .fluid_out(k_10_280), .air_in(c_11_0));
valve v_11_561 (.fluid_in(k_11_561), .fluid_out(k_10_280), .air_in(c_11_1));
valve v_11_562 (.fluid_in(k_11_562), .fluid_out(k_10_281), .air_in(c_11_0));
valve v_11_563 (.fluid_in(k_11_563), .fluid_out(k_10_281), .air_in(c_11_1));
valve v_11_564 (.fluid_in(k_11_564), .fluid_out(k_10_282), .air_in(c_11_0));
valve v_11_565 (.fluid_in(k_11_565), .fluid_out(k_10_282), .air_in(c_11_1));
valve v_11_566 (.fluid_in(k_11_566), .fluid_out(k_10_283), .air_in(c_11_0));
valve v_11_567 (.fluid_in(k_11_567), .fluid_out(k_10_283), .air_in(c_11_1));
valve v_11_568 (.fluid_in(k_11_568), .fluid_out(k_10_284), .air_in(c_11_0));
valve v_11_569 (.fluid_in(k_11_569), .fluid_out(k_10_284), .air_in(c_11_1));
valve v_11_570 (.fluid_in(k_11_570), .fluid_out(k_10_285), .air_in(c_11_0));
valve v_11_571 (.fluid_in(k_11_571), .fluid_out(k_10_285), .air_in(c_11_1));
valve v_11_572 (.fluid_in(k_11_572), .fluid_out(k_10_286), .air_in(c_11_0));
valve v_11_573 (.fluid_in(k_11_573), .fluid_out(k_10_286), .air_in(c_11_1));
valve v_11_574 (.fluid_in(k_11_574), .fluid_out(k_10_287), .air_in(c_11_0));
valve v_11_575 (.fluid_in(k_11_575), .fluid_out(k_10_287), .air_in(c_11_1));
valve v_11_576 (.fluid_in(k_11_576), .fluid_out(k_10_288), .air_in(c_11_0));
valve v_11_577 (.fluid_in(k_11_577), .fluid_out(k_10_288), .air_in(c_11_1));
valve v_11_578 (.fluid_in(k_11_578), .fluid_out(k_10_289), .air_in(c_11_0));
valve v_11_579 (.fluid_in(k_11_579), .fluid_out(k_10_289), .air_in(c_11_1));
valve v_11_580 (.fluid_in(k_11_580), .fluid_out(k_10_290), .air_in(c_11_0));
valve v_11_581 (.fluid_in(k_11_581), .fluid_out(k_10_290), .air_in(c_11_1));
valve v_11_582 (.fluid_in(k_11_582), .fluid_out(k_10_291), .air_in(c_11_0));
valve v_11_583 (.fluid_in(k_11_583), .fluid_out(k_10_291), .air_in(c_11_1));
valve v_11_584 (.fluid_in(k_11_584), .fluid_out(k_10_292), .air_in(c_11_0));
valve v_11_585 (.fluid_in(k_11_585), .fluid_out(k_10_292), .air_in(c_11_1));
valve v_11_586 (.fluid_in(k_11_586), .fluid_out(k_10_293), .air_in(c_11_0));
valve v_11_587 (.fluid_in(k_11_587), .fluid_out(k_10_293), .air_in(c_11_1));
valve v_11_588 (.fluid_in(k_11_588), .fluid_out(k_10_294), .air_in(c_11_0));
valve v_11_589 (.fluid_in(k_11_589), .fluid_out(k_10_294), .air_in(c_11_1));
valve v_11_590 (.fluid_in(k_11_590), .fluid_out(k_10_295), .air_in(c_11_0));
valve v_11_591 (.fluid_in(k_11_591), .fluid_out(k_10_295), .air_in(c_11_1));
valve v_11_592 (.fluid_in(k_11_592), .fluid_out(k_10_296), .air_in(c_11_0));
valve v_11_593 (.fluid_in(k_11_593), .fluid_out(k_10_296), .air_in(c_11_1));
valve v_11_594 (.fluid_in(k_11_594), .fluid_out(k_10_297), .air_in(c_11_0));
valve v_11_595 (.fluid_in(k_11_595), .fluid_out(k_10_297), .air_in(c_11_1));
valve v_11_596 (.fluid_in(k_11_596), .fluid_out(k_10_298), .air_in(c_11_0));
valve v_11_597 (.fluid_in(k_11_597), .fluid_out(k_10_298), .air_in(c_11_1));
valve v_11_598 (.fluid_in(k_11_598), .fluid_out(k_10_299), .air_in(c_11_0));
valve v_11_599 (.fluid_in(k_11_599), .fluid_out(k_10_299), .air_in(c_11_1));
valve v_11_600 (.fluid_in(k_11_600), .fluid_out(k_10_300), .air_in(c_11_0));
valve v_11_601 (.fluid_in(k_11_601), .fluid_out(k_10_300), .air_in(c_11_1));
valve v_11_602 (.fluid_in(k_11_602), .fluid_out(k_10_301), .air_in(c_11_0));
valve v_11_603 (.fluid_in(k_11_603), .fluid_out(k_10_301), .air_in(c_11_1));
valve v_11_604 (.fluid_in(k_11_604), .fluid_out(k_10_302), .air_in(c_11_0));
valve v_11_605 (.fluid_in(k_11_605), .fluid_out(k_10_302), .air_in(c_11_1));
valve v_11_606 (.fluid_in(k_11_606), .fluid_out(k_10_303), .air_in(c_11_0));
valve v_11_607 (.fluid_in(k_11_607), .fluid_out(k_10_303), .air_in(c_11_1));
valve v_11_608 (.fluid_in(k_11_608), .fluid_out(k_10_304), .air_in(c_11_0));
valve v_11_609 (.fluid_in(k_11_609), .fluid_out(k_10_304), .air_in(c_11_1));
valve v_11_610 (.fluid_in(k_11_610), .fluid_out(k_10_305), .air_in(c_11_0));
valve v_11_611 (.fluid_in(k_11_611), .fluid_out(k_10_305), .air_in(c_11_1));
valve v_11_612 (.fluid_in(k_11_612), .fluid_out(k_10_306), .air_in(c_11_0));
valve v_11_613 (.fluid_in(k_11_613), .fluid_out(k_10_306), .air_in(c_11_1));
valve v_11_614 (.fluid_in(k_11_614), .fluid_out(k_10_307), .air_in(c_11_0));
valve v_11_615 (.fluid_in(k_11_615), .fluid_out(k_10_307), .air_in(c_11_1));
valve v_11_616 (.fluid_in(k_11_616), .fluid_out(k_10_308), .air_in(c_11_0));
valve v_11_617 (.fluid_in(k_11_617), .fluid_out(k_10_308), .air_in(c_11_1));
valve v_11_618 (.fluid_in(k_11_618), .fluid_out(k_10_309), .air_in(c_11_0));
valve v_11_619 (.fluid_in(k_11_619), .fluid_out(k_10_309), .air_in(c_11_1));
valve v_11_620 (.fluid_in(k_11_620), .fluid_out(k_10_310), .air_in(c_11_0));
valve v_11_621 (.fluid_in(k_11_621), .fluid_out(k_10_310), .air_in(c_11_1));
valve v_11_622 (.fluid_in(k_11_622), .fluid_out(k_10_311), .air_in(c_11_0));
valve v_11_623 (.fluid_in(k_11_623), .fluid_out(k_10_311), .air_in(c_11_1));
valve v_11_624 (.fluid_in(k_11_624), .fluid_out(k_10_312), .air_in(c_11_0));
valve v_11_625 (.fluid_in(k_11_625), .fluid_out(k_10_312), .air_in(c_11_1));
valve v_11_626 (.fluid_in(k_11_626), .fluid_out(k_10_313), .air_in(c_11_0));
valve v_11_627 (.fluid_in(k_11_627), .fluid_out(k_10_313), .air_in(c_11_1));
valve v_11_628 (.fluid_in(k_11_628), .fluid_out(k_10_314), .air_in(c_11_0));
valve v_11_629 (.fluid_in(k_11_629), .fluid_out(k_10_314), .air_in(c_11_1));
valve v_11_630 (.fluid_in(k_11_630), .fluid_out(k_10_315), .air_in(c_11_0));
valve v_11_631 (.fluid_in(k_11_631), .fluid_out(k_10_315), .air_in(c_11_1));
valve v_11_632 (.fluid_in(k_11_632), .fluid_out(k_10_316), .air_in(c_11_0));
valve v_11_633 (.fluid_in(k_11_633), .fluid_out(k_10_316), .air_in(c_11_1));
valve v_11_634 (.fluid_in(k_11_634), .fluid_out(k_10_317), .air_in(c_11_0));
valve v_11_635 (.fluid_in(k_11_635), .fluid_out(k_10_317), .air_in(c_11_1));
valve v_11_636 (.fluid_in(k_11_636), .fluid_out(k_10_318), .air_in(c_11_0));
valve v_11_637 (.fluid_in(k_11_637), .fluid_out(k_10_318), .air_in(c_11_1));
valve v_11_638 (.fluid_in(k_11_638), .fluid_out(k_10_319), .air_in(c_11_0));
valve v_11_639 (.fluid_in(k_11_639), .fluid_out(k_10_319), .air_in(c_11_1));
valve v_11_640 (.fluid_in(k_11_640), .fluid_out(k_10_320), .air_in(c_11_0));
valve v_11_641 (.fluid_in(k_11_641), .fluid_out(k_10_320), .air_in(c_11_1));
valve v_11_642 (.fluid_in(k_11_642), .fluid_out(k_10_321), .air_in(c_11_0));
valve v_11_643 (.fluid_in(k_11_643), .fluid_out(k_10_321), .air_in(c_11_1));
valve v_11_644 (.fluid_in(k_11_644), .fluid_out(k_10_322), .air_in(c_11_0));
valve v_11_645 (.fluid_in(k_11_645), .fluid_out(k_10_322), .air_in(c_11_1));
valve v_11_646 (.fluid_in(k_11_646), .fluid_out(k_10_323), .air_in(c_11_0));
valve v_11_647 (.fluid_in(k_11_647), .fluid_out(k_10_323), .air_in(c_11_1));
valve v_11_648 (.fluid_in(k_11_648), .fluid_out(k_10_324), .air_in(c_11_0));
valve v_11_649 (.fluid_in(k_11_649), .fluid_out(k_10_324), .air_in(c_11_1));
valve v_11_650 (.fluid_in(k_11_650), .fluid_out(k_10_325), .air_in(c_11_0));
valve v_11_651 (.fluid_in(k_11_651), .fluid_out(k_10_325), .air_in(c_11_1));
valve v_11_652 (.fluid_in(k_11_652), .fluid_out(k_10_326), .air_in(c_11_0));
valve v_11_653 (.fluid_in(k_11_653), .fluid_out(k_10_326), .air_in(c_11_1));
valve v_11_654 (.fluid_in(k_11_654), .fluid_out(k_10_327), .air_in(c_11_0));
valve v_11_655 (.fluid_in(k_11_655), .fluid_out(k_10_327), .air_in(c_11_1));
valve v_11_656 (.fluid_in(k_11_656), .fluid_out(k_10_328), .air_in(c_11_0));
valve v_11_657 (.fluid_in(k_11_657), .fluid_out(k_10_328), .air_in(c_11_1));
valve v_11_658 (.fluid_in(k_11_658), .fluid_out(k_10_329), .air_in(c_11_0));
valve v_11_659 (.fluid_in(k_11_659), .fluid_out(k_10_329), .air_in(c_11_1));
valve v_11_660 (.fluid_in(k_11_660), .fluid_out(k_10_330), .air_in(c_11_0));
valve v_11_661 (.fluid_in(k_11_661), .fluid_out(k_10_330), .air_in(c_11_1));
valve v_11_662 (.fluid_in(k_11_662), .fluid_out(k_10_331), .air_in(c_11_0));
valve v_11_663 (.fluid_in(k_11_663), .fluid_out(k_10_331), .air_in(c_11_1));
valve v_11_664 (.fluid_in(k_11_664), .fluid_out(k_10_332), .air_in(c_11_0));
valve v_11_665 (.fluid_in(k_11_665), .fluid_out(k_10_332), .air_in(c_11_1));
valve v_11_666 (.fluid_in(k_11_666), .fluid_out(k_10_333), .air_in(c_11_0));
valve v_11_667 (.fluid_in(k_11_667), .fluid_out(k_10_333), .air_in(c_11_1));
valve v_11_668 (.fluid_in(k_11_668), .fluid_out(k_10_334), .air_in(c_11_0));
valve v_11_669 (.fluid_in(k_11_669), .fluid_out(k_10_334), .air_in(c_11_1));
valve v_11_670 (.fluid_in(k_11_670), .fluid_out(k_10_335), .air_in(c_11_0));
valve v_11_671 (.fluid_in(k_11_671), .fluid_out(k_10_335), .air_in(c_11_1));
valve v_11_672 (.fluid_in(k_11_672), .fluid_out(k_10_336), .air_in(c_11_0));
valve v_11_673 (.fluid_in(k_11_673), .fluid_out(k_10_336), .air_in(c_11_1));
valve v_11_674 (.fluid_in(k_11_674), .fluid_out(k_10_337), .air_in(c_11_0));
valve v_11_675 (.fluid_in(k_11_675), .fluid_out(k_10_337), .air_in(c_11_1));
valve v_11_676 (.fluid_in(k_11_676), .fluid_out(k_10_338), .air_in(c_11_0));
valve v_11_677 (.fluid_in(k_11_677), .fluid_out(k_10_338), .air_in(c_11_1));
valve v_11_678 (.fluid_in(k_11_678), .fluid_out(k_10_339), .air_in(c_11_0));
valve v_11_679 (.fluid_in(k_11_679), .fluid_out(k_10_339), .air_in(c_11_1));
valve v_11_680 (.fluid_in(k_11_680), .fluid_out(k_10_340), .air_in(c_11_0));
valve v_11_681 (.fluid_in(k_11_681), .fluid_out(k_10_340), .air_in(c_11_1));
valve v_11_682 (.fluid_in(k_11_682), .fluid_out(k_10_341), .air_in(c_11_0));
valve v_11_683 (.fluid_in(k_11_683), .fluid_out(k_10_341), .air_in(c_11_1));
valve v_11_684 (.fluid_in(k_11_684), .fluid_out(k_10_342), .air_in(c_11_0));
valve v_11_685 (.fluid_in(k_11_685), .fluid_out(k_10_342), .air_in(c_11_1));
valve v_11_686 (.fluid_in(k_11_686), .fluid_out(k_10_343), .air_in(c_11_0));
valve v_11_687 (.fluid_in(k_11_687), .fluid_out(k_10_343), .air_in(c_11_1));
valve v_11_688 (.fluid_in(k_11_688), .fluid_out(k_10_344), .air_in(c_11_0));
valve v_11_689 (.fluid_in(k_11_689), .fluid_out(k_10_344), .air_in(c_11_1));
valve v_11_690 (.fluid_in(k_11_690), .fluid_out(k_10_345), .air_in(c_11_0));
valve v_11_691 (.fluid_in(k_11_691), .fluid_out(k_10_345), .air_in(c_11_1));
valve v_11_692 (.fluid_in(k_11_692), .fluid_out(k_10_346), .air_in(c_11_0));
valve v_11_693 (.fluid_in(k_11_693), .fluid_out(k_10_346), .air_in(c_11_1));
valve v_11_694 (.fluid_in(k_11_694), .fluid_out(k_10_347), .air_in(c_11_0));
valve v_11_695 (.fluid_in(k_11_695), .fluid_out(k_10_347), .air_in(c_11_1));
valve v_11_696 (.fluid_in(k_11_696), .fluid_out(k_10_348), .air_in(c_11_0));
valve v_11_697 (.fluid_in(k_11_697), .fluid_out(k_10_348), .air_in(c_11_1));
valve v_11_698 (.fluid_in(k_11_698), .fluid_out(k_10_349), .air_in(c_11_0));
valve v_11_699 (.fluid_in(k_11_699), .fluid_out(k_10_349), .air_in(c_11_1));
valve v_11_700 (.fluid_in(k_11_700), .fluid_out(k_10_350), .air_in(c_11_0));
valve v_11_701 (.fluid_in(k_11_701), .fluid_out(k_10_350), .air_in(c_11_1));
valve v_11_702 (.fluid_in(k_11_702), .fluid_out(k_10_351), .air_in(c_11_0));
valve v_11_703 (.fluid_in(k_11_703), .fluid_out(k_10_351), .air_in(c_11_1));
valve v_11_704 (.fluid_in(k_11_704), .fluid_out(k_10_352), .air_in(c_11_0));
valve v_11_705 (.fluid_in(k_11_705), .fluid_out(k_10_352), .air_in(c_11_1));
valve v_11_706 (.fluid_in(k_11_706), .fluid_out(k_10_353), .air_in(c_11_0));
valve v_11_707 (.fluid_in(k_11_707), .fluid_out(k_10_353), .air_in(c_11_1));
valve v_11_708 (.fluid_in(k_11_708), .fluid_out(k_10_354), .air_in(c_11_0));
valve v_11_709 (.fluid_in(k_11_709), .fluid_out(k_10_354), .air_in(c_11_1));
valve v_11_710 (.fluid_in(k_11_710), .fluid_out(k_10_355), .air_in(c_11_0));
valve v_11_711 (.fluid_in(k_11_711), .fluid_out(k_10_355), .air_in(c_11_1));
valve v_11_712 (.fluid_in(k_11_712), .fluid_out(k_10_356), .air_in(c_11_0));
valve v_11_713 (.fluid_in(k_11_713), .fluid_out(k_10_356), .air_in(c_11_1));
valve v_11_714 (.fluid_in(k_11_714), .fluid_out(k_10_357), .air_in(c_11_0));
valve v_11_715 (.fluid_in(k_11_715), .fluid_out(k_10_357), .air_in(c_11_1));
valve v_11_716 (.fluid_in(k_11_716), .fluid_out(k_10_358), .air_in(c_11_0));
valve v_11_717 (.fluid_in(k_11_717), .fluid_out(k_10_358), .air_in(c_11_1));
valve v_11_718 (.fluid_in(k_11_718), .fluid_out(k_10_359), .air_in(c_11_0));
valve v_11_719 (.fluid_in(k_11_719), .fluid_out(k_10_359), .air_in(c_11_1));
valve v_11_720 (.fluid_in(k_11_720), .fluid_out(k_10_360), .air_in(c_11_0));
valve v_11_721 (.fluid_in(k_11_721), .fluid_out(k_10_360), .air_in(c_11_1));
valve v_11_722 (.fluid_in(k_11_722), .fluid_out(k_10_361), .air_in(c_11_0));
valve v_11_723 (.fluid_in(k_11_723), .fluid_out(k_10_361), .air_in(c_11_1));
valve v_11_724 (.fluid_in(k_11_724), .fluid_out(k_10_362), .air_in(c_11_0));
valve v_11_725 (.fluid_in(k_11_725), .fluid_out(k_10_362), .air_in(c_11_1));
valve v_11_726 (.fluid_in(k_11_726), .fluid_out(k_10_363), .air_in(c_11_0));
valve v_11_727 (.fluid_in(k_11_727), .fluid_out(k_10_363), .air_in(c_11_1));
valve v_11_728 (.fluid_in(k_11_728), .fluid_out(k_10_364), .air_in(c_11_0));
valve v_11_729 (.fluid_in(k_11_729), .fluid_out(k_10_364), .air_in(c_11_1));
valve v_11_730 (.fluid_in(k_11_730), .fluid_out(k_10_365), .air_in(c_11_0));
valve v_11_731 (.fluid_in(k_11_731), .fluid_out(k_10_365), .air_in(c_11_1));
valve v_11_732 (.fluid_in(k_11_732), .fluid_out(k_10_366), .air_in(c_11_0));
valve v_11_733 (.fluid_in(k_11_733), .fluid_out(k_10_366), .air_in(c_11_1));
valve v_11_734 (.fluid_in(k_11_734), .fluid_out(k_10_367), .air_in(c_11_0));
valve v_11_735 (.fluid_in(k_11_735), .fluid_out(k_10_367), .air_in(c_11_1));
valve v_11_736 (.fluid_in(k_11_736), .fluid_out(k_10_368), .air_in(c_11_0));
valve v_11_737 (.fluid_in(k_11_737), .fluid_out(k_10_368), .air_in(c_11_1));
valve v_11_738 (.fluid_in(k_11_738), .fluid_out(k_10_369), .air_in(c_11_0));
valve v_11_739 (.fluid_in(k_11_739), .fluid_out(k_10_369), .air_in(c_11_1));
valve v_11_740 (.fluid_in(k_11_740), .fluid_out(k_10_370), .air_in(c_11_0));
valve v_11_741 (.fluid_in(k_11_741), .fluid_out(k_10_370), .air_in(c_11_1));
valve v_11_742 (.fluid_in(k_11_742), .fluid_out(k_10_371), .air_in(c_11_0));
valve v_11_743 (.fluid_in(k_11_743), .fluid_out(k_10_371), .air_in(c_11_1));
valve v_11_744 (.fluid_in(k_11_744), .fluid_out(k_10_372), .air_in(c_11_0));
valve v_11_745 (.fluid_in(k_11_745), .fluid_out(k_10_372), .air_in(c_11_1));
valve v_11_746 (.fluid_in(k_11_746), .fluid_out(k_10_373), .air_in(c_11_0));
valve v_11_747 (.fluid_in(k_11_747), .fluid_out(k_10_373), .air_in(c_11_1));
valve v_11_748 (.fluid_in(k_11_748), .fluid_out(k_10_374), .air_in(c_11_0));
valve v_11_749 (.fluid_in(k_11_749), .fluid_out(k_10_374), .air_in(c_11_1));
valve v_11_750 (.fluid_in(k_11_750), .fluid_out(k_10_375), .air_in(c_11_0));
valve v_11_751 (.fluid_in(k_11_751), .fluid_out(k_10_375), .air_in(c_11_1));
valve v_11_752 (.fluid_in(k_11_752), .fluid_out(k_10_376), .air_in(c_11_0));
valve v_11_753 (.fluid_in(k_11_753), .fluid_out(k_10_376), .air_in(c_11_1));
valve v_11_754 (.fluid_in(k_11_754), .fluid_out(k_10_377), .air_in(c_11_0));
valve v_11_755 (.fluid_in(k_11_755), .fluid_out(k_10_377), .air_in(c_11_1));
valve v_11_756 (.fluid_in(k_11_756), .fluid_out(k_10_378), .air_in(c_11_0));
valve v_11_757 (.fluid_in(k_11_757), .fluid_out(k_10_378), .air_in(c_11_1));
valve v_11_758 (.fluid_in(k_11_758), .fluid_out(k_10_379), .air_in(c_11_0));
valve v_11_759 (.fluid_in(k_11_759), .fluid_out(k_10_379), .air_in(c_11_1));
valve v_11_760 (.fluid_in(k_11_760), .fluid_out(k_10_380), .air_in(c_11_0));
valve v_11_761 (.fluid_in(k_11_761), .fluid_out(k_10_380), .air_in(c_11_1));
valve v_11_762 (.fluid_in(k_11_762), .fluid_out(k_10_381), .air_in(c_11_0));
valve v_11_763 (.fluid_in(k_11_763), .fluid_out(k_10_381), .air_in(c_11_1));
valve v_11_764 (.fluid_in(k_11_764), .fluid_out(k_10_382), .air_in(c_11_0));
valve v_11_765 (.fluid_in(k_11_765), .fluid_out(k_10_382), .air_in(c_11_1));
valve v_11_766 (.fluid_in(k_11_766), .fluid_out(k_10_383), .air_in(c_11_0));
valve v_11_767 (.fluid_in(k_11_767), .fluid_out(k_10_383), .air_in(c_11_1));
valve v_11_768 (.fluid_in(k_11_768), .fluid_out(k_10_384), .air_in(c_11_0));
valve v_11_769 (.fluid_in(k_11_769), .fluid_out(k_10_384), .air_in(c_11_1));
valve v_11_770 (.fluid_in(k_11_770), .fluid_out(k_10_385), .air_in(c_11_0));
valve v_11_771 (.fluid_in(k_11_771), .fluid_out(k_10_385), .air_in(c_11_1));
valve v_11_772 (.fluid_in(k_11_772), .fluid_out(k_10_386), .air_in(c_11_0));
valve v_11_773 (.fluid_in(k_11_773), .fluid_out(k_10_386), .air_in(c_11_1));
valve v_11_774 (.fluid_in(k_11_774), .fluid_out(k_10_387), .air_in(c_11_0));
valve v_11_775 (.fluid_in(k_11_775), .fluid_out(k_10_387), .air_in(c_11_1));
valve v_11_776 (.fluid_in(k_11_776), .fluid_out(k_10_388), .air_in(c_11_0));
valve v_11_777 (.fluid_in(k_11_777), .fluid_out(k_10_388), .air_in(c_11_1));
valve v_11_778 (.fluid_in(k_11_778), .fluid_out(k_10_389), .air_in(c_11_0));
valve v_11_779 (.fluid_in(k_11_779), .fluid_out(k_10_389), .air_in(c_11_1));
valve v_11_780 (.fluid_in(k_11_780), .fluid_out(k_10_390), .air_in(c_11_0));
valve v_11_781 (.fluid_in(k_11_781), .fluid_out(k_10_390), .air_in(c_11_1));
valve v_11_782 (.fluid_in(k_11_782), .fluid_out(k_10_391), .air_in(c_11_0));
valve v_11_783 (.fluid_in(k_11_783), .fluid_out(k_10_391), .air_in(c_11_1));
valve v_11_784 (.fluid_in(k_11_784), .fluid_out(k_10_392), .air_in(c_11_0));
valve v_11_785 (.fluid_in(k_11_785), .fluid_out(k_10_392), .air_in(c_11_1));
valve v_11_786 (.fluid_in(k_11_786), .fluid_out(k_10_393), .air_in(c_11_0));
valve v_11_787 (.fluid_in(k_11_787), .fluid_out(k_10_393), .air_in(c_11_1));
valve v_11_788 (.fluid_in(k_11_788), .fluid_out(k_10_394), .air_in(c_11_0));
valve v_11_789 (.fluid_in(k_11_789), .fluid_out(k_10_394), .air_in(c_11_1));
valve v_11_790 (.fluid_in(k_11_790), .fluid_out(k_10_395), .air_in(c_11_0));
valve v_11_791 (.fluid_in(k_11_791), .fluid_out(k_10_395), .air_in(c_11_1));
valve v_11_792 (.fluid_in(k_11_792), .fluid_out(k_10_396), .air_in(c_11_0));
valve v_11_793 (.fluid_in(k_11_793), .fluid_out(k_10_396), .air_in(c_11_1));
valve v_11_794 (.fluid_in(k_11_794), .fluid_out(k_10_397), .air_in(c_11_0));
valve v_11_795 (.fluid_in(k_11_795), .fluid_out(k_10_397), .air_in(c_11_1));
valve v_11_796 (.fluid_in(k_11_796), .fluid_out(k_10_398), .air_in(c_11_0));
valve v_11_797 (.fluid_in(k_11_797), .fluid_out(k_10_398), .air_in(c_11_1));
valve v_11_798 (.fluid_in(k_11_798), .fluid_out(k_10_399), .air_in(c_11_0));
valve v_11_799 (.fluid_in(k_11_799), .fluid_out(k_10_399), .air_in(c_11_1));
valve v_11_800 (.fluid_in(k_11_800), .fluid_out(k_10_400), .air_in(c_11_0));
valve v_11_801 (.fluid_in(k_11_801), .fluid_out(k_10_400), .air_in(c_11_1));
valve v_11_802 (.fluid_in(k_11_802), .fluid_out(k_10_401), .air_in(c_11_0));
valve v_11_803 (.fluid_in(k_11_803), .fluid_out(k_10_401), .air_in(c_11_1));
valve v_11_804 (.fluid_in(k_11_804), .fluid_out(k_10_402), .air_in(c_11_0));
valve v_11_805 (.fluid_in(k_11_805), .fluid_out(k_10_402), .air_in(c_11_1));
valve v_11_806 (.fluid_in(k_11_806), .fluid_out(k_10_403), .air_in(c_11_0));
valve v_11_807 (.fluid_in(k_11_807), .fluid_out(k_10_403), .air_in(c_11_1));
valve v_11_808 (.fluid_in(k_11_808), .fluid_out(k_10_404), .air_in(c_11_0));
valve v_11_809 (.fluid_in(k_11_809), .fluid_out(k_10_404), .air_in(c_11_1));
valve v_11_810 (.fluid_in(k_11_810), .fluid_out(k_10_405), .air_in(c_11_0));
valve v_11_811 (.fluid_in(k_11_811), .fluid_out(k_10_405), .air_in(c_11_1));
valve v_11_812 (.fluid_in(k_11_812), .fluid_out(k_10_406), .air_in(c_11_0));
valve v_11_813 (.fluid_in(k_11_813), .fluid_out(k_10_406), .air_in(c_11_1));
valve v_11_814 (.fluid_in(k_11_814), .fluid_out(k_10_407), .air_in(c_11_0));
valve v_11_815 (.fluid_in(k_11_815), .fluid_out(k_10_407), .air_in(c_11_1));
valve v_11_816 (.fluid_in(k_11_816), .fluid_out(k_10_408), .air_in(c_11_0));
valve v_11_817 (.fluid_in(k_11_817), .fluid_out(k_10_408), .air_in(c_11_1));
valve v_11_818 (.fluid_in(k_11_818), .fluid_out(k_10_409), .air_in(c_11_0));
valve v_11_819 (.fluid_in(k_11_819), .fluid_out(k_10_409), .air_in(c_11_1));
valve v_11_820 (.fluid_in(k_11_820), .fluid_out(k_10_410), .air_in(c_11_0));
valve v_11_821 (.fluid_in(k_11_821), .fluid_out(k_10_410), .air_in(c_11_1));
valve v_11_822 (.fluid_in(k_11_822), .fluid_out(k_10_411), .air_in(c_11_0));
valve v_11_823 (.fluid_in(k_11_823), .fluid_out(k_10_411), .air_in(c_11_1));
valve v_11_824 (.fluid_in(k_11_824), .fluid_out(k_10_412), .air_in(c_11_0));
valve v_11_825 (.fluid_in(k_11_825), .fluid_out(k_10_412), .air_in(c_11_1));
valve v_11_826 (.fluid_in(k_11_826), .fluid_out(k_10_413), .air_in(c_11_0));
valve v_11_827 (.fluid_in(k_11_827), .fluid_out(k_10_413), .air_in(c_11_1));
valve v_11_828 (.fluid_in(k_11_828), .fluid_out(k_10_414), .air_in(c_11_0));
valve v_11_829 (.fluid_in(k_11_829), .fluid_out(k_10_414), .air_in(c_11_1));
valve v_11_830 (.fluid_in(k_11_830), .fluid_out(k_10_415), .air_in(c_11_0));
valve v_11_831 (.fluid_in(k_11_831), .fluid_out(k_10_415), .air_in(c_11_1));
valve v_11_832 (.fluid_in(k_11_832), .fluid_out(k_10_416), .air_in(c_11_0));
valve v_11_833 (.fluid_in(k_11_833), .fluid_out(k_10_416), .air_in(c_11_1));
valve v_11_834 (.fluid_in(k_11_834), .fluid_out(k_10_417), .air_in(c_11_0));
valve v_11_835 (.fluid_in(k_11_835), .fluid_out(k_10_417), .air_in(c_11_1));
valve v_11_836 (.fluid_in(k_11_836), .fluid_out(k_10_418), .air_in(c_11_0));
valve v_11_837 (.fluid_in(k_11_837), .fluid_out(k_10_418), .air_in(c_11_1));
valve v_11_838 (.fluid_in(k_11_838), .fluid_out(k_10_419), .air_in(c_11_0));
valve v_11_839 (.fluid_in(k_11_839), .fluid_out(k_10_419), .air_in(c_11_1));
valve v_11_840 (.fluid_in(k_11_840), .fluid_out(k_10_420), .air_in(c_11_0));
valve v_11_841 (.fluid_in(k_11_841), .fluid_out(k_10_420), .air_in(c_11_1));
valve v_11_842 (.fluid_in(k_11_842), .fluid_out(k_10_421), .air_in(c_11_0));
valve v_11_843 (.fluid_in(k_11_843), .fluid_out(k_10_421), .air_in(c_11_1));
valve v_11_844 (.fluid_in(k_11_844), .fluid_out(k_10_422), .air_in(c_11_0));
valve v_11_845 (.fluid_in(k_11_845), .fluid_out(k_10_422), .air_in(c_11_1));
valve v_11_846 (.fluid_in(k_11_846), .fluid_out(k_10_423), .air_in(c_11_0));
valve v_11_847 (.fluid_in(k_11_847), .fluid_out(k_10_423), .air_in(c_11_1));
valve v_11_848 (.fluid_in(k_11_848), .fluid_out(k_10_424), .air_in(c_11_0));
valve v_11_849 (.fluid_in(k_11_849), .fluid_out(k_10_424), .air_in(c_11_1));
valve v_11_850 (.fluid_in(k_11_850), .fluid_out(k_10_425), .air_in(c_11_0));
valve v_11_851 (.fluid_in(k_11_851), .fluid_out(k_10_425), .air_in(c_11_1));
valve v_11_852 (.fluid_in(k_11_852), .fluid_out(k_10_426), .air_in(c_11_0));
valve v_11_853 (.fluid_in(k_11_853), .fluid_out(k_10_426), .air_in(c_11_1));
valve v_11_854 (.fluid_in(k_11_854), .fluid_out(k_10_427), .air_in(c_11_0));
valve v_11_855 (.fluid_in(k_11_855), .fluid_out(k_10_427), .air_in(c_11_1));
valve v_11_856 (.fluid_in(k_11_856), .fluid_out(k_10_428), .air_in(c_11_0));
valve v_11_857 (.fluid_in(k_11_857), .fluid_out(k_10_428), .air_in(c_11_1));
valve v_11_858 (.fluid_in(k_11_858), .fluid_out(k_10_429), .air_in(c_11_0));
valve v_11_859 (.fluid_in(k_11_859), .fluid_out(k_10_429), .air_in(c_11_1));
valve v_11_860 (.fluid_in(k_11_860), .fluid_out(k_10_430), .air_in(c_11_0));
valve v_11_861 (.fluid_in(k_11_861), .fluid_out(k_10_430), .air_in(c_11_1));
valve v_11_862 (.fluid_in(k_11_862), .fluid_out(k_10_431), .air_in(c_11_0));
valve v_11_863 (.fluid_in(k_11_863), .fluid_out(k_10_431), .air_in(c_11_1));
valve v_11_864 (.fluid_in(k_11_864), .fluid_out(k_10_432), .air_in(c_11_0));
valve v_11_865 (.fluid_in(k_11_865), .fluid_out(k_10_432), .air_in(c_11_1));
valve v_11_866 (.fluid_in(k_11_866), .fluid_out(k_10_433), .air_in(c_11_0));
valve v_11_867 (.fluid_in(k_11_867), .fluid_out(k_10_433), .air_in(c_11_1));
valve v_11_868 (.fluid_in(k_11_868), .fluid_out(k_10_434), .air_in(c_11_0));
valve v_11_869 (.fluid_in(k_11_869), .fluid_out(k_10_434), .air_in(c_11_1));
valve v_11_870 (.fluid_in(k_11_870), .fluid_out(k_10_435), .air_in(c_11_0));
valve v_11_871 (.fluid_in(k_11_871), .fluid_out(k_10_435), .air_in(c_11_1));
valve v_11_872 (.fluid_in(k_11_872), .fluid_out(k_10_436), .air_in(c_11_0));
valve v_11_873 (.fluid_in(k_11_873), .fluid_out(k_10_436), .air_in(c_11_1));
valve v_11_874 (.fluid_in(k_11_874), .fluid_out(k_10_437), .air_in(c_11_0));
valve v_11_875 (.fluid_in(k_11_875), .fluid_out(k_10_437), .air_in(c_11_1));
valve v_11_876 (.fluid_in(k_11_876), .fluid_out(k_10_438), .air_in(c_11_0));
valve v_11_877 (.fluid_in(k_11_877), .fluid_out(k_10_438), .air_in(c_11_1));
valve v_11_878 (.fluid_in(k_11_878), .fluid_out(k_10_439), .air_in(c_11_0));
valve v_11_879 (.fluid_in(k_11_879), .fluid_out(k_10_439), .air_in(c_11_1));
valve v_11_880 (.fluid_in(k_11_880), .fluid_out(k_10_440), .air_in(c_11_0));
valve v_11_881 (.fluid_in(k_11_881), .fluid_out(k_10_440), .air_in(c_11_1));
valve v_11_882 (.fluid_in(k_11_882), .fluid_out(k_10_441), .air_in(c_11_0));
valve v_11_883 (.fluid_in(k_11_883), .fluid_out(k_10_441), .air_in(c_11_1));
valve v_11_884 (.fluid_in(k_11_884), .fluid_out(k_10_442), .air_in(c_11_0));
valve v_11_885 (.fluid_in(k_11_885), .fluid_out(k_10_442), .air_in(c_11_1));
valve v_11_886 (.fluid_in(k_11_886), .fluid_out(k_10_443), .air_in(c_11_0));
valve v_11_887 (.fluid_in(k_11_887), .fluid_out(k_10_443), .air_in(c_11_1));
valve v_11_888 (.fluid_in(k_11_888), .fluid_out(k_10_444), .air_in(c_11_0));
valve v_11_889 (.fluid_in(k_11_889), .fluid_out(k_10_444), .air_in(c_11_1));
valve v_11_890 (.fluid_in(k_11_890), .fluid_out(k_10_445), .air_in(c_11_0));
valve v_11_891 (.fluid_in(k_11_891), .fluid_out(k_10_445), .air_in(c_11_1));
valve v_11_892 (.fluid_in(k_11_892), .fluid_out(k_10_446), .air_in(c_11_0));
valve v_11_893 (.fluid_in(k_11_893), .fluid_out(k_10_446), .air_in(c_11_1));
valve v_11_894 (.fluid_in(k_11_894), .fluid_out(k_10_447), .air_in(c_11_0));
valve v_11_895 (.fluid_in(k_11_895), .fluid_out(k_10_447), .air_in(c_11_1));
valve v_11_896 (.fluid_in(k_11_896), .fluid_out(k_10_448), .air_in(c_11_0));
valve v_11_897 (.fluid_in(k_11_897), .fluid_out(k_10_448), .air_in(c_11_1));
valve v_11_898 (.fluid_in(k_11_898), .fluid_out(k_10_449), .air_in(c_11_0));
valve v_11_899 (.fluid_in(k_11_899), .fluid_out(k_10_449), .air_in(c_11_1));
valve v_11_900 (.fluid_in(k_11_900), .fluid_out(k_10_450), .air_in(c_11_0));
valve v_11_901 (.fluid_in(k_11_901), .fluid_out(k_10_450), .air_in(c_11_1));
valve v_11_902 (.fluid_in(k_11_902), .fluid_out(k_10_451), .air_in(c_11_0));
valve v_11_903 (.fluid_in(k_11_903), .fluid_out(k_10_451), .air_in(c_11_1));
valve v_11_904 (.fluid_in(k_11_904), .fluid_out(k_10_452), .air_in(c_11_0));
valve v_11_905 (.fluid_in(k_11_905), .fluid_out(k_10_452), .air_in(c_11_1));
valve v_11_906 (.fluid_in(k_11_906), .fluid_out(k_10_453), .air_in(c_11_0));
valve v_11_907 (.fluid_in(k_11_907), .fluid_out(k_10_453), .air_in(c_11_1));
valve v_11_908 (.fluid_in(k_11_908), .fluid_out(k_10_454), .air_in(c_11_0));
valve v_11_909 (.fluid_in(k_11_909), .fluid_out(k_10_454), .air_in(c_11_1));
valve v_11_910 (.fluid_in(k_11_910), .fluid_out(k_10_455), .air_in(c_11_0));
valve v_11_911 (.fluid_in(k_11_911), .fluid_out(k_10_455), .air_in(c_11_1));
valve v_11_912 (.fluid_in(k_11_912), .fluid_out(k_10_456), .air_in(c_11_0));
valve v_11_913 (.fluid_in(k_11_913), .fluid_out(k_10_456), .air_in(c_11_1));
valve v_11_914 (.fluid_in(k_11_914), .fluid_out(k_10_457), .air_in(c_11_0));
valve v_11_915 (.fluid_in(k_11_915), .fluid_out(k_10_457), .air_in(c_11_1));
valve v_11_916 (.fluid_in(k_11_916), .fluid_out(k_10_458), .air_in(c_11_0));
valve v_11_917 (.fluid_in(k_11_917), .fluid_out(k_10_458), .air_in(c_11_1));
valve v_11_918 (.fluid_in(k_11_918), .fluid_out(k_10_459), .air_in(c_11_0));
valve v_11_919 (.fluid_in(k_11_919), .fluid_out(k_10_459), .air_in(c_11_1));
valve v_11_920 (.fluid_in(k_11_920), .fluid_out(k_10_460), .air_in(c_11_0));
valve v_11_921 (.fluid_in(k_11_921), .fluid_out(k_10_460), .air_in(c_11_1));
valve v_11_922 (.fluid_in(k_11_922), .fluid_out(k_10_461), .air_in(c_11_0));
valve v_11_923 (.fluid_in(k_11_923), .fluid_out(k_10_461), .air_in(c_11_1));
valve v_11_924 (.fluid_in(k_11_924), .fluid_out(k_10_462), .air_in(c_11_0));
valve v_11_925 (.fluid_in(k_11_925), .fluid_out(k_10_462), .air_in(c_11_1));
valve v_11_926 (.fluid_in(k_11_926), .fluid_out(k_10_463), .air_in(c_11_0));
valve v_11_927 (.fluid_in(k_11_927), .fluid_out(k_10_463), .air_in(c_11_1));
valve v_11_928 (.fluid_in(k_11_928), .fluid_out(k_10_464), .air_in(c_11_0));
valve v_11_929 (.fluid_in(k_11_929), .fluid_out(k_10_464), .air_in(c_11_1));
valve v_11_930 (.fluid_in(k_11_930), .fluid_out(k_10_465), .air_in(c_11_0));
valve v_11_931 (.fluid_in(k_11_931), .fluid_out(k_10_465), .air_in(c_11_1));
valve v_11_932 (.fluid_in(k_11_932), .fluid_out(k_10_466), .air_in(c_11_0));
valve v_11_933 (.fluid_in(k_11_933), .fluid_out(k_10_466), .air_in(c_11_1));
valve v_11_934 (.fluid_in(k_11_934), .fluid_out(k_10_467), .air_in(c_11_0));
valve v_11_935 (.fluid_in(k_11_935), .fluid_out(k_10_467), .air_in(c_11_1));
valve v_11_936 (.fluid_in(k_11_936), .fluid_out(k_10_468), .air_in(c_11_0));
valve v_11_937 (.fluid_in(k_11_937), .fluid_out(k_10_468), .air_in(c_11_1));
valve v_11_938 (.fluid_in(k_11_938), .fluid_out(k_10_469), .air_in(c_11_0));
valve v_11_939 (.fluid_in(k_11_939), .fluid_out(k_10_469), .air_in(c_11_1));
valve v_11_940 (.fluid_in(k_11_940), .fluid_out(k_10_470), .air_in(c_11_0));
valve v_11_941 (.fluid_in(k_11_941), .fluid_out(k_10_470), .air_in(c_11_1));
valve v_11_942 (.fluid_in(k_11_942), .fluid_out(k_10_471), .air_in(c_11_0));
valve v_11_943 (.fluid_in(k_11_943), .fluid_out(k_10_471), .air_in(c_11_1));
valve v_11_944 (.fluid_in(k_11_944), .fluid_out(k_10_472), .air_in(c_11_0));
valve v_11_945 (.fluid_in(k_11_945), .fluid_out(k_10_472), .air_in(c_11_1));
valve v_11_946 (.fluid_in(k_11_946), .fluid_out(k_10_473), .air_in(c_11_0));
valve v_11_947 (.fluid_in(k_11_947), .fluid_out(k_10_473), .air_in(c_11_1));
valve v_11_948 (.fluid_in(k_11_948), .fluid_out(k_10_474), .air_in(c_11_0));
valve v_11_949 (.fluid_in(k_11_949), .fluid_out(k_10_474), .air_in(c_11_1));
valve v_11_950 (.fluid_in(k_11_950), .fluid_out(k_10_475), .air_in(c_11_0));
valve v_11_951 (.fluid_in(k_11_951), .fluid_out(k_10_475), .air_in(c_11_1));
valve v_11_952 (.fluid_in(k_11_952), .fluid_out(k_10_476), .air_in(c_11_0));
valve v_11_953 (.fluid_in(k_11_953), .fluid_out(k_10_476), .air_in(c_11_1));
valve v_11_954 (.fluid_in(k_11_954), .fluid_out(k_10_477), .air_in(c_11_0));
valve v_11_955 (.fluid_in(k_11_955), .fluid_out(k_10_477), .air_in(c_11_1));
valve v_11_956 (.fluid_in(k_11_956), .fluid_out(k_10_478), .air_in(c_11_0));
valve v_11_957 (.fluid_in(k_11_957), .fluid_out(k_10_478), .air_in(c_11_1));
valve v_11_958 (.fluid_in(k_11_958), .fluid_out(k_10_479), .air_in(c_11_0));
valve v_11_959 (.fluid_in(k_11_959), .fluid_out(k_10_479), .air_in(c_11_1));
valve v_11_960 (.fluid_in(k_11_960), .fluid_out(k_10_480), .air_in(c_11_0));
valve v_11_961 (.fluid_in(k_11_961), .fluid_out(k_10_480), .air_in(c_11_1));
valve v_11_962 (.fluid_in(k_11_962), .fluid_out(k_10_481), .air_in(c_11_0));
valve v_11_963 (.fluid_in(k_11_963), .fluid_out(k_10_481), .air_in(c_11_1));
valve v_11_964 (.fluid_in(k_11_964), .fluid_out(k_10_482), .air_in(c_11_0));
valve v_11_965 (.fluid_in(k_11_965), .fluid_out(k_10_482), .air_in(c_11_1));
valve v_11_966 (.fluid_in(k_11_966), .fluid_out(k_10_483), .air_in(c_11_0));
valve v_11_967 (.fluid_in(k_11_967), .fluid_out(k_10_483), .air_in(c_11_1));
valve v_11_968 (.fluid_in(k_11_968), .fluid_out(k_10_484), .air_in(c_11_0));
valve v_11_969 (.fluid_in(k_11_969), .fluid_out(k_10_484), .air_in(c_11_1));
valve v_11_970 (.fluid_in(k_11_970), .fluid_out(k_10_485), .air_in(c_11_0));
valve v_11_971 (.fluid_in(k_11_971), .fluid_out(k_10_485), .air_in(c_11_1));
valve v_11_972 (.fluid_in(k_11_972), .fluid_out(k_10_486), .air_in(c_11_0));
valve v_11_973 (.fluid_in(k_11_973), .fluid_out(k_10_486), .air_in(c_11_1));
valve v_11_974 (.fluid_in(k_11_974), .fluid_out(k_10_487), .air_in(c_11_0));
valve v_11_975 (.fluid_in(k_11_975), .fluid_out(k_10_487), .air_in(c_11_1));
valve v_11_976 (.fluid_in(k_11_976), .fluid_out(k_10_488), .air_in(c_11_0));
valve v_11_977 (.fluid_in(k_11_977), .fluid_out(k_10_488), .air_in(c_11_1));
valve v_11_978 (.fluid_in(k_11_978), .fluid_out(k_10_489), .air_in(c_11_0));
valve v_11_979 (.fluid_in(k_11_979), .fluid_out(k_10_489), .air_in(c_11_1));
valve v_11_980 (.fluid_in(k_11_980), .fluid_out(k_10_490), .air_in(c_11_0));
valve v_11_981 (.fluid_in(k_11_981), .fluid_out(k_10_490), .air_in(c_11_1));
valve v_11_982 (.fluid_in(k_11_982), .fluid_out(k_10_491), .air_in(c_11_0));
valve v_11_983 (.fluid_in(k_11_983), .fluid_out(k_10_491), .air_in(c_11_1));
valve v_11_984 (.fluid_in(k_11_984), .fluid_out(k_10_492), .air_in(c_11_0));
valve v_11_985 (.fluid_in(k_11_985), .fluid_out(k_10_492), .air_in(c_11_1));
valve v_11_986 (.fluid_in(k_11_986), .fluid_out(k_10_493), .air_in(c_11_0));
valve v_11_987 (.fluid_in(k_11_987), .fluid_out(k_10_493), .air_in(c_11_1));
valve v_11_988 (.fluid_in(k_11_988), .fluid_out(k_10_494), .air_in(c_11_0));
valve v_11_989 (.fluid_in(k_11_989), .fluid_out(k_10_494), .air_in(c_11_1));
valve v_11_990 (.fluid_in(k_11_990), .fluid_out(k_10_495), .air_in(c_11_0));
valve v_11_991 (.fluid_in(k_11_991), .fluid_out(k_10_495), .air_in(c_11_1));
valve v_11_992 (.fluid_in(k_11_992), .fluid_out(k_10_496), .air_in(c_11_0));
valve v_11_993 (.fluid_in(k_11_993), .fluid_out(k_10_496), .air_in(c_11_1));
valve v_11_994 (.fluid_in(k_11_994), .fluid_out(k_10_497), .air_in(c_11_0));
valve v_11_995 (.fluid_in(k_11_995), .fluid_out(k_10_497), .air_in(c_11_1));
valve v_11_996 (.fluid_in(k_11_996), .fluid_out(k_10_498), .air_in(c_11_0));
valve v_11_997 (.fluid_in(k_11_997), .fluid_out(k_10_498), .air_in(c_11_1));
valve v_11_998 (.fluid_in(k_11_998), .fluid_out(k_10_499), .air_in(c_11_0));
valve v_11_999 (.fluid_in(k_11_999), .fluid_out(k_10_499), .air_in(c_11_1));
valve v_11_1000 (.fluid_in(k_11_1000), .fluid_out(k_10_500), .air_in(c_11_0));
valve v_11_1001 (.fluid_in(k_11_1001), .fluid_out(k_10_500), .air_in(c_11_1));
valve v_11_1002 (.fluid_in(k_11_1002), .fluid_out(k_10_501), .air_in(c_11_0));
valve v_11_1003 (.fluid_in(k_11_1003), .fluid_out(k_10_501), .air_in(c_11_1));
valve v_11_1004 (.fluid_in(k_11_1004), .fluid_out(k_10_502), .air_in(c_11_0));
valve v_11_1005 (.fluid_in(k_11_1005), .fluid_out(k_10_502), .air_in(c_11_1));
valve v_11_1006 (.fluid_in(k_11_1006), .fluid_out(k_10_503), .air_in(c_11_0));
valve v_11_1007 (.fluid_in(k_11_1007), .fluid_out(k_10_503), .air_in(c_11_1));
valve v_11_1008 (.fluid_in(k_11_1008), .fluid_out(k_10_504), .air_in(c_11_0));
valve v_11_1009 (.fluid_in(k_11_1009), .fluid_out(k_10_504), .air_in(c_11_1));
valve v_11_1010 (.fluid_in(k_11_1010), .fluid_out(k_10_505), .air_in(c_11_0));
valve v_11_1011 (.fluid_in(k_11_1011), .fluid_out(k_10_505), .air_in(c_11_1));
valve v_11_1012 (.fluid_in(k_11_1012), .fluid_out(k_10_506), .air_in(c_11_0));
valve v_11_1013 (.fluid_in(k_11_1013), .fluid_out(k_10_506), .air_in(c_11_1));
valve v_11_1014 (.fluid_in(k_11_1014), .fluid_out(k_10_507), .air_in(c_11_0));
valve v_11_1015 (.fluid_in(k_11_1015), .fluid_out(k_10_507), .air_in(c_11_1));
valve v_11_1016 (.fluid_in(k_11_1016), .fluid_out(k_10_508), .air_in(c_11_0));
valve v_11_1017 (.fluid_in(k_11_1017), .fluid_out(k_10_508), .air_in(c_11_1));
valve v_11_1018 (.fluid_in(k_11_1018), .fluid_out(k_10_509), .air_in(c_11_0));
valve v_11_1019 (.fluid_in(k_11_1019), .fluid_out(k_10_509), .air_in(c_11_1));
valve v_11_1020 (.fluid_in(k_11_1020), .fluid_out(k_10_510), .air_in(c_11_0));
valve v_11_1021 (.fluid_in(k_11_1021), .fluid_out(k_10_510), .air_in(c_11_1));
valve v_11_1022 (.fluid_in(k_11_1022), .fluid_out(k_10_511), .air_in(c_11_0));
valve v_11_1023 (.fluid_in(k_11_1023), .fluid_out(k_10_511), .air_in(c_11_1));
valve v_11_1024 (.fluid_in(k_11_1024), .fluid_out(k_10_512), .air_in(c_11_0));
valve v_11_1025 (.fluid_in(k_11_1025), .fluid_out(k_10_512), .air_in(c_11_1));
valve v_11_1026 (.fluid_in(k_11_1026), .fluid_out(k_10_513), .air_in(c_11_0));
valve v_11_1027 (.fluid_in(k_11_1027), .fluid_out(k_10_513), .air_in(c_11_1));
valve v_11_1028 (.fluid_in(k_11_1028), .fluid_out(k_10_514), .air_in(c_11_0));
valve v_11_1029 (.fluid_in(k_11_1029), .fluid_out(k_10_514), .air_in(c_11_1));
valve v_11_1030 (.fluid_in(k_11_1030), .fluid_out(k_10_515), .air_in(c_11_0));
valve v_11_1031 (.fluid_in(k_11_1031), .fluid_out(k_10_515), .air_in(c_11_1));
valve v_11_1032 (.fluid_in(k_11_1032), .fluid_out(k_10_516), .air_in(c_11_0));
valve v_11_1033 (.fluid_in(k_11_1033), .fluid_out(k_10_516), .air_in(c_11_1));
valve v_11_1034 (.fluid_in(k_11_1034), .fluid_out(k_10_517), .air_in(c_11_0));
valve v_11_1035 (.fluid_in(k_11_1035), .fluid_out(k_10_517), .air_in(c_11_1));
valve v_11_1036 (.fluid_in(k_11_1036), .fluid_out(k_10_518), .air_in(c_11_0));
valve v_11_1037 (.fluid_in(k_11_1037), .fluid_out(k_10_518), .air_in(c_11_1));
valve v_11_1038 (.fluid_in(k_11_1038), .fluid_out(k_10_519), .air_in(c_11_0));
valve v_11_1039 (.fluid_in(k_11_1039), .fluid_out(k_10_519), .air_in(c_11_1));
valve v_11_1040 (.fluid_in(k_11_1040), .fluid_out(k_10_520), .air_in(c_11_0));
valve v_11_1041 (.fluid_in(k_11_1041), .fluid_out(k_10_520), .air_in(c_11_1));
valve v_11_1042 (.fluid_in(k_11_1042), .fluid_out(k_10_521), .air_in(c_11_0));
valve v_11_1043 (.fluid_in(k_11_1043), .fluid_out(k_10_521), .air_in(c_11_1));
valve v_11_1044 (.fluid_in(k_11_1044), .fluid_out(k_10_522), .air_in(c_11_0));
valve v_11_1045 (.fluid_in(k_11_1045), .fluid_out(k_10_522), .air_in(c_11_1));
valve v_11_1046 (.fluid_in(k_11_1046), .fluid_out(k_10_523), .air_in(c_11_0));
valve v_11_1047 (.fluid_in(k_11_1047), .fluid_out(k_10_523), .air_in(c_11_1));
valve v_11_1048 (.fluid_in(k_11_1048), .fluid_out(k_10_524), .air_in(c_11_0));
valve v_11_1049 (.fluid_in(k_11_1049), .fluid_out(k_10_524), .air_in(c_11_1));
valve v_11_1050 (.fluid_in(k_11_1050), .fluid_out(k_10_525), .air_in(c_11_0));
valve v_11_1051 (.fluid_in(k_11_1051), .fluid_out(k_10_525), .air_in(c_11_1));
valve v_11_1052 (.fluid_in(k_11_1052), .fluid_out(k_10_526), .air_in(c_11_0));
valve v_11_1053 (.fluid_in(k_11_1053), .fluid_out(k_10_526), .air_in(c_11_1));
valve v_11_1054 (.fluid_in(k_11_1054), .fluid_out(k_10_527), .air_in(c_11_0));
valve v_11_1055 (.fluid_in(k_11_1055), .fluid_out(k_10_527), .air_in(c_11_1));
valve v_11_1056 (.fluid_in(k_11_1056), .fluid_out(k_10_528), .air_in(c_11_0));
valve v_11_1057 (.fluid_in(k_11_1057), .fluid_out(k_10_528), .air_in(c_11_1));
valve v_11_1058 (.fluid_in(k_11_1058), .fluid_out(k_10_529), .air_in(c_11_0));
valve v_11_1059 (.fluid_in(k_11_1059), .fluid_out(k_10_529), .air_in(c_11_1));
valve v_11_1060 (.fluid_in(k_11_1060), .fluid_out(k_10_530), .air_in(c_11_0));
valve v_11_1061 (.fluid_in(k_11_1061), .fluid_out(k_10_530), .air_in(c_11_1));
valve v_11_1062 (.fluid_in(k_11_1062), .fluid_out(k_10_531), .air_in(c_11_0));
valve v_11_1063 (.fluid_in(k_11_1063), .fluid_out(k_10_531), .air_in(c_11_1));
valve v_11_1064 (.fluid_in(k_11_1064), .fluid_out(k_10_532), .air_in(c_11_0));
valve v_11_1065 (.fluid_in(k_11_1065), .fluid_out(k_10_532), .air_in(c_11_1));
valve v_11_1066 (.fluid_in(k_11_1066), .fluid_out(k_10_533), .air_in(c_11_0));
valve v_11_1067 (.fluid_in(k_11_1067), .fluid_out(k_10_533), .air_in(c_11_1));
valve v_11_1068 (.fluid_in(k_11_1068), .fluid_out(k_10_534), .air_in(c_11_0));
valve v_11_1069 (.fluid_in(k_11_1069), .fluid_out(k_10_534), .air_in(c_11_1));
valve v_11_1070 (.fluid_in(k_11_1070), .fluid_out(k_10_535), .air_in(c_11_0));
valve v_11_1071 (.fluid_in(k_11_1071), .fluid_out(k_10_535), .air_in(c_11_1));
valve v_11_1072 (.fluid_in(k_11_1072), .fluid_out(k_10_536), .air_in(c_11_0));
valve v_11_1073 (.fluid_in(k_11_1073), .fluid_out(k_10_536), .air_in(c_11_1));
valve v_11_1074 (.fluid_in(k_11_1074), .fluid_out(k_10_537), .air_in(c_11_0));
valve v_11_1075 (.fluid_in(k_11_1075), .fluid_out(k_10_537), .air_in(c_11_1));
valve v_11_1076 (.fluid_in(k_11_1076), .fluid_out(k_10_538), .air_in(c_11_0));
valve v_11_1077 (.fluid_in(k_11_1077), .fluid_out(k_10_538), .air_in(c_11_1));
valve v_11_1078 (.fluid_in(k_11_1078), .fluid_out(k_10_539), .air_in(c_11_0));
valve v_11_1079 (.fluid_in(k_11_1079), .fluid_out(k_10_539), .air_in(c_11_1));
valve v_11_1080 (.fluid_in(k_11_1080), .fluid_out(k_10_540), .air_in(c_11_0));
valve v_11_1081 (.fluid_in(k_11_1081), .fluid_out(k_10_540), .air_in(c_11_1));
valve v_11_1082 (.fluid_in(k_11_1082), .fluid_out(k_10_541), .air_in(c_11_0));
valve v_11_1083 (.fluid_in(k_11_1083), .fluid_out(k_10_541), .air_in(c_11_1));
valve v_11_1084 (.fluid_in(k_11_1084), .fluid_out(k_10_542), .air_in(c_11_0));
valve v_11_1085 (.fluid_in(k_11_1085), .fluid_out(k_10_542), .air_in(c_11_1));
valve v_11_1086 (.fluid_in(k_11_1086), .fluid_out(k_10_543), .air_in(c_11_0));
valve v_11_1087 (.fluid_in(k_11_1087), .fluid_out(k_10_543), .air_in(c_11_1));
valve v_11_1088 (.fluid_in(k_11_1088), .fluid_out(k_10_544), .air_in(c_11_0));
valve v_11_1089 (.fluid_in(k_11_1089), .fluid_out(k_10_544), .air_in(c_11_1));
valve v_11_1090 (.fluid_in(k_11_1090), .fluid_out(k_10_545), .air_in(c_11_0));
valve v_11_1091 (.fluid_in(k_11_1091), .fluid_out(k_10_545), .air_in(c_11_1));
valve v_11_1092 (.fluid_in(k_11_1092), .fluid_out(k_10_546), .air_in(c_11_0));
valve v_11_1093 (.fluid_in(k_11_1093), .fluid_out(k_10_546), .air_in(c_11_1));
valve v_11_1094 (.fluid_in(k_11_1094), .fluid_out(k_10_547), .air_in(c_11_0));
valve v_11_1095 (.fluid_in(k_11_1095), .fluid_out(k_10_547), .air_in(c_11_1));
valve v_11_1096 (.fluid_in(k_11_1096), .fluid_out(k_10_548), .air_in(c_11_0));
valve v_11_1097 (.fluid_in(k_11_1097), .fluid_out(k_10_548), .air_in(c_11_1));
valve v_11_1098 (.fluid_in(k_11_1098), .fluid_out(k_10_549), .air_in(c_11_0));
valve v_11_1099 (.fluid_in(k_11_1099), .fluid_out(k_10_549), .air_in(c_11_1));
valve v_11_1100 (.fluid_in(k_11_1100), .fluid_out(k_10_550), .air_in(c_11_0));
valve v_11_1101 (.fluid_in(k_11_1101), .fluid_out(k_10_550), .air_in(c_11_1));
valve v_11_1102 (.fluid_in(k_11_1102), .fluid_out(k_10_551), .air_in(c_11_0));
valve v_11_1103 (.fluid_in(k_11_1103), .fluid_out(k_10_551), .air_in(c_11_1));
valve v_11_1104 (.fluid_in(k_11_1104), .fluid_out(k_10_552), .air_in(c_11_0));
valve v_11_1105 (.fluid_in(k_11_1105), .fluid_out(k_10_552), .air_in(c_11_1));
valve v_11_1106 (.fluid_in(k_11_1106), .fluid_out(k_10_553), .air_in(c_11_0));
valve v_11_1107 (.fluid_in(k_11_1107), .fluid_out(k_10_553), .air_in(c_11_1));
valve v_11_1108 (.fluid_in(k_11_1108), .fluid_out(k_10_554), .air_in(c_11_0));
valve v_11_1109 (.fluid_in(k_11_1109), .fluid_out(k_10_554), .air_in(c_11_1));
valve v_11_1110 (.fluid_in(k_11_1110), .fluid_out(k_10_555), .air_in(c_11_0));
valve v_11_1111 (.fluid_in(k_11_1111), .fluid_out(k_10_555), .air_in(c_11_1));
valve v_11_1112 (.fluid_in(k_11_1112), .fluid_out(k_10_556), .air_in(c_11_0));
valve v_11_1113 (.fluid_in(k_11_1113), .fluid_out(k_10_556), .air_in(c_11_1));
valve v_11_1114 (.fluid_in(k_11_1114), .fluid_out(k_10_557), .air_in(c_11_0));
valve v_11_1115 (.fluid_in(k_11_1115), .fluid_out(k_10_557), .air_in(c_11_1));
valve v_11_1116 (.fluid_in(k_11_1116), .fluid_out(k_10_558), .air_in(c_11_0));
valve v_11_1117 (.fluid_in(k_11_1117), .fluid_out(k_10_558), .air_in(c_11_1));
valve v_11_1118 (.fluid_in(k_11_1118), .fluid_out(k_10_559), .air_in(c_11_0));
valve v_11_1119 (.fluid_in(k_11_1119), .fluid_out(k_10_559), .air_in(c_11_1));
valve v_11_1120 (.fluid_in(k_11_1120), .fluid_out(k_10_560), .air_in(c_11_0));
valve v_11_1121 (.fluid_in(k_11_1121), .fluid_out(k_10_560), .air_in(c_11_1));
valve v_11_1122 (.fluid_in(k_11_1122), .fluid_out(k_10_561), .air_in(c_11_0));
valve v_11_1123 (.fluid_in(k_11_1123), .fluid_out(k_10_561), .air_in(c_11_1));
valve v_11_1124 (.fluid_in(k_11_1124), .fluid_out(k_10_562), .air_in(c_11_0));
valve v_11_1125 (.fluid_in(k_11_1125), .fluid_out(k_10_562), .air_in(c_11_1));
valve v_11_1126 (.fluid_in(k_11_1126), .fluid_out(k_10_563), .air_in(c_11_0));
valve v_11_1127 (.fluid_in(k_11_1127), .fluid_out(k_10_563), .air_in(c_11_1));
valve v_11_1128 (.fluid_in(k_11_1128), .fluid_out(k_10_564), .air_in(c_11_0));
valve v_11_1129 (.fluid_in(k_11_1129), .fluid_out(k_10_564), .air_in(c_11_1));
valve v_11_1130 (.fluid_in(k_11_1130), .fluid_out(k_10_565), .air_in(c_11_0));
valve v_11_1131 (.fluid_in(k_11_1131), .fluid_out(k_10_565), .air_in(c_11_1));
valve v_11_1132 (.fluid_in(k_11_1132), .fluid_out(k_10_566), .air_in(c_11_0));
valve v_11_1133 (.fluid_in(k_11_1133), .fluid_out(k_10_566), .air_in(c_11_1));
valve v_11_1134 (.fluid_in(k_11_1134), .fluid_out(k_10_567), .air_in(c_11_0));
valve v_11_1135 (.fluid_in(k_11_1135), .fluid_out(k_10_567), .air_in(c_11_1));
valve v_11_1136 (.fluid_in(k_11_1136), .fluid_out(k_10_568), .air_in(c_11_0));
valve v_11_1137 (.fluid_in(k_11_1137), .fluid_out(k_10_568), .air_in(c_11_1));
valve v_11_1138 (.fluid_in(k_11_1138), .fluid_out(k_10_569), .air_in(c_11_0));
valve v_11_1139 (.fluid_in(k_11_1139), .fluid_out(k_10_569), .air_in(c_11_1));
valve v_11_1140 (.fluid_in(k_11_1140), .fluid_out(k_10_570), .air_in(c_11_0));
valve v_11_1141 (.fluid_in(k_11_1141), .fluid_out(k_10_570), .air_in(c_11_1));
valve v_11_1142 (.fluid_in(k_11_1142), .fluid_out(k_10_571), .air_in(c_11_0));
valve v_11_1143 (.fluid_in(k_11_1143), .fluid_out(k_10_571), .air_in(c_11_1));
valve v_11_1144 (.fluid_in(k_11_1144), .fluid_out(k_10_572), .air_in(c_11_0));
valve v_11_1145 (.fluid_in(k_11_1145), .fluid_out(k_10_572), .air_in(c_11_1));
valve v_11_1146 (.fluid_in(k_11_1146), .fluid_out(k_10_573), .air_in(c_11_0));
valve v_11_1147 (.fluid_in(k_11_1147), .fluid_out(k_10_573), .air_in(c_11_1));
valve v_11_1148 (.fluid_in(k_11_1148), .fluid_out(k_10_574), .air_in(c_11_0));
valve v_11_1149 (.fluid_in(k_11_1149), .fluid_out(k_10_574), .air_in(c_11_1));
valve v_11_1150 (.fluid_in(k_11_1150), .fluid_out(k_10_575), .air_in(c_11_0));
valve v_11_1151 (.fluid_in(k_11_1151), .fluid_out(k_10_575), .air_in(c_11_1));
valve v_11_1152 (.fluid_in(k_11_1152), .fluid_out(k_10_576), .air_in(c_11_0));
valve v_11_1153 (.fluid_in(k_11_1153), .fluid_out(k_10_576), .air_in(c_11_1));
valve v_11_1154 (.fluid_in(k_11_1154), .fluid_out(k_10_577), .air_in(c_11_0));
valve v_11_1155 (.fluid_in(k_11_1155), .fluid_out(k_10_577), .air_in(c_11_1));
valve v_11_1156 (.fluid_in(k_11_1156), .fluid_out(k_10_578), .air_in(c_11_0));
valve v_11_1157 (.fluid_in(k_11_1157), .fluid_out(k_10_578), .air_in(c_11_1));
valve v_11_1158 (.fluid_in(k_11_1158), .fluid_out(k_10_579), .air_in(c_11_0));
valve v_11_1159 (.fluid_in(k_11_1159), .fluid_out(k_10_579), .air_in(c_11_1));
valve v_11_1160 (.fluid_in(k_11_1160), .fluid_out(k_10_580), .air_in(c_11_0));
valve v_11_1161 (.fluid_in(k_11_1161), .fluid_out(k_10_580), .air_in(c_11_1));
valve v_11_1162 (.fluid_in(k_11_1162), .fluid_out(k_10_581), .air_in(c_11_0));
valve v_11_1163 (.fluid_in(k_11_1163), .fluid_out(k_10_581), .air_in(c_11_1));
valve v_11_1164 (.fluid_in(k_11_1164), .fluid_out(k_10_582), .air_in(c_11_0));
valve v_11_1165 (.fluid_in(k_11_1165), .fluid_out(k_10_582), .air_in(c_11_1));
valve v_11_1166 (.fluid_in(k_11_1166), .fluid_out(k_10_583), .air_in(c_11_0));
valve v_11_1167 (.fluid_in(k_11_1167), .fluid_out(k_10_583), .air_in(c_11_1));
valve v_11_1168 (.fluid_in(k_11_1168), .fluid_out(k_10_584), .air_in(c_11_0));
valve v_11_1169 (.fluid_in(k_11_1169), .fluid_out(k_10_584), .air_in(c_11_1));
valve v_11_1170 (.fluid_in(k_11_1170), .fluid_out(k_10_585), .air_in(c_11_0));
valve v_11_1171 (.fluid_in(k_11_1171), .fluid_out(k_10_585), .air_in(c_11_1));
valve v_11_1172 (.fluid_in(k_11_1172), .fluid_out(k_10_586), .air_in(c_11_0));
valve v_11_1173 (.fluid_in(k_11_1173), .fluid_out(k_10_586), .air_in(c_11_1));
valve v_11_1174 (.fluid_in(k_11_1174), .fluid_out(k_10_587), .air_in(c_11_0));
valve v_11_1175 (.fluid_in(k_11_1175), .fluid_out(k_10_587), .air_in(c_11_1));
valve v_11_1176 (.fluid_in(k_11_1176), .fluid_out(k_10_588), .air_in(c_11_0));
valve v_11_1177 (.fluid_in(k_11_1177), .fluid_out(k_10_588), .air_in(c_11_1));
valve v_11_1178 (.fluid_in(k_11_1178), .fluid_out(k_10_589), .air_in(c_11_0));
valve v_11_1179 (.fluid_in(k_11_1179), .fluid_out(k_10_589), .air_in(c_11_1));
valve v_11_1180 (.fluid_in(k_11_1180), .fluid_out(k_10_590), .air_in(c_11_0));
valve v_11_1181 (.fluid_in(k_11_1181), .fluid_out(k_10_590), .air_in(c_11_1));
valve v_11_1182 (.fluid_in(k_11_1182), .fluid_out(k_10_591), .air_in(c_11_0));
valve v_11_1183 (.fluid_in(k_11_1183), .fluid_out(k_10_591), .air_in(c_11_1));
valve v_11_1184 (.fluid_in(k_11_1184), .fluid_out(k_10_592), .air_in(c_11_0));
valve v_11_1185 (.fluid_in(k_11_1185), .fluid_out(k_10_592), .air_in(c_11_1));
valve v_11_1186 (.fluid_in(k_11_1186), .fluid_out(k_10_593), .air_in(c_11_0));
valve v_11_1187 (.fluid_in(k_11_1187), .fluid_out(k_10_593), .air_in(c_11_1));
valve v_11_1188 (.fluid_in(k_11_1188), .fluid_out(k_10_594), .air_in(c_11_0));
valve v_11_1189 (.fluid_in(k_11_1189), .fluid_out(k_10_594), .air_in(c_11_1));
valve v_11_1190 (.fluid_in(k_11_1190), .fluid_out(k_10_595), .air_in(c_11_0));
valve v_11_1191 (.fluid_in(k_11_1191), .fluid_out(k_10_595), .air_in(c_11_1));
valve v_11_1192 (.fluid_in(k_11_1192), .fluid_out(k_10_596), .air_in(c_11_0));
valve v_11_1193 (.fluid_in(k_11_1193), .fluid_out(k_10_596), .air_in(c_11_1));
valve v_11_1194 (.fluid_in(k_11_1194), .fluid_out(k_10_597), .air_in(c_11_0));
valve v_11_1195 (.fluid_in(k_11_1195), .fluid_out(k_10_597), .air_in(c_11_1));
valve v_11_1196 (.fluid_in(k_11_1196), .fluid_out(k_10_598), .air_in(c_11_0));
valve v_11_1197 (.fluid_in(k_11_1197), .fluid_out(k_10_598), .air_in(c_11_1));
valve v_11_1198 (.fluid_in(k_11_1198), .fluid_out(k_10_599), .air_in(c_11_0));
valve v_11_1199 (.fluid_in(k_11_1199), .fluid_out(k_10_599), .air_in(c_11_1));
valve v_11_1200 (.fluid_in(k_11_1200), .fluid_out(k_10_600), .air_in(c_11_0));
valve v_11_1201 (.fluid_in(k_11_1201), .fluid_out(k_10_600), .air_in(c_11_1));
valve v_11_1202 (.fluid_in(k_11_1202), .fluid_out(k_10_601), .air_in(c_11_0));
valve v_11_1203 (.fluid_in(k_11_1203), .fluid_out(k_10_601), .air_in(c_11_1));
valve v_11_1204 (.fluid_in(k_11_1204), .fluid_out(k_10_602), .air_in(c_11_0));
valve v_11_1205 (.fluid_in(k_11_1205), .fluid_out(k_10_602), .air_in(c_11_1));
valve v_11_1206 (.fluid_in(k_11_1206), .fluid_out(k_10_603), .air_in(c_11_0));
valve v_11_1207 (.fluid_in(k_11_1207), .fluid_out(k_10_603), .air_in(c_11_1));
valve v_11_1208 (.fluid_in(k_11_1208), .fluid_out(k_10_604), .air_in(c_11_0));
valve v_11_1209 (.fluid_in(k_11_1209), .fluid_out(k_10_604), .air_in(c_11_1));
valve v_11_1210 (.fluid_in(k_11_1210), .fluid_out(k_10_605), .air_in(c_11_0));
valve v_11_1211 (.fluid_in(k_11_1211), .fluid_out(k_10_605), .air_in(c_11_1));
valve v_11_1212 (.fluid_in(k_11_1212), .fluid_out(k_10_606), .air_in(c_11_0));
valve v_11_1213 (.fluid_in(k_11_1213), .fluid_out(k_10_606), .air_in(c_11_1));
valve v_11_1214 (.fluid_in(k_11_1214), .fluid_out(k_10_607), .air_in(c_11_0));
valve v_11_1215 (.fluid_in(k_11_1215), .fluid_out(k_10_607), .air_in(c_11_1));
valve v_11_1216 (.fluid_in(k_11_1216), .fluid_out(k_10_608), .air_in(c_11_0));
valve v_11_1217 (.fluid_in(k_11_1217), .fluid_out(k_10_608), .air_in(c_11_1));
valve v_11_1218 (.fluid_in(k_11_1218), .fluid_out(k_10_609), .air_in(c_11_0));
valve v_11_1219 (.fluid_in(k_11_1219), .fluid_out(k_10_609), .air_in(c_11_1));
valve v_11_1220 (.fluid_in(k_11_1220), .fluid_out(k_10_610), .air_in(c_11_0));
valve v_11_1221 (.fluid_in(k_11_1221), .fluid_out(k_10_610), .air_in(c_11_1));
valve v_11_1222 (.fluid_in(k_11_1222), .fluid_out(k_10_611), .air_in(c_11_0));
valve v_11_1223 (.fluid_in(k_11_1223), .fluid_out(k_10_611), .air_in(c_11_1));
valve v_11_1224 (.fluid_in(k_11_1224), .fluid_out(k_10_612), .air_in(c_11_0));
valve v_11_1225 (.fluid_in(k_11_1225), .fluid_out(k_10_612), .air_in(c_11_1));
valve v_11_1226 (.fluid_in(k_11_1226), .fluid_out(k_10_613), .air_in(c_11_0));
valve v_11_1227 (.fluid_in(k_11_1227), .fluid_out(k_10_613), .air_in(c_11_1));
valve v_11_1228 (.fluid_in(k_11_1228), .fluid_out(k_10_614), .air_in(c_11_0));
valve v_11_1229 (.fluid_in(k_11_1229), .fluid_out(k_10_614), .air_in(c_11_1));
valve v_11_1230 (.fluid_in(k_11_1230), .fluid_out(k_10_615), .air_in(c_11_0));
valve v_11_1231 (.fluid_in(k_11_1231), .fluid_out(k_10_615), .air_in(c_11_1));
valve v_11_1232 (.fluid_in(k_11_1232), .fluid_out(k_10_616), .air_in(c_11_0));
valve v_11_1233 (.fluid_in(k_11_1233), .fluid_out(k_10_616), .air_in(c_11_1));
valve v_11_1234 (.fluid_in(k_11_1234), .fluid_out(k_10_617), .air_in(c_11_0));
valve v_11_1235 (.fluid_in(k_11_1235), .fluid_out(k_10_617), .air_in(c_11_1));
valve v_11_1236 (.fluid_in(k_11_1236), .fluid_out(k_10_618), .air_in(c_11_0));
valve v_11_1237 (.fluid_in(k_11_1237), .fluid_out(k_10_618), .air_in(c_11_1));
valve v_11_1238 (.fluid_in(k_11_1238), .fluid_out(k_10_619), .air_in(c_11_0));
valve v_11_1239 (.fluid_in(k_11_1239), .fluid_out(k_10_619), .air_in(c_11_1));
valve v_11_1240 (.fluid_in(k_11_1240), .fluid_out(k_10_620), .air_in(c_11_0));
valve v_11_1241 (.fluid_in(k_11_1241), .fluid_out(k_10_620), .air_in(c_11_1));
valve v_11_1242 (.fluid_in(k_11_1242), .fluid_out(k_10_621), .air_in(c_11_0));
valve v_11_1243 (.fluid_in(k_11_1243), .fluid_out(k_10_621), .air_in(c_11_1));
valve v_11_1244 (.fluid_in(k_11_1244), .fluid_out(k_10_622), .air_in(c_11_0));
valve v_11_1245 (.fluid_in(k_11_1245), .fluid_out(k_10_622), .air_in(c_11_1));
valve v_11_1246 (.fluid_in(k_11_1246), .fluid_out(k_10_623), .air_in(c_11_0));
valve v_11_1247 (.fluid_in(k_11_1247), .fluid_out(k_10_623), .air_in(c_11_1));
valve v_11_1248 (.fluid_in(k_11_1248), .fluid_out(k_10_624), .air_in(c_11_0));
valve v_11_1249 (.fluid_in(k_11_1249), .fluid_out(k_10_624), .air_in(c_11_1));
valve v_11_1250 (.fluid_in(k_11_1250), .fluid_out(k_10_625), .air_in(c_11_0));
valve v_11_1251 (.fluid_in(k_11_1251), .fluid_out(k_10_625), .air_in(c_11_1));
valve v_11_1252 (.fluid_in(k_11_1252), .fluid_out(k_10_626), .air_in(c_11_0));
valve v_11_1253 (.fluid_in(k_11_1253), .fluid_out(k_10_626), .air_in(c_11_1));
valve v_11_1254 (.fluid_in(k_11_1254), .fluid_out(k_10_627), .air_in(c_11_0));
valve v_11_1255 (.fluid_in(k_11_1255), .fluid_out(k_10_627), .air_in(c_11_1));
valve v_11_1256 (.fluid_in(k_11_1256), .fluid_out(k_10_628), .air_in(c_11_0));
valve v_11_1257 (.fluid_in(k_11_1257), .fluid_out(k_10_628), .air_in(c_11_1));
valve v_11_1258 (.fluid_in(k_11_1258), .fluid_out(k_10_629), .air_in(c_11_0));
valve v_11_1259 (.fluid_in(k_11_1259), .fluid_out(k_10_629), .air_in(c_11_1));
valve v_11_1260 (.fluid_in(k_11_1260), .fluid_out(k_10_630), .air_in(c_11_0));
valve v_11_1261 (.fluid_in(k_11_1261), .fluid_out(k_10_630), .air_in(c_11_1));
valve v_11_1262 (.fluid_in(k_11_1262), .fluid_out(k_10_631), .air_in(c_11_0));
valve v_11_1263 (.fluid_in(k_11_1263), .fluid_out(k_10_631), .air_in(c_11_1));
valve v_11_1264 (.fluid_in(k_11_1264), .fluid_out(k_10_632), .air_in(c_11_0));
valve v_11_1265 (.fluid_in(k_11_1265), .fluid_out(k_10_632), .air_in(c_11_1));
valve v_11_1266 (.fluid_in(k_11_1266), .fluid_out(k_10_633), .air_in(c_11_0));
valve v_11_1267 (.fluid_in(k_11_1267), .fluid_out(k_10_633), .air_in(c_11_1));
valve v_11_1268 (.fluid_in(k_11_1268), .fluid_out(k_10_634), .air_in(c_11_0));
valve v_11_1269 (.fluid_in(k_11_1269), .fluid_out(k_10_634), .air_in(c_11_1));
valve v_11_1270 (.fluid_in(k_11_1270), .fluid_out(k_10_635), .air_in(c_11_0));
valve v_11_1271 (.fluid_in(k_11_1271), .fluid_out(k_10_635), .air_in(c_11_1));
valve v_11_1272 (.fluid_in(k_11_1272), .fluid_out(k_10_636), .air_in(c_11_0));
valve v_11_1273 (.fluid_in(k_11_1273), .fluid_out(k_10_636), .air_in(c_11_1));
valve v_11_1274 (.fluid_in(k_11_1274), .fluid_out(k_10_637), .air_in(c_11_0));
valve v_11_1275 (.fluid_in(k_11_1275), .fluid_out(k_10_637), .air_in(c_11_1));
valve v_11_1276 (.fluid_in(k_11_1276), .fluid_out(k_10_638), .air_in(c_11_0));
valve v_11_1277 (.fluid_in(k_11_1277), .fluid_out(k_10_638), .air_in(c_11_1));
valve v_11_1278 (.fluid_in(k_11_1278), .fluid_out(k_10_639), .air_in(c_11_0));
valve v_11_1279 (.fluid_in(k_11_1279), .fluid_out(k_10_639), .air_in(c_11_1));
valve v_11_1280 (.fluid_in(k_11_1280), .fluid_out(k_10_640), .air_in(c_11_0));
valve v_11_1281 (.fluid_in(k_11_1281), .fluid_out(k_10_640), .air_in(c_11_1));
valve v_11_1282 (.fluid_in(k_11_1282), .fluid_out(k_10_641), .air_in(c_11_0));
valve v_11_1283 (.fluid_in(k_11_1283), .fluid_out(k_10_641), .air_in(c_11_1));
valve v_11_1284 (.fluid_in(k_11_1284), .fluid_out(k_10_642), .air_in(c_11_0));
valve v_11_1285 (.fluid_in(k_11_1285), .fluid_out(k_10_642), .air_in(c_11_1));
valve v_11_1286 (.fluid_in(k_11_1286), .fluid_out(k_10_643), .air_in(c_11_0));
valve v_11_1287 (.fluid_in(k_11_1287), .fluid_out(k_10_643), .air_in(c_11_1));
valve v_11_1288 (.fluid_in(k_11_1288), .fluid_out(k_10_644), .air_in(c_11_0));
valve v_11_1289 (.fluid_in(k_11_1289), .fluid_out(k_10_644), .air_in(c_11_1));
valve v_11_1290 (.fluid_in(k_11_1290), .fluid_out(k_10_645), .air_in(c_11_0));
valve v_11_1291 (.fluid_in(k_11_1291), .fluid_out(k_10_645), .air_in(c_11_1));
valve v_11_1292 (.fluid_in(k_11_1292), .fluid_out(k_10_646), .air_in(c_11_0));
valve v_11_1293 (.fluid_in(k_11_1293), .fluid_out(k_10_646), .air_in(c_11_1));
valve v_11_1294 (.fluid_in(k_11_1294), .fluid_out(k_10_647), .air_in(c_11_0));
valve v_11_1295 (.fluid_in(k_11_1295), .fluid_out(k_10_647), .air_in(c_11_1));
valve v_11_1296 (.fluid_in(k_11_1296), .fluid_out(k_10_648), .air_in(c_11_0));
valve v_11_1297 (.fluid_in(k_11_1297), .fluid_out(k_10_648), .air_in(c_11_1));
valve v_11_1298 (.fluid_in(k_11_1298), .fluid_out(k_10_649), .air_in(c_11_0));
valve v_11_1299 (.fluid_in(k_11_1299), .fluid_out(k_10_649), .air_in(c_11_1));
valve v_11_1300 (.fluid_in(k_11_1300), .fluid_out(k_10_650), .air_in(c_11_0));
valve v_11_1301 (.fluid_in(k_11_1301), .fluid_out(k_10_650), .air_in(c_11_1));
valve v_11_1302 (.fluid_in(k_11_1302), .fluid_out(k_10_651), .air_in(c_11_0));
valve v_11_1303 (.fluid_in(k_11_1303), .fluid_out(k_10_651), .air_in(c_11_1));
valve v_11_1304 (.fluid_in(k_11_1304), .fluid_out(k_10_652), .air_in(c_11_0));
valve v_11_1305 (.fluid_in(k_11_1305), .fluid_out(k_10_652), .air_in(c_11_1));
valve v_11_1306 (.fluid_in(k_11_1306), .fluid_out(k_10_653), .air_in(c_11_0));
valve v_11_1307 (.fluid_in(k_11_1307), .fluid_out(k_10_653), .air_in(c_11_1));
valve v_11_1308 (.fluid_in(k_11_1308), .fluid_out(k_10_654), .air_in(c_11_0));
valve v_11_1309 (.fluid_in(k_11_1309), .fluid_out(k_10_654), .air_in(c_11_1));
valve v_11_1310 (.fluid_in(k_11_1310), .fluid_out(k_10_655), .air_in(c_11_0));
valve v_11_1311 (.fluid_in(k_11_1311), .fluid_out(k_10_655), .air_in(c_11_1));
valve v_11_1312 (.fluid_in(k_11_1312), .fluid_out(k_10_656), .air_in(c_11_0));
valve v_11_1313 (.fluid_in(k_11_1313), .fluid_out(k_10_656), .air_in(c_11_1));
valve v_11_1314 (.fluid_in(k_11_1314), .fluid_out(k_10_657), .air_in(c_11_0));
valve v_11_1315 (.fluid_in(k_11_1315), .fluid_out(k_10_657), .air_in(c_11_1));
valve v_11_1316 (.fluid_in(k_11_1316), .fluid_out(k_10_658), .air_in(c_11_0));
valve v_11_1317 (.fluid_in(k_11_1317), .fluid_out(k_10_658), .air_in(c_11_1));
valve v_11_1318 (.fluid_in(k_11_1318), .fluid_out(k_10_659), .air_in(c_11_0));
valve v_11_1319 (.fluid_in(k_11_1319), .fluid_out(k_10_659), .air_in(c_11_1));
valve v_11_1320 (.fluid_in(k_11_1320), .fluid_out(k_10_660), .air_in(c_11_0));
valve v_11_1321 (.fluid_in(k_11_1321), .fluid_out(k_10_660), .air_in(c_11_1));
valve v_11_1322 (.fluid_in(k_11_1322), .fluid_out(k_10_661), .air_in(c_11_0));
valve v_11_1323 (.fluid_in(k_11_1323), .fluid_out(k_10_661), .air_in(c_11_1));
valve v_11_1324 (.fluid_in(k_11_1324), .fluid_out(k_10_662), .air_in(c_11_0));
valve v_11_1325 (.fluid_in(k_11_1325), .fluid_out(k_10_662), .air_in(c_11_1));
valve v_11_1326 (.fluid_in(k_11_1326), .fluid_out(k_10_663), .air_in(c_11_0));
valve v_11_1327 (.fluid_in(k_11_1327), .fluid_out(k_10_663), .air_in(c_11_1));
valve v_11_1328 (.fluid_in(k_11_1328), .fluid_out(k_10_664), .air_in(c_11_0));
valve v_11_1329 (.fluid_in(k_11_1329), .fluid_out(k_10_664), .air_in(c_11_1));
valve v_11_1330 (.fluid_in(k_11_1330), .fluid_out(k_10_665), .air_in(c_11_0));
valve v_11_1331 (.fluid_in(k_11_1331), .fluid_out(k_10_665), .air_in(c_11_1));
valve v_11_1332 (.fluid_in(k_11_1332), .fluid_out(k_10_666), .air_in(c_11_0));
valve v_11_1333 (.fluid_in(k_11_1333), .fluid_out(k_10_666), .air_in(c_11_1));
valve v_11_1334 (.fluid_in(k_11_1334), .fluid_out(k_10_667), .air_in(c_11_0));
valve v_11_1335 (.fluid_in(k_11_1335), .fluid_out(k_10_667), .air_in(c_11_1));
valve v_11_1336 (.fluid_in(k_11_1336), .fluid_out(k_10_668), .air_in(c_11_0));
valve v_11_1337 (.fluid_in(k_11_1337), .fluid_out(k_10_668), .air_in(c_11_1));
valve v_11_1338 (.fluid_in(k_11_1338), .fluid_out(k_10_669), .air_in(c_11_0));
valve v_11_1339 (.fluid_in(k_11_1339), .fluid_out(k_10_669), .air_in(c_11_1));
valve v_11_1340 (.fluid_in(k_11_1340), .fluid_out(k_10_670), .air_in(c_11_0));
valve v_11_1341 (.fluid_in(k_11_1341), .fluid_out(k_10_670), .air_in(c_11_1));
valve v_11_1342 (.fluid_in(k_11_1342), .fluid_out(k_10_671), .air_in(c_11_0));
valve v_11_1343 (.fluid_in(k_11_1343), .fluid_out(k_10_671), .air_in(c_11_1));
valve v_11_1344 (.fluid_in(k_11_1344), .fluid_out(k_10_672), .air_in(c_11_0));
valve v_11_1345 (.fluid_in(k_11_1345), .fluid_out(k_10_672), .air_in(c_11_1));
valve v_11_1346 (.fluid_in(k_11_1346), .fluid_out(k_10_673), .air_in(c_11_0));
valve v_11_1347 (.fluid_in(k_11_1347), .fluid_out(k_10_673), .air_in(c_11_1));
valve v_11_1348 (.fluid_in(k_11_1348), .fluid_out(k_10_674), .air_in(c_11_0));
valve v_11_1349 (.fluid_in(k_11_1349), .fluid_out(k_10_674), .air_in(c_11_1));
valve v_11_1350 (.fluid_in(k_11_1350), .fluid_out(k_10_675), .air_in(c_11_0));
valve v_11_1351 (.fluid_in(k_11_1351), .fluid_out(k_10_675), .air_in(c_11_1));
valve v_11_1352 (.fluid_in(k_11_1352), .fluid_out(k_10_676), .air_in(c_11_0));
valve v_11_1353 (.fluid_in(k_11_1353), .fluid_out(k_10_676), .air_in(c_11_1));
valve v_11_1354 (.fluid_in(k_11_1354), .fluid_out(k_10_677), .air_in(c_11_0));
valve v_11_1355 (.fluid_in(k_11_1355), .fluid_out(k_10_677), .air_in(c_11_1));
valve v_11_1356 (.fluid_in(k_11_1356), .fluid_out(k_10_678), .air_in(c_11_0));
valve v_11_1357 (.fluid_in(k_11_1357), .fluid_out(k_10_678), .air_in(c_11_1));
valve v_11_1358 (.fluid_in(k_11_1358), .fluid_out(k_10_679), .air_in(c_11_0));
valve v_11_1359 (.fluid_in(k_11_1359), .fluid_out(k_10_679), .air_in(c_11_1));
valve v_11_1360 (.fluid_in(k_11_1360), .fluid_out(k_10_680), .air_in(c_11_0));
valve v_11_1361 (.fluid_in(k_11_1361), .fluid_out(k_10_680), .air_in(c_11_1));
valve v_11_1362 (.fluid_in(k_11_1362), .fluid_out(k_10_681), .air_in(c_11_0));
valve v_11_1363 (.fluid_in(k_11_1363), .fluid_out(k_10_681), .air_in(c_11_1));
valve v_11_1364 (.fluid_in(k_11_1364), .fluid_out(k_10_682), .air_in(c_11_0));
valve v_11_1365 (.fluid_in(k_11_1365), .fluid_out(k_10_682), .air_in(c_11_1));
valve v_11_1366 (.fluid_in(k_11_1366), .fluid_out(k_10_683), .air_in(c_11_0));
valve v_11_1367 (.fluid_in(k_11_1367), .fluid_out(k_10_683), .air_in(c_11_1));
valve v_11_1368 (.fluid_in(k_11_1368), .fluid_out(k_10_684), .air_in(c_11_0));
valve v_11_1369 (.fluid_in(k_11_1369), .fluid_out(k_10_684), .air_in(c_11_1));
valve v_11_1370 (.fluid_in(k_11_1370), .fluid_out(k_10_685), .air_in(c_11_0));
valve v_11_1371 (.fluid_in(k_11_1371), .fluid_out(k_10_685), .air_in(c_11_1));
valve v_11_1372 (.fluid_in(k_11_1372), .fluid_out(k_10_686), .air_in(c_11_0));
valve v_11_1373 (.fluid_in(k_11_1373), .fluid_out(k_10_686), .air_in(c_11_1));
valve v_11_1374 (.fluid_in(k_11_1374), .fluid_out(k_10_687), .air_in(c_11_0));
valve v_11_1375 (.fluid_in(k_11_1375), .fluid_out(k_10_687), .air_in(c_11_1));
valve v_11_1376 (.fluid_in(k_11_1376), .fluid_out(k_10_688), .air_in(c_11_0));
valve v_11_1377 (.fluid_in(k_11_1377), .fluid_out(k_10_688), .air_in(c_11_1));
valve v_11_1378 (.fluid_in(k_11_1378), .fluid_out(k_10_689), .air_in(c_11_0));
valve v_11_1379 (.fluid_in(k_11_1379), .fluid_out(k_10_689), .air_in(c_11_1));
valve v_11_1380 (.fluid_in(k_11_1380), .fluid_out(k_10_690), .air_in(c_11_0));
valve v_11_1381 (.fluid_in(k_11_1381), .fluid_out(k_10_690), .air_in(c_11_1));
valve v_11_1382 (.fluid_in(k_11_1382), .fluid_out(k_10_691), .air_in(c_11_0));
valve v_11_1383 (.fluid_in(k_11_1383), .fluid_out(k_10_691), .air_in(c_11_1));
valve v_11_1384 (.fluid_in(k_11_1384), .fluid_out(k_10_692), .air_in(c_11_0));
valve v_11_1385 (.fluid_in(k_11_1385), .fluid_out(k_10_692), .air_in(c_11_1));
valve v_11_1386 (.fluid_in(k_11_1386), .fluid_out(k_10_693), .air_in(c_11_0));
valve v_11_1387 (.fluid_in(k_11_1387), .fluid_out(k_10_693), .air_in(c_11_1));
valve v_11_1388 (.fluid_in(k_11_1388), .fluid_out(k_10_694), .air_in(c_11_0));
valve v_11_1389 (.fluid_in(k_11_1389), .fluid_out(k_10_694), .air_in(c_11_1));
valve v_11_1390 (.fluid_in(k_11_1390), .fluid_out(k_10_695), .air_in(c_11_0));
valve v_11_1391 (.fluid_in(k_11_1391), .fluid_out(k_10_695), .air_in(c_11_1));
valve v_11_1392 (.fluid_in(k_11_1392), .fluid_out(k_10_696), .air_in(c_11_0));
valve v_11_1393 (.fluid_in(k_11_1393), .fluid_out(k_10_696), .air_in(c_11_1));
valve v_11_1394 (.fluid_in(k_11_1394), .fluid_out(k_10_697), .air_in(c_11_0));
valve v_11_1395 (.fluid_in(k_11_1395), .fluid_out(k_10_697), .air_in(c_11_1));
valve v_11_1396 (.fluid_in(k_11_1396), .fluid_out(k_10_698), .air_in(c_11_0));
valve v_11_1397 (.fluid_in(k_11_1397), .fluid_out(k_10_698), .air_in(c_11_1));
valve v_11_1398 (.fluid_in(k_11_1398), .fluid_out(k_10_699), .air_in(c_11_0));
valve v_11_1399 (.fluid_in(k_11_1399), .fluid_out(k_10_699), .air_in(c_11_1));
valve v_11_1400 (.fluid_in(k_11_1400), .fluid_out(k_10_700), .air_in(c_11_0));
valve v_11_1401 (.fluid_in(k_11_1401), .fluid_out(k_10_700), .air_in(c_11_1));
valve v_11_1402 (.fluid_in(k_11_1402), .fluid_out(k_10_701), .air_in(c_11_0));
valve v_11_1403 (.fluid_in(k_11_1403), .fluid_out(k_10_701), .air_in(c_11_1));
valve v_11_1404 (.fluid_in(k_11_1404), .fluid_out(k_10_702), .air_in(c_11_0));
valve v_11_1405 (.fluid_in(k_11_1405), .fluid_out(k_10_702), .air_in(c_11_1));
valve v_11_1406 (.fluid_in(k_11_1406), .fluid_out(k_10_703), .air_in(c_11_0));
valve v_11_1407 (.fluid_in(k_11_1407), .fluid_out(k_10_703), .air_in(c_11_1));
valve v_11_1408 (.fluid_in(k_11_1408), .fluid_out(k_10_704), .air_in(c_11_0));
valve v_11_1409 (.fluid_in(k_11_1409), .fluid_out(k_10_704), .air_in(c_11_1));
valve v_11_1410 (.fluid_in(k_11_1410), .fluid_out(k_10_705), .air_in(c_11_0));
valve v_11_1411 (.fluid_in(k_11_1411), .fluid_out(k_10_705), .air_in(c_11_1));
valve v_11_1412 (.fluid_in(k_11_1412), .fluid_out(k_10_706), .air_in(c_11_0));
valve v_11_1413 (.fluid_in(k_11_1413), .fluid_out(k_10_706), .air_in(c_11_1));
valve v_11_1414 (.fluid_in(k_11_1414), .fluid_out(k_10_707), .air_in(c_11_0));
valve v_11_1415 (.fluid_in(k_11_1415), .fluid_out(k_10_707), .air_in(c_11_1));
valve v_11_1416 (.fluid_in(k_11_1416), .fluid_out(k_10_708), .air_in(c_11_0));
valve v_11_1417 (.fluid_in(k_11_1417), .fluid_out(k_10_708), .air_in(c_11_1));
valve v_11_1418 (.fluid_in(k_11_1418), .fluid_out(k_10_709), .air_in(c_11_0));
valve v_11_1419 (.fluid_in(k_11_1419), .fluid_out(k_10_709), .air_in(c_11_1));
valve v_11_1420 (.fluid_in(k_11_1420), .fluid_out(k_10_710), .air_in(c_11_0));
valve v_11_1421 (.fluid_in(k_11_1421), .fluid_out(k_10_710), .air_in(c_11_1));
valve v_11_1422 (.fluid_in(k_11_1422), .fluid_out(k_10_711), .air_in(c_11_0));
valve v_11_1423 (.fluid_in(k_11_1423), .fluid_out(k_10_711), .air_in(c_11_1));
valve v_11_1424 (.fluid_in(k_11_1424), .fluid_out(k_10_712), .air_in(c_11_0));
valve v_11_1425 (.fluid_in(k_11_1425), .fluid_out(k_10_712), .air_in(c_11_1));
valve v_11_1426 (.fluid_in(k_11_1426), .fluid_out(k_10_713), .air_in(c_11_0));
valve v_11_1427 (.fluid_in(k_11_1427), .fluid_out(k_10_713), .air_in(c_11_1));
valve v_11_1428 (.fluid_in(k_11_1428), .fluid_out(k_10_714), .air_in(c_11_0));
valve v_11_1429 (.fluid_in(k_11_1429), .fluid_out(k_10_714), .air_in(c_11_1));
valve v_11_1430 (.fluid_in(k_11_1430), .fluid_out(k_10_715), .air_in(c_11_0));
valve v_11_1431 (.fluid_in(k_11_1431), .fluid_out(k_10_715), .air_in(c_11_1));
valve v_11_1432 (.fluid_in(k_11_1432), .fluid_out(k_10_716), .air_in(c_11_0));
valve v_11_1433 (.fluid_in(k_11_1433), .fluid_out(k_10_716), .air_in(c_11_1));
valve v_11_1434 (.fluid_in(k_11_1434), .fluid_out(k_10_717), .air_in(c_11_0));
valve v_11_1435 (.fluid_in(k_11_1435), .fluid_out(k_10_717), .air_in(c_11_1));
valve v_11_1436 (.fluid_in(k_11_1436), .fluid_out(k_10_718), .air_in(c_11_0));
valve v_11_1437 (.fluid_in(k_11_1437), .fluid_out(k_10_718), .air_in(c_11_1));
valve v_11_1438 (.fluid_in(k_11_1438), .fluid_out(k_10_719), .air_in(c_11_0));
valve v_11_1439 (.fluid_in(k_11_1439), .fluid_out(k_10_719), .air_in(c_11_1));
valve v_11_1440 (.fluid_in(k_11_1440), .fluid_out(k_10_720), .air_in(c_11_0));
valve v_11_1441 (.fluid_in(k_11_1441), .fluid_out(k_10_720), .air_in(c_11_1));
valve v_11_1442 (.fluid_in(k_11_1442), .fluid_out(k_10_721), .air_in(c_11_0));
valve v_11_1443 (.fluid_in(k_11_1443), .fluid_out(k_10_721), .air_in(c_11_1));
valve v_11_1444 (.fluid_in(k_11_1444), .fluid_out(k_10_722), .air_in(c_11_0));
valve v_11_1445 (.fluid_in(k_11_1445), .fluid_out(k_10_722), .air_in(c_11_1));
valve v_11_1446 (.fluid_in(k_11_1446), .fluid_out(k_10_723), .air_in(c_11_0));
valve v_11_1447 (.fluid_in(k_11_1447), .fluid_out(k_10_723), .air_in(c_11_1));
valve v_11_1448 (.fluid_in(k_11_1448), .fluid_out(k_10_724), .air_in(c_11_0));
valve v_11_1449 (.fluid_in(k_11_1449), .fluid_out(k_10_724), .air_in(c_11_1));
valve v_11_1450 (.fluid_in(k_11_1450), .fluid_out(k_10_725), .air_in(c_11_0));
valve v_11_1451 (.fluid_in(k_11_1451), .fluid_out(k_10_725), .air_in(c_11_1));
valve v_11_1452 (.fluid_in(k_11_1452), .fluid_out(k_10_726), .air_in(c_11_0));
valve v_11_1453 (.fluid_in(k_11_1453), .fluid_out(k_10_726), .air_in(c_11_1));
valve v_11_1454 (.fluid_in(k_11_1454), .fluid_out(k_10_727), .air_in(c_11_0));
valve v_11_1455 (.fluid_in(k_11_1455), .fluid_out(k_10_727), .air_in(c_11_1));
valve v_11_1456 (.fluid_in(k_11_1456), .fluid_out(k_10_728), .air_in(c_11_0));
valve v_11_1457 (.fluid_in(k_11_1457), .fluid_out(k_10_728), .air_in(c_11_1));
valve v_11_1458 (.fluid_in(k_11_1458), .fluid_out(k_10_729), .air_in(c_11_0));
valve v_11_1459 (.fluid_in(k_11_1459), .fluid_out(k_10_729), .air_in(c_11_1));
valve v_11_1460 (.fluid_in(k_11_1460), .fluid_out(k_10_730), .air_in(c_11_0));
valve v_11_1461 (.fluid_in(k_11_1461), .fluid_out(k_10_730), .air_in(c_11_1));
valve v_11_1462 (.fluid_in(k_11_1462), .fluid_out(k_10_731), .air_in(c_11_0));
valve v_11_1463 (.fluid_in(k_11_1463), .fluid_out(k_10_731), .air_in(c_11_1));
valve v_11_1464 (.fluid_in(k_11_1464), .fluid_out(k_10_732), .air_in(c_11_0));
valve v_11_1465 (.fluid_in(k_11_1465), .fluid_out(k_10_732), .air_in(c_11_1));
valve v_11_1466 (.fluid_in(k_11_1466), .fluid_out(k_10_733), .air_in(c_11_0));
valve v_11_1467 (.fluid_in(k_11_1467), .fluid_out(k_10_733), .air_in(c_11_1));
valve v_11_1468 (.fluid_in(k_11_1468), .fluid_out(k_10_734), .air_in(c_11_0));
valve v_11_1469 (.fluid_in(k_11_1469), .fluid_out(k_10_734), .air_in(c_11_1));
valve v_11_1470 (.fluid_in(k_11_1470), .fluid_out(k_10_735), .air_in(c_11_0));
valve v_11_1471 (.fluid_in(k_11_1471), .fluid_out(k_10_735), .air_in(c_11_1));
valve v_11_1472 (.fluid_in(k_11_1472), .fluid_out(k_10_736), .air_in(c_11_0));
valve v_11_1473 (.fluid_in(k_11_1473), .fluid_out(k_10_736), .air_in(c_11_1));
valve v_11_1474 (.fluid_in(k_11_1474), .fluid_out(k_10_737), .air_in(c_11_0));
valve v_11_1475 (.fluid_in(k_11_1475), .fluid_out(k_10_737), .air_in(c_11_1));
valve v_11_1476 (.fluid_in(k_11_1476), .fluid_out(k_10_738), .air_in(c_11_0));
valve v_11_1477 (.fluid_in(k_11_1477), .fluid_out(k_10_738), .air_in(c_11_1));
valve v_11_1478 (.fluid_in(k_11_1478), .fluid_out(k_10_739), .air_in(c_11_0));
valve v_11_1479 (.fluid_in(k_11_1479), .fluid_out(k_10_739), .air_in(c_11_1));
valve v_11_1480 (.fluid_in(k_11_1480), .fluid_out(k_10_740), .air_in(c_11_0));
valve v_11_1481 (.fluid_in(k_11_1481), .fluid_out(k_10_740), .air_in(c_11_1));
valve v_11_1482 (.fluid_in(k_11_1482), .fluid_out(k_10_741), .air_in(c_11_0));
valve v_11_1483 (.fluid_in(k_11_1483), .fluid_out(k_10_741), .air_in(c_11_1));
valve v_11_1484 (.fluid_in(k_11_1484), .fluid_out(k_10_742), .air_in(c_11_0));
valve v_11_1485 (.fluid_in(k_11_1485), .fluid_out(k_10_742), .air_in(c_11_1));
valve v_11_1486 (.fluid_in(k_11_1486), .fluid_out(k_10_743), .air_in(c_11_0));
valve v_11_1487 (.fluid_in(k_11_1487), .fluid_out(k_10_743), .air_in(c_11_1));
valve v_11_1488 (.fluid_in(k_11_1488), .fluid_out(k_10_744), .air_in(c_11_0));
valve v_11_1489 (.fluid_in(k_11_1489), .fluid_out(k_10_744), .air_in(c_11_1));
valve v_11_1490 (.fluid_in(k_11_1490), .fluid_out(k_10_745), .air_in(c_11_0));
valve v_11_1491 (.fluid_in(k_11_1491), .fluid_out(k_10_745), .air_in(c_11_1));
valve v_11_1492 (.fluid_in(k_11_1492), .fluid_out(k_10_746), .air_in(c_11_0));
valve v_11_1493 (.fluid_in(k_11_1493), .fluid_out(k_10_746), .air_in(c_11_1));
valve v_11_1494 (.fluid_in(k_11_1494), .fluid_out(k_10_747), .air_in(c_11_0));
valve v_11_1495 (.fluid_in(k_11_1495), .fluid_out(k_10_747), .air_in(c_11_1));
valve v_11_1496 (.fluid_in(k_11_1496), .fluid_out(k_10_748), .air_in(c_11_0));
valve v_11_1497 (.fluid_in(k_11_1497), .fluid_out(k_10_748), .air_in(c_11_1));
valve v_11_1498 (.fluid_in(k_11_1498), .fluid_out(k_10_749), .air_in(c_11_0));
valve v_11_1499 (.fluid_in(k_11_1499), .fluid_out(k_10_749), .air_in(c_11_1));
valve v_11_1500 (.fluid_in(k_11_1500), .fluid_out(k_10_750), .air_in(c_11_0));
valve v_11_1501 (.fluid_in(k_11_1501), .fluid_out(k_10_750), .air_in(c_11_1));
valve v_11_1502 (.fluid_in(k_11_1502), .fluid_out(k_10_751), .air_in(c_11_0));
valve v_11_1503 (.fluid_in(k_11_1503), .fluid_out(k_10_751), .air_in(c_11_1));
valve v_11_1504 (.fluid_in(k_11_1504), .fluid_out(k_10_752), .air_in(c_11_0));
valve v_11_1505 (.fluid_in(k_11_1505), .fluid_out(k_10_752), .air_in(c_11_1));
valve v_11_1506 (.fluid_in(k_11_1506), .fluid_out(k_10_753), .air_in(c_11_0));
valve v_11_1507 (.fluid_in(k_11_1507), .fluid_out(k_10_753), .air_in(c_11_1));
valve v_11_1508 (.fluid_in(k_11_1508), .fluid_out(k_10_754), .air_in(c_11_0));
valve v_11_1509 (.fluid_in(k_11_1509), .fluid_out(k_10_754), .air_in(c_11_1));
valve v_11_1510 (.fluid_in(k_11_1510), .fluid_out(k_10_755), .air_in(c_11_0));
valve v_11_1511 (.fluid_in(k_11_1511), .fluid_out(k_10_755), .air_in(c_11_1));
valve v_11_1512 (.fluid_in(k_11_1512), .fluid_out(k_10_756), .air_in(c_11_0));
valve v_11_1513 (.fluid_in(k_11_1513), .fluid_out(k_10_756), .air_in(c_11_1));
valve v_11_1514 (.fluid_in(k_11_1514), .fluid_out(k_10_757), .air_in(c_11_0));
valve v_11_1515 (.fluid_in(k_11_1515), .fluid_out(k_10_757), .air_in(c_11_1));
valve v_11_1516 (.fluid_in(k_11_1516), .fluid_out(k_10_758), .air_in(c_11_0));
valve v_11_1517 (.fluid_in(k_11_1517), .fluid_out(k_10_758), .air_in(c_11_1));
valve v_11_1518 (.fluid_in(k_11_1518), .fluid_out(k_10_759), .air_in(c_11_0));
valve v_11_1519 (.fluid_in(k_11_1519), .fluid_out(k_10_759), .air_in(c_11_1));
valve v_11_1520 (.fluid_in(k_11_1520), .fluid_out(k_10_760), .air_in(c_11_0));
valve v_11_1521 (.fluid_in(k_11_1521), .fluid_out(k_10_760), .air_in(c_11_1));
valve v_11_1522 (.fluid_in(k_11_1522), .fluid_out(k_10_761), .air_in(c_11_0));
valve v_11_1523 (.fluid_in(k_11_1523), .fluid_out(k_10_761), .air_in(c_11_1));
valve v_11_1524 (.fluid_in(k_11_1524), .fluid_out(k_10_762), .air_in(c_11_0));
valve v_11_1525 (.fluid_in(k_11_1525), .fluid_out(k_10_762), .air_in(c_11_1));
valve v_11_1526 (.fluid_in(k_11_1526), .fluid_out(k_10_763), .air_in(c_11_0));
valve v_11_1527 (.fluid_in(k_11_1527), .fluid_out(k_10_763), .air_in(c_11_1));
valve v_11_1528 (.fluid_in(k_11_1528), .fluid_out(k_10_764), .air_in(c_11_0));
valve v_11_1529 (.fluid_in(k_11_1529), .fluid_out(k_10_764), .air_in(c_11_1));
valve v_11_1530 (.fluid_in(k_11_1530), .fluid_out(k_10_765), .air_in(c_11_0));
valve v_11_1531 (.fluid_in(k_11_1531), .fluid_out(k_10_765), .air_in(c_11_1));
valve v_11_1532 (.fluid_in(k_11_1532), .fluid_out(k_10_766), .air_in(c_11_0));
valve v_11_1533 (.fluid_in(k_11_1533), .fluid_out(k_10_766), .air_in(c_11_1));
valve v_11_1534 (.fluid_in(k_11_1534), .fluid_out(k_10_767), .air_in(c_11_0));
valve v_11_1535 (.fluid_in(k_11_1535), .fluid_out(k_10_767), .air_in(c_11_1));
valve v_11_1536 (.fluid_in(k_11_1536), .fluid_out(k_10_768), .air_in(c_11_0));
valve v_11_1537 (.fluid_in(k_11_1537), .fluid_out(k_10_768), .air_in(c_11_1));
valve v_11_1538 (.fluid_in(k_11_1538), .fluid_out(k_10_769), .air_in(c_11_0));
valve v_11_1539 (.fluid_in(k_11_1539), .fluid_out(k_10_769), .air_in(c_11_1));
valve v_11_1540 (.fluid_in(k_11_1540), .fluid_out(k_10_770), .air_in(c_11_0));
valve v_11_1541 (.fluid_in(k_11_1541), .fluid_out(k_10_770), .air_in(c_11_1));
valve v_11_1542 (.fluid_in(k_11_1542), .fluid_out(k_10_771), .air_in(c_11_0));
valve v_11_1543 (.fluid_in(k_11_1543), .fluid_out(k_10_771), .air_in(c_11_1));
valve v_11_1544 (.fluid_in(k_11_1544), .fluid_out(k_10_772), .air_in(c_11_0));
valve v_11_1545 (.fluid_in(k_11_1545), .fluid_out(k_10_772), .air_in(c_11_1));
valve v_11_1546 (.fluid_in(k_11_1546), .fluid_out(k_10_773), .air_in(c_11_0));
valve v_11_1547 (.fluid_in(k_11_1547), .fluid_out(k_10_773), .air_in(c_11_1));
valve v_11_1548 (.fluid_in(k_11_1548), .fluid_out(k_10_774), .air_in(c_11_0));
valve v_11_1549 (.fluid_in(k_11_1549), .fluid_out(k_10_774), .air_in(c_11_1));
valve v_11_1550 (.fluid_in(k_11_1550), .fluid_out(k_10_775), .air_in(c_11_0));
valve v_11_1551 (.fluid_in(k_11_1551), .fluid_out(k_10_775), .air_in(c_11_1));
valve v_11_1552 (.fluid_in(k_11_1552), .fluid_out(k_10_776), .air_in(c_11_0));
valve v_11_1553 (.fluid_in(k_11_1553), .fluid_out(k_10_776), .air_in(c_11_1));
valve v_11_1554 (.fluid_in(k_11_1554), .fluid_out(k_10_777), .air_in(c_11_0));
valve v_11_1555 (.fluid_in(k_11_1555), .fluid_out(k_10_777), .air_in(c_11_1));
valve v_11_1556 (.fluid_in(k_11_1556), .fluid_out(k_10_778), .air_in(c_11_0));
valve v_11_1557 (.fluid_in(k_11_1557), .fluid_out(k_10_778), .air_in(c_11_1));
valve v_11_1558 (.fluid_in(k_11_1558), .fluid_out(k_10_779), .air_in(c_11_0));
valve v_11_1559 (.fluid_in(k_11_1559), .fluid_out(k_10_779), .air_in(c_11_1));
valve v_11_1560 (.fluid_in(k_11_1560), .fluid_out(k_10_780), .air_in(c_11_0));
valve v_11_1561 (.fluid_in(k_11_1561), .fluid_out(k_10_780), .air_in(c_11_1));
valve v_11_1562 (.fluid_in(k_11_1562), .fluid_out(k_10_781), .air_in(c_11_0));
valve v_11_1563 (.fluid_in(k_11_1563), .fluid_out(k_10_781), .air_in(c_11_1));
valve v_11_1564 (.fluid_in(k_11_1564), .fluid_out(k_10_782), .air_in(c_11_0));
valve v_11_1565 (.fluid_in(k_11_1565), .fluid_out(k_10_782), .air_in(c_11_1));
valve v_11_1566 (.fluid_in(k_11_1566), .fluid_out(k_10_783), .air_in(c_11_0));
valve v_11_1567 (.fluid_in(k_11_1567), .fluid_out(k_10_783), .air_in(c_11_1));
valve v_11_1568 (.fluid_in(k_11_1568), .fluid_out(k_10_784), .air_in(c_11_0));
valve v_11_1569 (.fluid_in(k_11_1569), .fluid_out(k_10_784), .air_in(c_11_1));
valve v_11_1570 (.fluid_in(k_11_1570), .fluid_out(k_10_785), .air_in(c_11_0));
valve v_11_1571 (.fluid_in(k_11_1571), .fluid_out(k_10_785), .air_in(c_11_1));
valve v_11_1572 (.fluid_in(k_11_1572), .fluid_out(k_10_786), .air_in(c_11_0));
valve v_11_1573 (.fluid_in(k_11_1573), .fluid_out(k_10_786), .air_in(c_11_1));
valve v_11_1574 (.fluid_in(k_11_1574), .fluid_out(k_10_787), .air_in(c_11_0));
valve v_11_1575 (.fluid_in(k_11_1575), .fluid_out(k_10_787), .air_in(c_11_1));
valve v_11_1576 (.fluid_in(k_11_1576), .fluid_out(k_10_788), .air_in(c_11_0));
valve v_11_1577 (.fluid_in(k_11_1577), .fluid_out(k_10_788), .air_in(c_11_1));
valve v_11_1578 (.fluid_in(k_11_1578), .fluid_out(k_10_789), .air_in(c_11_0));
valve v_11_1579 (.fluid_in(k_11_1579), .fluid_out(k_10_789), .air_in(c_11_1));
valve v_11_1580 (.fluid_in(k_11_1580), .fluid_out(k_10_790), .air_in(c_11_0));
valve v_11_1581 (.fluid_in(k_11_1581), .fluid_out(k_10_790), .air_in(c_11_1));
valve v_11_1582 (.fluid_in(k_11_1582), .fluid_out(k_10_791), .air_in(c_11_0));
valve v_11_1583 (.fluid_in(k_11_1583), .fluid_out(k_10_791), .air_in(c_11_1));
valve v_11_1584 (.fluid_in(k_11_1584), .fluid_out(k_10_792), .air_in(c_11_0));
valve v_11_1585 (.fluid_in(k_11_1585), .fluid_out(k_10_792), .air_in(c_11_1));
valve v_11_1586 (.fluid_in(k_11_1586), .fluid_out(k_10_793), .air_in(c_11_0));
valve v_11_1587 (.fluid_in(k_11_1587), .fluid_out(k_10_793), .air_in(c_11_1));
valve v_11_1588 (.fluid_in(k_11_1588), .fluid_out(k_10_794), .air_in(c_11_0));
valve v_11_1589 (.fluid_in(k_11_1589), .fluid_out(k_10_794), .air_in(c_11_1));
valve v_11_1590 (.fluid_in(k_11_1590), .fluid_out(k_10_795), .air_in(c_11_0));
valve v_11_1591 (.fluid_in(k_11_1591), .fluid_out(k_10_795), .air_in(c_11_1));
valve v_11_1592 (.fluid_in(k_11_1592), .fluid_out(k_10_796), .air_in(c_11_0));
valve v_11_1593 (.fluid_in(k_11_1593), .fluid_out(k_10_796), .air_in(c_11_1));
valve v_11_1594 (.fluid_in(k_11_1594), .fluid_out(k_10_797), .air_in(c_11_0));
valve v_11_1595 (.fluid_in(k_11_1595), .fluid_out(k_10_797), .air_in(c_11_1));
valve v_11_1596 (.fluid_in(k_11_1596), .fluid_out(k_10_798), .air_in(c_11_0));
valve v_11_1597 (.fluid_in(k_11_1597), .fluid_out(k_10_798), .air_in(c_11_1));
valve v_11_1598 (.fluid_in(k_11_1598), .fluid_out(k_10_799), .air_in(c_11_0));
valve v_11_1599 (.fluid_in(k_11_1599), .fluid_out(k_10_799), .air_in(c_11_1));
valve v_11_1600 (.fluid_in(k_11_1600), .fluid_out(k_10_800), .air_in(c_11_0));
valve v_11_1601 (.fluid_in(k_11_1601), .fluid_out(k_10_800), .air_in(c_11_1));
valve v_11_1602 (.fluid_in(k_11_1602), .fluid_out(k_10_801), .air_in(c_11_0));
valve v_11_1603 (.fluid_in(k_11_1603), .fluid_out(k_10_801), .air_in(c_11_1));
valve v_11_1604 (.fluid_in(k_11_1604), .fluid_out(k_10_802), .air_in(c_11_0));
valve v_11_1605 (.fluid_in(k_11_1605), .fluid_out(k_10_802), .air_in(c_11_1));
valve v_11_1606 (.fluid_in(k_11_1606), .fluid_out(k_10_803), .air_in(c_11_0));
valve v_11_1607 (.fluid_in(k_11_1607), .fluid_out(k_10_803), .air_in(c_11_1));
valve v_11_1608 (.fluid_in(k_11_1608), .fluid_out(k_10_804), .air_in(c_11_0));
valve v_11_1609 (.fluid_in(k_11_1609), .fluid_out(k_10_804), .air_in(c_11_1));
valve v_11_1610 (.fluid_in(k_11_1610), .fluid_out(k_10_805), .air_in(c_11_0));
valve v_11_1611 (.fluid_in(k_11_1611), .fluid_out(k_10_805), .air_in(c_11_1));
valve v_11_1612 (.fluid_in(k_11_1612), .fluid_out(k_10_806), .air_in(c_11_0));
valve v_11_1613 (.fluid_in(k_11_1613), .fluid_out(k_10_806), .air_in(c_11_1));
valve v_11_1614 (.fluid_in(k_11_1614), .fluid_out(k_10_807), .air_in(c_11_0));
valve v_11_1615 (.fluid_in(k_11_1615), .fluid_out(k_10_807), .air_in(c_11_1));
valve v_11_1616 (.fluid_in(k_11_1616), .fluid_out(k_10_808), .air_in(c_11_0));
valve v_11_1617 (.fluid_in(k_11_1617), .fluid_out(k_10_808), .air_in(c_11_1));
valve v_11_1618 (.fluid_in(k_11_1618), .fluid_out(k_10_809), .air_in(c_11_0));
valve v_11_1619 (.fluid_in(k_11_1619), .fluid_out(k_10_809), .air_in(c_11_1));
valve v_11_1620 (.fluid_in(k_11_1620), .fluid_out(k_10_810), .air_in(c_11_0));
valve v_11_1621 (.fluid_in(k_11_1621), .fluid_out(k_10_810), .air_in(c_11_1));
valve v_11_1622 (.fluid_in(k_11_1622), .fluid_out(k_10_811), .air_in(c_11_0));
valve v_11_1623 (.fluid_in(k_11_1623), .fluid_out(k_10_811), .air_in(c_11_1));
valve v_11_1624 (.fluid_in(k_11_1624), .fluid_out(k_10_812), .air_in(c_11_0));
valve v_11_1625 (.fluid_in(k_11_1625), .fluid_out(k_10_812), .air_in(c_11_1));
valve v_11_1626 (.fluid_in(k_11_1626), .fluid_out(k_10_813), .air_in(c_11_0));
valve v_11_1627 (.fluid_in(k_11_1627), .fluid_out(k_10_813), .air_in(c_11_1));
valve v_11_1628 (.fluid_in(k_11_1628), .fluid_out(k_10_814), .air_in(c_11_0));
valve v_11_1629 (.fluid_in(k_11_1629), .fluid_out(k_10_814), .air_in(c_11_1));
valve v_11_1630 (.fluid_in(k_11_1630), .fluid_out(k_10_815), .air_in(c_11_0));
valve v_11_1631 (.fluid_in(k_11_1631), .fluid_out(k_10_815), .air_in(c_11_1));
valve v_11_1632 (.fluid_in(k_11_1632), .fluid_out(k_10_816), .air_in(c_11_0));
valve v_11_1633 (.fluid_in(k_11_1633), .fluid_out(k_10_816), .air_in(c_11_1));
valve v_11_1634 (.fluid_in(k_11_1634), .fluid_out(k_10_817), .air_in(c_11_0));
valve v_11_1635 (.fluid_in(k_11_1635), .fluid_out(k_10_817), .air_in(c_11_1));
valve v_11_1636 (.fluid_in(k_11_1636), .fluid_out(k_10_818), .air_in(c_11_0));
valve v_11_1637 (.fluid_in(k_11_1637), .fluid_out(k_10_818), .air_in(c_11_1));
valve v_11_1638 (.fluid_in(k_11_1638), .fluid_out(k_10_819), .air_in(c_11_0));
valve v_11_1639 (.fluid_in(k_11_1639), .fluid_out(k_10_819), .air_in(c_11_1));
valve v_11_1640 (.fluid_in(k_11_1640), .fluid_out(k_10_820), .air_in(c_11_0));
valve v_11_1641 (.fluid_in(k_11_1641), .fluid_out(k_10_820), .air_in(c_11_1));
valve v_11_1642 (.fluid_in(k_11_1642), .fluid_out(k_10_821), .air_in(c_11_0));
valve v_11_1643 (.fluid_in(k_11_1643), .fluid_out(k_10_821), .air_in(c_11_1));
valve v_11_1644 (.fluid_in(k_11_1644), .fluid_out(k_10_822), .air_in(c_11_0));
valve v_11_1645 (.fluid_in(k_11_1645), .fluid_out(k_10_822), .air_in(c_11_1));
valve v_11_1646 (.fluid_in(k_11_1646), .fluid_out(k_10_823), .air_in(c_11_0));
valve v_11_1647 (.fluid_in(k_11_1647), .fluid_out(k_10_823), .air_in(c_11_1));
valve v_11_1648 (.fluid_in(k_11_1648), .fluid_out(k_10_824), .air_in(c_11_0));
valve v_11_1649 (.fluid_in(k_11_1649), .fluid_out(k_10_824), .air_in(c_11_1));
valve v_11_1650 (.fluid_in(k_11_1650), .fluid_out(k_10_825), .air_in(c_11_0));
valve v_11_1651 (.fluid_in(k_11_1651), .fluid_out(k_10_825), .air_in(c_11_1));
valve v_11_1652 (.fluid_in(k_11_1652), .fluid_out(k_10_826), .air_in(c_11_0));
valve v_11_1653 (.fluid_in(k_11_1653), .fluid_out(k_10_826), .air_in(c_11_1));
valve v_11_1654 (.fluid_in(k_11_1654), .fluid_out(k_10_827), .air_in(c_11_0));
valve v_11_1655 (.fluid_in(k_11_1655), .fluid_out(k_10_827), .air_in(c_11_1));
valve v_11_1656 (.fluid_in(k_11_1656), .fluid_out(k_10_828), .air_in(c_11_0));
valve v_11_1657 (.fluid_in(k_11_1657), .fluid_out(k_10_828), .air_in(c_11_1));
valve v_11_1658 (.fluid_in(k_11_1658), .fluid_out(k_10_829), .air_in(c_11_0));
valve v_11_1659 (.fluid_in(k_11_1659), .fluid_out(k_10_829), .air_in(c_11_1));
valve v_11_1660 (.fluid_in(k_11_1660), .fluid_out(k_10_830), .air_in(c_11_0));
valve v_11_1661 (.fluid_in(k_11_1661), .fluid_out(k_10_830), .air_in(c_11_1));
valve v_11_1662 (.fluid_in(k_11_1662), .fluid_out(k_10_831), .air_in(c_11_0));
valve v_11_1663 (.fluid_in(k_11_1663), .fluid_out(k_10_831), .air_in(c_11_1));
valve v_11_1664 (.fluid_in(k_11_1664), .fluid_out(k_10_832), .air_in(c_11_0));
valve v_11_1665 (.fluid_in(k_11_1665), .fluid_out(k_10_832), .air_in(c_11_1));
valve v_11_1666 (.fluid_in(k_11_1666), .fluid_out(k_10_833), .air_in(c_11_0));
valve v_11_1667 (.fluid_in(k_11_1667), .fluid_out(k_10_833), .air_in(c_11_1));
valve v_11_1668 (.fluid_in(k_11_1668), .fluid_out(k_10_834), .air_in(c_11_0));
valve v_11_1669 (.fluid_in(k_11_1669), .fluid_out(k_10_834), .air_in(c_11_1));
valve v_11_1670 (.fluid_in(k_11_1670), .fluid_out(k_10_835), .air_in(c_11_0));
valve v_11_1671 (.fluid_in(k_11_1671), .fluid_out(k_10_835), .air_in(c_11_1));
valve v_11_1672 (.fluid_in(k_11_1672), .fluid_out(k_10_836), .air_in(c_11_0));
valve v_11_1673 (.fluid_in(k_11_1673), .fluid_out(k_10_836), .air_in(c_11_1));
valve v_11_1674 (.fluid_in(k_11_1674), .fluid_out(k_10_837), .air_in(c_11_0));
valve v_11_1675 (.fluid_in(k_11_1675), .fluid_out(k_10_837), .air_in(c_11_1));
valve v_11_1676 (.fluid_in(k_11_1676), .fluid_out(k_10_838), .air_in(c_11_0));
valve v_11_1677 (.fluid_in(k_11_1677), .fluid_out(k_10_838), .air_in(c_11_1));
valve v_11_1678 (.fluid_in(k_11_1678), .fluid_out(k_10_839), .air_in(c_11_0));
valve v_11_1679 (.fluid_in(k_11_1679), .fluid_out(k_10_839), .air_in(c_11_1));
valve v_11_1680 (.fluid_in(k_11_1680), .fluid_out(k_10_840), .air_in(c_11_0));
valve v_11_1681 (.fluid_in(k_11_1681), .fluid_out(k_10_840), .air_in(c_11_1));
valve v_11_1682 (.fluid_in(k_11_1682), .fluid_out(k_10_841), .air_in(c_11_0));
valve v_11_1683 (.fluid_in(k_11_1683), .fluid_out(k_10_841), .air_in(c_11_1));
valve v_11_1684 (.fluid_in(k_11_1684), .fluid_out(k_10_842), .air_in(c_11_0));
valve v_11_1685 (.fluid_in(k_11_1685), .fluid_out(k_10_842), .air_in(c_11_1));
valve v_11_1686 (.fluid_in(k_11_1686), .fluid_out(k_10_843), .air_in(c_11_0));
valve v_11_1687 (.fluid_in(k_11_1687), .fluid_out(k_10_843), .air_in(c_11_1));
valve v_11_1688 (.fluid_in(k_11_1688), .fluid_out(k_10_844), .air_in(c_11_0));
valve v_11_1689 (.fluid_in(k_11_1689), .fluid_out(k_10_844), .air_in(c_11_1));
valve v_11_1690 (.fluid_in(k_11_1690), .fluid_out(k_10_845), .air_in(c_11_0));
valve v_11_1691 (.fluid_in(k_11_1691), .fluid_out(k_10_845), .air_in(c_11_1));
valve v_11_1692 (.fluid_in(k_11_1692), .fluid_out(k_10_846), .air_in(c_11_0));
valve v_11_1693 (.fluid_in(k_11_1693), .fluid_out(k_10_846), .air_in(c_11_1));
valve v_11_1694 (.fluid_in(k_11_1694), .fluid_out(k_10_847), .air_in(c_11_0));
valve v_11_1695 (.fluid_in(k_11_1695), .fluid_out(k_10_847), .air_in(c_11_1));
valve v_11_1696 (.fluid_in(k_11_1696), .fluid_out(k_10_848), .air_in(c_11_0));
valve v_11_1697 (.fluid_in(k_11_1697), .fluid_out(k_10_848), .air_in(c_11_1));
valve v_11_1698 (.fluid_in(k_11_1698), .fluid_out(k_10_849), .air_in(c_11_0));
valve v_11_1699 (.fluid_in(k_11_1699), .fluid_out(k_10_849), .air_in(c_11_1));
valve v_11_1700 (.fluid_in(k_11_1700), .fluid_out(k_10_850), .air_in(c_11_0));
valve v_11_1701 (.fluid_in(k_11_1701), .fluid_out(k_10_850), .air_in(c_11_1));
valve v_11_1702 (.fluid_in(k_11_1702), .fluid_out(k_10_851), .air_in(c_11_0));
valve v_11_1703 (.fluid_in(k_11_1703), .fluid_out(k_10_851), .air_in(c_11_1));
valve v_11_1704 (.fluid_in(k_11_1704), .fluid_out(k_10_852), .air_in(c_11_0));
valve v_11_1705 (.fluid_in(k_11_1705), .fluid_out(k_10_852), .air_in(c_11_1));
valve v_11_1706 (.fluid_in(k_11_1706), .fluid_out(k_10_853), .air_in(c_11_0));
valve v_11_1707 (.fluid_in(k_11_1707), .fluid_out(k_10_853), .air_in(c_11_1));
valve v_11_1708 (.fluid_in(k_11_1708), .fluid_out(k_10_854), .air_in(c_11_0));
valve v_11_1709 (.fluid_in(k_11_1709), .fluid_out(k_10_854), .air_in(c_11_1));
valve v_11_1710 (.fluid_in(k_11_1710), .fluid_out(k_10_855), .air_in(c_11_0));
valve v_11_1711 (.fluid_in(k_11_1711), .fluid_out(k_10_855), .air_in(c_11_1));
valve v_11_1712 (.fluid_in(k_11_1712), .fluid_out(k_10_856), .air_in(c_11_0));
valve v_11_1713 (.fluid_in(k_11_1713), .fluid_out(k_10_856), .air_in(c_11_1));
valve v_11_1714 (.fluid_in(k_11_1714), .fluid_out(k_10_857), .air_in(c_11_0));
valve v_11_1715 (.fluid_in(k_11_1715), .fluid_out(k_10_857), .air_in(c_11_1));
valve v_11_1716 (.fluid_in(k_11_1716), .fluid_out(k_10_858), .air_in(c_11_0));
valve v_11_1717 (.fluid_in(k_11_1717), .fluid_out(k_10_858), .air_in(c_11_1));
valve v_11_1718 (.fluid_in(k_11_1718), .fluid_out(k_10_859), .air_in(c_11_0));
valve v_11_1719 (.fluid_in(k_11_1719), .fluid_out(k_10_859), .air_in(c_11_1));
valve v_11_1720 (.fluid_in(k_11_1720), .fluid_out(k_10_860), .air_in(c_11_0));
valve v_11_1721 (.fluid_in(k_11_1721), .fluid_out(k_10_860), .air_in(c_11_1));
valve v_11_1722 (.fluid_in(k_11_1722), .fluid_out(k_10_861), .air_in(c_11_0));
valve v_11_1723 (.fluid_in(k_11_1723), .fluid_out(k_10_861), .air_in(c_11_1));
valve v_11_1724 (.fluid_in(k_11_1724), .fluid_out(k_10_862), .air_in(c_11_0));
valve v_11_1725 (.fluid_in(k_11_1725), .fluid_out(k_10_862), .air_in(c_11_1));
valve v_11_1726 (.fluid_in(k_11_1726), .fluid_out(k_10_863), .air_in(c_11_0));
valve v_11_1727 (.fluid_in(k_11_1727), .fluid_out(k_10_863), .air_in(c_11_1));
valve v_11_1728 (.fluid_in(k_11_1728), .fluid_out(k_10_864), .air_in(c_11_0));
valve v_11_1729 (.fluid_in(k_11_1729), .fluid_out(k_10_864), .air_in(c_11_1));
valve v_11_1730 (.fluid_in(k_11_1730), .fluid_out(k_10_865), .air_in(c_11_0));
valve v_11_1731 (.fluid_in(k_11_1731), .fluid_out(k_10_865), .air_in(c_11_1));
valve v_11_1732 (.fluid_in(k_11_1732), .fluid_out(k_10_866), .air_in(c_11_0));
valve v_11_1733 (.fluid_in(k_11_1733), .fluid_out(k_10_866), .air_in(c_11_1));
valve v_11_1734 (.fluid_in(k_11_1734), .fluid_out(k_10_867), .air_in(c_11_0));
valve v_11_1735 (.fluid_in(k_11_1735), .fluid_out(k_10_867), .air_in(c_11_1));
valve v_11_1736 (.fluid_in(k_11_1736), .fluid_out(k_10_868), .air_in(c_11_0));
valve v_11_1737 (.fluid_in(k_11_1737), .fluid_out(k_10_868), .air_in(c_11_1));
valve v_11_1738 (.fluid_in(k_11_1738), .fluid_out(k_10_869), .air_in(c_11_0));
valve v_11_1739 (.fluid_in(k_11_1739), .fluid_out(k_10_869), .air_in(c_11_1));
valve v_11_1740 (.fluid_in(k_11_1740), .fluid_out(k_10_870), .air_in(c_11_0));
valve v_11_1741 (.fluid_in(k_11_1741), .fluid_out(k_10_870), .air_in(c_11_1));
valve v_11_1742 (.fluid_in(k_11_1742), .fluid_out(k_10_871), .air_in(c_11_0));
valve v_11_1743 (.fluid_in(k_11_1743), .fluid_out(k_10_871), .air_in(c_11_1));
valve v_11_1744 (.fluid_in(k_11_1744), .fluid_out(k_10_872), .air_in(c_11_0));
valve v_11_1745 (.fluid_in(k_11_1745), .fluid_out(k_10_872), .air_in(c_11_1));
valve v_11_1746 (.fluid_in(k_11_1746), .fluid_out(k_10_873), .air_in(c_11_0));
valve v_11_1747 (.fluid_in(k_11_1747), .fluid_out(k_10_873), .air_in(c_11_1));
valve v_11_1748 (.fluid_in(k_11_1748), .fluid_out(k_10_874), .air_in(c_11_0));
valve v_11_1749 (.fluid_in(k_11_1749), .fluid_out(k_10_874), .air_in(c_11_1));
valve v_11_1750 (.fluid_in(k_11_1750), .fluid_out(k_10_875), .air_in(c_11_0));
valve v_11_1751 (.fluid_in(k_11_1751), .fluid_out(k_10_875), .air_in(c_11_1));
valve v_11_1752 (.fluid_in(k_11_1752), .fluid_out(k_10_876), .air_in(c_11_0));
valve v_11_1753 (.fluid_in(k_11_1753), .fluid_out(k_10_876), .air_in(c_11_1));
valve v_11_1754 (.fluid_in(k_11_1754), .fluid_out(k_10_877), .air_in(c_11_0));
valve v_11_1755 (.fluid_in(k_11_1755), .fluid_out(k_10_877), .air_in(c_11_1));
valve v_11_1756 (.fluid_in(k_11_1756), .fluid_out(k_10_878), .air_in(c_11_0));
valve v_11_1757 (.fluid_in(k_11_1757), .fluid_out(k_10_878), .air_in(c_11_1));
valve v_11_1758 (.fluid_in(k_11_1758), .fluid_out(k_10_879), .air_in(c_11_0));
valve v_11_1759 (.fluid_in(k_11_1759), .fluid_out(k_10_879), .air_in(c_11_1));
valve v_11_1760 (.fluid_in(k_11_1760), .fluid_out(k_10_880), .air_in(c_11_0));
valve v_11_1761 (.fluid_in(k_11_1761), .fluid_out(k_10_880), .air_in(c_11_1));
valve v_11_1762 (.fluid_in(k_11_1762), .fluid_out(k_10_881), .air_in(c_11_0));
valve v_11_1763 (.fluid_in(k_11_1763), .fluid_out(k_10_881), .air_in(c_11_1));
valve v_11_1764 (.fluid_in(k_11_1764), .fluid_out(k_10_882), .air_in(c_11_0));
valve v_11_1765 (.fluid_in(k_11_1765), .fluid_out(k_10_882), .air_in(c_11_1));
valve v_11_1766 (.fluid_in(k_11_1766), .fluid_out(k_10_883), .air_in(c_11_0));
valve v_11_1767 (.fluid_in(k_11_1767), .fluid_out(k_10_883), .air_in(c_11_1));
valve v_11_1768 (.fluid_in(k_11_1768), .fluid_out(k_10_884), .air_in(c_11_0));
valve v_11_1769 (.fluid_in(k_11_1769), .fluid_out(k_10_884), .air_in(c_11_1));
valve v_11_1770 (.fluid_in(k_11_1770), .fluid_out(k_10_885), .air_in(c_11_0));
valve v_11_1771 (.fluid_in(k_11_1771), .fluid_out(k_10_885), .air_in(c_11_1));
valve v_11_1772 (.fluid_in(k_11_1772), .fluid_out(k_10_886), .air_in(c_11_0));
valve v_11_1773 (.fluid_in(k_11_1773), .fluid_out(k_10_886), .air_in(c_11_1));
valve v_11_1774 (.fluid_in(k_11_1774), .fluid_out(k_10_887), .air_in(c_11_0));
valve v_11_1775 (.fluid_in(k_11_1775), .fluid_out(k_10_887), .air_in(c_11_1));
valve v_11_1776 (.fluid_in(k_11_1776), .fluid_out(k_10_888), .air_in(c_11_0));
valve v_11_1777 (.fluid_in(k_11_1777), .fluid_out(k_10_888), .air_in(c_11_1));
valve v_11_1778 (.fluid_in(k_11_1778), .fluid_out(k_10_889), .air_in(c_11_0));
valve v_11_1779 (.fluid_in(k_11_1779), .fluid_out(k_10_889), .air_in(c_11_1));
valve v_11_1780 (.fluid_in(k_11_1780), .fluid_out(k_10_890), .air_in(c_11_0));
valve v_11_1781 (.fluid_in(k_11_1781), .fluid_out(k_10_890), .air_in(c_11_1));
valve v_11_1782 (.fluid_in(k_11_1782), .fluid_out(k_10_891), .air_in(c_11_0));
valve v_11_1783 (.fluid_in(k_11_1783), .fluid_out(k_10_891), .air_in(c_11_1));
valve v_11_1784 (.fluid_in(k_11_1784), .fluid_out(k_10_892), .air_in(c_11_0));
valve v_11_1785 (.fluid_in(k_11_1785), .fluid_out(k_10_892), .air_in(c_11_1));
valve v_11_1786 (.fluid_in(k_11_1786), .fluid_out(k_10_893), .air_in(c_11_0));
valve v_11_1787 (.fluid_in(k_11_1787), .fluid_out(k_10_893), .air_in(c_11_1));
valve v_11_1788 (.fluid_in(k_11_1788), .fluid_out(k_10_894), .air_in(c_11_0));
valve v_11_1789 (.fluid_in(k_11_1789), .fluid_out(k_10_894), .air_in(c_11_1));
valve v_11_1790 (.fluid_in(k_11_1790), .fluid_out(k_10_895), .air_in(c_11_0));
valve v_11_1791 (.fluid_in(k_11_1791), .fluid_out(k_10_895), .air_in(c_11_1));
valve v_11_1792 (.fluid_in(k_11_1792), .fluid_out(k_10_896), .air_in(c_11_0));
valve v_11_1793 (.fluid_in(k_11_1793), .fluid_out(k_10_896), .air_in(c_11_1));
valve v_11_1794 (.fluid_in(k_11_1794), .fluid_out(k_10_897), .air_in(c_11_0));
valve v_11_1795 (.fluid_in(k_11_1795), .fluid_out(k_10_897), .air_in(c_11_1));
valve v_11_1796 (.fluid_in(k_11_1796), .fluid_out(k_10_898), .air_in(c_11_0));
valve v_11_1797 (.fluid_in(k_11_1797), .fluid_out(k_10_898), .air_in(c_11_1));
valve v_11_1798 (.fluid_in(k_11_1798), .fluid_out(k_10_899), .air_in(c_11_0));
valve v_11_1799 (.fluid_in(k_11_1799), .fluid_out(k_10_899), .air_in(c_11_1));
valve v_11_1800 (.fluid_in(k_11_1800), .fluid_out(k_10_900), .air_in(c_11_0));
valve v_11_1801 (.fluid_in(k_11_1801), .fluid_out(k_10_900), .air_in(c_11_1));
valve v_11_1802 (.fluid_in(k_11_1802), .fluid_out(k_10_901), .air_in(c_11_0));
valve v_11_1803 (.fluid_in(k_11_1803), .fluid_out(k_10_901), .air_in(c_11_1));
valve v_11_1804 (.fluid_in(k_11_1804), .fluid_out(k_10_902), .air_in(c_11_0));
valve v_11_1805 (.fluid_in(k_11_1805), .fluid_out(k_10_902), .air_in(c_11_1));
valve v_11_1806 (.fluid_in(k_11_1806), .fluid_out(k_10_903), .air_in(c_11_0));
valve v_11_1807 (.fluid_in(k_11_1807), .fluid_out(k_10_903), .air_in(c_11_1));
valve v_11_1808 (.fluid_in(k_11_1808), .fluid_out(k_10_904), .air_in(c_11_0));
valve v_11_1809 (.fluid_in(k_11_1809), .fluid_out(k_10_904), .air_in(c_11_1));
valve v_11_1810 (.fluid_in(k_11_1810), .fluid_out(k_10_905), .air_in(c_11_0));
valve v_11_1811 (.fluid_in(k_11_1811), .fluid_out(k_10_905), .air_in(c_11_1));
valve v_11_1812 (.fluid_in(k_11_1812), .fluid_out(k_10_906), .air_in(c_11_0));
valve v_11_1813 (.fluid_in(k_11_1813), .fluid_out(k_10_906), .air_in(c_11_1));
valve v_11_1814 (.fluid_in(k_11_1814), .fluid_out(k_10_907), .air_in(c_11_0));
valve v_11_1815 (.fluid_in(k_11_1815), .fluid_out(k_10_907), .air_in(c_11_1));
valve v_11_1816 (.fluid_in(k_11_1816), .fluid_out(k_10_908), .air_in(c_11_0));
valve v_11_1817 (.fluid_in(k_11_1817), .fluid_out(k_10_908), .air_in(c_11_1));
valve v_11_1818 (.fluid_in(k_11_1818), .fluid_out(k_10_909), .air_in(c_11_0));
valve v_11_1819 (.fluid_in(k_11_1819), .fluid_out(k_10_909), .air_in(c_11_1));
valve v_11_1820 (.fluid_in(k_11_1820), .fluid_out(k_10_910), .air_in(c_11_0));
valve v_11_1821 (.fluid_in(k_11_1821), .fluid_out(k_10_910), .air_in(c_11_1));
valve v_11_1822 (.fluid_in(k_11_1822), .fluid_out(k_10_911), .air_in(c_11_0));
valve v_11_1823 (.fluid_in(k_11_1823), .fluid_out(k_10_911), .air_in(c_11_1));
valve v_11_1824 (.fluid_in(k_11_1824), .fluid_out(k_10_912), .air_in(c_11_0));
valve v_11_1825 (.fluid_in(k_11_1825), .fluid_out(k_10_912), .air_in(c_11_1));
valve v_11_1826 (.fluid_in(k_11_1826), .fluid_out(k_10_913), .air_in(c_11_0));
valve v_11_1827 (.fluid_in(k_11_1827), .fluid_out(k_10_913), .air_in(c_11_1));
valve v_11_1828 (.fluid_in(k_11_1828), .fluid_out(k_10_914), .air_in(c_11_0));
valve v_11_1829 (.fluid_in(k_11_1829), .fluid_out(k_10_914), .air_in(c_11_1));
valve v_11_1830 (.fluid_in(k_11_1830), .fluid_out(k_10_915), .air_in(c_11_0));
valve v_11_1831 (.fluid_in(k_11_1831), .fluid_out(k_10_915), .air_in(c_11_1));
valve v_11_1832 (.fluid_in(k_11_1832), .fluid_out(k_10_916), .air_in(c_11_0));
valve v_11_1833 (.fluid_in(k_11_1833), .fluid_out(k_10_916), .air_in(c_11_1));
valve v_11_1834 (.fluid_in(k_11_1834), .fluid_out(k_10_917), .air_in(c_11_0));
valve v_11_1835 (.fluid_in(k_11_1835), .fluid_out(k_10_917), .air_in(c_11_1));
valve v_11_1836 (.fluid_in(k_11_1836), .fluid_out(k_10_918), .air_in(c_11_0));
valve v_11_1837 (.fluid_in(k_11_1837), .fluid_out(k_10_918), .air_in(c_11_1));
valve v_11_1838 (.fluid_in(k_11_1838), .fluid_out(k_10_919), .air_in(c_11_0));
valve v_11_1839 (.fluid_in(k_11_1839), .fluid_out(k_10_919), .air_in(c_11_1));
valve v_11_1840 (.fluid_in(k_11_1840), .fluid_out(k_10_920), .air_in(c_11_0));
valve v_11_1841 (.fluid_in(k_11_1841), .fluid_out(k_10_920), .air_in(c_11_1));
valve v_11_1842 (.fluid_in(k_11_1842), .fluid_out(k_10_921), .air_in(c_11_0));
valve v_11_1843 (.fluid_in(k_11_1843), .fluid_out(k_10_921), .air_in(c_11_1));
valve v_11_1844 (.fluid_in(k_11_1844), .fluid_out(k_10_922), .air_in(c_11_0));
valve v_11_1845 (.fluid_in(k_11_1845), .fluid_out(k_10_922), .air_in(c_11_1));
valve v_11_1846 (.fluid_in(k_11_1846), .fluid_out(k_10_923), .air_in(c_11_0));
valve v_11_1847 (.fluid_in(k_11_1847), .fluid_out(k_10_923), .air_in(c_11_1));
valve v_11_1848 (.fluid_in(k_11_1848), .fluid_out(k_10_924), .air_in(c_11_0));
valve v_11_1849 (.fluid_in(k_11_1849), .fluid_out(k_10_924), .air_in(c_11_1));
valve v_11_1850 (.fluid_in(k_11_1850), .fluid_out(k_10_925), .air_in(c_11_0));
valve v_11_1851 (.fluid_in(k_11_1851), .fluid_out(k_10_925), .air_in(c_11_1));
valve v_11_1852 (.fluid_in(k_11_1852), .fluid_out(k_10_926), .air_in(c_11_0));
valve v_11_1853 (.fluid_in(k_11_1853), .fluid_out(k_10_926), .air_in(c_11_1));
valve v_11_1854 (.fluid_in(k_11_1854), .fluid_out(k_10_927), .air_in(c_11_0));
valve v_11_1855 (.fluid_in(k_11_1855), .fluid_out(k_10_927), .air_in(c_11_1));
valve v_11_1856 (.fluid_in(k_11_1856), .fluid_out(k_10_928), .air_in(c_11_0));
valve v_11_1857 (.fluid_in(k_11_1857), .fluid_out(k_10_928), .air_in(c_11_1));
valve v_11_1858 (.fluid_in(k_11_1858), .fluid_out(k_10_929), .air_in(c_11_0));
valve v_11_1859 (.fluid_in(k_11_1859), .fluid_out(k_10_929), .air_in(c_11_1));
valve v_11_1860 (.fluid_in(k_11_1860), .fluid_out(k_10_930), .air_in(c_11_0));
valve v_11_1861 (.fluid_in(k_11_1861), .fluid_out(k_10_930), .air_in(c_11_1));
valve v_11_1862 (.fluid_in(k_11_1862), .fluid_out(k_10_931), .air_in(c_11_0));
valve v_11_1863 (.fluid_in(k_11_1863), .fluid_out(k_10_931), .air_in(c_11_1));
valve v_11_1864 (.fluid_in(k_11_1864), .fluid_out(k_10_932), .air_in(c_11_0));
valve v_11_1865 (.fluid_in(k_11_1865), .fluid_out(k_10_932), .air_in(c_11_1));
valve v_11_1866 (.fluid_in(k_11_1866), .fluid_out(k_10_933), .air_in(c_11_0));
valve v_11_1867 (.fluid_in(k_11_1867), .fluid_out(k_10_933), .air_in(c_11_1));
valve v_11_1868 (.fluid_in(k_11_1868), .fluid_out(k_10_934), .air_in(c_11_0));
valve v_11_1869 (.fluid_in(k_11_1869), .fluid_out(k_10_934), .air_in(c_11_1));
valve v_11_1870 (.fluid_in(k_11_1870), .fluid_out(k_10_935), .air_in(c_11_0));
valve v_11_1871 (.fluid_in(k_11_1871), .fluid_out(k_10_935), .air_in(c_11_1));
valve v_11_1872 (.fluid_in(k_11_1872), .fluid_out(k_10_936), .air_in(c_11_0));
valve v_11_1873 (.fluid_in(k_11_1873), .fluid_out(k_10_936), .air_in(c_11_1));
valve v_11_1874 (.fluid_in(k_11_1874), .fluid_out(k_10_937), .air_in(c_11_0));
valve v_11_1875 (.fluid_in(k_11_1875), .fluid_out(k_10_937), .air_in(c_11_1));
valve v_11_1876 (.fluid_in(k_11_1876), .fluid_out(k_10_938), .air_in(c_11_0));
valve v_11_1877 (.fluid_in(k_11_1877), .fluid_out(k_10_938), .air_in(c_11_1));
valve v_11_1878 (.fluid_in(k_11_1878), .fluid_out(k_10_939), .air_in(c_11_0));
valve v_11_1879 (.fluid_in(k_11_1879), .fluid_out(k_10_939), .air_in(c_11_1));
valve v_11_1880 (.fluid_in(k_11_1880), .fluid_out(k_10_940), .air_in(c_11_0));
valve v_11_1881 (.fluid_in(k_11_1881), .fluid_out(k_10_940), .air_in(c_11_1));
valve v_11_1882 (.fluid_in(k_11_1882), .fluid_out(k_10_941), .air_in(c_11_0));
valve v_11_1883 (.fluid_in(k_11_1883), .fluid_out(k_10_941), .air_in(c_11_1));
valve v_11_1884 (.fluid_in(k_11_1884), .fluid_out(k_10_942), .air_in(c_11_0));
valve v_11_1885 (.fluid_in(k_11_1885), .fluid_out(k_10_942), .air_in(c_11_1));
valve v_11_1886 (.fluid_in(k_11_1886), .fluid_out(k_10_943), .air_in(c_11_0));
valve v_11_1887 (.fluid_in(k_11_1887), .fluid_out(k_10_943), .air_in(c_11_1));
valve v_11_1888 (.fluid_in(k_11_1888), .fluid_out(k_10_944), .air_in(c_11_0));
valve v_11_1889 (.fluid_in(k_11_1889), .fluid_out(k_10_944), .air_in(c_11_1));
valve v_11_1890 (.fluid_in(k_11_1890), .fluid_out(k_10_945), .air_in(c_11_0));
valve v_11_1891 (.fluid_in(k_11_1891), .fluid_out(k_10_945), .air_in(c_11_1));
valve v_11_1892 (.fluid_in(k_11_1892), .fluid_out(k_10_946), .air_in(c_11_0));
valve v_11_1893 (.fluid_in(k_11_1893), .fluid_out(k_10_946), .air_in(c_11_1));
valve v_11_1894 (.fluid_in(k_11_1894), .fluid_out(k_10_947), .air_in(c_11_0));
valve v_11_1895 (.fluid_in(k_11_1895), .fluid_out(k_10_947), .air_in(c_11_1));
valve v_11_1896 (.fluid_in(k_11_1896), .fluid_out(k_10_948), .air_in(c_11_0));
valve v_11_1897 (.fluid_in(k_11_1897), .fluid_out(k_10_948), .air_in(c_11_1));
valve v_11_1898 (.fluid_in(k_11_1898), .fluid_out(k_10_949), .air_in(c_11_0));
valve v_11_1899 (.fluid_in(k_11_1899), .fluid_out(k_10_949), .air_in(c_11_1));
valve v_11_1900 (.fluid_in(k_11_1900), .fluid_out(k_10_950), .air_in(c_11_0));
valve v_11_1901 (.fluid_in(k_11_1901), .fluid_out(k_10_950), .air_in(c_11_1));
valve v_11_1902 (.fluid_in(k_11_1902), .fluid_out(k_10_951), .air_in(c_11_0));
valve v_11_1903 (.fluid_in(k_11_1903), .fluid_out(k_10_951), .air_in(c_11_1));
valve v_11_1904 (.fluid_in(k_11_1904), .fluid_out(k_10_952), .air_in(c_11_0));
valve v_11_1905 (.fluid_in(k_11_1905), .fluid_out(k_10_952), .air_in(c_11_1));
valve v_11_1906 (.fluid_in(k_11_1906), .fluid_out(k_10_953), .air_in(c_11_0));
valve v_11_1907 (.fluid_in(k_11_1907), .fluid_out(k_10_953), .air_in(c_11_1));
valve v_11_1908 (.fluid_in(k_11_1908), .fluid_out(k_10_954), .air_in(c_11_0));
valve v_11_1909 (.fluid_in(k_11_1909), .fluid_out(k_10_954), .air_in(c_11_1));
valve v_11_1910 (.fluid_in(k_11_1910), .fluid_out(k_10_955), .air_in(c_11_0));
valve v_11_1911 (.fluid_in(k_11_1911), .fluid_out(k_10_955), .air_in(c_11_1));
valve v_11_1912 (.fluid_in(k_11_1912), .fluid_out(k_10_956), .air_in(c_11_0));
valve v_11_1913 (.fluid_in(k_11_1913), .fluid_out(k_10_956), .air_in(c_11_1));
valve v_11_1914 (.fluid_in(k_11_1914), .fluid_out(k_10_957), .air_in(c_11_0));
valve v_11_1915 (.fluid_in(k_11_1915), .fluid_out(k_10_957), .air_in(c_11_1));
valve v_11_1916 (.fluid_in(k_11_1916), .fluid_out(k_10_958), .air_in(c_11_0));
valve v_11_1917 (.fluid_in(k_11_1917), .fluid_out(k_10_958), .air_in(c_11_1));
valve v_11_1918 (.fluid_in(k_11_1918), .fluid_out(k_10_959), .air_in(c_11_0));
valve v_11_1919 (.fluid_in(k_11_1919), .fluid_out(k_10_959), .air_in(c_11_1));
valve v_11_1920 (.fluid_in(k_11_1920), .fluid_out(k_10_960), .air_in(c_11_0));
valve v_11_1921 (.fluid_in(k_11_1921), .fluid_out(k_10_960), .air_in(c_11_1));
valve v_11_1922 (.fluid_in(k_11_1922), .fluid_out(k_10_961), .air_in(c_11_0));
valve v_11_1923 (.fluid_in(k_11_1923), .fluid_out(k_10_961), .air_in(c_11_1));
valve v_11_1924 (.fluid_in(k_11_1924), .fluid_out(k_10_962), .air_in(c_11_0));
valve v_11_1925 (.fluid_in(k_11_1925), .fluid_out(k_10_962), .air_in(c_11_1));
valve v_11_1926 (.fluid_in(k_11_1926), .fluid_out(k_10_963), .air_in(c_11_0));
valve v_11_1927 (.fluid_in(k_11_1927), .fluid_out(k_10_963), .air_in(c_11_1));
valve v_11_1928 (.fluid_in(k_11_1928), .fluid_out(k_10_964), .air_in(c_11_0));
valve v_11_1929 (.fluid_in(k_11_1929), .fluid_out(k_10_964), .air_in(c_11_1));
valve v_11_1930 (.fluid_in(k_11_1930), .fluid_out(k_10_965), .air_in(c_11_0));
valve v_11_1931 (.fluid_in(k_11_1931), .fluid_out(k_10_965), .air_in(c_11_1));
valve v_11_1932 (.fluid_in(k_11_1932), .fluid_out(k_10_966), .air_in(c_11_0));
valve v_11_1933 (.fluid_in(k_11_1933), .fluid_out(k_10_966), .air_in(c_11_1));
valve v_11_1934 (.fluid_in(k_11_1934), .fluid_out(k_10_967), .air_in(c_11_0));
valve v_11_1935 (.fluid_in(k_11_1935), .fluid_out(k_10_967), .air_in(c_11_1));
valve v_11_1936 (.fluid_in(k_11_1936), .fluid_out(k_10_968), .air_in(c_11_0));
valve v_11_1937 (.fluid_in(k_11_1937), .fluid_out(k_10_968), .air_in(c_11_1));
valve v_11_1938 (.fluid_in(k_11_1938), .fluid_out(k_10_969), .air_in(c_11_0));
valve v_11_1939 (.fluid_in(k_11_1939), .fluid_out(k_10_969), .air_in(c_11_1));
valve v_11_1940 (.fluid_in(k_11_1940), .fluid_out(k_10_970), .air_in(c_11_0));
valve v_11_1941 (.fluid_in(k_11_1941), .fluid_out(k_10_970), .air_in(c_11_1));
valve v_11_1942 (.fluid_in(k_11_1942), .fluid_out(k_10_971), .air_in(c_11_0));
valve v_11_1943 (.fluid_in(k_11_1943), .fluid_out(k_10_971), .air_in(c_11_1));
valve v_11_1944 (.fluid_in(k_11_1944), .fluid_out(k_10_972), .air_in(c_11_0));
valve v_11_1945 (.fluid_in(k_11_1945), .fluid_out(k_10_972), .air_in(c_11_1));
valve v_11_1946 (.fluid_in(k_11_1946), .fluid_out(k_10_973), .air_in(c_11_0));
valve v_11_1947 (.fluid_in(k_11_1947), .fluid_out(k_10_973), .air_in(c_11_1));
valve v_11_1948 (.fluid_in(k_11_1948), .fluid_out(k_10_974), .air_in(c_11_0));
valve v_11_1949 (.fluid_in(k_11_1949), .fluid_out(k_10_974), .air_in(c_11_1));
valve v_11_1950 (.fluid_in(k_11_1950), .fluid_out(k_10_975), .air_in(c_11_0));
valve v_11_1951 (.fluid_in(k_11_1951), .fluid_out(k_10_975), .air_in(c_11_1));
valve v_11_1952 (.fluid_in(k_11_1952), .fluid_out(k_10_976), .air_in(c_11_0));
valve v_11_1953 (.fluid_in(k_11_1953), .fluid_out(k_10_976), .air_in(c_11_1));
valve v_11_1954 (.fluid_in(k_11_1954), .fluid_out(k_10_977), .air_in(c_11_0));
valve v_11_1955 (.fluid_in(k_11_1955), .fluid_out(k_10_977), .air_in(c_11_1));
valve v_11_1956 (.fluid_in(k_11_1956), .fluid_out(k_10_978), .air_in(c_11_0));
valve v_11_1957 (.fluid_in(k_11_1957), .fluid_out(k_10_978), .air_in(c_11_1));
valve v_11_1958 (.fluid_in(k_11_1958), .fluid_out(k_10_979), .air_in(c_11_0));
valve v_11_1959 (.fluid_in(k_11_1959), .fluid_out(k_10_979), .air_in(c_11_1));
valve v_11_1960 (.fluid_in(k_11_1960), .fluid_out(k_10_980), .air_in(c_11_0));
valve v_11_1961 (.fluid_in(k_11_1961), .fluid_out(k_10_980), .air_in(c_11_1));
valve v_11_1962 (.fluid_in(k_11_1962), .fluid_out(k_10_981), .air_in(c_11_0));
valve v_11_1963 (.fluid_in(k_11_1963), .fluid_out(k_10_981), .air_in(c_11_1));
valve v_11_1964 (.fluid_in(k_11_1964), .fluid_out(k_10_982), .air_in(c_11_0));
valve v_11_1965 (.fluid_in(k_11_1965), .fluid_out(k_10_982), .air_in(c_11_1));
valve v_11_1966 (.fluid_in(k_11_1966), .fluid_out(k_10_983), .air_in(c_11_0));
valve v_11_1967 (.fluid_in(k_11_1967), .fluid_out(k_10_983), .air_in(c_11_1));
valve v_11_1968 (.fluid_in(k_11_1968), .fluid_out(k_10_984), .air_in(c_11_0));
valve v_11_1969 (.fluid_in(k_11_1969), .fluid_out(k_10_984), .air_in(c_11_1));
valve v_11_1970 (.fluid_in(k_11_1970), .fluid_out(k_10_985), .air_in(c_11_0));
valve v_11_1971 (.fluid_in(k_11_1971), .fluid_out(k_10_985), .air_in(c_11_1));
valve v_11_1972 (.fluid_in(k_11_1972), .fluid_out(k_10_986), .air_in(c_11_0));
valve v_11_1973 (.fluid_in(k_11_1973), .fluid_out(k_10_986), .air_in(c_11_1));
valve v_11_1974 (.fluid_in(k_11_1974), .fluid_out(k_10_987), .air_in(c_11_0));
valve v_11_1975 (.fluid_in(k_11_1975), .fluid_out(k_10_987), .air_in(c_11_1));
valve v_11_1976 (.fluid_in(k_11_1976), .fluid_out(k_10_988), .air_in(c_11_0));
valve v_11_1977 (.fluid_in(k_11_1977), .fluid_out(k_10_988), .air_in(c_11_1));
valve v_11_1978 (.fluid_in(k_11_1978), .fluid_out(k_10_989), .air_in(c_11_0));
valve v_11_1979 (.fluid_in(k_11_1979), .fluid_out(k_10_989), .air_in(c_11_1));
valve v_11_1980 (.fluid_in(k_11_1980), .fluid_out(k_10_990), .air_in(c_11_0));
valve v_11_1981 (.fluid_in(k_11_1981), .fluid_out(k_10_990), .air_in(c_11_1));
valve v_11_1982 (.fluid_in(k_11_1982), .fluid_out(k_10_991), .air_in(c_11_0));
valve v_11_1983 (.fluid_in(k_11_1983), .fluid_out(k_10_991), .air_in(c_11_1));
valve v_11_1984 (.fluid_in(k_11_1984), .fluid_out(k_10_992), .air_in(c_11_0));
valve v_11_1985 (.fluid_in(k_11_1985), .fluid_out(k_10_992), .air_in(c_11_1));
valve v_11_1986 (.fluid_in(k_11_1986), .fluid_out(k_10_993), .air_in(c_11_0));
valve v_11_1987 (.fluid_in(k_11_1987), .fluid_out(k_10_993), .air_in(c_11_1));
valve v_11_1988 (.fluid_in(k_11_1988), .fluid_out(k_10_994), .air_in(c_11_0));
valve v_11_1989 (.fluid_in(k_11_1989), .fluid_out(k_10_994), .air_in(c_11_1));
valve v_11_1990 (.fluid_in(k_11_1990), .fluid_out(k_10_995), .air_in(c_11_0));
valve v_11_1991 (.fluid_in(k_11_1991), .fluid_out(k_10_995), .air_in(c_11_1));
valve v_11_1992 (.fluid_in(k_11_1992), .fluid_out(k_10_996), .air_in(c_11_0));
valve v_11_1993 (.fluid_in(k_11_1993), .fluid_out(k_10_996), .air_in(c_11_1));
valve v_11_1994 (.fluid_in(k_11_1994), .fluid_out(k_10_997), .air_in(c_11_0));
valve v_11_1995 (.fluid_in(k_11_1995), .fluid_out(k_10_997), .air_in(c_11_1));
valve v_11_1996 (.fluid_in(k_11_1996), .fluid_out(k_10_998), .air_in(c_11_0));
valve v_11_1997 (.fluid_in(k_11_1997), .fluid_out(k_10_998), .air_in(c_11_1));
valve v_11_1998 (.fluid_in(k_11_1998), .fluid_out(k_10_999), .air_in(c_11_0));
valve v_11_1999 (.fluid_in(k_11_1999), .fluid_out(k_10_999), .air_in(c_11_1));
valve v_11_2000 (.fluid_in(k_11_2000), .fluid_out(k_10_1000), .air_in(c_11_0));
valve v_11_2001 (.fluid_in(k_11_2001), .fluid_out(k_10_1000), .air_in(c_11_1));
valve v_11_2002 (.fluid_in(k_11_2002), .fluid_out(k_10_1001), .air_in(c_11_0));
valve v_11_2003 (.fluid_in(k_11_2003), .fluid_out(k_10_1001), .air_in(c_11_1));
valve v_11_2004 (.fluid_in(k_11_2004), .fluid_out(k_10_1002), .air_in(c_11_0));
valve v_11_2005 (.fluid_in(k_11_2005), .fluid_out(k_10_1002), .air_in(c_11_1));
valve v_11_2006 (.fluid_in(k_11_2006), .fluid_out(k_10_1003), .air_in(c_11_0));
valve v_11_2007 (.fluid_in(k_11_2007), .fluid_out(k_10_1003), .air_in(c_11_1));
valve v_11_2008 (.fluid_in(k_11_2008), .fluid_out(k_10_1004), .air_in(c_11_0));
valve v_11_2009 (.fluid_in(k_11_2009), .fluid_out(k_10_1004), .air_in(c_11_1));
valve v_11_2010 (.fluid_in(k_11_2010), .fluid_out(k_10_1005), .air_in(c_11_0));
valve v_11_2011 (.fluid_in(k_11_2011), .fluid_out(k_10_1005), .air_in(c_11_1));
valve v_11_2012 (.fluid_in(k_11_2012), .fluid_out(k_10_1006), .air_in(c_11_0));
valve v_11_2013 (.fluid_in(k_11_2013), .fluid_out(k_10_1006), .air_in(c_11_1));
valve v_11_2014 (.fluid_in(k_11_2014), .fluid_out(k_10_1007), .air_in(c_11_0));
valve v_11_2015 (.fluid_in(k_11_2015), .fluid_out(k_10_1007), .air_in(c_11_1));
valve v_11_2016 (.fluid_in(k_11_2016), .fluid_out(k_10_1008), .air_in(c_11_0));
valve v_11_2017 (.fluid_in(k_11_2017), .fluid_out(k_10_1008), .air_in(c_11_1));
valve v_11_2018 (.fluid_in(k_11_2018), .fluid_out(k_10_1009), .air_in(c_11_0));
valve v_11_2019 (.fluid_in(k_11_2019), .fluid_out(k_10_1009), .air_in(c_11_1));
valve v_11_2020 (.fluid_in(k_11_2020), .fluid_out(k_10_1010), .air_in(c_11_0));
valve v_11_2021 (.fluid_in(k_11_2021), .fluid_out(k_10_1010), .air_in(c_11_1));
valve v_11_2022 (.fluid_in(k_11_2022), .fluid_out(k_10_1011), .air_in(c_11_0));
valve v_11_2023 (.fluid_in(k_11_2023), .fluid_out(k_10_1011), .air_in(c_11_1));
valve v_11_2024 (.fluid_in(k_11_2024), .fluid_out(k_10_1012), .air_in(c_11_0));
valve v_11_2025 (.fluid_in(k_11_2025), .fluid_out(k_10_1012), .air_in(c_11_1));
valve v_11_2026 (.fluid_in(k_11_2026), .fluid_out(k_10_1013), .air_in(c_11_0));
valve v_11_2027 (.fluid_in(k_11_2027), .fluid_out(k_10_1013), .air_in(c_11_1));
valve v_11_2028 (.fluid_in(k_11_2028), .fluid_out(k_10_1014), .air_in(c_11_0));
valve v_11_2029 (.fluid_in(k_11_2029), .fluid_out(k_10_1014), .air_in(c_11_1));
valve v_11_2030 (.fluid_in(k_11_2030), .fluid_out(k_10_1015), .air_in(c_11_0));
valve v_11_2031 (.fluid_in(k_11_2031), .fluid_out(k_10_1015), .air_in(c_11_1));
valve v_11_2032 (.fluid_in(k_11_2032), .fluid_out(k_10_1016), .air_in(c_11_0));
valve v_11_2033 (.fluid_in(k_11_2033), .fluid_out(k_10_1016), .air_in(c_11_1));
valve v_11_2034 (.fluid_in(k_11_2034), .fluid_out(k_10_1017), .air_in(c_11_0));
valve v_11_2035 (.fluid_in(k_11_2035), .fluid_out(k_10_1017), .air_in(c_11_1));
valve v_11_2036 (.fluid_in(k_11_2036), .fluid_out(k_10_1018), .air_in(c_11_0));
valve v_11_2037 (.fluid_in(k_11_2037), .fluid_out(k_10_1018), .air_in(c_11_1));
valve v_11_2038 (.fluid_in(k_11_2038), .fluid_out(k_10_1019), .air_in(c_11_0));
valve v_11_2039 (.fluid_in(k_11_2039), .fluid_out(k_10_1019), .air_in(c_11_1));
valve v_11_2040 (.fluid_in(k_11_2040), .fluid_out(k_10_1020), .air_in(c_11_0));
valve v_11_2041 (.fluid_in(k_11_2041), .fluid_out(k_10_1020), .air_in(c_11_1));
valve v_11_2042 (.fluid_in(k_11_2042), .fluid_out(k_10_1021), .air_in(c_11_0));
valve v_11_2043 (.fluid_in(k_11_2043), .fluid_out(k_10_1021), .air_in(c_11_1));
valve v_11_2044 (.fluid_in(k_11_2044), .fluid_out(k_10_1022), .air_in(c_11_0));
valve v_11_2045 (.fluid_in(k_11_2045), .fluid_out(k_10_1022), .air_in(c_11_1));
valve v_11_2046 (.fluid_in(k_11_2046), .fluid_out(k_10_1023), .air_in(c_11_0));
valve v_11_2047 (.fluid_in(k_11_2047), .fluid_out(k_10_1023), .air_in(c_11_1));
valve v_12_0 (.fluid_in(k_12_0), .fluid_out(k_11_0), .air_in(c_12_0));
valve v_12_1 (.fluid_in(k_12_1), .fluid_out(k_11_0), .air_in(c_12_1));
valve v_12_2 (.fluid_in(k_12_2), .fluid_out(k_11_1), .air_in(c_12_0));
valve v_12_3 (.fluid_in(k_12_3), .fluid_out(k_11_1), .air_in(c_12_1));
valve v_12_4 (.fluid_in(k_12_4), .fluid_out(k_11_2), .air_in(c_12_0));
valve v_12_5 (.fluid_in(k_12_5), .fluid_out(k_11_2), .air_in(c_12_1));
valve v_12_6 (.fluid_in(k_12_6), .fluid_out(k_11_3), .air_in(c_12_0));
valve v_12_7 (.fluid_in(k_12_7), .fluid_out(k_11_3), .air_in(c_12_1));
valve v_12_8 (.fluid_in(k_12_8), .fluid_out(k_11_4), .air_in(c_12_0));
valve v_12_9 (.fluid_in(k_12_9), .fluid_out(k_11_4), .air_in(c_12_1));
valve v_12_10 (.fluid_in(k_12_10), .fluid_out(k_11_5), .air_in(c_12_0));
valve v_12_11 (.fluid_in(k_12_11), .fluid_out(k_11_5), .air_in(c_12_1));
valve v_12_12 (.fluid_in(k_12_12), .fluid_out(k_11_6), .air_in(c_12_0));
valve v_12_13 (.fluid_in(k_12_13), .fluid_out(k_11_6), .air_in(c_12_1));
valve v_12_14 (.fluid_in(k_12_14), .fluid_out(k_11_7), .air_in(c_12_0));
valve v_12_15 (.fluid_in(k_12_15), .fluid_out(k_11_7), .air_in(c_12_1));
valve v_12_16 (.fluid_in(k_12_16), .fluid_out(k_11_8), .air_in(c_12_0));
valve v_12_17 (.fluid_in(k_12_17), .fluid_out(k_11_8), .air_in(c_12_1));
valve v_12_18 (.fluid_in(k_12_18), .fluid_out(k_11_9), .air_in(c_12_0));
valve v_12_19 (.fluid_in(k_12_19), .fluid_out(k_11_9), .air_in(c_12_1));
valve v_12_20 (.fluid_in(k_12_20), .fluid_out(k_11_10), .air_in(c_12_0));
valve v_12_21 (.fluid_in(k_12_21), .fluid_out(k_11_10), .air_in(c_12_1));
valve v_12_22 (.fluid_in(k_12_22), .fluid_out(k_11_11), .air_in(c_12_0));
valve v_12_23 (.fluid_in(k_12_23), .fluid_out(k_11_11), .air_in(c_12_1));
valve v_12_24 (.fluid_in(k_12_24), .fluid_out(k_11_12), .air_in(c_12_0));
valve v_12_25 (.fluid_in(k_12_25), .fluid_out(k_11_12), .air_in(c_12_1));
valve v_12_26 (.fluid_in(k_12_26), .fluid_out(k_11_13), .air_in(c_12_0));
valve v_12_27 (.fluid_in(k_12_27), .fluid_out(k_11_13), .air_in(c_12_1));
valve v_12_28 (.fluid_in(k_12_28), .fluid_out(k_11_14), .air_in(c_12_0));
valve v_12_29 (.fluid_in(k_12_29), .fluid_out(k_11_14), .air_in(c_12_1));
valve v_12_30 (.fluid_in(k_12_30), .fluid_out(k_11_15), .air_in(c_12_0));
valve v_12_31 (.fluid_in(k_12_31), .fluid_out(k_11_15), .air_in(c_12_1));
valve v_12_32 (.fluid_in(k_12_32), .fluid_out(k_11_16), .air_in(c_12_0));
valve v_12_33 (.fluid_in(k_12_33), .fluid_out(k_11_16), .air_in(c_12_1));
valve v_12_34 (.fluid_in(k_12_34), .fluid_out(k_11_17), .air_in(c_12_0));
valve v_12_35 (.fluid_in(k_12_35), .fluid_out(k_11_17), .air_in(c_12_1));
valve v_12_36 (.fluid_in(k_12_36), .fluid_out(k_11_18), .air_in(c_12_0));
valve v_12_37 (.fluid_in(k_12_37), .fluid_out(k_11_18), .air_in(c_12_1));
valve v_12_38 (.fluid_in(k_12_38), .fluid_out(k_11_19), .air_in(c_12_0));
valve v_12_39 (.fluid_in(k_12_39), .fluid_out(k_11_19), .air_in(c_12_1));
valve v_12_40 (.fluid_in(k_12_40), .fluid_out(k_11_20), .air_in(c_12_0));
valve v_12_41 (.fluid_in(k_12_41), .fluid_out(k_11_20), .air_in(c_12_1));
valve v_12_42 (.fluid_in(k_12_42), .fluid_out(k_11_21), .air_in(c_12_0));
valve v_12_43 (.fluid_in(k_12_43), .fluid_out(k_11_21), .air_in(c_12_1));
valve v_12_44 (.fluid_in(k_12_44), .fluid_out(k_11_22), .air_in(c_12_0));
valve v_12_45 (.fluid_in(k_12_45), .fluid_out(k_11_22), .air_in(c_12_1));
valve v_12_46 (.fluid_in(k_12_46), .fluid_out(k_11_23), .air_in(c_12_0));
valve v_12_47 (.fluid_in(k_12_47), .fluid_out(k_11_23), .air_in(c_12_1));
valve v_12_48 (.fluid_in(k_12_48), .fluid_out(k_11_24), .air_in(c_12_0));
valve v_12_49 (.fluid_in(k_12_49), .fluid_out(k_11_24), .air_in(c_12_1));
valve v_12_50 (.fluid_in(k_12_50), .fluid_out(k_11_25), .air_in(c_12_0));
valve v_12_51 (.fluid_in(k_12_51), .fluid_out(k_11_25), .air_in(c_12_1));
valve v_12_52 (.fluid_in(k_12_52), .fluid_out(k_11_26), .air_in(c_12_0));
valve v_12_53 (.fluid_in(k_12_53), .fluid_out(k_11_26), .air_in(c_12_1));
valve v_12_54 (.fluid_in(k_12_54), .fluid_out(k_11_27), .air_in(c_12_0));
valve v_12_55 (.fluid_in(k_12_55), .fluid_out(k_11_27), .air_in(c_12_1));
valve v_12_56 (.fluid_in(k_12_56), .fluid_out(k_11_28), .air_in(c_12_0));
valve v_12_57 (.fluid_in(k_12_57), .fluid_out(k_11_28), .air_in(c_12_1));
valve v_12_58 (.fluid_in(k_12_58), .fluid_out(k_11_29), .air_in(c_12_0));
valve v_12_59 (.fluid_in(k_12_59), .fluid_out(k_11_29), .air_in(c_12_1));
valve v_12_60 (.fluid_in(k_12_60), .fluid_out(k_11_30), .air_in(c_12_0));
valve v_12_61 (.fluid_in(k_12_61), .fluid_out(k_11_30), .air_in(c_12_1));
valve v_12_62 (.fluid_in(k_12_62), .fluid_out(k_11_31), .air_in(c_12_0));
valve v_12_63 (.fluid_in(k_12_63), .fluid_out(k_11_31), .air_in(c_12_1));
valve v_12_64 (.fluid_in(k_12_64), .fluid_out(k_11_32), .air_in(c_12_0));
valve v_12_65 (.fluid_in(k_12_65), .fluid_out(k_11_32), .air_in(c_12_1));
valve v_12_66 (.fluid_in(k_12_66), .fluid_out(k_11_33), .air_in(c_12_0));
valve v_12_67 (.fluid_in(k_12_67), .fluid_out(k_11_33), .air_in(c_12_1));
valve v_12_68 (.fluid_in(k_12_68), .fluid_out(k_11_34), .air_in(c_12_0));
valve v_12_69 (.fluid_in(k_12_69), .fluid_out(k_11_34), .air_in(c_12_1));
valve v_12_70 (.fluid_in(k_12_70), .fluid_out(k_11_35), .air_in(c_12_0));
valve v_12_71 (.fluid_in(k_12_71), .fluid_out(k_11_35), .air_in(c_12_1));
valve v_12_72 (.fluid_in(k_12_72), .fluid_out(k_11_36), .air_in(c_12_0));
valve v_12_73 (.fluid_in(k_12_73), .fluid_out(k_11_36), .air_in(c_12_1));
valve v_12_74 (.fluid_in(k_12_74), .fluid_out(k_11_37), .air_in(c_12_0));
valve v_12_75 (.fluid_in(k_12_75), .fluid_out(k_11_37), .air_in(c_12_1));
valve v_12_76 (.fluid_in(k_12_76), .fluid_out(k_11_38), .air_in(c_12_0));
valve v_12_77 (.fluid_in(k_12_77), .fluid_out(k_11_38), .air_in(c_12_1));
valve v_12_78 (.fluid_in(k_12_78), .fluid_out(k_11_39), .air_in(c_12_0));
valve v_12_79 (.fluid_in(k_12_79), .fluid_out(k_11_39), .air_in(c_12_1));
valve v_12_80 (.fluid_in(k_12_80), .fluid_out(k_11_40), .air_in(c_12_0));
valve v_12_81 (.fluid_in(k_12_81), .fluid_out(k_11_40), .air_in(c_12_1));
valve v_12_82 (.fluid_in(k_12_82), .fluid_out(k_11_41), .air_in(c_12_0));
valve v_12_83 (.fluid_in(k_12_83), .fluid_out(k_11_41), .air_in(c_12_1));
valve v_12_84 (.fluid_in(k_12_84), .fluid_out(k_11_42), .air_in(c_12_0));
valve v_12_85 (.fluid_in(k_12_85), .fluid_out(k_11_42), .air_in(c_12_1));
valve v_12_86 (.fluid_in(k_12_86), .fluid_out(k_11_43), .air_in(c_12_0));
valve v_12_87 (.fluid_in(k_12_87), .fluid_out(k_11_43), .air_in(c_12_1));
valve v_12_88 (.fluid_in(k_12_88), .fluid_out(k_11_44), .air_in(c_12_0));
valve v_12_89 (.fluid_in(k_12_89), .fluid_out(k_11_44), .air_in(c_12_1));
valve v_12_90 (.fluid_in(k_12_90), .fluid_out(k_11_45), .air_in(c_12_0));
valve v_12_91 (.fluid_in(k_12_91), .fluid_out(k_11_45), .air_in(c_12_1));
valve v_12_92 (.fluid_in(k_12_92), .fluid_out(k_11_46), .air_in(c_12_0));
valve v_12_93 (.fluid_in(k_12_93), .fluid_out(k_11_46), .air_in(c_12_1));
valve v_12_94 (.fluid_in(k_12_94), .fluid_out(k_11_47), .air_in(c_12_0));
valve v_12_95 (.fluid_in(k_12_95), .fluid_out(k_11_47), .air_in(c_12_1));
valve v_12_96 (.fluid_in(k_12_96), .fluid_out(k_11_48), .air_in(c_12_0));
valve v_12_97 (.fluid_in(k_12_97), .fluid_out(k_11_48), .air_in(c_12_1));
valve v_12_98 (.fluid_in(k_12_98), .fluid_out(k_11_49), .air_in(c_12_0));
valve v_12_99 (.fluid_in(k_12_99), .fluid_out(k_11_49), .air_in(c_12_1));
valve v_12_100 (.fluid_in(k_12_100), .fluid_out(k_11_50), .air_in(c_12_0));
valve v_12_101 (.fluid_in(k_12_101), .fluid_out(k_11_50), .air_in(c_12_1));
valve v_12_102 (.fluid_in(k_12_102), .fluid_out(k_11_51), .air_in(c_12_0));
valve v_12_103 (.fluid_in(k_12_103), .fluid_out(k_11_51), .air_in(c_12_1));
valve v_12_104 (.fluid_in(k_12_104), .fluid_out(k_11_52), .air_in(c_12_0));
valve v_12_105 (.fluid_in(k_12_105), .fluid_out(k_11_52), .air_in(c_12_1));
valve v_12_106 (.fluid_in(k_12_106), .fluid_out(k_11_53), .air_in(c_12_0));
valve v_12_107 (.fluid_in(k_12_107), .fluid_out(k_11_53), .air_in(c_12_1));
valve v_12_108 (.fluid_in(k_12_108), .fluid_out(k_11_54), .air_in(c_12_0));
valve v_12_109 (.fluid_in(k_12_109), .fluid_out(k_11_54), .air_in(c_12_1));
valve v_12_110 (.fluid_in(k_12_110), .fluid_out(k_11_55), .air_in(c_12_0));
valve v_12_111 (.fluid_in(k_12_111), .fluid_out(k_11_55), .air_in(c_12_1));
valve v_12_112 (.fluid_in(k_12_112), .fluid_out(k_11_56), .air_in(c_12_0));
valve v_12_113 (.fluid_in(k_12_113), .fluid_out(k_11_56), .air_in(c_12_1));
valve v_12_114 (.fluid_in(k_12_114), .fluid_out(k_11_57), .air_in(c_12_0));
valve v_12_115 (.fluid_in(k_12_115), .fluid_out(k_11_57), .air_in(c_12_1));
valve v_12_116 (.fluid_in(k_12_116), .fluid_out(k_11_58), .air_in(c_12_0));
valve v_12_117 (.fluid_in(k_12_117), .fluid_out(k_11_58), .air_in(c_12_1));
valve v_12_118 (.fluid_in(k_12_118), .fluid_out(k_11_59), .air_in(c_12_0));
valve v_12_119 (.fluid_in(k_12_119), .fluid_out(k_11_59), .air_in(c_12_1));
valve v_12_120 (.fluid_in(k_12_120), .fluid_out(k_11_60), .air_in(c_12_0));
valve v_12_121 (.fluid_in(k_12_121), .fluid_out(k_11_60), .air_in(c_12_1));
valve v_12_122 (.fluid_in(k_12_122), .fluid_out(k_11_61), .air_in(c_12_0));
valve v_12_123 (.fluid_in(k_12_123), .fluid_out(k_11_61), .air_in(c_12_1));
valve v_12_124 (.fluid_in(k_12_124), .fluid_out(k_11_62), .air_in(c_12_0));
valve v_12_125 (.fluid_in(k_12_125), .fluid_out(k_11_62), .air_in(c_12_1));
valve v_12_126 (.fluid_in(k_12_126), .fluid_out(k_11_63), .air_in(c_12_0));
valve v_12_127 (.fluid_in(k_12_127), .fluid_out(k_11_63), .air_in(c_12_1));
valve v_12_128 (.fluid_in(k_12_128), .fluid_out(k_11_64), .air_in(c_12_0));
valve v_12_129 (.fluid_in(k_12_129), .fluid_out(k_11_64), .air_in(c_12_1));
valve v_12_130 (.fluid_in(k_12_130), .fluid_out(k_11_65), .air_in(c_12_0));
valve v_12_131 (.fluid_in(k_12_131), .fluid_out(k_11_65), .air_in(c_12_1));
valve v_12_132 (.fluid_in(k_12_132), .fluid_out(k_11_66), .air_in(c_12_0));
valve v_12_133 (.fluid_in(k_12_133), .fluid_out(k_11_66), .air_in(c_12_1));
valve v_12_134 (.fluid_in(k_12_134), .fluid_out(k_11_67), .air_in(c_12_0));
valve v_12_135 (.fluid_in(k_12_135), .fluid_out(k_11_67), .air_in(c_12_1));
valve v_12_136 (.fluid_in(k_12_136), .fluid_out(k_11_68), .air_in(c_12_0));
valve v_12_137 (.fluid_in(k_12_137), .fluid_out(k_11_68), .air_in(c_12_1));
valve v_12_138 (.fluid_in(k_12_138), .fluid_out(k_11_69), .air_in(c_12_0));
valve v_12_139 (.fluid_in(k_12_139), .fluid_out(k_11_69), .air_in(c_12_1));
valve v_12_140 (.fluid_in(k_12_140), .fluid_out(k_11_70), .air_in(c_12_0));
valve v_12_141 (.fluid_in(k_12_141), .fluid_out(k_11_70), .air_in(c_12_1));
valve v_12_142 (.fluid_in(k_12_142), .fluid_out(k_11_71), .air_in(c_12_0));
valve v_12_143 (.fluid_in(k_12_143), .fluid_out(k_11_71), .air_in(c_12_1));
valve v_12_144 (.fluid_in(k_12_144), .fluid_out(k_11_72), .air_in(c_12_0));
valve v_12_145 (.fluid_in(k_12_145), .fluid_out(k_11_72), .air_in(c_12_1));
valve v_12_146 (.fluid_in(k_12_146), .fluid_out(k_11_73), .air_in(c_12_0));
valve v_12_147 (.fluid_in(k_12_147), .fluid_out(k_11_73), .air_in(c_12_1));
valve v_12_148 (.fluid_in(k_12_148), .fluid_out(k_11_74), .air_in(c_12_0));
valve v_12_149 (.fluid_in(k_12_149), .fluid_out(k_11_74), .air_in(c_12_1));
valve v_12_150 (.fluid_in(k_12_150), .fluid_out(k_11_75), .air_in(c_12_0));
valve v_12_151 (.fluid_in(k_12_151), .fluid_out(k_11_75), .air_in(c_12_1));
valve v_12_152 (.fluid_in(k_12_152), .fluid_out(k_11_76), .air_in(c_12_0));
valve v_12_153 (.fluid_in(k_12_153), .fluid_out(k_11_76), .air_in(c_12_1));
valve v_12_154 (.fluid_in(k_12_154), .fluid_out(k_11_77), .air_in(c_12_0));
valve v_12_155 (.fluid_in(k_12_155), .fluid_out(k_11_77), .air_in(c_12_1));
valve v_12_156 (.fluid_in(k_12_156), .fluid_out(k_11_78), .air_in(c_12_0));
valve v_12_157 (.fluid_in(k_12_157), .fluid_out(k_11_78), .air_in(c_12_1));
valve v_12_158 (.fluid_in(k_12_158), .fluid_out(k_11_79), .air_in(c_12_0));
valve v_12_159 (.fluid_in(k_12_159), .fluid_out(k_11_79), .air_in(c_12_1));
valve v_12_160 (.fluid_in(k_12_160), .fluid_out(k_11_80), .air_in(c_12_0));
valve v_12_161 (.fluid_in(k_12_161), .fluid_out(k_11_80), .air_in(c_12_1));
valve v_12_162 (.fluid_in(k_12_162), .fluid_out(k_11_81), .air_in(c_12_0));
valve v_12_163 (.fluid_in(k_12_163), .fluid_out(k_11_81), .air_in(c_12_1));
valve v_12_164 (.fluid_in(k_12_164), .fluid_out(k_11_82), .air_in(c_12_0));
valve v_12_165 (.fluid_in(k_12_165), .fluid_out(k_11_82), .air_in(c_12_1));
valve v_12_166 (.fluid_in(k_12_166), .fluid_out(k_11_83), .air_in(c_12_0));
valve v_12_167 (.fluid_in(k_12_167), .fluid_out(k_11_83), .air_in(c_12_1));
valve v_12_168 (.fluid_in(k_12_168), .fluid_out(k_11_84), .air_in(c_12_0));
valve v_12_169 (.fluid_in(k_12_169), .fluid_out(k_11_84), .air_in(c_12_1));
valve v_12_170 (.fluid_in(k_12_170), .fluid_out(k_11_85), .air_in(c_12_0));
valve v_12_171 (.fluid_in(k_12_171), .fluid_out(k_11_85), .air_in(c_12_1));
valve v_12_172 (.fluid_in(k_12_172), .fluid_out(k_11_86), .air_in(c_12_0));
valve v_12_173 (.fluid_in(k_12_173), .fluid_out(k_11_86), .air_in(c_12_1));
valve v_12_174 (.fluid_in(k_12_174), .fluid_out(k_11_87), .air_in(c_12_0));
valve v_12_175 (.fluid_in(k_12_175), .fluid_out(k_11_87), .air_in(c_12_1));
valve v_12_176 (.fluid_in(k_12_176), .fluid_out(k_11_88), .air_in(c_12_0));
valve v_12_177 (.fluid_in(k_12_177), .fluid_out(k_11_88), .air_in(c_12_1));
valve v_12_178 (.fluid_in(k_12_178), .fluid_out(k_11_89), .air_in(c_12_0));
valve v_12_179 (.fluid_in(k_12_179), .fluid_out(k_11_89), .air_in(c_12_1));
valve v_12_180 (.fluid_in(k_12_180), .fluid_out(k_11_90), .air_in(c_12_0));
valve v_12_181 (.fluid_in(k_12_181), .fluid_out(k_11_90), .air_in(c_12_1));
valve v_12_182 (.fluid_in(k_12_182), .fluid_out(k_11_91), .air_in(c_12_0));
valve v_12_183 (.fluid_in(k_12_183), .fluid_out(k_11_91), .air_in(c_12_1));
valve v_12_184 (.fluid_in(k_12_184), .fluid_out(k_11_92), .air_in(c_12_0));
valve v_12_185 (.fluid_in(k_12_185), .fluid_out(k_11_92), .air_in(c_12_1));
valve v_12_186 (.fluid_in(k_12_186), .fluid_out(k_11_93), .air_in(c_12_0));
valve v_12_187 (.fluid_in(k_12_187), .fluid_out(k_11_93), .air_in(c_12_1));
valve v_12_188 (.fluid_in(k_12_188), .fluid_out(k_11_94), .air_in(c_12_0));
valve v_12_189 (.fluid_in(k_12_189), .fluid_out(k_11_94), .air_in(c_12_1));
valve v_12_190 (.fluid_in(k_12_190), .fluid_out(k_11_95), .air_in(c_12_0));
valve v_12_191 (.fluid_in(k_12_191), .fluid_out(k_11_95), .air_in(c_12_1));
valve v_12_192 (.fluid_in(k_12_192), .fluid_out(k_11_96), .air_in(c_12_0));
valve v_12_193 (.fluid_in(k_12_193), .fluid_out(k_11_96), .air_in(c_12_1));
valve v_12_194 (.fluid_in(k_12_194), .fluid_out(k_11_97), .air_in(c_12_0));
valve v_12_195 (.fluid_in(k_12_195), .fluid_out(k_11_97), .air_in(c_12_1));
valve v_12_196 (.fluid_in(k_12_196), .fluid_out(k_11_98), .air_in(c_12_0));
valve v_12_197 (.fluid_in(k_12_197), .fluid_out(k_11_98), .air_in(c_12_1));
valve v_12_198 (.fluid_in(k_12_198), .fluid_out(k_11_99), .air_in(c_12_0));
valve v_12_199 (.fluid_in(k_12_199), .fluid_out(k_11_99), .air_in(c_12_1));
valve v_12_200 (.fluid_in(k_12_200), .fluid_out(k_11_100), .air_in(c_12_0));
valve v_12_201 (.fluid_in(k_12_201), .fluid_out(k_11_100), .air_in(c_12_1));
valve v_12_202 (.fluid_in(k_12_202), .fluid_out(k_11_101), .air_in(c_12_0));
valve v_12_203 (.fluid_in(k_12_203), .fluid_out(k_11_101), .air_in(c_12_1));
valve v_12_204 (.fluid_in(k_12_204), .fluid_out(k_11_102), .air_in(c_12_0));
valve v_12_205 (.fluid_in(k_12_205), .fluid_out(k_11_102), .air_in(c_12_1));
valve v_12_206 (.fluid_in(k_12_206), .fluid_out(k_11_103), .air_in(c_12_0));
valve v_12_207 (.fluid_in(k_12_207), .fluid_out(k_11_103), .air_in(c_12_1));
valve v_12_208 (.fluid_in(k_12_208), .fluid_out(k_11_104), .air_in(c_12_0));
valve v_12_209 (.fluid_in(k_12_209), .fluid_out(k_11_104), .air_in(c_12_1));
valve v_12_210 (.fluid_in(k_12_210), .fluid_out(k_11_105), .air_in(c_12_0));
valve v_12_211 (.fluid_in(k_12_211), .fluid_out(k_11_105), .air_in(c_12_1));
valve v_12_212 (.fluid_in(k_12_212), .fluid_out(k_11_106), .air_in(c_12_0));
valve v_12_213 (.fluid_in(k_12_213), .fluid_out(k_11_106), .air_in(c_12_1));
valve v_12_214 (.fluid_in(k_12_214), .fluid_out(k_11_107), .air_in(c_12_0));
valve v_12_215 (.fluid_in(k_12_215), .fluid_out(k_11_107), .air_in(c_12_1));
valve v_12_216 (.fluid_in(k_12_216), .fluid_out(k_11_108), .air_in(c_12_0));
valve v_12_217 (.fluid_in(k_12_217), .fluid_out(k_11_108), .air_in(c_12_1));
valve v_12_218 (.fluid_in(k_12_218), .fluid_out(k_11_109), .air_in(c_12_0));
valve v_12_219 (.fluid_in(k_12_219), .fluid_out(k_11_109), .air_in(c_12_1));
valve v_12_220 (.fluid_in(k_12_220), .fluid_out(k_11_110), .air_in(c_12_0));
valve v_12_221 (.fluid_in(k_12_221), .fluid_out(k_11_110), .air_in(c_12_1));
valve v_12_222 (.fluid_in(k_12_222), .fluid_out(k_11_111), .air_in(c_12_0));
valve v_12_223 (.fluid_in(k_12_223), .fluid_out(k_11_111), .air_in(c_12_1));
valve v_12_224 (.fluid_in(k_12_224), .fluid_out(k_11_112), .air_in(c_12_0));
valve v_12_225 (.fluid_in(k_12_225), .fluid_out(k_11_112), .air_in(c_12_1));
valve v_12_226 (.fluid_in(k_12_226), .fluid_out(k_11_113), .air_in(c_12_0));
valve v_12_227 (.fluid_in(k_12_227), .fluid_out(k_11_113), .air_in(c_12_1));
valve v_12_228 (.fluid_in(k_12_228), .fluid_out(k_11_114), .air_in(c_12_0));
valve v_12_229 (.fluid_in(k_12_229), .fluid_out(k_11_114), .air_in(c_12_1));
valve v_12_230 (.fluid_in(k_12_230), .fluid_out(k_11_115), .air_in(c_12_0));
valve v_12_231 (.fluid_in(k_12_231), .fluid_out(k_11_115), .air_in(c_12_1));
valve v_12_232 (.fluid_in(k_12_232), .fluid_out(k_11_116), .air_in(c_12_0));
valve v_12_233 (.fluid_in(k_12_233), .fluid_out(k_11_116), .air_in(c_12_1));
valve v_12_234 (.fluid_in(k_12_234), .fluid_out(k_11_117), .air_in(c_12_0));
valve v_12_235 (.fluid_in(k_12_235), .fluid_out(k_11_117), .air_in(c_12_1));
valve v_12_236 (.fluid_in(k_12_236), .fluid_out(k_11_118), .air_in(c_12_0));
valve v_12_237 (.fluid_in(k_12_237), .fluid_out(k_11_118), .air_in(c_12_1));
valve v_12_238 (.fluid_in(k_12_238), .fluid_out(k_11_119), .air_in(c_12_0));
valve v_12_239 (.fluid_in(k_12_239), .fluid_out(k_11_119), .air_in(c_12_1));
valve v_12_240 (.fluid_in(k_12_240), .fluid_out(k_11_120), .air_in(c_12_0));
valve v_12_241 (.fluid_in(k_12_241), .fluid_out(k_11_120), .air_in(c_12_1));
valve v_12_242 (.fluid_in(k_12_242), .fluid_out(k_11_121), .air_in(c_12_0));
valve v_12_243 (.fluid_in(k_12_243), .fluid_out(k_11_121), .air_in(c_12_1));
valve v_12_244 (.fluid_in(k_12_244), .fluid_out(k_11_122), .air_in(c_12_0));
valve v_12_245 (.fluid_in(k_12_245), .fluid_out(k_11_122), .air_in(c_12_1));
valve v_12_246 (.fluid_in(k_12_246), .fluid_out(k_11_123), .air_in(c_12_0));
valve v_12_247 (.fluid_in(k_12_247), .fluid_out(k_11_123), .air_in(c_12_1));
valve v_12_248 (.fluid_in(k_12_248), .fluid_out(k_11_124), .air_in(c_12_0));
valve v_12_249 (.fluid_in(k_12_249), .fluid_out(k_11_124), .air_in(c_12_1));
valve v_12_250 (.fluid_in(k_12_250), .fluid_out(k_11_125), .air_in(c_12_0));
valve v_12_251 (.fluid_in(k_12_251), .fluid_out(k_11_125), .air_in(c_12_1));
valve v_12_252 (.fluid_in(k_12_252), .fluid_out(k_11_126), .air_in(c_12_0));
valve v_12_253 (.fluid_in(k_12_253), .fluid_out(k_11_126), .air_in(c_12_1));
valve v_12_254 (.fluid_in(k_12_254), .fluid_out(k_11_127), .air_in(c_12_0));
valve v_12_255 (.fluid_in(k_12_255), .fluid_out(k_11_127), .air_in(c_12_1));
valve v_12_256 (.fluid_in(k_12_256), .fluid_out(k_11_128), .air_in(c_12_0));
valve v_12_257 (.fluid_in(k_12_257), .fluid_out(k_11_128), .air_in(c_12_1));
valve v_12_258 (.fluid_in(k_12_258), .fluid_out(k_11_129), .air_in(c_12_0));
valve v_12_259 (.fluid_in(k_12_259), .fluid_out(k_11_129), .air_in(c_12_1));
valve v_12_260 (.fluid_in(k_12_260), .fluid_out(k_11_130), .air_in(c_12_0));
valve v_12_261 (.fluid_in(k_12_261), .fluid_out(k_11_130), .air_in(c_12_1));
valve v_12_262 (.fluid_in(k_12_262), .fluid_out(k_11_131), .air_in(c_12_0));
valve v_12_263 (.fluid_in(k_12_263), .fluid_out(k_11_131), .air_in(c_12_1));
valve v_12_264 (.fluid_in(k_12_264), .fluid_out(k_11_132), .air_in(c_12_0));
valve v_12_265 (.fluid_in(k_12_265), .fluid_out(k_11_132), .air_in(c_12_1));
valve v_12_266 (.fluid_in(k_12_266), .fluid_out(k_11_133), .air_in(c_12_0));
valve v_12_267 (.fluid_in(k_12_267), .fluid_out(k_11_133), .air_in(c_12_1));
valve v_12_268 (.fluid_in(k_12_268), .fluid_out(k_11_134), .air_in(c_12_0));
valve v_12_269 (.fluid_in(k_12_269), .fluid_out(k_11_134), .air_in(c_12_1));
valve v_12_270 (.fluid_in(k_12_270), .fluid_out(k_11_135), .air_in(c_12_0));
valve v_12_271 (.fluid_in(k_12_271), .fluid_out(k_11_135), .air_in(c_12_1));
valve v_12_272 (.fluid_in(k_12_272), .fluid_out(k_11_136), .air_in(c_12_0));
valve v_12_273 (.fluid_in(k_12_273), .fluid_out(k_11_136), .air_in(c_12_1));
valve v_12_274 (.fluid_in(k_12_274), .fluid_out(k_11_137), .air_in(c_12_0));
valve v_12_275 (.fluid_in(k_12_275), .fluid_out(k_11_137), .air_in(c_12_1));
valve v_12_276 (.fluid_in(k_12_276), .fluid_out(k_11_138), .air_in(c_12_0));
valve v_12_277 (.fluid_in(k_12_277), .fluid_out(k_11_138), .air_in(c_12_1));
valve v_12_278 (.fluid_in(k_12_278), .fluid_out(k_11_139), .air_in(c_12_0));
valve v_12_279 (.fluid_in(k_12_279), .fluid_out(k_11_139), .air_in(c_12_1));
valve v_12_280 (.fluid_in(k_12_280), .fluid_out(k_11_140), .air_in(c_12_0));
valve v_12_281 (.fluid_in(k_12_281), .fluid_out(k_11_140), .air_in(c_12_1));
valve v_12_282 (.fluid_in(k_12_282), .fluid_out(k_11_141), .air_in(c_12_0));
valve v_12_283 (.fluid_in(k_12_283), .fluid_out(k_11_141), .air_in(c_12_1));
valve v_12_284 (.fluid_in(k_12_284), .fluid_out(k_11_142), .air_in(c_12_0));
valve v_12_285 (.fluid_in(k_12_285), .fluid_out(k_11_142), .air_in(c_12_1));
valve v_12_286 (.fluid_in(k_12_286), .fluid_out(k_11_143), .air_in(c_12_0));
valve v_12_287 (.fluid_in(k_12_287), .fluid_out(k_11_143), .air_in(c_12_1));
valve v_12_288 (.fluid_in(k_12_288), .fluid_out(k_11_144), .air_in(c_12_0));
valve v_12_289 (.fluid_in(k_12_289), .fluid_out(k_11_144), .air_in(c_12_1));
valve v_12_290 (.fluid_in(k_12_290), .fluid_out(k_11_145), .air_in(c_12_0));
valve v_12_291 (.fluid_in(k_12_291), .fluid_out(k_11_145), .air_in(c_12_1));
valve v_12_292 (.fluid_in(k_12_292), .fluid_out(k_11_146), .air_in(c_12_0));
valve v_12_293 (.fluid_in(k_12_293), .fluid_out(k_11_146), .air_in(c_12_1));
valve v_12_294 (.fluid_in(k_12_294), .fluid_out(k_11_147), .air_in(c_12_0));
valve v_12_295 (.fluid_in(k_12_295), .fluid_out(k_11_147), .air_in(c_12_1));
valve v_12_296 (.fluid_in(k_12_296), .fluid_out(k_11_148), .air_in(c_12_0));
valve v_12_297 (.fluid_in(k_12_297), .fluid_out(k_11_148), .air_in(c_12_1));
valve v_12_298 (.fluid_in(k_12_298), .fluid_out(k_11_149), .air_in(c_12_0));
valve v_12_299 (.fluid_in(k_12_299), .fluid_out(k_11_149), .air_in(c_12_1));
valve v_12_300 (.fluid_in(k_12_300), .fluid_out(k_11_150), .air_in(c_12_0));
valve v_12_301 (.fluid_in(k_12_301), .fluid_out(k_11_150), .air_in(c_12_1));
valve v_12_302 (.fluid_in(k_12_302), .fluid_out(k_11_151), .air_in(c_12_0));
valve v_12_303 (.fluid_in(k_12_303), .fluid_out(k_11_151), .air_in(c_12_1));
valve v_12_304 (.fluid_in(k_12_304), .fluid_out(k_11_152), .air_in(c_12_0));
valve v_12_305 (.fluid_in(k_12_305), .fluid_out(k_11_152), .air_in(c_12_1));
valve v_12_306 (.fluid_in(k_12_306), .fluid_out(k_11_153), .air_in(c_12_0));
valve v_12_307 (.fluid_in(k_12_307), .fluid_out(k_11_153), .air_in(c_12_1));
valve v_12_308 (.fluid_in(k_12_308), .fluid_out(k_11_154), .air_in(c_12_0));
valve v_12_309 (.fluid_in(k_12_309), .fluid_out(k_11_154), .air_in(c_12_1));
valve v_12_310 (.fluid_in(k_12_310), .fluid_out(k_11_155), .air_in(c_12_0));
valve v_12_311 (.fluid_in(k_12_311), .fluid_out(k_11_155), .air_in(c_12_1));
valve v_12_312 (.fluid_in(k_12_312), .fluid_out(k_11_156), .air_in(c_12_0));
valve v_12_313 (.fluid_in(k_12_313), .fluid_out(k_11_156), .air_in(c_12_1));
valve v_12_314 (.fluid_in(k_12_314), .fluid_out(k_11_157), .air_in(c_12_0));
valve v_12_315 (.fluid_in(k_12_315), .fluid_out(k_11_157), .air_in(c_12_1));
valve v_12_316 (.fluid_in(k_12_316), .fluid_out(k_11_158), .air_in(c_12_0));
valve v_12_317 (.fluid_in(k_12_317), .fluid_out(k_11_158), .air_in(c_12_1));
valve v_12_318 (.fluid_in(k_12_318), .fluid_out(k_11_159), .air_in(c_12_0));
valve v_12_319 (.fluid_in(k_12_319), .fluid_out(k_11_159), .air_in(c_12_1));
valve v_12_320 (.fluid_in(k_12_320), .fluid_out(k_11_160), .air_in(c_12_0));
valve v_12_321 (.fluid_in(k_12_321), .fluid_out(k_11_160), .air_in(c_12_1));
valve v_12_322 (.fluid_in(k_12_322), .fluid_out(k_11_161), .air_in(c_12_0));
valve v_12_323 (.fluid_in(k_12_323), .fluid_out(k_11_161), .air_in(c_12_1));
valve v_12_324 (.fluid_in(k_12_324), .fluid_out(k_11_162), .air_in(c_12_0));
valve v_12_325 (.fluid_in(k_12_325), .fluid_out(k_11_162), .air_in(c_12_1));
valve v_12_326 (.fluid_in(k_12_326), .fluid_out(k_11_163), .air_in(c_12_0));
valve v_12_327 (.fluid_in(k_12_327), .fluid_out(k_11_163), .air_in(c_12_1));
valve v_12_328 (.fluid_in(k_12_328), .fluid_out(k_11_164), .air_in(c_12_0));
valve v_12_329 (.fluid_in(k_12_329), .fluid_out(k_11_164), .air_in(c_12_1));
valve v_12_330 (.fluid_in(k_12_330), .fluid_out(k_11_165), .air_in(c_12_0));
valve v_12_331 (.fluid_in(k_12_331), .fluid_out(k_11_165), .air_in(c_12_1));
valve v_12_332 (.fluid_in(k_12_332), .fluid_out(k_11_166), .air_in(c_12_0));
valve v_12_333 (.fluid_in(k_12_333), .fluid_out(k_11_166), .air_in(c_12_1));
valve v_12_334 (.fluid_in(k_12_334), .fluid_out(k_11_167), .air_in(c_12_0));
valve v_12_335 (.fluid_in(k_12_335), .fluid_out(k_11_167), .air_in(c_12_1));
valve v_12_336 (.fluid_in(k_12_336), .fluid_out(k_11_168), .air_in(c_12_0));
valve v_12_337 (.fluid_in(k_12_337), .fluid_out(k_11_168), .air_in(c_12_1));
valve v_12_338 (.fluid_in(k_12_338), .fluid_out(k_11_169), .air_in(c_12_0));
valve v_12_339 (.fluid_in(k_12_339), .fluid_out(k_11_169), .air_in(c_12_1));
valve v_12_340 (.fluid_in(k_12_340), .fluid_out(k_11_170), .air_in(c_12_0));
valve v_12_341 (.fluid_in(k_12_341), .fluid_out(k_11_170), .air_in(c_12_1));
valve v_12_342 (.fluid_in(k_12_342), .fluid_out(k_11_171), .air_in(c_12_0));
valve v_12_343 (.fluid_in(k_12_343), .fluid_out(k_11_171), .air_in(c_12_1));
valve v_12_344 (.fluid_in(k_12_344), .fluid_out(k_11_172), .air_in(c_12_0));
valve v_12_345 (.fluid_in(k_12_345), .fluid_out(k_11_172), .air_in(c_12_1));
valve v_12_346 (.fluid_in(k_12_346), .fluid_out(k_11_173), .air_in(c_12_0));
valve v_12_347 (.fluid_in(k_12_347), .fluid_out(k_11_173), .air_in(c_12_1));
valve v_12_348 (.fluid_in(k_12_348), .fluid_out(k_11_174), .air_in(c_12_0));
valve v_12_349 (.fluid_in(k_12_349), .fluid_out(k_11_174), .air_in(c_12_1));
valve v_12_350 (.fluid_in(k_12_350), .fluid_out(k_11_175), .air_in(c_12_0));
valve v_12_351 (.fluid_in(k_12_351), .fluid_out(k_11_175), .air_in(c_12_1));
valve v_12_352 (.fluid_in(k_12_352), .fluid_out(k_11_176), .air_in(c_12_0));
valve v_12_353 (.fluid_in(k_12_353), .fluid_out(k_11_176), .air_in(c_12_1));
valve v_12_354 (.fluid_in(k_12_354), .fluid_out(k_11_177), .air_in(c_12_0));
valve v_12_355 (.fluid_in(k_12_355), .fluid_out(k_11_177), .air_in(c_12_1));
valve v_12_356 (.fluid_in(k_12_356), .fluid_out(k_11_178), .air_in(c_12_0));
valve v_12_357 (.fluid_in(k_12_357), .fluid_out(k_11_178), .air_in(c_12_1));
valve v_12_358 (.fluid_in(k_12_358), .fluid_out(k_11_179), .air_in(c_12_0));
valve v_12_359 (.fluid_in(k_12_359), .fluid_out(k_11_179), .air_in(c_12_1));
valve v_12_360 (.fluid_in(k_12_360), .fluid_out(k_11_180), .air_in(c_12_0));
valve v_12_361 (.fluid_in(k_12_361), .fluid_out(k_11_180), .air_in(c_12_1));
valve v_12_362 (.fluid_in(k_12_362), .fluid_out(k_11_181), .air_in(c_12_0));
valve v_12_363 (.fluid_in(k_12_363), .fluid_out(k_11_181), .air_in(c_12_1));
valve v_12_364 (.fluid_in(k_12_364), .fluid_out(k_11_182), .air_in(c_12_0));
valve v_12_365 (.fluid_in(k_12_365), .fluid_out(k_11_182), .air_in(c_12_1));
valve v_12_366 (.fluid_in(k_12_366), .fluid_out(k_11_183), .air_in(c_12_0));
valve v_12_367 (.fluid_in(k_12_367), .fluid_out(k_11_183), .air_in(c_12_1));
valve v_12_368 (.fluid_in(k_12_368), .fluid_out(k_11_184), .air_in(c_12_0));
valve v_12_369 (.fluid_in(k_12_369), .fluid_out(k_11_184), .air_in(c_12_1));
valve v_12_370 (.fluid_in(k_12_370), .fluid_out(k_11_185), .air_in(c_12_0));
valve v_12_371 (.fluid_in(k_12_371), .fluid_out(k_11_185), .air_in(c_12_1));
valve v_12_372 (.fluid_in(k_12_372), .fluid_out(k_11_186), .air_in(c_12_0));
valve v_12_373 (.fluid_in(k_12_373), .fluid_out(k_11_186), .air_in(c_12_1));
valve v_12_374 (.fluid_in(k_12_374), .fluid_out(k_11_187), .air_in(c_12_0));
valve v_12_375 (.fluid_in(k_12_375), .fluid_out(k_11_187), .air_in(c_12_1));
valve v_12_376 (.fluid_in(k_12_376), .fluid_out(k_11_188), .air_in(c_12_0));
valve v_12_377 (.fluid_in(k_12_377), .fluid_out(k_11_188), .air_in(c_12_1));
valve v_12_378 (.fluid_in(k_12_378), .fluid_out(k_11_189), .air_in(c_12_0));
valve v_12_379 (.fluid_in(k_12_379), .fluid_out(k_11_189), .air_in(c_12_1));
valve v_12_380 (.fluid_in(k_12_380), .fluid_out(k_11_190), .air_in(c_12_0));
valve v_12_381 (.fluid_in(k_12_381), .fluid_out(k_11_190), .air_in(c_12_1));
valve v_12_382 (.fluid_in(k_12_382), .fluid_out(k_11_191), .air_in(c_12_0));
valve v_12_383 (.fluid_in(k_12_383), .fluid_out(k_11_191), .air_in(c_12_1));
valve v_12_384 (.fluid_in(k_12_384), .fluid_out(k_11_192), .air_in(c_12_0));
valve v_12_385 (.fluid_in(k_12_385), .fluid_out(k_11_192), .air_in(c_12_1));
valve v_12_386 (.fluid_in(k_12_386), .fluid_out(k_11_193), .air_in(c_12_0));
valve v_12_387 (.fluid_in(k_12_387), .fluid_out(k_11_193), .air_in(c_12_1));
valve v_12_388 (.fluid_in(k_12_388), .fluid_out(k_11_194), .air_in(c_12_0));
valve v_12_389 (.fluid_in(k_12_389), .fluid_out(k_11_194), .air_in(c_12_1));
valve v_12_390 (.fluid_in(k_12_390), .fluid_out(k_11_195), .air_in(c_12_0));
valve v_12_391 (.fluid_in(k_12_391), .fluid_out(k_11_195), .air_in(c_12_1));
valve v_12_392 (.fluid_in(k_12_392), .fluid_out(k_11_196), .air_in(c_12_0));
valve v_12_393 (.fluid_in(k_12_393), .fluid_out(k_11_196), .air_in(c_12_1));
valve v_12_394 (.fluid_in(k_12_394), .fluid_out(k_11_197), .air_in(c_12_0));
valve v_12_395 (.fluid_in(k_12_395), .fluid_out(k_11_197), .air_in(c_12_1));
valve v_12_396 (.fluid_in(k_12_396), .fluid_out(k_11_198), .air_in(c_12_0));
valve v_12_397 (.fluid_in(k_12_397), .fluid_out(k_11_198), .air_in(c_12_1));
valve v_12_398 (.fluid_in(k_12_398), .fluid_out(k_11_199), .air_in(c_12_0));
valve v_12_399 (.fluid_in(k_12_399), .fluid_out(k_11_199), .air_in(c_12_1));
valve v_12_400 (.fluid_in(k_12_400), .fluid_out(k_11_200), .air_in(c_12_0));
valve v_12_401 (.fluid_in(k_12_401), .fluid_out(k_11_200), .air_in(c_12_1));
valve v_12_402 (.fluid_in(k_12_402), .fluid_out(k_11_201), .air_in(c_12_0));
valve v_12_403 (.fluid_in(k_12_403), .fluid_out(k_11_201), .air_in(c_12_1));
valve v_12_404 (.fluid_in(k_12_404), .fluid_out(k_11_202), .air_in(c_12_0));
valve v_12_405 (.fluid_in(k_12_405), .fluid_out(k_11_202), .air_in(c_12_1));
valve v_12_406 (.fluid_in(k_12_406), .fluid_out(k_11_203), .air_in(c_12_0));
valve v_12_407 (.fluid_in(k_12_407), .fluid_out(k_11_203), .air_in(c_12_1));
valve v_12_408 (.fluid_in(k_12_408), .fluid_out(k_11_204), .air_in(c_12_0));
valve v_12_409 (.fluid_in(k_12_409), .fluid_out(k_11_204), .air_in(c_12_1));
valve v_12_410 (.fluid_in(k_12_410), .fluid_out(k_11_205), .air_in(c_12_0));
valve v_12_411 (.fluid_in(k_12_411), .fluid_out(k_11_205), .air_in(c_12_1));
valve v_12_412 (.fluid_in(k_12_412), .fluid_out(k_11_206), .air_in(c_12_0));
valve v_12_413 (.fluid_in(k_12_413), .fluid_out(k_11_206), .air_in(c_12_1));
valve v_12_414 (.fluid_in(k_12_414), .fluid_out(k_11_207), .air_in(c_12_0));
valve v_12_415 (.fluid_in(k_12_415), .fluid_out(k_11_207), .air_in(c_12_1));
valve v_12_416 (.fluid_in(k_12_416), .fluid_out(k_11_208), .air_in(c_12_0));
valve v_12_417 (.fluid_in(k_12_417), .fluid_out(k_11_208), .air_in(c_12_1));
valve v_12_418 (.fluid_in(k_12_418), .fluid_out(k_11_209), .air_in(c_12_0));
valve v_12_419 (.fluid_in(k_12_419), .fluid_out(k_11_209), .air_in(c_12_1));
valve v_12_420 (.fluid_in(k_12_420), .fluid_out(k_11_210), .air_in(c_12_0));
valve v_12_421 (.fluid_in(k_12_421), .fluid_out(k_11_210), .air_in(c_12_1));
valve v_12_422 (.fluid_in(k_12_422), .fluid_out(k_11_211), .air_in(c_12_0));
valve v_12_423 (.fluid_in(k_12_423), .fluid_out(k_11_211), .air_in(c_12_1));
valve v_12_424 (.fluid_in(k_12_424), .fluid_out(k_11_212), .air_in(c_12_0));
valve v_12_425 (.fluid_in(k_12_425), .fluid_out(k_11_212), .air_in(c_12_1));
valve v_12_426 (.fluid_in(k_12_426), .fluid_out(k_11_213), .air_in(c_12_0));
valve v_12_427 (.fluid_in(k_12_427), .fluid_out(k_11_213), .air_in(c_12_1));
valve v_12_428 (.fluid_in(k_12_428), .fluid_out(k_11_214), .air_in(c_12_0));
valve v_12_429 (.fluid_in(k_12_429), .fluid_out(k_11_214), .air_in(c_12_1));
valve v_12_430 (.fluid_in(k_12_430), .fluid_out(k_11_215), .air_in(c_12_0));
valve v_12_431 (.fluid_in(k_12_431), .fluid_out(k_11_215), .air_in(c_12_1));
valve v_12_432 (.fluid_in(k_12_432), .fluid_out(k_11_216), .air_in(c_12_0));
valve v_12_433 (.fluid_in(k_12_433), .fluid_out(k_11_216), .air_in(c_12_1));
valve v_12_434 (.fluid_in(k_12_434), .fluid_out(k_11_217), .air_in(c_12_0));
valve v_12_435 (.fluid_in(k_12_435), .fluid_out(k_11_217), .air_in(c_12_1));
valve v_12_436 (.fluid_in(k_12_436), .fluid_out(k_11_218), .air_in(c_12_0));
valve v_12_437 (.fluid_in(k_12_437), .fluid_out(k_11_218), .air_in(c_12_1));
valve v_12_438 (.fluid_in(k_12_438), .fluid_out(k_11_219), .air_in(c_12_0));
valve v_12_439 (.fluid_in(k_12_439), .fluid_out(k_11_219), .air_in(c_12_1));
valve v_12_440 (.fluid_in(k_12_440), .fluid_out(k_11_220), .air_in(c_12_0));
valve v_12_441 (.fluid_in(k_12_441), .fluid_out(k_11_220), .air_in(c_12_1));
valve v_12_442 (.fluid_in(k_12_442), .fluid_out(k_11_221), .air_in(c_12_0));
valve v_12_443 (.fluid_in(k_12_443), .fluid_out(k_11_221), .air_in(c_12_1));
valve v_12_444 (.fluid_in(k_12_444), .fluid_out(k_11_222), .air_in(c_12_0));
valve v_12_445 (.fluid_in(k_12_445), .fluid_out(k_11_222), .air_in(c_12_1));
valve v_12_446 (.fluid_in(k_12_446), .fluid_out(k_11_223), .air_in(c_12_0));
valve v_12_447 (.fluid_in(k_12_447), .fluid_out(k_11_223), .air_in(c_12_1));
valve v_12_448 (.fluid_in(k_12_448), .fluid_out(k_11_224), .air_in(c_12_0));
valve v_12_449 (.fluid_in(k_12_449), .fluid_out(k_11_224), .air_in(c_12_1));
valve v_12_450 (.fluid_in(k_12_450), .fluid_out(k_11_225), .air_in(c_12_0));
valve v_12_451 (.fluid_in(k_12_451), .fluid_out(k_11_225), .air_in(c_12_1));
valve v_12_452 (.fluid_in(k_12_452), .fluid_out(k_11_226), .air_in(c_12_0));
valve v_12_453 (.fluid_in(k_12_453), .fluid_out(k_11_226), .air_in(c_12_1));
valve v_12_454 (.fluid_in(k_12_454), .fluid_out(k_11_227), .air_in(c_12_0));
valve v_12_455 (.fluid_in(k_12_455), .fluid_out(k_11_227), .air_in(c_12_1));
valve v_12_456 (.fluid_in(k_12_456), .fluid_out(k_11_228), .air_in(c_12_0));
valve v_12_457 (.fluid_in(k_12_457), .fluid_out(k_11_228), .air_in(c_12_1));
valve v_12_458 (.fluid_in(k_12_458), .fluid_out(k_11_229), .air_in(c_12_0));
valve v_12_459 (.fluid_in(k_12_459), .fluid_out(k_11_229), .air_in(c_12_1));
valve v_12_460 (.fluid_in(k_12_460), .fluid_out(k_11_230), .air_in(c_12_0));
valve v_12_461 (.fluid_in(k_12_461), .fluid_out(k_11_230), .air_in(c_12_1));
valve v_12_462 (.fluid_in(k_12_462), .fluid_out(k_11_231), .air_in(c_12_0));
valve v_12_463 (.fluid_in(k_12_463), .fluid_out(k_11_231), .air_in(c_12_1));
valve v_12_464 (.fluid_in(k_12_464), .fluid_out(k_11_232), .air_in(c_12_0));
valve v_12_465 (.fluid_in(k_12_465), .fluid_out(k_11_232), .air_in(c_12_1));
valve v_12_466 (.fluid_in(k_12_466), .fluid_out(k_11_233), .air_in(c_12_0));
valve v_12_467 (.fluid_in(k_12_467), .fluid_out(k_11_233), .air_in(c_12_1));
valve v_12_468 (.fluid_in(k_12_468), .fluid_out(k_11_234), .air_in(c_12_0));
valve v_12_469 (.fluid_in(k_12_469), .fluid_out(k_11_234), .air_in(c_12_1));
valve v_12_470 (.fluid_in(k_12_470), .fluid_out(k_11_235), .air_in(c_12_0));
valve v_12_471 (.fluid_in(k_12_471), .fluid_out(k_11_235), .air_in(c_12_1));
valve v_12_472 (.fluid_in(k_12_472), .fluid_out(k_11_236), .air_in(c_12_0));
valve v_12_473 (.fluid_in(k_12_473), .fluid_out(k_11_236), .air_in(c_12_1));
valve v_12_474 (.fluid_in(k_12_474), .fluid_out(k_11_237), .air_in(c_12_0));
valve v_12_475 (.fluid_in(k_12_475), .fluid_out(k_11_237), .air_in(c_12_1));
valve v_12_476 (.fluid_in(k_12_476), .fluid_out(k_11_238), .air_in(c_12_0));
valve v_12_477 (.fluid_in(k_12_477), .fluid_out(k_11_238), .air_in(c_12_1));
valve v_12_478 (.fluid_in(k_12_478), .fluid_out(k_11_239), .air_in(c_12_0));
valve v_12_479 (.fluid_in(k_12_479), .fluid_out(k_11_239), .air_in(c_12_1));
valve v_12_480 (.fluid_in(k_12_480), .fluid_out(k_11_240), .air_in(c_12_0));
valve v_12_481 (.fluid_in(k_12_481), .fluid_out(k_11_240), .air_in(c_12_1));
valve v_12_482 (.fluid_in(k_12_482), .fluid_out(k_11_241), .air_in(c_12_0));
valve v_12_483 (.fluid_in(k_12_483), .fluid_out(k_11_241), .air_in(c_12_1));
valve v_12_484 (.fluid_in(k_12_484), .fluid_out(k_11_242), .air_in(c_12_0));
valve v_12_485 (.fluid_in(k_12_485), .fluid_out(k_11_242), .air_in(c_12_1));
valve v_12_486 (.fluid_in(k_12_486), .fluid_out(k_11_243), .air_in(c_12_0));
valve v_12_487 (.fluid_in(k_12_487), .fluid_out(k_11_243), .air_in(c_12_1));
valve v_12_488 (.fluid_in(k_12_488), .fluid_out(k_11_244), .air_in(c_12_0));
valve v_12_489 (.fluid_in(k_12_489), .fluid_out(k_11_244), .air_in(c_12_1));
valve v_12_490 (.fluid_in(k_12_490), .fluid_out(k_11_245), .air_in(c_12_0));
valve v_12_491 (.fluid_in(k_12_491), .fluid_out(k_11_245), .air_in(c_12_1));
valve v_12_492 (.fluid_in(k_12_492), .fluid_out(k_11_246), .air_in(c_12_0));
valve v_12_493 (.fluid_in(k_12_493), .fluid_out(k_11_246), .air_in(c_12_1));
valve v_12_494 (.fluid_in(k_12_494), .fluid_out(k_11_247), .air_in(c_12_0));
valve v_12_495 (.fluid_in(k_12_495), .fluid_out(k_11_247), .air_in(c_12_1));
valve v_12_496 (.fluid_in(k_12_496), .fluid_out(k_11_248), .air_in(c_12_0));
valve v_12_497 (.fluid_in(k_12_497), .fluid_out(k_11_248), .air_in(c_12_1));
valve v_12_498 (.fluid_in(k_12_498), .fluid_out(k_11_249), .air_in(c_12_0));
valve v_12_499 (.fluid_in(k_12_499), .fluid_out(k_11_249), .air_in(c_12_1));
valve v_12_500 (.fluid_in(k_12_500), .fluid_out(k_11_250), .air_in(c_12_0));
valve v_12_501 (.fluid_in(k_12_501), .fluid_out(k_11_250), .air_in(c_12_1));
valve v_12_502 (.fluid_in(k_12_502), .fluid_out(k_11_251), .air_in(c_12_0));
valve v_12_503 (.fluid_in(k_12_503), .fluid_out(k_11_251), .air_in(c_12_1));
valve v_12_504 (.fluid_in(k_12_504), .fluid_out(k_11_252), .air_in(c_12_0));
valve v_12_505 (.fluid_in(k_12_505), .fluid_out(k_11_252), .air_in(c_12_1));
valve v_12_506 (.fluid_in(k_12_506), .fluid_out(k_11_253), .air_in(c_12_0));
valve v_12_507 (.fluid_in(k_12_507), .fluid_out(k_11_253), .air_in(c_12_1));
valve v_12_508 (.fluid_in(k_12_508), .fluid_out(k_11_254), .air_in(c_12_0));
valve v_12_509 (.fluid_in(k_12_509), .fluid_out(k_11_254), .air_in(c_12_1));
valve v_12_510 (.fluid_in(k_12_510), .fluid_out(k_11_255), .air_in(c_12_0));
valve v_12_511 (.fluid_in(k_12_511), .fluid_out(k_11_255), .air_in(c_12_1));
valve v_12_512 (.fluid_in(k_12_512), .fluid_out(k_11_256), .air_in(c_12_0));
valve v_12_513 (.fluid_in(k_12_513), .fluid_out(k_11_256), .air_in(c_12_1));
valve v_12_514 (.fluid_in(k_12_514), .fluid_out(k_11_257), .air_in(c_12_0));
valve v_12_515 (.fluid_in(k_12_515), .fluid_out(k_11_257), .air_in(c_12_1));
valve v_12_516 (.fluid_in(k_12_516), .fluid_out(k_11_258), .air_in(c_12_0));
valve v_12_517 (.fluid_in(k_12_517), .fluid_out(k_11_258), .air_in(c_12_1));
valve v_12_518 (.fluid_in(k_12_518), .fluid_out(k_11_259), .air_in(c_12_0));
valve v_12_519 (.fluid_in(k_12_519), .fluid_out(k_11_259), .air_in(c_12_1));
valve v_12_520 (.fluid_in(k_12_520), .fluid_out(k_11_260), .air_in(c_12_0));
valve v_12_521 (.fluid_in(k_12_521), .fluid_out(k_11_260), .air_in(c_12_1));
valve v_12_522 (.fluid_in(k_12_522), .fluid_out(k_11_261), .air_in(c_12_0));
valve v_12_523 (.fluid_in(k_12_523), .fluid_out(k_11_261), .air_in(c_12_1));
valve v_12_524 (.fluid_in(k_12_524), .fluid_out(k_11_262), .air_in(c_12_0));
valve v_12_525 (.fluid_in(k_12_525), .fluid_out(k_11_262), .air_in(c_12_1));
valve v_12_526 (.fluid_in(k_12_526), .fluid_out(k_11_263), .air_in(c_12_0));
valve v_12_527 (.fluid_in(k_12_527), .fluid_out(k_11_263), .air_in(c_12_1));
valve v_12_528 (.fluid_in(k_12_528), .fluid_out(k_11_264), .air_in(c_12_0));
valve v_12_529 (.fluid_in(k_12_529), .fluid_out(k_11_264), .air_in(c_12_1));
valve v_12_530 (.fluid_in(k_12_530), .fluid_out(k_11_265), .air_in(c_12_0));
valve v_12_531 (.fluid_in(k_12_531), .fluid_out(k_11_265), .air_in(c_12_1));
valve v_12_532 (.fluid_in(k_12_532), .fluid_out(k_11_266), .air_in(c_12_0));
valve v_12_533 (.fluid_in(k_12_533), .fluid_out(k_11_266), .air_in(c_12_1));
valve v_12_534 (.fluid_in(k_12_534), .fluid_out(k_11_267), .air_in(c_12_0));
valve v_12_535 (.fluid_in(k_12_535), .fluid_out(k_11_267), .air_in(c_12_1));
valve v_12_536 (.fluid_in(k_12_536), .fluid_out(k_11_268), .air_in(c_12_0));
valve v_12_537 (.fluid_in(k_12_537), .fluid_out(k_11_268), .air_in(c_12_1));
valve v_12_538 (.fluid_in(k_12_538), .fluid_out(k_11_269), .air_in(c_12_0));
valve v_12_539 (.fluid_in(k_12_539), .fluid_out(k_11_269), .air_in(c_12_1));
valve v_12_540 (.fluid_in(k_12_540), .fluid_out(k_11_270), .air_in(c_12_0));
valve v_12_541 (.fluid_in(k_12_541), .fluid_out(k_11_270), .air_in(c_12_1));
valve v_12_542 (.fluid_in(k_12_542), .fluid_out(k_11_271), .air_in(c_12_0));
valve v_12_543 (.fluid_in(k_12_543), .fluid_out(k_11_271), .air_in(c_12_1));
valve v_12_544 (.fluid_in(k_12_544), .fluid_out(k_11_272), .air_in(c_12_0));
valve v_12_545 (.fluid_in(k_12_545), .fluid_out(k_11_272), .air_in(c_12_1));
valve v_12_546 (.fluid_in(k_12_546), .fluid_out(k_11_273), .air_in(c_12_0));
valve v_12_547 (.fluid_in(k_12_547), .fluid_out(k_11_273), .air_in(c_12_1));
valve v_12_548 (.fluid_in(k_12_548), .fluid_out(k_11_274), .air_in(c_12_0));
valve v_12_549 (.fluid_in(k_12_549), .fluid_out(k_11_274), .air_in(c_12_1));
valve v_12_550 (.fluid_in(k_12_550), .fluid_out(k_11_275), .air_in(c_12_0));
valve v_12_551 (.fluid_in(k_12_551), .fluid_out(k_11_275), .air_in(c_12_1));
valve v_12_552 (.fluid_in(k_12_552), .fluid_out(k_11_276), .air_in(c_12_0));
valve v_12_553 (.fluid_in(k_12_553), .fluid_out(k_11_276), .air_in(c_12_1));
valve v_12_554 (.fluid_in(k_12_554), .fluid_out(k_11_277), .air_in(c_12_0));
valve v_12_555 (.fluid_in(k_12_555), .fluid_out(k_11_277), .air_in(c_12_1));
valve v_12_556 (.fluid_in(k_12_556), .fluid_out(k_11_278), .air_in(c_12_0));
valve v_12_557 (.fluid_in(k_12_557), .fluid_out(k_11_278), .air_in(c_12_1));
valve v_12_558 (.fluid_in(k_12_558), .fluid_out(k_11_279), .air_in(c_12_0));
valve v_12_559 (.fluid_in(k_12_559), .fluid_out(k_11_279), .air_in(c_12_1));
valve v_12_560 (.fluid_in(k_12_560), .fluid_out(k_11_280), .air_in(c_12_0));
valve v_12_561 (.fluid_in(k_12_561), .fluid_out(k_11_280), .air_in(c_12_1));
valve v_12_562 (.fluid_in(k_12_562), .fluid_out(k_11_281), .air_in(c_12_0));
valve v_12_563 (.fluid_in(k_12_563), .fluid_out(k_11_281), .air_in(c_12_1));
valve v_12_564 (.fluid_in(k_12_564), .fluid_out(k_11_282), .air_in(c_12_0));
valve v_12_565 (.fluid_in(k_12_565), .fluid_out(k_11_282), .air_in(c_12_1));
valve v_12_566 (.fluid_in(k_12_566), .fluid_out(k_11_283), .air_in(c_12_0));
valve v_12_567 (.fluid_in(k_12_567), .fluid_out(k_11_283), .air_in(c_12_1));
valve v_12_568 (.fluid_in(k_12_568), .fluid_out(k_11_284), .air_in(c_12_0));
valve v_12_569 (.fluid_in(k_12_569), .fluid_out(k_11_284), .air_in(c_12_1));
valve v_12_570 (.fluid_in(k_12_570), .fluid_out(k_11_285), .air_in(c_12_0));
valve v_12_571 (.fluid_in(k_12_571), .fluid_out(k_11_285), .air_in(c_12_1));
valve v_12_572 (.fluid_in(k_12_572), .fluid_out(k_11_286), .air_in(c_12_0));
valve v_12_573 (.fluid_in(k_12_573), .fluid_out(k_11_286), .air_in(c_12_1));
valve v_12_574 (.fluid_in(k_12_574), .fluid_out(k_11_287), .air_in(c_12_0));
valve v_12_575 (.fluid_in(k_12_575), .fluid_out(k_11_287), .air_in(c_12_1));
valve v_12_576 (.fluid_in(k_12_576), .fluid_out(k_11_288), .air_in(c_12_0));
valve v_12_577 (.fluid_in(k_12_577), .fluid_out(k_11_288), .air_in(c_12_1));
valve v_12_578 (.fluid_in(k_12_578), .fluid_out(k_11_289), .air_in(c_12_0));
valve v_12_579 (.fluid_in(k_12_579), .fluid_out(k_11_289), .air_in(c_12_1));
valve v_12_580 (.fluid_in(k_12_580), .fluid_out(k_11_290), .air_in(c_12_0));
valve v_12_581 (.fluid_in(k_12_581), .fluid_out(k_11_290), .air_in(c_12_1));
valve v_12_582 (.fluid_in(k_12_582), .fluid_out(k_11_291), .air_in(c_12_0));
valve v_12_583 (.fluid_in(k_12_583), .fluid_out(k_11_291), .air_in(c_12_1));
valve v_12_584 (.fluid_in(k_12_584), .fluid_out(k_11_292), .air_in(c_12_0));
valve v_12_585 (.fluid_in(k_12_585), .fluid_out(k_11_292), .air_in(c_12_1));
valve v_12_586 (.fluid_in(k_12_586), .fluid_out(k_11_293), .air_in(c_12_0));
valve v_12_587 (.fluid_in(k_12_587), .fluid_out(k_11_293), .air_in(c_12_1));
valve v_12_588 (.fluid_in(k_12_588), .fluid_out(k_11_294), .air_in(c_12_0));
valve v_12_589 (.fluid_in(k_12_589), .fluid_out(k_11_294), .air_in(c_12_1));
valve v_12_590 (.fluid_in(k_12_590), .fluid_out(k_11_295), .air_in(c_12_0));
valve v_12_591 (.fluid_in(k_12_591), .fluid_out(k_11_295), .air_in(c_12_1));
valve v_12_592 (.fluid_in(k_12_592), .fluid_out(k_11_296), .air_in(c_12_0));
valve v_12_593 (.fluid_in(k_12_593), .fluid_out(k_11_296), .air_in(c_12_1));
valve v_12_594 (.fluid_in(k_12_594), .fluid_out(k_11_297), .air_in(c_12_0));
valve v_12_595 (.fluid_in(k_12_595), .fluid_out(k_11_297), .air_in(c_12_1));
valve v_12_596 (.fluid_in(k_12_596), .fluid_out(k_11_298), .air_in(c_12_0));
valve v_12_597 (.fluid_in(k_12_597), .fluid_out(k_11_298), .air_in(c_12_1));
valve v_12_598 (.fluid_in(k_12_598), .fluid_out(k_11_299), .air_in(c_12_0));
valve v_12_599 (.fluid_in(k_12_599), .fluid_out(k_11_299), .air_in(c_12_1));
valve v_12_600 (.fluid_in(k_12_600), .fluid_out(k_11_300), .air_in(c_12_0));
valve v_12_601 (.fluid_in(k_12_601), .fluid_out(k_11_300), .air_in(c_12_1));
valve v_12_602 (.fluid_in(k_12_602), .fluid_out(k_11_301), .air_in(c_12_0));
valve v_12_603 (.fluid_in(k_12_603), .fluid_out(k_11_301), .air_in(c_12_1));
valve v_12_604 (.fluid_in(k_12_604), .fluid_out(k_11_302), .air_in(c_12_0));
valve v_12_605 (.fluid_in(k_12_605), .fluid_out(k_11_302), .air_in(c_12_1));
valve v_12_606 (.fluid_in(k_12_606), .fluid_out(k_11_303), .air_in(c_12_0));
valve v_12_607 (.fluid_in(k_12_607), .fluid_out(k_11_303), .air_in(c_12_1));
valve v_12_608 (.fluid_in(k_12_608), .fluid_out(k_11_304), .air_in(c_12_0));
valve v_12_609 (.fluid_in(k_12_609), .fluid_out(k_11_304), .air_in(c_12_1));
valve v_12_610 (.fluid_in(k_12_610), .fluid_out(k_11_305), .air_in(c_12_0));
valve v_12_611 (.fluid_in(k_12_611), .fluid_out(k_11_305), .air_in(c_12_1));
valve v_12_612 (.fluid_in(k_12_612), .fluid_out(k_11_306), .air_in(c_12_0));
valve v_12_613 (.fluid_in(k_12_613), .fluid_out(k_11_306), .air_in(c_12_1));
valve v_12_614 (.fluid_in(k_12_614), .fluid_out(k_11_307), .air_in(c_12_0));
valve v_12_615 (.fluid_in(k_12_615), .fluid_out(k_11_307), .air_in(c_12_1));
valve v_12_616 (.fluid_in(k_12_616), .fluid_out(k_11_308), .air_in(c_12_0));
valve v_12_617 (.fluid_in(k_12_617), .fluid_out(k_11_308), .air_in(c_12_1));
valve v_12_618 (.fluid_in(k_12_618), .fluid_out(k_11_309), .air_in(c_12_0));
valve v_12_619 (.fluid_in(k_12_619), .fluid_out(k_11_309), .air_in(c_12_1));
valve v_12_620 (.fluid_in(k_12_620), .fluid_out(k_11_310), .air_in(c_12_0));
valve v_12_621 (.fluid_in(k_12_621), .fluid_out(k_11_310), .air_in(c_12_1));
valve v_12_622 (.fluid_in(k_12_622), .fluid_out(k_11_311), .air_in(c_12_0));
valve v_12_623 (.fluid_in(k_12_623), .fluid_out(k_11_311), .air_in(c_12_1));
valve v_12_624 (.fluid_in(k_12_624), .fluid_out(k_11_312), .air_in(c_12_0));
valve v_12_625 (.fluid_in(k_12_625), .fluid_out(k_11_312), .air_in(c_12_1));
valve v_12_626 (.fluid_in(k_12_626), .fluid_out(k_11_313), .air_in(c_12_0));
valve v_12_627 (.fluid_in(k_12_627), .fluid_out(k_11_313), .air_in(c_12_1));
valve v_12_628 (.fluid_in(k_12_628), .fluid_out(k_11_314), .air_in(c_12_0));
valve v_12_629 (.fluid_in(k_12_629), .fluid_out(k_11_314), .air_in(c_12_1));
valve v_12_630 (.fluid_in(k_12_630), .fluid_out(k_11_315), .air_in(c_12_0));
valve v_12_631 (.fluid_in(k_12_631), .fluid_out(k_11_315), .air_in(c_12_1));
valve v_12_632 (.fluid_in(k_12_632), .fluid_out(k_11_316), .air_in(c_12_0));
valve v_12_633 (.fluid_in(k_12_633), .fluid_out(k_11_316), .air_in(c_12_1));
valve v_12_634 (.fluid_in(k_12_634), .fluid_out(k_11_317), .air_in(c_12_0));
valve v_12_635 (.fluid_in(k_12_635), .fluid_out(k_11_317), .air_in(c_12_1));
valve v_12_636 (.fluid_in(k_12_636), .fluid_out(k_11_318), .air_in(c_12_0));
valve v_12_637 (.fluid_in(k_12_637), .fluid_out(k_11_318), .air_in(c_12_1));
valve v_12_638 (.fluid_in(k_12_638), .fluid_out(k_11_319), .air_in(c_12_0));
valve v_12_639 (.fluid_in(k_12_639), .fluid_out(k_11_319), .air_in(c_12_1));
valve v_12_640 (.fluid_in(k_12_640), .fluid_out(k_11_320), .air_in(c_12_0));
valve v_12_641 (.fluid_in(k_12_641), .fluid_out(k_11_320), .air_in(c_12_1));
valve v_12_642 (.fluid_in(k_12_642), .fluid_out(k_11_321), .air_in(c_12_0));
valve v_12_643 (.fluid_in(k_12_643), .fluid_out(k_11_321), .air_in(c_12_1));
valve v_12_644 (.fluid_in(k_12_644), .fluid_out(k_11_322), .air_in(c_12_0));
valve v_12_645 (.fluid_in(k_12_645), .fluid_out(k_11_322), .air_in(c_12_1));
valve v_12_646 (.fluid_in(k_12_646), .fluid_out(k_11_323), .air_in(c_12_0));
valve v_12_647 (.fluid_in(k_12_647), .fluid_out(k_11_323), .air_in(c_12_1));
valve v_12_648 (.fluid_in(k_12_648), .fluid_out(k_11_324), .air_in(c_12_0));
valve v_12_649 (.fluid_in(k_12_649), .fluid_out(k_11_324), .air_in(c_12_1));
valve v_12_650 (.fluid_in(k_12_650), .fluid_out(k_11_325), .air_in(c_12_0));
valve v_12_651 (.fluid_in(k_12_651), .fluid_out(k_11_325), .air_in(c_12_1));
valve v_12_652 (.fluid_in(k_12_652), .fluid_out(k_11_326), .air_in(c_12_0));
valve v_12_653 (.fluid_in(k_12_653), .fluid_out(k_11_326), .air_in(c_12_1));
valve v_12_654 (.fluid_in(k_12_654), .fluid_out(k_11_327), .air_in(c_12_0));
valve v_12_655 (.fluid_in(k_12_655), .fluid_out(k_11_327), .air_in(c_12_1));
valve v_12_656 (.fluid_in(k_12_656), .fluid_out(k_11_328), .air_in(c_12_0));
valve v_12_657 (.fluid_in(k_12_657), .fluid_out(k_11_328), .air_in(c_12_1));
valve v_12_658 (.fluid_in(k_12_658), .fluid_out(k_11_329), .air_in(c_12_0));
valve v_12_659 (.fluid_in(k_12_659), .fluid_out(k_11_329), .air_in(c_12_1));
valve v_12_660 (.fluid_in(k_12_660), .fluid_out(k_11_330), .air_in(c_12_0));
valve v_12_661 (.fluid_in(k_12_661), .fluid_out(k_11_330), .air_in(c_12_1));
valve v_12_662 (.fluid_in(k_12_662), .fluid_out(k_11_331), .air_in(c_12_0));
valve v_12_663 (.fluid_in(k_12_663), .fluid_out(k_11_331), .air_in(c_12_1));
valve v_12_664 (.fluid_in(k_12_664), .fluid_out(k_11_332), .air_in(c_12_0));
valve v_12_665 (.fluid_in(k_12_665), .fluid_out(k_11_332), .air_in(c_12_1));
valve v_12_666 (.fluid_in(k_12_666), .fluid_out(k_11_333), .air_in(c_12_0));
valve v_12_667 (.fluid_in(k_12_667), .fluid_out(k_11_333), .air_in(c_12_1));
valve v_12_668 (.fluid_in(k_12_668), .fluid_out(k_11_334), .air_in(c_12_0));
valve v_12_669 (.fluid_in(k_12_669), .fluid_out(k_11_334), .air_in(c_12_1));
valve v_12_670 (.fluid_in(k_12_670), .fluid_out(k_11_335), .air_in(c_12_0));
valve v_12_671 (.fluid_in(k_12_671), .fluid_out(k_11_335), .air_in(c_12_1));
valve v_12_672 (.fluid_in(k_12_672), .fluid_out(k_11_336), .air_in(c_12_0));
valve v_12_673 (.fluid_in(k_12_673), .fluid_out(k_11_336), .air_in(c_12_1));
valve v_12_674 (.fluid_in(k_12_674), .fluid_out(k_11_337), .air_in(c_12_0));
valve v_12_675 (.fluid_in(k_12_675), .fluid_out(k_11_337), .air_in(c_12_1));
valve v_12_676 (.fluid_in(k_12_676), .fluid_out(k_11_338), .air_in(c_12_0));
valve v_12_677 (.fluid_in(k_12_677), .fluid_out(k_11_338), .air_in(c_12_1));
valve v_12_678 (.fluid_in(k_12_678), .fluid_out(k_11_339), .air_in(c_12_0));
valve v_12_679 (.fluid_in(k_12_679), .fluid_out(k_11_339), .air_in(c_12_1));
valve v_12_680 (.fluid_in(k_12_680), .fluid_out(k_11_340), .air_in(c_12_0));
valve v_12_681 (.fluid_in(k_12_681), .fluid_out(k_11_340), .air_in(c_12_1));
valve v_12_682 (.fluid_in(k_12_682), .fluid_out(k_11_341), .air_in(c_12_0));
valve v_12_683 (.fluid_in(k_12_683), .fluid_out(k_11_341), .air_in(c_12_1));
valve v_12_684 (.fluid_in(k_12_684), .fluid_out(k_11_342), .air_in(c_12_0));
valve v_12_685 (.fluid_in(k_12_685), .fluid_out(k_11_342), .air_in(c_12_1));
valve v_12_686 (.fluid_in(k_12_686), .fluid_out(k_11_343), .air_in(c_12_0));
valve v_12_687 (.fluid_in(k_12_687), .fluid_out(k_11_343), .air_in(c_12_1));
valve v_12_688 (.fluid_in(k_12_688), .fluid_out(k_11_344), .air_in(c_12_0));
valve v_12_689 (.fluid_in(k_12_689), .fluid_out(k_11_344), .air_in(c_12_1));
valve v_12_690 (.fluid_in(k_12_690), .fluid_out(k_11_345), .air_in(c_12_0));
valve v_12_691 (.fluid_in(k_12_691), .fluid_out(k_11_345), .air_in(c_12_1));
valve v_12_692 (.fluid_in(k_12_692), .fluid_out(k_11_346), .air_in(c_12_0));
valve v_12_693 (.fluid_in(k_12_693), .fluid_out(k_11_346), .air_in(c_12_1));
valve v_12_694 (.fluid_in(k_12_694), .fluid_out(k_11_347), .air_in(c_12_0));
valve v_12_695 (.fluid_in(k_12_695), .fluid_out(k_11_347), .air_in(c_12_1));
valve v_12_696 (.fluid_in(k_12_696), .fluid_out(k_11_348), .air_in(c_12_0));
valve v_12_697 (.fluid_in(k_12_697), .fluid_out(k_11_348), .air_in(c_12_1));
valve v_12_698 (.fluid_in(k_12_698), .fluid_out(k_11_349), .air_in(c_12_0));
valve v_12_699 (.fluid_in(k_12_699), .fluid_out(k_11_349), .air_in(c_12_1));
valve v_12_700 (.fluid_in(k_12_700), .fluid_out(k_11_350), .air_in(c_12_0));
valve v_12_701 (.fluid_in(k_12_701), .fluid_out(k_11_350), .air_in(c_12_1));
valve v_12_702 (.fluid_in(k_12_702), .fluid_out(k_11_351), .air_in(c_12_0));
valve v_12_703 (.fluid_in(k_12_703), .fluid_out(k_11_351), .air_in(c_12_1));
valve v_12_704 (.fluid_in(k_12_704), .fluid_out(k_11_352), .air_in(c_12_0));
valve v_12_705 (.fluid_in(k_12_705), .fluid_out(k_11_352), .air_in(c_12_1));
valve v_12_706 (.fluid_in(k_12_706), .fluid_out(k_11_353), .air_in(c_12_0));
valve v_12_707 (.fluid_in(k_12_707), .fluid_out(k_11_353), .air_in(c_12_1));
valve v_12_708 (.fluid_in(k_12_708), .fluid_out(k_11_354), .air_in(c_12_0));
valve v_12_709 (.fluid_in(k_12_709), .fluid_out(k_11_354), .air_in(c_12_1));
valve v_12_710 (.fluid_in(k_12_710), .fluid_out(k_11_355), .air_in(c_12_0));
valve v_12_711 (.fluid_in(k_12_711), .fluid_out(k_11_355), .air_in(c_12_1));
valve v_12_712 (.fluid_in(k_12_712), .fluid_out(k_11_356), .air_in(c_12_0));
valve v_12_713 (.fluid_in(k_12_713), .fluid_out(k_11_356), .air_in(c_12_1));
valve v_12_714 (.fluid_in(k_12_714), .fluid_out(k_11_357), .air_in(c_12_0));
valve v_12_715 (.fluid_in(k_12_715), .fluid_out(k_11_357), .air_in(c_12_1));
valve v_12_716 (.fluid_in(k_12_716), .fluid_out(k_11_358), .air_in(c_12_0));
valve v_12_717 (.fluid_in(k_12_717), .fluid_out(k_11_358), .air_in(c_12_1));
valve v_12_718 (.fluid_in(k_12_718), .fluid_out(k_11_359), .air_in(c_12_0));
valve v_12_719 (.fluid_in(k_12_719), .fluid_out(k_11_359), .air_in(c_12_1));
valve v_12_720 (.fluid_in(k_12_720), .fluid_out(k_11_360), .air_in(c_12_0));
valve v_12_721 (.fluid_in(k_12_721), .fluid_out(k_11_360), .air_in(c_12_1));
valve v_12_722 (.fluid_in(k_12_722), .fluid_out(k_11_361), .air_in(c_12_0));
valve v_12_723 (.fluid_in(k_12_723), .fluid_out(k_11_361), .air_in(c_12_1));
valve v_12_724 (.fluid_in(k_12_724), .fluid_out(k_11_362), .air_in(c_12_0));
valve v_12_725 (.fluid_in(k_12_725), .fluid_out(k_11_362), .air_in(c_12_1));
valve v_12_726 (.fluid_in(k_12_726), .fluid_out(k_11_363), .air_in(c_12_0));
valve v_12_727 (.fluid_in(k_12_727), .fluid_out(k_11_363), .air_in(c_12_1));
valve v_12_728 (.fluid_in(k_12_728), .fluid_out(k_11_364), .air_in(c_12_0));
valve v_12_729 (.fluid_in(k_12_729), .fluid_out(k_11_364), .air_in(c_12_1));
valve v_12_730 (.fluid_in(k_12_730), .fluid_out(k_11_365), .air_in(c_12_0));
valve v_12_731 (.fluid_in(k_12_731), .fluid_out(k_11_365), .air_in(c_12_1));
valve v_12_732 (.fluid_in(k_12_732), .fluid_out(k_11_366), .air_in(c_12_0));
valve v_12_733 (.fluid_in(k_12_733), .fluid_out(k_11_366), .air_in(c_12_1));
valve v_12_734 (.fluid_in(k_12_734), .fluid_out(k_11_367), .air_in(c_12_0));
valve v_12_735 (.fluid_in(k_12_735), .fluid_out(k_11_367), .air_in(c_12_1));
valve v_12_736 (.fluid_in(k_12_736), .fluid_out(k_11_368), .air_in(c_12_0));
valve v_12_737 (.fluid_in(k_12_737), .fluid_out(k_11_368), .air_in(c_12_1));
valve v_12_738 (.fluid_in(k_12_738), .fluid_out(k_11_369), .air_in(c_12_0));
valve v_12_739 (.fluid_in(k_12_739), .fluid_out(k_11_369), .air_in(c_12_1));
valve v_12_740 (.fluid_in(k_12_740), .fluid_out(k_11_370), .air_in(c_12_0));
valve v_12_741 (.fluid_in(k_12_741), .fluid_out(k_11_370), .air_in(c_12_1));
valve v_12_742 (.fluid_in(k_12_742), .fluid_out(k_11_371), .air_in(c_12_0));
valve v_12_743 (.fluid_in(k_12_743), .fluid_out(k_11_371), .air_in(c_12_1));
valve v_12_744 (.fluid_in(k_12_744), .fluid_out(k_11_372), .air_in(c_12_0));
valve v_12_745 (.fluid_in(k_12_745), .fluid_out(k_11_372), .air_in(c_12_1));
valve v_12_746 (.fluid_in(k_12_746), .fluid_out(k_11_373), .air_in(c_12_0));
valve v_12_747 (.fluid_in(k_12_747), .fluid_out(k_11_373), .air_in(c_12_1));
valve v_12_748 (.fluid_in(k_12_748), .fluid_out(k_11_374), .air_in(c_12_0));
valve v_12_749 (.fluid_in(k_12_749), .fluid_out(k_11_374), .air_in(c_12_1));
valve v_12_750 (.fluid_in(k_12_750), .fluid_out(k_11_375), .air_in(c_12_0));
valve v_12_751 (.fluid_in(k_12_751), .fluid_out(k_11_375), .air_in(c_12_1));
valve v_12_752 (.fluid_in(k_12_752), .fluid_out(k_11_376), .air_in(c_12_0));
valve v_12_753 (.fluid_in(k_12_753), .fluid_out(k_11_376), .air_in(c_12_1));
valve v_12_754 (.fluid_in(k_12_754), .fluid_out(k_11_377), .air_in(c_12_0));
valve v_12_755 (.fluid_in(k_12_755), .fluid_out(k_11_377), .air_in(c_12_1));
valve v_12_756 (.fluid_in(k_12_756), .fluid_out(k_11_378), .air_in(c_12_0));
valve v_12_757 (.fluid_in(k_12_757), .fluid_out(k_11_378), .air_in(c_12_1));
valve v_12_758 (.fluid_in(k_12_758), .fluid_out(k_11_379), .air_in(c_12_0));
valve v_12_759 (.fluid_in(k_12_759), .fluid_out(k_11_379), .air_in(c_12_1));
valve v_12_760 (.fluid_in(k_12_760), .fluid_out(k_11_380), .air_in(c_12_0));
valve v_12_761 (.fluid_in(k_12_761), .fluid_out(k_11_380), .air_in(c_12_1));
valve v_12_762 (.fluid_in(k_12_762), .fluid_out(k_11_381), .air_in(c_12_0));
valve v_12_763 (.fluid_in(k_12_763), .fluid_out(k_11_381), .air_in(c_12_1));
valve v_12_764 (.fluid_in(k_12_764), .fluid_out(k_11_382), .air_in(c_12_0));
valve v_12_765 (.fluid_in(k_12_765), .fluid_out(k_11_382), .air_in(c_12_1));
valve v_12_766 (.fluid_in(k_12_766), .fluid_out(k_11_383), .air_in(c_12_0));
valve v_12_767 (.fluid_in(k_12_767), .fluid_out(k_11_383), .air_in(c_12_1));
valve v_12_768 (.fluid_in(k_12_768), .fluid_out(k_11_384), .air_in(c_12_0));
valve v_12_769 (.fluid_in(k_12_769), .fluid_out(k_11_384), .air_in(c_12_1));
valve v_12_770 (.fluid_in(k_12_770), .fluid_out(k_11_385), .air_in(c_12_0));
valve v_12_771 (.fluid_in(k_12_771), .fluid_out(k_11_385), .air_in(c_12_1));
valve v_12_772 (.fluid_in(k_12_772), .fluid_out(k_11_386), .air_in(c_12_0));
valve v_12_773 (.fluid_in(k_12_773), .fluid_out(k_11_386), .air_in(c_12_1));
valve v_12_774 (.fluid_in(k_12_774), .fluid_out(k_11_387), .air_in(c_12_0));
valve v_12_775 (.fluid_in(k_12_775), .fluid_out(k_11_387), .air_in(c_12_1));
valve v_12_776 (.fluid_in(k_12_776), .fluid_out(k_11_388), .air_in(c_12_0));
valve v_12_777 (.fluid_in(k_12_777), .fluid_out(k_11_388), .air_in(c_12_1));
valve v_12_778 (.fluid_in(k_12_778), .fluid_out(k_11_389), .air_in(c_12_0));
valve v_12_779 (.fluid_in(k_12_779), .fluid_out(k_11_389), .air_in(c_12_1));
valve v_12_780 (.fluid_in(k_12_780), .fluid_out(k_11_390), .air_in(c_12_0));
valve v_12_781 (.fluid_in(k_12_781), .fluid_out(k_11_390), .air_in(c_12_1));
valve v_12_782 (.fluid_in(k_12_782), .fluid_out(k_11_391), .air_in(c_12_0));
valve v_12_783 (.fluid_in(k_12_783), .fluid_out(k_11_391), .air_in(c_12_1));
valve v_12_784 (.fluid_in(k_12_784), .fluid_out(k_11_392), .air_in(c_12_0));
valve v_12_785 (.fluid_in(k_12_785), .fluid_out(k_11_392), .air_in(c_12_1));
valve v_12_786 (.fluid_in(k_12_786), .fluid_out(k_11_393), .air_in(c_12_0));
valve v_12_787 (.fluid_in(k_12_787), .fluid_out(k_11_393), .air_in(c_12_1));
valve v_12_788 (.fluid_in(k_12_788), .fluid_out(k_11_394), .air_in(c_12_0));
valve v_12_789 (.fluid_in(k_12_789), .fluid_out(k_11_394), .air_in(c_12_1));
valve v_12_790 (.fluid_in(k_12_790), .fluid_out(k_11_395), .air_in(c_12_0));
valve v_12_791 (.fluid_in(k_12_791), .fluid_out(k_11_395), .air_in(c_12_1));
valve v_12_792 (.fluid_in(k_12_792), .fluid_out(k_11_396), .air_in(c_12_0));
valve v_12_793 (.fluid_in(k_12_793), .fluid_out(k_11_396), .air_in(c_12_1));
valve v_12_794 (.fluid_in(k_12_794), .fluid_out(k_11_397), .air_in(c_12_0));
valve v_12_795 (.fluid_in(k_12_795), .fluid_out(k_11_397), .air_in(c_12_1));
valve v_12_796 (.fluid_in(k_12_796), .fluid_out(k_11_398), .air_in(c_12_0));
valve v_12_797 (.fluid_in(k_12_797), .fluid_out(k_11_398), .air_in(c_12_1));
valve v_12_798 (.fluid_in(k_12_798), .fluid_out(k_11_399), .air_in(c_12_0));
valve v_12_799 (.fluid_in(k_12_799), .fluid_out(k_11_399), .air_in(c_12_1));
valve v_12_800 (.fluid_in(k_12_800), .fluid_out(k_11_400), .air_in(c_12_0));
valve v_12_801 (.fluid_in(k_12_801), .fluid_out(k_11_400), .air_in(c_12_1));
valve v_12_802 (.fluid_in(k_12_802), .fluid_out(k_11_401), .air_in(c_12_0));
valve v_12_803 (.fluid_in(k_12_803), .fluid_out(k_11_401), .air_in(c_12_1));
valve v_12_804 (.fluid_in(k_12_804), .fluid_out(k_11_402), .air_in(c_12_0));
valve v_12_805 (.fluid_in(k_12_805), .fluid_out(k_11_402), .air_in(c_12_1));
valve v_12_806 (.fluid_in(k_12_806), .fluid_out(k_11_403), .air_in(c_12_0));
valve v_12_807 (.fluid_in(k_12_807), .fluid_out(k_11_403), .air_in(c_12_1));
valve v_12_808 (.fluid_in(k_12_808), .fluid_out(k_11_404), .air_in(c_12_0));
valve v_12_809 (.fluid_in(k_12_809), .fluid_out(k_11_404), .air_in(c_12_1));
valve v_12_810 (.fluid_in(k_12_810), .fluid_out(k_11_405), .air_in(c_12_0));
valve v_12_811 (.fluid_in(k_12_811), .fluid_out(k_11_405), .air_in(c_12_1));
valve v_12_812 (.fluid_in(k_12_812), .fluid_out(k_11_406), .air_in(c_12_0));
valve v_12_813 (.fluid_in(k_12_813), .fluid_out(k_11_406), .air_in(c_12_1));
valve v_12_814 (.fluid_in(k_12_814), .fluid_out(k_11_407), .air_in(c_12_0));
valve v_12_815 (.fluid_in(k_12_815), .fluid_out(k_11_407), .air_in(c_12_1));
valve v_12_816 (.fluid_in(k_12_816), .fluid_out(k_11_408), .air_in(c_12_0));
valve v_12_817 (.fluid_in(k_12_817), .fluid_out(k_11_408), .air_in(c_12_1));
valve v_12_818 (.fluid_in(k_12_818), .fluid_out(k_11_409), .air_in(c_12_0));
valve v_12_819 (.fluid_in(k_12_819), .fluid_out(k_11_409), .air_in(c_12_1));
valve v_12_820 (.fluid_in(k_12_820), .fluid_out(k_11_410), .air_in(c_12_0));
valve v_12_821 (.fluid_in(k_12_821), .fluid_out(k_11_410), .air_in(c_12_1));
valve v_12_822 (.fluid_in(k_12_822), .fluid_out(k_11_411), .air_in(c_12_0));
valve v_12_823 (.fluid_in(k_12_823), .fluid_out(k_11_411), .air_in(c_12_1));
valve v_12_824 (.fluid_in(k_12_824), .fluid_out(k_11_412), .air_in(c_12_0));
valve v_12_825 (.fluid_in(k_12_825), .fluid_out(k_11_412), .air_in(c_12_1));
valve v_12_826 (.fluid_in(k_12_826), .fluid_out(k_11_413), .air_in(c_12_0));
valve v_12_827 (.fluid_in(k_12_827), .fluid_out(k_11_413), .air_in(c_12_1));
valve v_12_828 (.fluid_in(k_12_828), .fluid_out(k_11_414), .air_in(c_12_0));
valve v_12_829 (.fluid_in(k_12_829), .fluid_out(k_11_414), .air_in(c_12_1));
valve v_12_830 (.fluid_in(k_12_830), .fluid_out(k_11_415), .air_in(c_12_0));
valve v_12_831 (.fluid_in(k_12_831), .fluid_out(k_11_415), .air_in(c_12_1));
valve v_12_832 (.fluid_in(k_12_832), .fluid_out(k_11_416), .air_in(c_12_0));
valve v_12_833 (.fluid_in(k_12_833), .fluid_out(k_11_416), .air_in(c_12_1));
valve v_12_834 (.fluid_in(k_12_834), .fluid_out(k_11_417), .air_in(c_12_0));
valve v_12_835 (.fluid_in(k_12_835), .fluid_out(k_11_417), .air_in(c_12_1));
valve v_12_836 (.fluid_in(k_12_836), .fluid_out(k_11_418), .air_in(c_12_0));
valve v_12_837 (.fluid_in(k_12_837), .fluid_out(k_11_418), .air_in(c_12_1));
valve v_12_838 (.fluid_in(k_12_838), .fluid_out(k_11_419), .air_in(c_12_0));
valve v_12_839 (.fluid_in(k_12_839), .fluid_out(k_11_419), .air_in(c_12_1));
valve v_12_840 (.fluid_in(k_12_840), .fluid_out(k_11_420), .air_in(c_12_0));
valve v_12_841 (.fluid_in(k_12_841), .fluid_out(k_11_420), .air_in(c_12_1));
valve v_12_842 (.fluid_in(k_12_842), .fluid_out(k_11_421), .air_in(c_12_0));
valve v_12_843 (.fluid_in(k_12_843), .fluid_out(k_11_421), .air_in(c_12_1));
valve v_12_844 (.fluid_in(k_12_844), .fluid_out(k_11_422), .air_in(c_12_0));
valve v_12_845 (.fluid_in(k_12_845), .fluid_out(k_11_422), .air_in(c_12_1));
valve v_12_846 (.fluid_in(k_12_846), .fluid_out(k_11_423), .air_in(c_12_0));
valve v_12_847 (.fluid_in(k_12_847), .fluid_out(k_11_423), .air_in(c_12_1));
valve v_12_848 (.fluid_in(k_12_848), .fluid_out(k_11_424), .air_in(c_12_0));
valve v_12_849 (.fluid_in(k_12_849), .fluid_out(k_11_424), .air_in(c_12_1));
valve v_12_850 (.fluid_in(k_12_850), .fluid_out(k_11_425), .air_in(c_12_0));
valve v_12_851 (.fluid_in(k_12_851), .fluid_out(k_11_425), .air_in(c_12_1));
valve v_12_852 (.fluid_in(k_12_852), .fluid_out(k_11_426), .air_in(c_12_0));
valve v_12_853 (.fluid_in(k_12_853), .fluid_out(k_11_426), .air_in(c_12_1));
valve v_12_854 (.fluid_in(k_12_854), .fluid_out(k_11_427), .air_in(c_12_0));
valve v_12_855 (.fluid_in(k_12_855), .fluid_out(k_11_427), .air_in(c_12_1));
valve v_12_856 (.fluid_in(k_12_856), .fluid_out(k_11_428), .air_in(c_12_0));
valve v_12_857 (.fluid_in(k_12_857), .fluid_out(k_11_428), .air_in(c_12_1));
valve v_12_858 (.fluid_in(k_12_858), .fluid_out(k_11_429), .air_in(c_12_0));
valve v_12_859 (.fluid_in(k_12_859), .fluid_out(k_11_429), .air_in(c_12_1));
valve v_12_860 (.fluid_in(k_12_860), .fluid_out(k_11_430), .air_in(c_12_0));
valve v_12_861 (.fluid_in(k_12_861), .fluid_out(k_11_430), .air_in(c_12_1));
valve v_12_862 (.fluid_in(k_12_862), .fluid_out(k_11_431), .air_in(c_12_0));
valve v_12_863 (.fluid_in(k_12_863), .fluid_out(k_11_431), .air_in(c_12_1));
valve v_12_864 (.fluid_in(k_12_864), .fluid_out(k_11_432), .air_in(c_12_0));
valve v_12_865 (.fluid_in(k_12_865), .fluid_out(k_11_432), .air_in(c_12_1));
valve v_12_866 (.fluid_in(k_12_866), .fluid_out(k_11_433), .air_in(c_12_0));
valve v_12_867 (.fluid_in(k_12_867), .fluid_out(k_11_433), .air_in(c_12_1));
valve v_12_868 (.fluid_in(k_12_868), .fluid_out(k_11_434), .air_in(c_12_0));
valve v_12_869 (.fluid_in(k_12_869), .fluid_out(k_11_434), .air_in(c_12_1));
valve v_12_870 (.fluid_in(k_12_870), .fluid_out(k_11_435), .air_in(c_12_0));
valve v_12_871 (.fluid_in(k_12_871), .fluid_out(k_11_435), .air_in(c_12_1));
valve v_12_872 (.fluid_in(k_12_872), .fluid_out(k_11_436), .air_in(c_12_0));
valve v_12_873 (.fluid_in(k_12_873), .fluid_out(k_11_436), .air_in(c_12_1));
valve v_12_874 (.fluid_in(k_12_874), .fluid_out(k_11_437), .air_in(c_12_0));
valve v_12_875 (.fluid_in(k_12_875), .fluid_out(k_11_437), .air_in(c_12_1));
valve v_12_876 (.fluid_in(k_12_876), .fluid_out(k_11_438), .air_in(c_12_0));
valve v_12_877 (.fluid_in(k_12_877), .fluid_out(k_11_438), .air_in(c_12_1));
valve v_12_878 (.fluid_in(k_12_878), .fluid_out(k_11_439), .air_in(c_12_0));
valve v_12_879 (.fluid_in(k_12_879), .fluid_out(k_11_439), .air_in(c_12_1));
valve v_12_880 (.fluid_in(k_12_880), .fluid_out(k_11_440), .air_in(c_12_0));
valve v_12_881 (.fluid_in(k_12_881), .fluid_out(k_11_440), .air_in(c_12_1));
valve v_12_882 (.fluid_in(k_12_882), .fluid_out(k_11_441), .air_in(c_12_0));
valve v_12_883 (.fluid_in(k_12_883), .fluid_out(k_11_441), .air_in(c_12_1));
valve v_12_884 (.fluid_in(k_12_884), .fluid_out(k_11_442), .air_in(c_12_0));
valve v_12_885 (.fluid_in(k_12_885), .fluid_out(k_11_442), .air_in(c_12_1));
valve v_12_886 (.fluid_in(k_12_886), .fluid_out(k_11_443), .air_in(c_12_0));
valve v_12_887 (.fluid_in(k_12_887), .fluid_out(k_11_443), .air_in(c_12_1));
valve v_12_888 (.fluid_in(k_12_888), .fluid_out(k_11_444), .air_in(c_12_0));
valve v_12_889 (.fluid_in(k_12_889), .fluid_out(k_11_444), .air_in(c_12_1));
valve v_12_890 (.fluid_in(k_12_890), .fluid_out(k_11_445), .air_in(c_12_0));
valve v_12_891 (.fluid_in(k_12_891), .fluid_out(k_11_445), .air_in(c_12_1));
valve v_12_892 (.fluid_in(k_12_892), .fluid_out(k_11_446), .air_in(c_12_0));
valve v_12_893 (.fluid_in(k_12_893), .fluid_out(k_11_446), .air_in(c_12_1));
valve v_12_894 (.fluid_in(k_12_894), .fluid_out(k_11_447), .air_in(c_12_0));
valve v_12_895 (.fluid_in(k_12_895), .fluid_out(k_11_447), .air_in(c_12_1));
valve v_12_896 (.fluid_in(k_12_896), .fluid_out(k_11_448), .air_in(c_12_0));
valve v_12_897 (.fluid_in(k_12_897), .fluid_out(k_11_448), .air_in(c_12_1));
valve v_12_898 (.fluid_in(k_12_898), .fluid_out(k_11_449), .air_in(c_12_0));
valve v_12_899 (.fluid_in(k_12_899), .fluid_out(k_11_449), .air_in(c_12_1));
valve v_12_900 (.fluid_in(k_12_900), .fluid_out(k_11_450), .air_in(c_12_0));
valve v_12_901 (.fluid_in(k_12_901), .fluid_out(k_11_450), .air_in(c_12_1));
valve v_12_902 (.fluid_in(k_12_902), .fluid_out(k_11_451), .air_in(c_12_0));
valve v_12_903 (.fluid_in(k_12_903), .fluid_out(k_11_451), .air_in(c_12_1));
valve v_12_904 (.fluid_in(k_12_904), .fluid_out(k_11_452), .air_in(c_12_0));
valve v_12_905 (.fluid_in(k_12_905), .fluid_out(k_11_452), .air_in(c_12_1));
valve v_12_906 (.fluid_in(k_12_906), .fluid_out(k_11_453), .air_in(c_12_0));
valve v_12_907 (.fluid_in(k_12_907), .fluid_out(k_11_453), .air_in(c_12_1));
valve v_12_908 (.fluid_in(k_12_908), .fluid_out(k_11_454), .air_in(c_12_0));
valve v_12_909 (.fluid_in(k_12_909), .fluid_out(k_11_454), .air_in(c_12_1));
valve v_12_910 (.fluid_in(k_12_910), .fluid_out(k_11_455), .air_in(c_12_0));
valve v_12_911 (.fluid_in(k_12_911), .fluid_out(k_11_455), .air_in(c_12_1));
valve v_12_912 (.fluid_in(k_12_912), .fluid_out(k_11_456), .air_in(c_12_0));
valve v_12_913 (.fluid_in(k_12_913), .fluid_out(k_11_456), .air_in(c_12_1));
valve v_12_914 (.fluid_in(k_12_914), .fluid_out(k_11_457), .air_in(c_12_0));
valve v_12_915 (.fluid_in(k_12_915), .fluid_out(k_11_457), .air_in(c_12_1));
valve v_12_916 (.fluid_in(k_12_916), .fluid_out(k_11_458), .air_in(c_12_0));
valve v_12_917 (.fluid_in(k_12_917), .fluid_out(k_11_458), .air_in(c_12_1));
valve v_12_918 (.fluid_in(k_12_918), .fluid_out(k_11_459), .air_in(c_12_0));
valve v_12_919 (.fluid_in(k_12_919), .fluid_out(k_11_459), .air_in(c_12_1));
valve v_12_920 (.fluid_in(k_12_920), .fluid_out(k_11_460), .air_in(c_12_0));
valve v_12_921 (.fluid_in(k_12_921), .fluid_out(k_11_460), .air_in(c_12_1));
valve v_12_922 (.fluid_in(k_12_922), .fluid_out(k_11_461), .air_in(c_12_0));
valve v_12_923 (.fluid_in(k_12_923), .fluid_out(k_11_461), .air_in(c_12_1));
valve v_12_924 (.fluid_in(k_12_924), .fluid_out(k_11_462), .air_in(c_12_0));
valve v_12_925 (.fluid_in(k_12_925), .fluid_out(k_11_462), .air_in(c_12_1));
valve v_12_926 (.fluid_in(k_12_926), .fluid_out(k_11_463), .air_in(c_12_0));
valve v_12_927 (.fluid_in(k_12_927), .fluid_out(k_11_463), .air_in(c_12_1));
valve v_12_928 (.fluid_in(k_12_928), .fluid_out(k_11_464), .air_in(c_12_0));
valve v_12_929 (.fluid_in(k_12_929), .fluid_out(k_11_464), .air_in(c_12_1));
valve v_12_930 (.fluid_in(k_12_930), .fluid_out(k_11_465), .air_in(c_12_0));
valve v_12_931 (.fluid_in(k_12_931), .fluid_out(k_11_465), .air_in(c_12_1));
valve v_12_932 (.fluid_in(k_12_932), .fluid_out(k_11_466), .air_in(c_12_0));
valve v_12_933 (.fluid_in(k_12_933), .fluid_out(k_11_466), .air_in(c_12_1));
valve v_12_934 (.fluid_in(k_12_934), .fluid_out(k_11_467), .air_in(c_12_0));
valve v_12_935 (.fluid_in(k_12_935), .fluid_out(k_11_467), .air_in(c_12_1));
valve v_12_936 (.fluid_in(k_12_936), .fluid_out(k_11_468), .air_in(c_12_0));
valve v_12_937 (.fluid_in(k_12_937), .fluid_out(k_11_468), .air_in(c_12_1));
valve v_12_938 (.fluid_in(k_12_938), .fluid_out(k_11_469), .air_in(c_12_0));
valve v_12_939 (.fluid_in(k_12_939), .fluid_out(k_11_469), .air_in(c_12_1));
valve v_12_940 (.fluid_in(k_12_940), .fluid_out(k_11_470), .air_in(c_12_0));
valve v_12_941 (.fluid_in(k_12_941), .fluid_out(k_11_470), .air_in(c_12_1));
valve v_12_942 (.fluid_in(k_12_942), .fluid_out(k_11_471), .air_in(c_12_0));
valve v_12_943 (.fluid_in(k_12_943), .fluid_out(k_11_471), .air_in(c_12_1));
valve v_12_944 (.fluid_in(k_12_944), .fluid_out(k_11_472), .air_in(c_12_0));
valve v_12_945 (.fluid_in(k_12_945), .fluid_out(k_11_472), .air_in(c_12_1));
valve v_12_946 (.fluid_in(k_12_946), .fluid_out(k_11_473), .air_in(c_12_0));
valve v_12_947 (.fluid_in(k_12_947), .fluid_out(k_11_473), .air_in(c_12_1));
valve v_12_948 (.fluid_in(k_12_948), .fluid_out(k_11_474), .air_in(c_12_0));
valve v_12_949 (.fluid_in(k_12_949), .fluid_out(k_11_474), .air_in(c_12_1));
valve v_12_950 (.fluid_in(k_12_950), .fluid_out(k_11_475), .air_in(c_12_0));
valve v_12_951 (.fluid_in(k_12_951), .fluid_out(k_11_475), .air_in(c_12_1));
valve v_12_952 (.fluid_in(k_12_952), .fluid_out(k_11_476), .air_in(c_12_0));
valve v_12_953 (.fluid_in(k_12_953), .fluid_out(k_11_476), .air_in(c_12_1));
valve v_12_954 (.fluid_in(k_12_954), .fluid_out(k_11_477), .air_in(c_12_0));
valve v_12_955 (.fluid_in(k_12_955), .fluid_out(k_11_477), .air_in(c_12_1));
valve v_12_956 (.fluid_in(k_12_956), .fluid_out(k_11_478), .air_in(c_12_0));
valve v_12_957 (.fluid_in(k_12_957), .fluid_out(k_11_478), .air_in(c_12_1));
valve v_12_958 (.fluid_in(k_12_958), .fluid_out(k_11_479), .air_in(c_12_0));
valve v_12_959 (.fluid_in(k_12_959), .fluid_out(k_11_479), .air_in(c_12_1));
valve v_12_960 (.fluid_in(k_12_960), .fluid_out(k_11_480), .air_in(c_12_0));
valve v_12_961 (.fluid_in(k_12_961), .fluid_out(k_11_480), .air_in(c_12_1));
valve v_12_962 (.fluid_in(k_12_962), .fluid_out(k_11_481), .air_in(c_12_0));
valve v_12_963 (.fluid_in(k_12_963), .fluid_out(k_11_481), .air_in(c_12_1));
valve v_12_964 (.fluid_in(k_12_964), .fluid_out(k_11_482), .air_in(c_12_0));
valve v_12_965 (.fluid_in(k_12_965), .fluid_out(k_11_482), .air_in(c_12_1));
valve v_12_966 (.fluid_in(k_12_966), .fluid_out(k_11_483), .air_in(c_12_0));
valve v_12_967 (.fluid_in(k_12_967), .fluid_out(k_11_483), .air_in(c_12_1));
valve v_12_968 (.fluid_in(k_12_968), .fluid_out(k_11_484), .air_in(c_12_0));
valve v_12_969 (.fluid_in(k_12_969), .fluid_out(k_11_484), .air_in(c_12_1));
valve v_12_970 (.fluid_in(k_12_970), .fluid_out(k_11_485), .air_in(c_12_0));
valve v_12_971 (.fluid_in(k_12_971), .fluid_out(k_11_485), .air_in(c_12_1));
valve v_12_972 (.fluid_in(k_12_972), .fluid_out(k_11_486), .air_in(c_12_0));
valve v_12_973 (.fluid_in(k_12_973), .fluid_out(k_11_486), .air_in(c_12_1));
valve v_12_974 (.fluid_in(k_12_974), .fluid_out(k_11_487), .air_in(c_12_0));
valve v_12_975 (.fluid_in(k_12_975), .fluid_out(k_11_487), .air_in(c_12_1));
valve v_12_976 (.fluid_in(k_12_976), .fluid_out(k_11_488), .air_in(c_12_0));
valve v_12_977 (.fluid_in(k_12_977), .fluid_out(k_11_488), .air_in(c_12_1));
valve v_12_978 (.fluid_in(k_12_978), .fluid_out(k_11_489), .air_in(c_12_0));
valve v_12_979 (.fluid_in(k_12_979), .fluid_out(k_11_489), .air_in(c_12_1));
valve v_12_980 (.fluid_in(k_12_980), .fluid_out(k_11_490), .air_in(c_12_0));
valve v_12_981 (.fluid_in(k_12_981), .fluid_out(k_11_490), .air_in(c_12_1));
valve v_12_982 (.fluid_in(k_12_982), .fluid_out(k_11_491), .air_in(c_12_0));
valve v_12_983 (.fluid_in(k_12_983), .fluid_out(k_11_491), .air_in(c_12_1));
valve v_12_984 (.fluid_in(k_12_984), .fluid_out(k_11_492), .air_in(c_12_0));
valve v_12_985 (.fluid_in(k_12_985), .fluid_out(k_11_492), .air_in(c_12_1));
valve v_12_986 (.fluid_in(k_12_986), .fluid_out(k_11_493), .air_in(c_12_0));
valve v_12_987 (.fluid_in(k_12_987), .fluid_out(k_11_493), .air_in(c_12_1));
valve v_12_988 (.fluid_in(k_12_988), .fluid_out(k_11_494), .air_in(c_12_0));
valve v_12_989 (.fluid_in(k_12_989), .fluid_out(k_11_494), .air_in(c_12_1));
valve v_12_990 (.fluid_in(k_12_990), .fluid_out(k_11_495), .air_in(c_12_0));
valve v_12_991 (.fluid_in(k_12_991), .fluid_out(k_11_495), .air_in(c_12_1));
valve v_12_992 (.fluid_in(k_12_992), .fluid_out(k_11_496), .air_in(c_12_0));
valve v_12_993 (.fluid_in(k_12_993), .fluid_out(k_11_496), .air_in(c_12_1));
valve v_12_994 (.fluid_in(k_12_994), .fluid_out(k_11_497), .air_in(c_12_0));
valve v_12_995 (.fluid_in(k_12_995), .fluid_out(k_11_497), .air_in(c_12_1));
valve v_12_996 (.fluid_in(k_12_996), .fluid_out(k_11_498), .air_in(c_12_0));
valve v_12_997 (.fluid_in(k_12_997), .fluid_out(k_11_498), .air_in(c_12_1));
valve v_12_998 (.fluid_in(k_12_998), .fluid_out(k_11_499), .air_in(c_12_0));
valve v_12_999 (.fluid_in(k_12_999), .fluid_out(k_11_499), .air_in(c_12_1));
valve v_12_1000 (.fluid_in(k_12_1000), .fluid_out(k_11_500), .air_in(c_12_0));
valve v_12_1001 (.fluid_in(k_12_1001), .fluid_out(k_11_500), .air_in(c_12_1));
valve v_12_1002 (.fluid_in(k_12_1002), .fluid_out(k_11_501), .air_in(c_12_0));
valve v_12_1003 (.fluid_in(k_12_1003), .fluid_out(k_11_501), .air_in(c_12_1));
valve v_12_1004 (.fluid_in(k_12_1004), .fluid_out(k_11_502), .air_in(c_12_0));
valve v_12_1005 (.fluid_in(k_12_1005), .fluid_out(k_11_502), .air_in(c_12_1));
valve v_12_1006 (.fluid_in(k_12_1006), .fluid_out(k_11_503), .air_in(c_12_0));
valve v_12_1007 (.fluid_in(k_12_1007), .fluid_out(k_11_503), .air_in(c_12_1));
valve v_12_1008 (.fluid_in(k_12_1008), .fluid_out(k_11_504), .air_in(c_12_0));
valve v_12_1009 (.fluid_in(k_12_1009), .fluid_out(k_11_504), .air_in(c_12_1));
valve v_12_1010 (.fluid_in(k_12_1010), .fluid_out(k_11_505), .air_in(c_12_0));
valve v_12_1011 (.fluid_in(k_12_1011), .fluid_out(k_11_505), .air_in(c_12_1));
valve v_12_1012 (.fluid_in(k_12_1012), .fluid_out(k_11_506), .air_in(c_12_0));
valve v_12_1013 (.fluid_in(k_12_1013), .fluid_out(k_11_506), .air_in(c_12_1));
valve v_12_1014 (.fluid_in(k_12_1014), .fluid_out(k_11_507), .air_in(c_12_0));
valve v_12_1015 (.fluid_in(k_12_1015), .fluid_out(k_11_507), .air_in(c_12_1));
valve v_12_1016 (.fluid_in(k_12_1016), .fluid_out(k_11_508), .air_in(c_12_0));
valve v_12_1017 (.fluid_in(k_12_1017), .fluid_out(k_11_508), .air_in(c_12_1));
valve v_12_1018 (.fluid_in(k_12_1018), .fluid_out(k_11_509), .air_in(c_12_0));
valve v_12_1019 (.fluid_in(k_12_1019), .fluid_out(k_11_509), .air_in(c_12_1));
valve v_12_1020 (.fluid_in(k_12_1020), .fluid_out(k_11_510), .air_in(c_12_0));
valve v_12_1021 (.fluid_in(k_12_1021), .fluid_out(k_11_510), .air_in(c_12_1));
valve v_12_1022 (.fluid_in(k_12_1022), .fluid_out(k_11_511), .air_in(c_12_0));
valve v_12_1023 (.fluid_in(k_12_1023), .fluid_out(k_11_511), .air_in(c_12_1));
valve v_12_1024 (.fluid_in(k_12_1024), .fluid_out(k_11_512), .air_in(c_12_0));
valve v_12_1025 (.fluid_in(k_12_1025), .fluid_out(k_11_512), .air_in(c_12_1));
valve v_12_1026 (.fluid_in(k_12_1026), .fluid_out(k_11_513), .air_in(c_12_0));
valve v_12_1027 (.fluid_in(k_12_1027), .fluid_out(k_11_513), .air_in(c_12_1));
valve v_12_1028 (.fluid_in(k_12_1028), .fluid_out(k_11_514), .air_in(c_12_0));
valve v_12_1029 (.fluid_in(k_12_1029), .fluid_out(k_11_514), .air_in(c_12_1));
valve v_12_1030 (.fluid_in(k_12_1030), .fluid_out(k_11_515), .air_in(c_12_0));
valve v_12_1031 (.fluid_in(k_12_1031), .fluid_out(k_11_515), .air_in(c_12_1));
valve v_12_1032 (.fluid_in(k_12_1032), .fluid_out(k_11_516), .air_in(c_12_0));
valve v_12_1033 (.fluid_in(k_12_1033), .fluid_out(k_11_516), .air_in(c_12_1));
valve v_12_1034 (.fluid_in(k_12_1034), .fluid_out(k_11_517), .air_in(c_12_0));
valve v_12_1035 (.fluid_in(k_12_1035), .fluid_out(k_11_517), .air_in(c_12_1));
valve v_12_1036 (.fluid_in(k_12_1036), .fluid_out(k_11_518), .air_in(c_12_0));
valve v_12_1037 (.fluid_in(k_12_1037), .fluid_out(k_11_518), .air_in(c_12_1));
valve v_12_1038 (.fluid_in(k_12_1038), .fluid_out(k_11_519), .air_in(c_12_0));
valve v_12_1039 (.fluid_in(k_12_1039), .fluid_out(k_11_519), .air_in(c_12_1));
valve v_12_1040 (.fluid_in(k_12_1040), .fluid_out(k_11_520), .air_in(c_12_0));
valve v_12_1041 (.fluid_in(k_12_1041), .fluid_out(k_11_520), .air_in(c_12_1));
valve v_12_1042 (.fluid_in(k_12_1042), .fluid_out(k_11_521), .air_in(c_12_0));
valve v_12_1043 (.fluid_in(k_12_1043), .fluid_out(k_11_521), .air_in(c_12_1));
valve v_12_1044 (.fluid_in(k_12_1044), .fluid_out(k_11_522), .air_in(c_12_0));
valve v_12_1045 (.fluid_in(k_12_1045), .fluid_out(k_11_522), .air_in(c_12_1));
valve v_12_1046 (.fluid_in(k_12_1046), .fluid_out(k_11_523), .air_in(c_12_0));
valve v_12_1047 (.fluid_in(k_12_1047), .fluid_out(k_11_523), .air_in(c_12_1));
valve v_12_1048 (.fluid_in(k_12_1048), .fluid_out(k_11_524), .air_in(c_12_0));
valve v_12_1049 (.fluid_in(k_12_1049), .fluid_out(k_11_524), .air_in(c_12_1));
valve v_12_1050 (.fluid_in(k_12_1050), .fluid_out(k_11_525), .air_in(c_12_0));
valve v_12_1051 (.fluid_in(k_12_1051), .fluid_out(k_11_525), .air_in(c_12_1));
valve v_12_1052 (.fluid_in(k_12_1052), .fluid_out(k_11_526), .air_in(c_12_0));
valve v_12_1053 (.fluid_in(k_12_1053), .fluid_out(k_11_526), .air_in(c_12_1));
valve v_12_1054 (.fluid_in(k_12_1054), .fluid_out(k_11_527), .air_in(c_12_0));
valve v_12_1055 (.fluid_in(k_12_1055), .fluid_out(k_11_527), .air_in(c_12_1));
valve v_12_1056 (.fluid_in(k_12_1056), .fluid_out(k_11_528), .air_in(c_12_0));
valve v_12_1057 (.fluid_in(k_12_1057), .fluid_out(k_11_528), .air_in(c_12_1));
valve v_12_1058 (.fluid_in(k_12_1058), .fluid_out(k_11_529), .air_in(c_12_0));
valve v_12_1059 (.fluid_in(k_12_1059), .fluid_out(k_11_529), .air_in(c_12_1));
valve v_12_1060 (.fluid_in(k_12_1060), .fluid_out(k_11_530), .air_in(c_12_0));
valve v_12_1061 (.fluid_in(k_12_1061), .fluid_out(k_11_530), .air_in(c_12_1));
valve v_12_1062 (.fluid_in(k_12_1062), .fluid_out(k_11_531), .air_in(c_12_0));
valve v_12_1063 (.fluid_in(k_12_1063), .fluid_out(k_11_531), .air_in(c_12_1));
valve v_12_1064 (.fluid_in(k_12_1064), .fluid_out(k_11_532), .air_in(c_12_0));
valve v_12_1065 (.fluid_in(k_12_1065), .fluid_out(k_11_532), .air_in(c_12_1));
valve v_12_1066 (.fluid_in(k_12_1066), .fluid_out(k_11_533), .air_in(c_12_0));
valve v_12_1067 (.fluid_in(k_12_1067), .fluid_out(k_11_533), .air_in(c_12_1));
valve v_12_1068 (.fluid_in(k_12_1068), .fluid_out(k_11_534), .air_in(c_12_0));
valve v_12_1069 (.fluid_in(k_12_1069), .fluid_out(k_11_534), .air_in(c_12_1));
valve v_12_1070 (.fluid_in(k_12_1070), .fluid_out(k_11_535), .air_in(c_12_0));
valve v_12_1071 (.fluid_in(k_12_1071), .fluid_out(k_11_535), .air_in(c_12_1));
valve v_12_1072 (.fluid_in(k_12_1072), .fluid_out(k_11_536), .air_in(c_12_0));
valve v_12_1073 (.fluid_in(k_12_1073), .fluid_out(k_11_536), .air_in(c_12_1));
valve v_12_1074 (.fluid_in(k_12_1074), .fluid_out(k_11_537), .air_in(c_12_0));
valve v_12_1075 (.fluid_in(k_12_1075), .fluid_out(k_11_537), .air_in(c_12_1));
valve v_12_1076 (.fluid_in(k_12_1076), .fluid_out(k_11_538), .air_in(c_12_0));
valve v_12_1077 (.fluid_in(k_12_1077), .fluid_out(k_11_538), .air_in(c_12_1));
valve v_12_1078 (.fluid_in(k_12_1078), .fluid_out(k_11_539), .air_in(c_12_0));
valve v_12_1079 (.fluid_in(k_12_1079), .fluid_out(k_11_539), .air_in(c_12_1));
valve v_12_1080 (.fluid_in(k_12_1080), .fluid_out(k_11_540), .air_in(c_12_0));
valve v_12_1081 (.fluid_in(k_12_1081), .fluid_out(k_11_540), .air_in(c_12_1));
valve v_12_1082 (.fluid_in(k_12_1082), .fluid_out(k_11_541), .air_in(c_12_0));
valve v_12_1083 (.fluid_in(k_12_1083), .fluid_out(k_11_541), .air_in(c_12_1));
valve v_12_1084 (.fluid_in(k_12_1084), .fluid_out(k_11_542), .air_in(c_12_0));
valve v_12_1085 (.fluid_in(k_12_1085), .fluid_out(k_11_542), .air_in(c_12_1));
valve v_12_1086 (.fluid_in(k_12_1086), .fluid_out(k_11_543), .air_in(c_12_0));
valve v_12_1087 (.fluid_in(k_12_1087), .fluid_out(k_11_543), .air_in(c_12_1));
valve v_12_1088 (.fluid_in(k_12_1088), .fluid_out(k_11_544), .air_in(c_12_0));
valve v_12_1089 (.fluid_in(k_12_1089), .fluid_out(k_11_544), .air_in(c_12_1));
valve v_12_1090 (.fluid_in(k_12_1090), .fluid_out(k_11_545), .air_in(c_12_0));
valve v_12_1091 (.fluid_in(k_12_1091), .fluid_out(k_11_545), .air_in(c_12_1));
valve v_12_1092 (.fluid_in(k_12_1092), .fluid_out(k_11_546), .air_in(c_12_0));
valve v_12_1093 (.fluid_in(k_12_1093), .fluid_out(k_11_546), .air_in(c_12_1));
valve v_12_1094 (.fluid_in(k_12_1094), .fluid_out(k_11_547), .air_in(c_12_0));
valve v_12_1095 (.fluid_in(k_12_1095), .fluid_out(k_11_547), .air_in(c_12_1));
valve v_12_1096 (.fluid_in(k_12_1096), .fluid_out(k_11_548), .air_in(c_12_0));
valve v_12_1097 (.fluid_in(k_12_1097), .fluid_out(k_11_548), .air_in(c_12_1));
valve v_12_1098 (.fluid_in(k_12_1098), .fluid_out(k_11_549), .air_in(c_12_0));
valve v_12_1099 (.fluid_in(k_12_1099), .fluid_out(k_11_549), .air_in(c_12_1));
valve v_12_1100 (.fluid_in(k_12_1100), .fluid_out(k_11_550), .air_in(c_12_0));
valve v_12_1101 (.fluid_in(k_12_1101), .fluid_out(k_11_550), .air_in(c_12_1));
valve v_12_1102 (.fluid_in(k_12_1102), .fluid_out(k_11_551), .air_in(c_12_0));
valve v_12_1103 (.fluid_in(k_12_1103), .fluid_out(k_11_551), .air_in(c_12_1));
valve v_12_1104 (.fluid_in(k_12_1104), .fluid_out(k_11_552), .air_in(c_12_0));
valve v_12_1105 (.fluid_in(k_12_1105), .fluid_out(k_11_552), .air_in(c_12_1));
valve v_12_1106 (.fluid_in(k_12_1106), .fluid_out(k_11_553), .air_in(c_12_0));
valve v_12_1107 (.fluid_in(k_12_1107), .fluid_out(k_11_553), .air_in(c_12_1));
valve v_12_1108 (.fluid_in(k_12_1108), .fluid_out(k_11_554), .air_in(c_12_0));
valve v_12_1109 (.fluid_in(k_12_1109), .fluid_out(k_11_554), .air_in(c_12_1));
valve v_12_1110 (.fluid_in(k_12_1110), .fluid_out(k_11_555), .air_in(c_12_0));
valve v_12_1111 (.fluid_in(k_12_1111), .fluid_out(k_11_555), .air_in(c_12_1));
valve v_12_1112 (.fluid_in(k_12_1112), .fluid_out(k_11_556), .air_in(c_12_0));
valve v_12_1113 (.fluid_in(k_12_1113), .fluid_out(k_11_556), .air_in(c_12_1));
valve v_12_1114 (.fluid_in(k_12_1114), .fluid_out(k_11_557), .air_in(c_12_0));
valve v_12_1115 (.fluid_in(k_12_1115), .fluid_out(k_11_557), .air_in(c_12_1));
valve v_12_1116 (.fluid_in(k_12_1116), .fluid_out(k_11_558), .air_in(c_12_0));
valve v_12_1117 (.fluid_in(k_12_1117), .fluid_out(k_11_558), .air_in(c_12_1));
valve v_12_1118 (.fluid_in(k_12_1118), .fluid_out(k_11_559), .air_in(c_12_0));
valve v_12_1119 (.fluid_in(k_12_1119), .fluid_out(k_11_559), .air_in(c_12_1));
valve v_12_1120 (.fluid_in(k_12_1120), .fluid_out(k_11_560), .air_in(c_12_0));
valve v_12_1121 (.fluid_in(k_12_1121), .fluid_out(k_11_560), .air_in(c_12_1));
valve v_12_1122 (.fluid_in(k_12_1122), .fluid_out(k_11_561), .air_in(c_12_0));
valve v_12_1123 (.fluid_in(k_12_1123), .fluid_out(k_11_561), .air_in(c_12_1));
valve v_12_1124 (.fluid_in(k_12_1124), .fluid_out(k_11_562), .air_in(c_12_0));
valve v_12_1125 (.fluid_in(k_12_1125), .fluid_out(k_11_562), .air_in(c_12_1));
valve v_12_1126 (.fluid_in(k_12_1126), .fluid_out(k_11_563), .air_in(c_12_0));
valve v_12_1127 (.fluid_in(k_12_1127), .fluid_out(k_11_563), .air_in(c_12_1));
valve v_12_1128 (.fluid_in(k_12_1128), .fluid_out(k_11_564), .air_in(c_12_0));
valve v_12_1129 (.fluid_in(k_12_1129), .fluid_out(k_11_564), .air_in(c_12_1));
valve v_12_1130 (.fluid_in(k_12_1130), .fluid_out(k_11_565), .air_in(c_12_0));
valve v_12_1131 (.fluid_in(k_12_1131), .fluid_out(k_11_565), .air_in(c_12_1));
valve v_12_1132 (.fluid_in(k_12_1132), .fluid_out(k_11_566), .air_in(c_12_0));
valve v_12_1133 (.fluid_in(k_12_1133), .fluid_out(k_11_566), .air_in(c_12_1));
valve v_12_1134 (.fluid_in(k_12_1134), .fluid_out(k_11_567), .air_in(c_12_0));
valve v_12_1135 (.fluid_in(k_12_1135), .fluid_out(k_11_567), .air_in(c_12_1));
valve v_12_1136 (.fluid_in(k_12_1136), .fluid_out(k_11_568), .air_in(c_12_0));
valve v_12_1137 (.fluid_in(k_12_1137), .fluid_out(k_11_568), .air_in(c_12_1));
valve v_12_1138 (.fluid_in(k_12_1138), .fluid_out(k_11_569), .air_in(c_12_0));
valve v_12_1139 (.fluid_in(k_12_1139), .fluid_out(k_11_569), .air_in(c_12_1));
valve v_12_1140 (.fluid_in(k_12_1140), .fluid_out(k_11_570), .air_in(c_12_0));
valve v_12_1141 (.fluid_in(k_12_1141), .fluid_out(k_11_570), .air_in(c_12_1));
valve v_12_1142 (.fluid_in(k_12_1142), .fluid_out(k_11_571), .air_in(c_12_0));
valve v_12_1143 (.fluid_in(k_12_1143), .fluid_out(k_11_571), .air_in(c_12_1));
valve v_12_1144 (.fluid_in(k_12_1144), .fluid_out(k_11_572), .air_in(c_12_0));
valve v_12_1145 (.fluid_in(k_12_1145), .fluid_out(k_11_572), .air_in(c_12_1));
valve v_12_1146 (.fluid_in(k_12_1146), .fluid_out(k_11_573), .air_in(c_12_0));
valve v_12_1147 (.fluid_in(k_12_1147), .fluid_out(k_11_573), .air_in(c_12_1));
valve v_12_1148 (.fluid_in(k_12_1148), .fluid_out(k_11_574), .air_in(c_12_0));
valve v_12_1149 (.fluid_in(k_12_1149), .fluid_out(k_11_574), .air_in(c_12_1));
valve v_12_1150 (.fluid_in(k_12_1150), .fluid_out(k_11_575), .air_in(c_12_0));
valve v_12_1151 (.fluid_in(k_12_1151), .fluid_out(k_11_575), .air_in(c_12_1));
valve v_12_1152 (.fluid_in(k_12_1152), .fluid_out(k_11_576), .air_in(c_12_0));
valve v_12_1153 (.fluid_in(k_12_1153), .fluid_out(k_11_576), .air_in(c_12_1));
valve v_12_1154 (.fluid_in(k_12_1154), .fluid_out(k_11_577), .air_in(c_12_0));
valve v_12_1155 (.fluid_in(k_12_1155), .fluid_out(k_11_577), .air_in(c_12_1));
valve v_12_1156 (.fluid_in(k_12_1156), .fluid_out(k_11_578), .air_in(c_12_0));
valve v_12_1157 (.fluid_in(k_12_1157), .fluid_out(k_11_578), .air_in(c_12_1));
valve v_12_1158 (.fluid_in(k_12_1158), .fluid_out(k_11_579), .air_in(c_12_0));
valve v_12_1159 (.fluid_in(k_12_1159), .fluid_out(k_11_579), .air_in(c_12_1));
valve v_12_1160 (.fluid_in(k_12_1160), .fluid_out(k_11_580), .air_in(c_12_0));
valve v_12_1161 (.fluid_in(k_12_1161), .fluid_out(k_11_580), .air_in(c_12_1));
valve v_12_1162 (.fluid_in(k_12_1162), .fluid_out(k_11_581), .air_in(c_12_0));
valve v_12_1163 (.fluid_in(k_12_1163), .fluid_out(k_11_581), .air_in(c_12_1));
valve v_12_1164 (.fluid_in(k_12_1164), .fluid_out(k_11_582), .air_in(c_12_0));
valve v_12_1165 (.fluid_in(k_12_1165), .fluid_out(k_11_582), .air_in(c_12_1));
valve v_12_1166 (.fluid_in(k_12_1166), .fluid_out(k_11_583), .air_in(c_12_0));
valve v_12_1167 (.fluid_in(k_12_1167), .fluid_out(k_11_583), .air_in(c_12_1));
valve v_12_1168 (.fluid_in(k_12_1168), .fluid_out(k_11_584), .air_in(c_12_0));
valve v_12_1169 (.fluid_in(k_12_1169), .fluid_out(k_11_584), .air_in(c_12_1));
valve v_12_1170 (.fluid_in(k_12_1170), .fluid_out(k_11_585), .air_in(c_12_0));
valve v_12_1171 (.fluid_in(k_12_1171), .fluid_out(k_11_585), .air_in(c_12_1));
valve v_12_1172 (.fluid_in(k_12_1172), .fluid_out(k_11_586), .air_in(c_12_0));
valve v_12_1173 (.fluid_in(k_12_1173), .fluid_out(k_11_586), .air_in(c_12_1));
valve v_12_1174 (.fluid_in(k_12_1174), .fluid_out(k_11_587), .air_in(c_12_0));
valve v_12_1175 (.fluid_in(k_12_1175), .fluid_out(k_11_587), .air_in(c_12_1));
valve v_12_1176 (.fluid_in(k_12_1176), .fluid_out(k_11_588), .air_in(c_12_0));
valve v_12_1177 (.fluid_in(k_12_1177), .fluid_out(k_11_588), .air_in(c_12_1));
valve v_12_1178 (.fluid_in(k_12_1178), .fluid_out(k_11_589), .air_in(c_12_0));
valve v_12_1179 (.fluid_in(k_12_1179), .fluid_out(k_11_589), .air_in(c_12_1));
valve v_12_1180 (.fluid_in(k_12_1180), .fluid_out(k_11_590), .air_in(c_12_0));
valve v_12_1181 (.fluid_in(k_12_1181), .fluid_out(k_11_590), .air_in(c_12_1));
valve v_12_1182 (.fluid_in(k_12_1182), .fluid_out(k_11_591), .air_in(c_12_0));
valve v_12_1183 (.fluid_in(k_12_1183), .fluid_out(k_11_591), .air_in(c_12_1));
valve v_12_1184 (.fluid_in(k_12_1184), .fluid_out(k_11_592), .air_in(c_12_0));
valve v_12_1185 (.fluid_in(k_12_1185), .fluid_out(k_11_592), .air_in(c_12_1));
valve v_12_1186 (.fluid_in(k_12_1186), .fluid_out(k_11_593), .air_in(c_12_0));
valve v_12_1187 (.fluid_in(k_12_1187), .fluid_out(k_11_593), .air_in(c_12_1));
valve v_12_1188 (.fluid_in(k_12_1188), .fluid_out(k_11_594), .air_in(c_12_0));
valve v_12_1189 (.fluid_in(k_12_1189), .fluid_out(k_11_594), .air_in(c_12_1));
valve v_12_1190 (.fluid_in(k_12_1190), .fluid_out(k_11_595), .air_in(c_12_0));
valve v_12_1191 (.fluid_in(k_12_1191), .fluid_out(k_11_595), .air_in(c_12_1));
valve v_12_1192 (.fluid_in(k_12_1192), .fluid_out(k_11_596), .air_in(c_12_0));
valve v_12_1193 (.fluid_in(k_12_1193), .fluid_out(k_11_596), .air_in(c_12_1));
valve v_12_1194 (.fluid_in(k_12_1194), .fluid_out(k_11_597), .air_in(c_12_0));
valve v_12_1195 (.fluid_in(k_12_1195), .fluid_out(k_11_597), .air_in(c_12_1));
valve v_12_1196 (.fluid_in(k_12_1196), .fluid_out(k_11_598), .air_in(c_12_0));
valve v_12_1197 (.fluid_in(k_12_1197), .fluid_out(k_11_598), .air_in(c_12_1));
valve v_12_1198 (.fluid_in(k_12_1198), .fluid_out(k_11_599), .air_in(c_12_0));
valve v_12_1199 (.fluid_in(k_12_1199), .fluid_out(k_11_599), .air_in(c_12_1));
valve v_12_1200 (.fluid_in(k_12_1200), .fluid_out(k_11_600), .air_in(c_12_0));
valve v_12_1201 (.fluid_in(k_12_1201), .fluid_out(k_11_600), .air_in(c_12_1));
valve v_12_1202 (.fluid_in(k_12_1202), .fluid_out(k_11_601), .air_in(c_12_0));
valve v_12_1203 (.fluid_in(k_12_1203), .fluid_out(k_11_601), .air_in(c_12_1));
valve v_12_1204 (.fluid_in(k_12_1204), .fluid_out(k_11_602), .air_in(c_12_0));
valve v_12_1205 (.fluid_in(k_12_1205), .fluid_out(k_11_602), .air_in(c_12_1));
valve v_12_1206 (.fluid_in(k_12_1206), .fluid_out(k_11_603), .air_in(c_12_0));
valve v_12_1207 (.fluid_in(k_12_1207), .fluid_out(k_11_603), .air_in(c_12_1));
valve v_12_1208 (.fluid_in(k_12_1208), .fluid_out(k_11_604), .air_in(c_12_0));
valve v_12_1209 (.fluid_in(k_12_1209), .fluid_out(k_11_604), .air_in(c_12_1));
valve v_12_1210 (.fluid_in(k_12_1210), .fluid_out(k_11_605), .air_in(c_12_0));
valve v_12_1211 (.fluid_in(k_12_1211), .fluid_out(k_11_605), .air_in(c_12_1));
valve v_12_1212 (.fluid_in(k_12_1212), .fluid_out(k_11_606), .air_in(c_12_0));
valve v_12_1213 (.fluid_in(k_12_1213), .fluid_out(k_11_606), .air_in(c_12_1));
valve v_12_1214 (.fluid_in(k_12_1214), .fluid_out(k_11_607), .air_in(c_12_0));
valve v_12_1215 (.fluid_in(k_12_1215), .fluid_out(k_11_607), .air_in(c_12_1));
valve v_12_1216 (.fluid_in(k_12_1216), .fluid_out(k_11_608), .air_in(c_12_0));
valve v_12_1217 (.fluid_in(k_12_1217), .fluid_out(k_11_608), .air_in(c_12_1));
valve v_12_1218 (.fluid_in(k_12_1218), .fluid_out(k_11_609), .air_in(c_12_0));
valve v_12_1219 (.fluid_in(k_12_1219), .fluid_out(k_11_609), .air_in(c_12_1));
valve v_12_1220 (.fluid_in(k_12_1220), .fluid_out(k_11_610), .air_in(c_12_0));
valve v_12_1221 (.fluid_in(k_12_1221), .fluid_out(k_11_610), .air_in(c_12_1));
valve v_12_1222 (.fluid_in(k_12_1222), .fluid_out(k_11_611), .air_in(c_12_0));
valve v_12_1223 (.fluid_in(k_12_1223), .fluid_out(k_11_611), .air_in(c_12_1));
valve v_12_1224 (.fluid_in(k_12_1224), .fluid_out(k_11_612), .air_in(c_12_0));
valve v_12_1225 (.fluid_in(k_12_1225), .fluid_out(k_11_612), .air_in(c_12_1));
valve v_12_1226 (.fluid_in(k_12_1226), .fluid_out(k_11_613), .air_in(c_12_0));
valve v_12_1227 (.fluid_in(k_12_1227), .fluid_out(k_11_613), .air_in(c_12_1));
valve v_12_1228 (.fluid_in(k_12_1228), .fluid_out(k_11_614), .air_in(c_12_0));
valve v_12_1229 (.fluid_in(k_12_1229), .fluid_out(k_11_614), .air_in(c_12_1));
valve v_12_1230 (.fluid_in(k_12_1230), .fluid_out(k_11_615), .air_in(c_12_0));
valve v_12_1231 (.fluid_in(k_12_1231), .fluid_out(k_11_615), .air_in(c_12_1));
valve v_12_1232 (.fluid_in(k_12_1232), .fluid_out(k_11_616), .air_in(c_12_0));
valve v_12_1233 (.fluid_in(k_12_1233), .fluid_out(k_11_616), .air_in(c_12_1));
valve v_12_1234 (.fluid_in(k_12_1234), .fluid_out(k_11_617), .air_in(c_12_0));
valve v_12_1235 (.fluid_in(k_12_1235), .fluid_out(k_11_617), .air_in(c_12_1));
valve v_12_1236 (.fluid_in(k_12_1236), .fluid_out(k_11_618), .air_in(c_12_0));
valve v_12_1237 (.fluid_in(k_12_1237), .fluid_out(k_11_618), .air_in(c_12_1));
valve v_12_1238 (.fluid_in(k_12_1238), .fluid_out(k_11_619), .air_in(c_12_0));
valve v_12_1239 (.fluid_in(k_12_1239), .fluid_out(k_11_619), .air_in(c_12_1));
valve v_12_1240 (.fluid_in(k_12_1240), .fluid_out(k_11_620), .air_in(c_12_0));
valve v_12_1241 (.fluid_in(k_12_1241), .fluid_out(k_11_620), .air_in(c_12_1));
valve v_12_1242 (.fluid_in(k_12_1242), .fluid_out(k_11_621), .air_in(c_12_0));
valve v_12_1243 (.fluid_in(k_12_1243), .fluid_out(k_11_621), .air_in(c_12_1));
valve v_12_1244 (.fluid_in(k_12_1244), .fluid_out(k_11_622), .air_in(c_12_0));
valve v_12_1245 (.fluid_in(k_12_1245), .fluid_out(k_11_622), .air_in(c_12_1));
valve v_12_1246 (.fluid_in(k_12_1246), .fluid_out(k_11_623), .air_in(c_12_0));
valve v_12_1247 (.fluid_in(k_12_1247), .fluid_out(k_11_623), .air_in(c_12_1));
valve v_12_1248 (.fluid_in(k_12_1248), .fluid_out(k_11_624), .air_in(c_12_0));
valve v_12_1249 (.fluid_in(k_12_1249), .fluid_out(k_11_624), .air_in(c_12_1));
valve v_12_1250 (.fluid_in(k_12_1250), .fluid_out(k_11_625), .air_in(c_12_0));
valve v_12_1251 (.fluid_in(k_12_1251), .fluid_out(k_11_625), .air_in(c_12_1));
valve v_12_1252 (.fluid_in(k_12_1252), .fluid_out(k_11_626), .air_in(c_12_0));
valve v_12_1253 (.fluid_in(k_12_1253), .fluid_out(k_11_626), .air_in(c_12_1));
valve v_12_1254 (.fluid_in(k_12_1254), .fluid_out(k_11_627), .air_in(c_12_0));
valve v_12_1255 (.fluid_in(k_12_1255), .fluid_out(k_11_627), .air_in(c_12_1));
valve v_12_1256 (.fluid_in(k_12_1256), .fluid_out(k_11_628), .air_in(c_12_0));
valve v_12_1257 (.fluid_in(k_12_1257), .fluid_out(k_11_628), .air_in(c_12_1));
valve v_12_1258 (.fluid_in(k_12_1258), .fluid_out(k_11_629), .air_in(c_12_0));
valve v_12_1259 (.fluid_in(k_12_1259), .fluid_out(k_11_629), .air_in(c_12_1));
valve v_12_1260 (.fluid_in(k_12_1260), .fluid_out(k_11_630), .air_in(c_12_0));
valve v_12_1261 (.fluid_in(k_12_1261), .fluid_out(k_11_630), .air_in(c_12_1));
valve v_12_1262 (.fluid_in(k_12_1262), .fluid_out(k_11_631), .air_in(c_12_0));
valve v_12_1263 (.fluid_in(k_12_1263), .fluid_out(k_11_631), .air_in(c_12_1));
valve v_12_1264 (.fluid_in(k_12_1264), .fluid_out(k_11_632), .air_in(c_12_0));
valve v_12_1265 (.fluid_in(k_12_1265), .fluid_out(k_11_632), .air_in(c_12_1));
valve v_12_1266 (.fluid_in(k_12_1266), .fluid_out(k_11_633), .air_in(c_12_0));
valve v_12_1267 (.fluid_in(k_12_1267), .fluid_out(k_11_633), .air_in(c_12_1));
valve v_12_1268 (.fluid_in(k_12_1268), .fluid_out(k_11_634), .air_in(c_12_0));
valve v_12_1269 (.fluid_in(k_12_1269), .fluid_out(k_11_634), .air_in(c_12_1));
valve v_12_1270 (.fluid_in(k_12_1270), .fluid_out(k_11_635), .air_in(c_12_0));
valve v_12_1271 (.fluid_in(k_12_1271), .fluid_out(k_11_635), .air_in(c_12_1));
valve v_12_1272 (.fluid_in(k_12_1272), .fluid_out(k_11_636), .air_in(c_12_0));
valve v_12_1273 (.fluid_in(k_12_1273), .fluid_out(k_11_636), .air_in(c_12_1));
valve v_12_1274 (.fluid_in(k_12_1274), .fluid_out(k_11_637), .air_in(c_12_0));
valve v_12_1275 (.fluid_in(k_12_1275), .fluid_out(k_11_637), .air_in(c_12_1));
valve v_12_1276 (.fluid_in(k_12_1276), .fluid_out(k_11_638), .air_in(c_12_0));
valve v_12_1277 (.fluid_in(k_12_1277), .fluid_out(k_11_638), .air_in(c_12_1));
valve v_12_1278 (.fluid_in(k_12_1278), .fluid_out(k_11_639), .air_in(c_12_0));
valve v_12_1279 (.fluid_in(k_12_1279), .fluid_out(k_11_639), .air_in(c_12_1));
valve v_12_1280 (.fluid_in(k_12_1280), .fluid_out(k_11_640), .air_in(c_12_0));
valve v_12_1281 (.fluid_in(k_12_1281), .fluid_out(k_11_640), .air_in(c_12_1));
valve v_12_1282 (.fluid_in(k_12_1282), .fluid_out(k_11_641), .air_in(c_12_0));
valve v_12_1283 (.fluid_in(k_12_1283), .fluid_out(k_11_641), .air_in(c_12_1));
valve v_12_1284 (.fluid_in(k_12_1284), .fluid_out(k_11_642), .air_in(c_12_0));
valve v_12_1285 (.fluid_in(k_12_1285), .fluid_out(k_11_642), .air_in(c_12_1));
valve v_12_1286 (.fluid_in(k_12_1286), .fluid_out(k_11_643), .air_in(c_12_0));
valve v_12_1287 (.fluid_in(k_12_1287), .fluid_out(k_11_643), .air_in(c_12_1));
valve v_12_1288 (.fluid_in(k_12_1288), .fluid_out(k_11_644), .air_in(c_12_0));
valve v_12_1289 (.fluid_in(k_12_1289), .fluid_out(k_11_644), .air_in(c_12_1));
valve v_12_1290 (.fluid_in(k_12_1290), .fluid_out(k_11_645), .air_in(c_12_0));
valve v_12_1291 (.fluid_in(k_12_1291), .fluid_out(k_11_645), .air_in(c_12_1));
valve v_12_1292 (.fluid_in(k_12_1292), .fluid_out(k_11_646), .air_in(c_12_0));
valve v_12_1293 (.fluid_in(k_12_1293), .fluid_out(k_11_646), .air_in(c_12_1));
valve v_12_1294 (.fluid_in(k_12_1294), .fluid_out(k_11_647), .air_in(c_12_0));
valve v_12_1295 (.fluid_in(k_12_1295), .fluid_out(k_11_647), .air_in(c_12_1));
valve v_12_1296 (.fluid_in(k_12_1296), .fluid_out(k_11_648), .air_in(c_12_0));
valve v_12_1297 (.fluid_in(k_12_1297), .fluid_out(k_11_648), .air_in(c_12_1));
valve v_12_1298 (.fluid_in(k_12_1298), .fluid_out(k_11_649), .air_in(c_12_0));
valve v_12_1299 (.fluid_in(k_12_1299), .fluid_out(k_11_649), .air_in(c_12_1));
valve v_12_1300 (.fluid_in(k_12_1300), .fluid_out(k_11_650), .air_in(c_12_0));
valve v_12_1301 (.fluid_in(k_12_1301), .fluid_out(k_11_650), .air_in(c_12_1));
valve v_12_1302 (.fluid_in(k_12_1302), .fluid_out(k_11_651), .air_in(c_12_0));
valve v_12_1303 (.fluid_in(k_12_1303), .fluid_out(k_11_651), .air_in(c_12_1));
valve v_12_1304 (.fluid_in(k_12_1304), .fluid_out(k_11_652), .air_in(c_12_0));
valve v_12_1305 (.fluid_in(k_12_1305), .fluid_out(k_11_652), .air_in(c_12_1));
valve v_12_1306 (.fluid_in(k_12_1306), .fluid_out(k_11_653), .air_in(c_12_0));
valve v_12_1307 (.fluid_in(k_12_1307), .fluid_out(k_11_653), .air_in(c_12_1));
valve v_12_1308 (.fluid_in(k_12_1308), .fluid_out(k_11_654), .air_in(c_12_0));
valve v_12_1309 (.fluid_in(k_12_1309), .fluid_out(k_11_654), .air_in(c_12_1));
valve v_12_1310 (.fluid_in(k_12_1310), .fluid_out(k_11_655), .air_in(c_12_0));
valve v_12_1311 (.fluid_in(k_12_1311), .fluid_out(k_11_655), .air_in(c_12_1));
valve v_12_1312 (.fluid_in(k_12_1312), .fluid_out(k_11_656), .air_in(c_12_0));
valve v_12_1313 (.fluid_in(k_12_1313), .fluid_out(k_11_656), .air_in(c_12_1));
valve v_12_1314 (.fluid_in(k_12_1314), .fluid_out(k_11_657), .air_in(c_12_0));
valve v_12_1315 (.fluid_in(k_12_1315), .fluid_out(k_11_657), .air_in(c_12_1));
valve v_12_1316 (.fluid_in(k_12_1316), .fluid_out(k_11_658), .air_in(c_12_0));
valve v_12_1317 (.fluid_in(k_12_1317), .fluid_out(k_11_658), .air_in(c_12_1));
valve v_12_1318 (.fluid_in(k_12_1318), .fluid_out(k_11_659), .air_in(c_12_0));
valve v_12_1319 (.fluid_in(k_12_1319), .fluid_out(k_11_659), .air_in(c_12_1));
valve v_12_1320 (.fluid_in(k_12_1320), .fluid_out(k_11_660), .air_in(c_12_0));
valve v_12_1321 (.fluid_in(k_12_1321), .fluid_out(k_11_660), .air_in(c_12_1));
valve v_12_1322 (.fluid_in(k_12_1322), .fluid_out(k_11_661), .air_in(c_12_0));
valve v_12_1323 (.fluid_in(k_12_1323), .fluid_out(k_11_661), .air_in(c_12_1));
valve v_12_1324 (.fluid_in(k_12_1324), .fluid_out(k_11_662), .air_in(c_12_0));
valve v_12_1325 (.fluid_in(k_12_1325), .fluid_out(k_11_662), .air_in(c_12_1));
valve v_12_1326 (.fluid_in(k_12_1326), .fluid_out(k_11_663), .air_in(c_12_0));
valve v_12_1327 (.fluid_in(k_12_1327), .fluid_out(k_11_663), .air_in(c_12_1));
valve v_12_1328 (.fluid_in(k_12_1328), .fluid_out(k_11_664), .air_in(c_12_0));
valve v_12_1329 (.fluid_in(k_12_1329), .fluid_out(k_11_664), .air_in(c_12_1));
valve v_12_1330 (.fluid_in(k_12_1330), .fluid_out(k_11_665), .air_in(c_12_0));
valve v_12_1331 (.fluid_in(k_12_1331), .fluid_out(k_11_665), .air_in(c_12_1));
valve v_12_1332 (.fluid_in(k_12_1332), .fluid_out(k_11_666), .air_in(c_12_0));
valve v_12_1333 (.fluid_in(k_12_1333), .fluid_out(k_11_666), .air_in(c_12_1));
valve v_12_1334 (.fluid_in(k_12_1334), .fluid_out(k_11_667), .air_in(c_12_0));
valve v_12_1335 (.fluid_in(k_12_1335), .fluid_out(k_11_667), .air_in(c_12_1));
valve v_12_1336 (.fluid_in(k_12_1336), .fluid_out(k_11_668), .air_in(c_12_0));
valve v_12_1337 (.fluid_in(k_12_1337), .fluid_out(k_11_668), .air_in(c_12_1));
valve v_12_1338 (.fluid_in(k_12_1338), .fluid_out(k_11_669), .air_in(c_12_0));
valve v_12_1339 (.fluid_in(k_12_1339), .fluid_out(k_11_669), .air_in(c_12_1));
valve v_12_1340 (.fluid_in(k_12_1340), .fluid_out(k_11_670), .air_in(c_12_0));
valve v_12_1341 (.fluid_in(k_12_1341), .fluid_out(k_11_670), .air_in(c_12_1));
valve v_12_1342 (.fluid_in(k_12_1342), .fluid_out(k_11_671), .air_in(c_12_0));
valve v_12_1343 (.fluid_in(k_12_1343), .fluid_out(k_11_671), .air_in(c_12_1));
valve v_12_1344 (.fluid_in(k_12_1344), .fluid_out(k_11_672), .air_in(c_12_0));
valve v_12_1345 (.fluid_in(k_12_1345), .fluid_out(k_11_672), .air_in(c_12_1));
valve v_12_1346 (.fluid_in(k_12_1346), .fluid_out(k_11_673), .air_in(c_12_0));
valve v_12_1347 (.fluid_in(k_12_1347), .fluid_out(k_11_673), .air_in(c_12_1));
valve v_12_1348 (.fluid_in(k_12_1348), .fluid_out(k_11_674), .air_in(c_12_0));
valve v_12_1349 (.fluid_in(k_12_1349), .fluid_out(k_11_674), .air_in(c_12_1));
valve v_12_1350 (.fluid_in(k_12_1350), .fluid_out(k_11_675), .air_in(c_12_0));
valve v_12_1351 (.fluid_in(k_12_1351), .fluid_out(k_11_675), .air_in(c_12_1));
valve v_12_1352 (.fluid_in(k_12_1352), .fluid_out(k_11_676), .air_in(c_12_0));
valve v_12_1353 (.fluid_in(k_12_1353), .fluid_out(k_11_676), .air_in(c_12_1));
valve v_12_1354 (.fluid_in(k_12_1354), .fluid_out(k_11_677), .air_in(c_12_0));
valve v_12_1355 (.fluid_in(k_12_1355), .fluid_out(k_11_677), .air_in(c_12_1));
valve v_12_1356 (.fluid_in(k_12_1356), .fluid_out(k_11_678), .air_in(c_12_0));
valve v_12_1357 (.fluid_in(k_12_1357), .fluid_out(k_11_678), .air_in(c_12_1));
valve v_12_1358 (.fluid_in(k_12_1358), .fluid_out(k_11_679), .air_in(c_12_0));
valve v_12_1359 (.fluid_in(k_12_1359), .fluid_out(k_11_679), .air_in(c_12_1));
valve v_12_1360 (.fluid_in(k_12_1360), .fluid_out(k_11_680), .air_in(c_12_0));
valve v_12_1361 (.fluid_in(k_12_1361), .fluid_out(k_11_680), .air_in(c_12_1));
valve v_12_1362 (.fluid_in(k_12_1362), .fluid_out(k_11_681), .air_in(c_12_0));
valve v_12_1363 (.fluid_in(k_12_1363), .fluid_out(k_11_681), .air_in(c_12_1));
valve v_12_1364 (.fluid_in(k_12_1364), .fluid_out(k_11_682), .air_in(c_12_0));
valve v_12_1365 (.fluid_in(k_12_1365), .fluid_out(k_11_682), .air_in(c_12_1));
valve v_12_1366 (.fluid_in(k_12_1366), .fluid_out(k_11_683), .air_in(c_12_0));
valve v_12_1367 (.fluid_in(k_12_1367), .fluid_out(k_11_683), .air_in(c_12_1));
valve v_12_1368 (.fluid_in(k_12_1368), .fluid_out(k_11_684), .air_in(c_12_0));
valve v_12_1369 (.fluid_in(k_12_1369), .fluid_out(k_11_684), .air_in(c_12_1));
valve v_12_1370 (.fluid_in(k_12_1370), .fluid_out(k_11_685), .air_in(c_12_0));
valve v_12_1371 (.fluid_in(k_12_1371), .fluid_out(k_11_685), .air_in(c_12_1));
valve v_12_1372 (.fluid_in(k_12_1372), .fluid_out(k_11_686), .air_in(c_12_0));
valve v_12_1373 (.fluid_in(k_12_1373), .fluid_out(k_11_686), .air_in(c_12_1));
valve v_12_1374 (.fluid_in(k_12_1374), .fluid_out(k_11_687), .air_in(c_12_0));
valve v_12_1375 (.fluid_in(k_12_1375), .fluid_out(k_11_687), .air_in(c_12_1));
valve v_12_1376 (.fluid_in(k_12_1376), .fluid_out(k_11_688), .air_in(c_12_0));
valve v_12_1377 (.fluid_in(k_12_1377), .fluid_out(k_11_688), .air_in(c_12_1));
valve v_12_1378 (.fluid_in(k_12_1378), .fluid_out(k_11_689), .air_in(c_12_0));
valve v_12_1379 (.fluid_in(k_12_1379), .fluid_out(k_11_689), .air_in(c_12_1));
valve v_12_1380 (.fluid_in(k_12_1380), .fluid_out(k_11_690), .air_in(c_12_0));
valve v_12_1381 (.fluid_in(k_12_1381), .fluid_out(k_11_690), .air_in(c_12_1));
valve v_12_1382 (.fluid_in(k_12_1382), .fluid_out(k_11_691), .air_in(c_12_0));
valve v_12_1383 (.fluid_in(k_12_1383), .fluid_out(k_11_691), .air_in(c_12_1));
valve v_12_1384 (.fluid_in(k_12_1384), .fluid_out(k_11_692), .air_in(c_12_0));
valve v_12_1385 (.fluid_in(k_12_1385), .fluid_out(k_11_692), .air_in(c_12_1));
valve v_12_1386 (.fluid_in(k_12_1386), .fluid_out(k_11_693), .air_in(c_12_0));
valve v_12_1387 (.fluid_in(k_12_1387), .fluid_out(k_11_693), .air_in(c_12_1));
valve v_12_1388 (.fluid_in(k_12_1388), .fluid_out(k_11_694), .air_in(c_12_0));
valve v_12_1389 (.fluid_in(k_12_1389), .fluid_out(k_11_694), .air_in(c_12_1));
valve v_12_1390 (.fluid_in(k_12_1390), .fluid_out(k_11_695), .air_in(c_12_0));
valve v_12_1391 (.fluid_in(k_12_1391), .fluid_out(k_11_695), .air_in(c_12_1));
valve v_12_1392 (.fluid_in(k_12_1392), .fluid_out(k_11_696), .air_in(c_12_0));
valve v_12_1393 (.fluid_in(k_12_1393), .fluid_out(k_11_696), .air_in(c_12_1));
valve v_12_1394 (.fluid_in(k_12_1394), .fluid_out(k_11_697), .air_in(c_12_0));
valve v_12_1395 (.fluid_in(k_12_1395), .fluid_out(k_11_697), .air_in(c_12_1));
valve v_12_1396 (.fluid_in(k_12_1396), .fluid_out(k_11_698), .air_in(c_12_0));
valve v_12_1397 (.fluid_in(k_12_1397), .fluid_out(k_11_698), .air_in(c_12_1));
valve v_12_1398 (.fluid_in(k_12_1398), .fluid_out(k_11_699), .air_in(c_12_0));
valve v_12_1399 (.fluid_in(k_12_1399), .fluid_out(k_11_699), .air_in(c_12_1));
valve v_12_1400 (.fluid_in(k_12_1400), .fluid_out(k_11_700), .air_in(c_12_0));
valve v_12_1401 (.fluid_in(k_12_1401), .fluid_out(k_11_700), .air_in(c_12_1));
valve v_12_1402 (.fluid_in(k_12_1402), .fluid_out(k_11_701), .air_in(c_12_0));
valve v_12_1403 (.fluid_in(k_12_1403), .fluid_out(k_11_701), .air_in(c_12_1));
valve v_12_1404 (.fluid_in(k_12_1404), .fluid_out(k_11_702), .air_in(c_12_0));
valve v_12_1405 (.fluid_in(k_12_1405), .fluid_out(k_11_702), .air_in(c_12_1));
valve v_12_1406 (.fluid_in(k_12_1406), .fluid_out(k_11_703), .air_in(c_12_0));
valve v_12_1407 (.fluid_in(k_12_1407), .fluid_out(k_11_703), .air_in(c_12_1));
valve v_12_1408 (.fluid_in(k_12_1408), .fluid_out(k_11_704), .air_in(c_12_0));
valve v_12_1409 (.fluid_in(k_12_1409), .fluid_out(k_11_704), .air_in(c_12_1));
valve v_12_1410 (.fluid_in(k_12_1410), .fluid_out(k_11_705), .air_in(c_12_0));
valve v_12_1411 (.fluid_in(k_12_1411), .fluid_out(k_11_705), .air_in(c_12_1));
valve v_12_1412 (.fluid_in(k_12_1412), .fluid_out(k_11_706), .air_in(c_12_0));
valve v_12_1413 (.fluid_in(k_12_1413), .fluid_out(k_11_706), .air_in(c_12_1));
valve v_12_1414 (.fluid_in(k_12_1414), .fluid_out(k_11_707), .air_in(c_12_0));
valve v_12_1415 (.fluid_in(k_12_1415), .fluid_out(k_11_707), .air_in(c_12_1));
valve v_12_1416 (.fluid_in(k_12_1416), .fluid_out(k_11_708), .air_in(c_12_0));
valve v_12_1417 (.fluid_in(k_12_1417), .fluid_out(k_11_708), .air_in(c_12_1));
valve v_12_1418 (.fluid_in(k_12_1418), .fluid_out(k_11_709), .air_in(c_12_0));
valve v_12_1419 (.fluid_in(k_12_1419), .fluid_out(k_11_709), .air_in(c_12_1));
valve v_12_1420 (.fluid_in(k_12_1420), .fluid_out(k_11_710), .air_in(c_12_0));
valve v_12_1421 (.fluid_in(k_12_1421), .fluid_out(k_11_710), .air_in(c_12_1));
valve v_12_1422 (.fluid_in(k_12_1422), .fluid_out(k_11_711), .air_in(c_12_0));
valve v_12_1423 (.fluid_in(k_12_1423), .fluid_out(k_11_711), .air_in(c_12_1));
valve v_12_1424 (.fluid_in(k_12_1424), .fluid_out(k_11_712), .air_in(c_12_0));
valve v_12_1425 (.fluid_in(k_12_1425), .fluid_out(k_11_712), .air_in(c_12_1));
valve v_12_1426 (.fluid_in(k_12_1426), .fluid_out(k_11_713), .air_in(c_12_0));
valve v_12_1427 (.fluid_in(k_12_1427), .fluid_out(k_11_713), .air_in(c_12_1));
valve v_12_1428 (.fluid_in(k_12_1428), .fluid_out(k_11_714), .air_in(c_12_0));
valve v_12_1429 (.fluid_in(k_12_1429), .fluid_out(k_11_714), .air_in(c_12_1));
valve v_12_1430 (.fluid_in(k_12_1430), .fluid_out(k_11_715), .air_in(c_12_0));
valve v_12_1431 (.fluid_in(k_12_1431), .fluid_out(k_11_715), .air_in(c_12_1));
valve v_12_1432 (.fluid_in(k_12_1432), .fluid_out(k_11_716), .air_in(c_12_0));
valve v_12_1433 (.fluid_in(k_12_1433), .fluid_out(k_11_716), .air_in(c_12_1));
valve v_12_1434 (.fluid_in(k_12_1434), .fluid_out(k_11_717), .air_in(c_12_0));
valve v_12_1435 (.fluid_in(k_12_1435), .fluid_out(k_11_717), .air_in(c_12_1));
valve v_12_1436 (.fluid_in(k_12_1436), .fluid_out(k_11_718), .air_in(c_12_0));
valve v_12_1437 (.fluid_in(k_12_1437), .fluid_out(k_11_718), .air_in(c_12_1));
valve v_12_1438 (.fluid_in(k_12_1438), .fluid_out(k_11_719), .air_in(c_12_0));
valve v_12_1439 (.fluid_in(k_12_1439), .fluid_out(k_11_719), .air_in(c_12_1));
valve v_12_1440 (.fluid_in(k_12_1440), .fluid_out(k_11_720), .air_in(c_12_0));
valve v_12_1441 (.fluid_in(k_12_1441), .fluid_out(k_11_720), .air_in(c_12_1));
valve v_12_1442 (.fluid_in(k_12_1442), .fluid_out(k_11_721), .air_in(c_12_0));
valve v_12_1443 (.fluid_in(k_12_1443), .fluid_out(k_11_721), .air_in(c_12_1));
valve v_12_1444 (.fluid_in(k_12_1444), .fluid_out(k_11_722), .air_in(c_12_0));
valve v_12_1445 (.fluid_in(k_12_1445), .fluid_out(k_11_722), .air_in(c_12_1));
valve v_12_1446 (.fluid_in(k_12_1446), .fluid_out(k_11_723), .air_in(c_12_0));
valve v_12_1447 (.fluid_in(k_12_1447), .fluid_out(k_11_723), .air_in(c_12_1));
valve v_12_1448 (.fluid_in(k_12_1448), .fluid_out(k_11_724), .air_in(c_12_0));
valve v_12_1449 (.fluid_in(k_12_1449), .fluid_out(k_11_724), .air_in(c_12_1));
valve v_12_1450 (.fluid_in(k_12_1450), .fluid_out(k_11_725), .air_in(c_12_0));
valve v_12_1451 (.fluid_in(k_12_1451), .fluid_out(k_11_725), .air_in(c_12_1));
valve v_12_1452 (.fluid_in(k_12_1452), .fluid_out(k_11_726), .air_in(c_12_0));
valve v_12_1453 (.fluid_in(k_12_1453), .fluid_out(k_11_726), .air_in(c_12_1));
valve v_12_1454 (.fluid_in(k_12_1454), .fluid_out(k_11_727), .air_in(c_12_0));
valve v_12_1455 (.fluid_in(k_12_1455), .fluid_out(k_11_727), .air_in(c_12_1));
valve v_12_1456 (.fluid_in(k_12_1456), .fluid_out(k_11_728), .air_in(c_12_0));
valve v_12_1457 (.fluid_in(k_12_1457), .fluid_out(k_11_728), .air_in(c_12_1));
valve v_12_1458 (.fluid_in(k_12_1458), .fluid_out(k_11_729), .air_in(c_12_0));
valve v_12_1459 (.fluid_in(k_12_1459), .fluid_out(k_11_729), .air_in(c_12_1));
valve v_12_1460 (.fluid_in(k_12_1460), .fluid_out(k_11_730), .air_in(c_12_0));
valve v_12_1461 (.fluid_in(k_12_1461), .fluid_out(k_11_730), .air_in(c_12_1));
valve v_12_1462 (.fluid_in(k_12_1462), .fluid_out(k_11_731), .air_in(c_12_0));
valve v_12_1463 (.fluid_in(k_12_1463), .fluid_out(k_11_731), .air_in(c_12_1));
valve v_12_1464 (.fluid_in(k_12_1464), .fluid_out(k_11_732), .air_in(c_12_0));
valve v_12_1465 (.fluid_in(k_12_1465), .fluid_out(k_11_732), .air_in(c_12_1));
valve v_12_1466 (.fluid_in(k_12_1466), .fluid_out(k_11_733), .air_in(c_12_0));
valve v_12_1467 (.fluid_in(k_12_1467), .fluid_out(k_11_733), .air_in(c_12_1));
valve v_12_1468 (.fluid_in(k_12_1468), .fluid_out(k_11_734), .air_in(c_12_0));
valve v_12_1469 (.fluid_in(k_12_1469), .fluid_out(k_11_734), .air_in(c_12_1));
valve v_12_1470 (.fluid_in(k_12_1470), .fluid_out(k_11_735), .air_in(c_12_0));
valve v_12_1471 (.fluid_in(k_12_1471), .fluid_out(k_11_735), .air_in(c_12_1));
valve v_12_1472 (.fluid_in(k_12_1472), .fluid_out(k_11_736), .air_in(c_12_0));
valve v_12_1473 (.fluid_in(k_12_1473), .fluid_out(k_11_736), .air_in(c_12_1));
valve v_12_1474 (.fluid_in(k_12_1474), .fluid_out(k_11_737), .air_in(c_12_0));
valve v_12_1475 (.fluid_in(k_12_1475), .fluid_out(k_11_737), .air_in(c_12_1));
valve v_12_1476 (.fluid_in(k_12_1476), .fluid_out(k_11_738), .air_in(c_12_0));
valve v_12_1477 (.fluid_in(k_12_1477), .fluid_out(k_11_738), .air_in(c_12_1));
valve v_12_1478 (.fluid_in(k_12_1478), .fluid_out(k_11_739), .air_in(c_12_0));
valve v_12_1479 (.fluid_in(k_12_1479), .fluid_out(k_11_739), .air_in(c_12_1));
valve v_12_1480 (.fluid_in(k_12_1480), .fluid_out(k_11_740), .air_in(c_12_0));
valve v_12_1481 (.fluid_in(k_12_1481), .fluid_out(k_11_740), .air_in(c_12_1));
valve v_12_1482 (.fluid_in(k_12_1482), .fluid_out(k_11_741), .air_in(c_12_0));
valve v_12_1483 (.fluid_in(k_12_1483), .fluid_out(k_11_741), .air_in(c_12_1));
valve v_12_1484 (.fluid_in(k_12_1484), .fluid_out(k_11_742), .air_in(c_12_0));
valve v_12_1485 (.fluid_in(k_12_1485), .fluid_out(k_11_742), .air_in(c_12_1));
valve v_12_1486 (.fluid_in(k_12_1486), .fluid_out(k_11_743), .air_in(c_12_0));
valve v_12_1487 (.fluid_in(k_12_1487), .fluid_out(k_11_743), .air_in(c_12_1));
valve v_12_1488 (.fluid_in(k_12_1488), .fluid_out(k_11_744), .air_in(c_12_0));
valve v_12_1489 (.fluid_in(k_12_1489), .fluid_out(k_11_744), .air_in(c_12_1));
valve v_12_1490 (.fluid_in(k_12_1490), .fluid_out(k_11_745), .air_in(c_12_0));
valve v_12_1491 (.fluid_in(k_12_1491), .fluid_out(k_11_745), .air_in(c_12_1));
valve v_12_1492 (.fluid_in(k_12_1492), .fluid_out(k_11_746), .air_in(c_12_0));
valve v_12_1493 (.fluid_in(k_12_1493), .fluid_out(k_11_746), .air_in(c_12_1));
valve v_12_1494 (.fluid_in(k_12_1494), .fluid_out(k_11_747), .air_in(c_12_0));
valve v_12_1495 (.fluid_in(k_12_1495), .fluid_out(k_11_747), .air_in(c_12_1));
valve v_12_1496 (.fluid_in(k_12_1496), .fluid_out(k_11_748), .air_in(c_12_0));
valve v_12_1497 (.fluid_in(k_12_1497), .fluid_out(k_11_748), .air_in(c_12_1));
valve v_12_1498 (.fluid_in(k_12_1498), .fluid_out(k_11_749), .air_in(c_12_0));
valve v_12_1499 (.fluid_in(k_12_1499), .fluid_out(k_11_749), .air_in(c_12_1));
valve v_12_1500 (.fluid_in(k_12_1500), .fluid_out(k_11_750), .air_in(c_12_0));
valve v_12_1501 (.fluid_in(k_12_1501), .fluid_out(k_11_750), .air_in(c_12_1));
valve v_12_1502 (.fluid_in(k_12_1502), .fluid_out(k_11_751), .air_in(c_12_0));
valve v_12_1503 (.fluid_in(k_12_1503), .fluid_out(k_11_751), .air_in(c_12_1));
valve v_12_1504 (.fluid_in(k_12_1504), .fluid_out(k_11_752), .air_in(c_12_0));
valve v_12_1505 (.fluid_in(k_12_1505), .fluid_out(k_11_752), .air_in(c_12_1));
valve v_12_1506 (.fluid_in(k_12_1506), .fluid_out(k_11_753), .air_in(c_12_0));
valve v_12_1507 (.fluid_in(k_12_1507), .fluid_out(k_11_753), .air_in(c_12_1));
valve v_12_1508 (.fluid_in(k_12_1508), .fluid_out(k_11_754), .air_in(c_12_0));
valve v_12_1509 (.fluid_in(k_12_1509), .fluid_out(k_11_754), .air_in(c_12_1));
valve v_12_1510 (.fluid_in(k_12_1510), .fluid_out(k_11_755), .air_in(c_12_0));
valve v_12_1511 (.fluid_in(k_12_1511), .fluid_out(k_11_755), .air_in(c_12_1));
valve v_12_1512 (.fluid_in(k_12_1512), .fluid_out(k_11_756), .air_in(c_12_0));
valve v_12_1513 (.fluid_in(k_12_1513), .fluid_out(k_11_756), .air_in(c_12_1));
valve v_12_1514 (.fluid_in(k_12_1514), .fluid_out(k_11_757), .air_in(c_12_0));
valve v_12_1515 (.fluid_in(k_12_1515), .fluid_out(k_11_757), .air_in(c_12_1));
valve v_12_1516 (.fluid_in(k_12_1516), .fluid_out(k_11_758), .air_in(c_12_0));
valve v_12_1517 (.fluid_in(k_12_1517), .fluid_out(k_11_758), .air_in(c_12_1));
valve v_12_1518 (.fluid_in(k_12_1518), .fluid_out(k_11_759), .air_in(c_12_0));
valve v_12_1519 (.fluid_in(k_12_1519), .fluid_out(k_11_759), .air_in(c_12_1));
valve v_12_1520 (.fluid_in(k_12_1520), .fluid_out(k_11_760), .air_in(c_12_0));
valve v_12_1521 (.fluid_in(k_12_1521), .fluid_out(k_11_760), .air_in(c_12_1));
valve v_12_1522 (.fluid_in(k_12_1522), .fluid_out(k_11_761), .air_in(c_12_0));
valve v_12_1523 (.fluid_in(k_12_1523), .fluid_out(k_11_761), .air_in(c_12_1));
valve v_12_1524 (.fluid_in(k_12_1524), .fluid_out(k_11_762), .air_in(c_12_0));
valve v_12_1525 (.fluid_in(k_12_1525), .fluid_out(k_11_762), .air_in(c_12_1));
valve v_12_1526 (.fluid_in(k_12_1526), .fluid_out(k_11_763), .air_in(c_12_0));
valve v_12_1527 (.fluid_in(k_12_1527), .fluid_out(k_11_763), .air_in(c_12_1));
valve v_12_1528 (.fluid_in(k_12_1528), .fluid_out(k_11_764), .air_in(c_12_0));
valve v_12_1529 (.fluid_in(k_12_1529), .fluid_out(k_11_764), .air_in(c_12_1));
valve v_12_1530 (.fluid_in(k_12_1530), .fluid_out(k_11_765), .air_in(c_12_0));
valve v_12_1531 (.fluid_in(k_12_1531), .fluid_out(k_11_765), .air_in(c_12_1));
valve v_12_1532 (.fluid_in(k_12_1532), .fluid_out(k_11_766), .air_in(c_12_0));
valve v_12_1533 (.fluid_in(k_12_1533), .fluid_out(k_11_766), .air_in(c_12_1));
valve v_12_1534 (.fluid_in(k_12_1534), .fluid_out(k_11_767), .air_in(c_12_0));
valve v_12_1535 (.fluid_in(k_12_1535), .fluid_out(k_11_767), .air_in(c_12_1));
valve v_12_1536 (.fluid_in(k_12_1536), .fluid_out(k_11_768), .air_in(c_12_0));
valve v_12_1537 (.fluid_in(k_12_1537), .fluid_out(k_11_768), .air_in(c_12_1));
valve v_12_1538 (.fluid_in(k_12_1538), .fluid_out(k_11_769), .air_in(c_12_0));
valve v_12_1539 (.fluid_in(k_12_1539), .fluid_out(k_11_769), .air_in(c_12_1));
valve v_12_1540 (.fluid_in(k_12_1540), .fluid_out(k_11_770), .air_in(c_12_0));
valve v_12_1541 (.fluid_in(k_12_1541), .fluid_out(k_11_770), .air_in(c_12_1));
valve v_12_1542 (.fluid_in(k_12_1542), .fluid_out(k_11_771), .air_in(c_12_0));
valve v_12_1543 (.fluid_in(k_12_1543), .fluid_out(k_11_771), .air_in(c_12_1));
valve v_12_1544 (.fluid_in(k_12_1544), .fluid_out(k_11_772), .air_in(c_12_0));
valve v_12_1545 (.fluid_in(k_12_1545), .fluid_out(k_11_772), .air_in(c_12_1));
valve v_12_1546 (.fluid_in(k_12_1546), .fluid_out(k_11_773), .air_in(c_12_0));
valve v_12_1547 (.fluid_in(k_12_1547), .fluid_out(k_11_773), .air_in(c_12_1));
valve v_12_1548 (.fluid_in(k_12_1548), .fluid_out(k_11_774), .air_in(c_12_0));
valve v_12_1549 (.fluid_in(k_12_1549), .fluid_out(k_11_774), .air_in(c_12_1));
valve v_12_1550 (.fluid_in(k_12_1550), .fluid_out(k_11_775), .air_in(c_12_0));
valve v_12_1551 (.fluid_in(k_12_1551), .fluid_out(k_11_775), .air_in(c_12_1));
valve v_12_1552 (.fluid_in(k_12_1552), .fluid_out(k_11_776), .air_in(c_12_0));
valve v_12_1553 (.fluid_in(k_12_1553), .fluid_out(k_11_776), .air_in(c_12_1));
valve v_12_1554 (.fluid_in(k_12_1554), .fluid_out(k_11_777), .air_in(c_12_0));
valve v_12_1555 (.fluid_in(k_12_1555), .fluid_out(k_11_777), .air_in(c_12_1));
valve v_12_1556 (.fluid_in(k_12_1556), .fluid_out(k_11_778), .air_in(c_12_0));
valve v_12_1557 (.fluid_in(k_12_1557), .fluid_out(k_11_778), .air_in(c_12_1));
valve v_12_1558 (.fluid_in(k_12_1558), .fluid_out(k_11_779), .air_in(c_12_0));
valve v_12_1559 (.fluid_in(k_12_1559), .fluid_out(k_11_779), .air_in(c_12_1));
valve v_12_1560 (.fluid_in(k_12_1560), .fluid_out(k_11_780), .air_in(c_12_0));
valve v_12_1561 (.fluid_in(k_12_1561), .fluid_out(k_11_780), .air_in(c_12_1));
valve v_12_1562 (.fluid_in(k_12_1562), .fluid_out(k_11_781), .air_in(c_12_0));
valve v_12_1563 (.fluid_in(k_12_1563), .fluid_out(k_11_781), .air_in(c_12_1));
valve v_12_1564 (.fluid_in(k_12_1564), .fluid_out(k_11_782), .air_in(c_12_0));
valve v_12_1565 (.fluid_in(k_12_1565), .fluid_out(k_11_782), .air_in(c_12_1));
valve v_12_1566 (.fluid_in(k_12_1566), .fluid_out(k_11_783), .air_in(c_12_0));
valve v_12_1567 (.fluid_in(k_12_1567), .fluid_out(k_11_783), .air_in(c_12_1));
valve v_12_1568 (.fluid_in(k_12_1568), .fluid_out(k_11_784), .air_in(c_12_0));
valve v_12_1569 (.fluid_in(k_12_1569), .fluid_out(k_11_784), .air_in(c_12_1));
valve v_12_1570 (.fluid_in(k_12_1570), .fluid_out(k_11_785), .air_in(c_12_0));
valve v_12_1571 (.fluid_in(k_12_1571), .fluid_out(k_11_785), .air_in(c_12_1));
valve v_12_1572 (.fluid_in(k_12_1572), .fluid_out(k_11_786), .air_in(c_12_0));
valve v_12_1573 (.fluid_in(k_12_1573), .fluid_out(k_11_786), .air_in(c_12_1));
valve v_12_1574 (.fluid_in(k_12_1574), .fluid_out(k_11_787), .air_in(c_12_0));
valve v_12_1575 (.fluid_in(k_12_1575), .fluid_out(k_11_787), .air_in(c_12_1));
valve v_12_1576 (.fluid_in(k_12_1576), .fluid_out(k_11_788), .air_in(c_12_0));
valve v_12_1577 (.fluid_in(k_12_1577), .fluid_out(k_11_788), .air_in(c_12_1));
valve v_12_1578 (.fluid_in(k_12_1578), .fluid_out(k_11_789), .air_in(c_12_0));
valve v_12_1579 (.fluid_in(k_12_1579), .fluid_out(k_11_789), .air_in(c_12_1));
valve v_12_1580 (.fluid_in(k_12_1580), .fluid_out(k_11_790), .air_in(c_12_0));
valve v_12_1581 (.fluid_in(k_12_1581), .fluid_out(k_11_790), .air_in(c_12_1));
valve v_12_1582 (.fluid_in(k_12_1582), .fluid_out(k_11_791), .air_in(c_12_0));
valve v_12_1583 (.fluid_in(k_12_1583), .fluid_out(k_11_791), .air_in(c_12_1));
valve v_12_1584 (.fluid_in(k_12_1584), .fluid_out(k_11_792), .air_in(c_12_0));
valve v_12_1585 (.fluid_in(k_12_1585), .fluid_out(k_11_792), .air_in(c_12_1));
valve v_12_1586 (.fluid_in(k_12_1586), .fluid_out(k_11_793), .air_in(c_12_0));
valve v_12_1587 (.fluid_in(k_12_1587), .fluid_out(k_11_793), .air_in(c_12_1));
valve v_12_1588 (.fluid_in(k_12_1588), .fluid_out(k_11_794), .air_in(c_12_0));
valve v_12_1589 (.fluid_in(k_12_1589), .fluid_out(k_11_794), .air_in(c_12_1));
valve v_12_1590 (.fluid_in(k_12_1590), .fluid_out(k_11_795), .air_in(c_12_0));
valve v_12_1591 (.fluid_in(k_12_1591), .fluid_out(k_11_795), .air_in(c_12_1));
valve v_12_1592 (.fluid_in(k_12_1592), .fluid_out(k_11_796), .air_in(c_12_0));
valve v_12_1593 (.fluid_in(k_12_1593), .fluid_out(k_11_796), .air_in(c_12_1));
valve v_12_1594 (.fluid_in(k_12_1594), .fluid_out(k_11_797), .air_in(c_12_0));
valve v_12_1595 (.fluid_in(k_12_1595), .fluid_out(k_11_797), .air_in(c_12_1));
valve v_12_1596 (.fluid_in(k_12_1596), .fluid_out(k_11_798), .air_in(c_12_0));
valve v_12_1597 (.fluid_in(k_12_1597), .fluid_out(k_11_798), .air_in(c_12_1));
valve v_12_1598 (.fluid_in(k_12_1598), .fluid_out(k_11_799), .air_in(c_12_0));
valve v_12_1599 (.fluid_in(k_12_1599), .fluid_out(k_11_799), .air_in(c_12_1));
valve v_12_1600 (.fluid_in(k_12_1600), .fluid_out(k_11_800), .air_in(c_12_0));
valve v_12_1601 (.fluid_in(k_12_1601), .fluid_out(k_11_800), .air_in(c_12_1));
valve v_12_1602 (.fluid_in(k_12_1602), .fluid_out(k_11_801), .air_in(c_12_0));
valve v_12_1603 (.fluid_in(k_12_1603), .fluid_out(k_11_801), .air_in(c_12_1));
valve v_12_1604 (.fluid_in(k_12_1604), .fluid_out(k_11_802), .air_in(c_12_0));
valve v_12_1605 (.fluid_in(k_12_1605), .fluid_out(k_11_802), .air_in(c_12_1));
valve v_12_1606 (.fluid_in(k_12_1606), .fluid_out(k_11_803), .air_in(c_12_0));
valve v_12_1607 (.fluid_in(k_12_1607), .fluid_out(k_11_803), .air_in(c_12_1));
valve v_12_1608 (.fluid_in(k_12_1608), .fluid_out(k_11_804), .air_in(c_12_0));
valve v_12_1609 (.fluid_in(k_12_1609), .fluid_out(k_11_804), .air_in(c_12_1));
valve v_12_1610 (.fluid_in(k_12_1610), .fluid_out(k_11_805), .air_in(c_12_0));
valve v_12_1611 (.fluid_in(k_12_1611), .fluid_out(k_11_805), .air_in(c_12_1));
valve v_12_1612 (.fluid_in(k_12_1612), .fluid_out(k_11_806), .air_in(c_12_0));
valve v_12_1613 (.fluid_in(k_12_1613), .fluid_out(k_11_806), .air_in(c_12_1));
valve v_12_1614 (.fluid_in(k_12_1614), .fluid_out(k_11_807), .air_in(c_12_0));
valve v_12_1615 (.fluid_in(k_12_1615), .fluid_out(k_11_807), .air_in(c_12_1));
valve v_12_1616 (.fluid_in(k_12_1616), .fluid_out(k_11_808), .air_in(c_12_0));
valve v_12_1617 (.fluid_in(k_12_1617), .fluid_out(k_11_808), .air_in(c_12_1));
valve v_12_1618 (.fluid_in(k_12_1618), .fluid_out(k_11_809), .air_in(c_12_0));
valve v_12_1619 (.fluid_in(k_12_1619), .fluid_out(k_11_809), .air_in(c_12_1));
valve v_12_1620 (.fluid_in(k_12_1620), .fluid_out(k_11_810), .air_in(c_12_0));
valve v_12_1621 (.fluid_in(k_12_1621), .fluid_out(k_11_810), .air_in(c_12_1));
valve v_12_1622 (.fluid_in(k_12_1622), .fluid_out(k_11_811), .air_in(c_12_0));
valve v_12_1623 (.fluid_in(k_12_1623), .fluid_out(k_11_811), .air_in(c_12_1));
valve v_12_1624 (.fluid_in(k_12_1624), .fluid_out(k_11_812), .air_in(c_12_0));
valve v_12_1625 (.fluid_in(k_12_1625), .fluid_out(k_11_812), .air_in(c_12_1));
valve v_12_1626 (.fluid_in(k_12_1626), .fluid_out(k_11_813), .air_in(c_12_0));
valve v_12_1627 (.fluid_in(k_12_1627), .fluid_out(k_11_813), .air_in(c_12_1));
valve v_12_1628 (.fluid_in(k_12_1628), .fluid_out(k_11_814), .air_in(c_12_0));
valve v_12_1629 (.fluid_in(k_12_1629), .fluid_out(k_11_814), .air_in(c_12_1));
valve v_12_1630 (.fluid_in(k_12_1630), .fluid_out(k_11_815), .air_in(c_12_0));
valve v_12_1631 (.fluid_in(k_12_1631), .fluid_out(k_11_815), .air_in(c_12_1));
valve v_12_1632 (.fluid_in(k_12_1632), .fluid_out(k_11_816), .air_in(c_12_0));
valve v_12_1633 (.fluid_in(k_12_1633), .fluid_out(k_11_816), .air_in(c_12_1));
valve v_12_1634 (.fluid_in(k_12_1634), .fluid_out(k_11_817), .air_in(c_12_0));
valve v_12_1635 (.fluid_in(k_12_1635), .fluid_out(k_11_817), .air_in(c_12_1));
valve v_12_1636 (.fluid_in(k_12_1636), .fluid_out(k_11_818), .air_in(c_12_0));
valve v_12_1637 (.fluid_in(k_12_1637), .fluid_out(k_11_818), .air_in(c_12_1));
valve v_12_1638 (.fluid_in(k_12_1638), .fluid_out(k_11_819), .air_in(c_12_0));
valve v_12_1639 (.fluid_in(k_12_1639), .fluid_out(k_11_819), .air_in(c_12_1));
valve v_12_1640 (.fluid_in(k_12_1640), .fluid_out(k_11_820), .air_in(c_12_0));
valve v_12_1641 (.fluid_in(k_12_1641), .fluid_out(k_11_820), .air_in(c_12_1));
valve v_12_1642 (.fluid_in(k_12_1642), .fluid_out(k_11_821), .air_in(c_12_0));
valve v_12_1643 (.fluid_in(k_12_1643), .fluid_out(k_11_821), .air_in(c_12_1));
valve v_12_1644 (.fluid_in(k_12_1644), .fluid_out(k_11_822), .air_in(c_12_0));
valve v_12_1645 (.fluid_in(k_12_1645), .fluid_out(k_11_822), .air_in(c_12_1));
valve v_12_1646 (.fluid_in(k_12_1646), .fluid_out(k_11_823), .air_in(c_12_0));
valve v_12_1647 (.fluid_in(k_12_1647), .fluid_out(k_11_823), .air_in(c_12_1));
valve v_12_1648 (.fluid_in(k_12_1648), .fluid_out(k_11_824), .air_in(c_12_0));
valve v_12_1649 (.fluid_in(k_12_1649), .fluid_out(k_11_824), .air_in(c_12_1));
valve v_12_1650 (.fluid_in(k_12_1650), .fluid_out(k_11_825), .air_in(c_12_0));
valve v_12_1651 (.fluid_in(k_12_1651), .fluid_out(k_11_825), .air_in(c_12_1));
valve v_12_1652 (.fluid_in(k_12_1652), .fluid_out(k_11_826), .air_in(c_12_0));
valve v_12_1653 (.fluid_in(k_12_1653), .fluid_out(k_11_826), .air_in(c_12_1));
valve v_12_1654 (.fluid_in(k_12_1654), .fluid_out(k_11_827), .air_in(c_12_0));
valve v_12_1655 (.fluid_in(k_12_1655), .fluid_out(k_11_827), .air_in(c_12_1));
valve v_12_1656 (.fluid_in(k_12_1656), .fluid_out(k_11_828), .air_in(c_12_0));
valve v_12_1657 (.fluid_in(k_12_1657), .fluid_out(k_11_828), .air_in(c_12_1));
valve v_12_1658 (.fluid_in(k_12_1658), .fluid_out(k_11_829), .air_in(c_12_0));
valve v_12_1659 (.fluid_in(k_12_1659), .fluid_out(k_11_829), .air_in(c_12_1));
valve v_12_1660 (.fluid_in(k_12_1660), .fluid_out(k_11_830), .air_in(c_12_0));
valve v_12_1661 (.fluid_in(k_12_1661), .fluid_out(k_11_830), .air_in(c_12_1));
valve v_12_1662 (.fluid_in(k_12_1662), .fluid_out(k_11_831), .air_in(c_12_0));
valve v_12_1663 (.fluid_in(k_12_1663), .fluid_out(k_11_831), .air_in(c_12_1));
valve v_12_1664 (.fluid_in(k_12_1664), .fluid_out(k_11_832), .air_in(c_12_0));
valve v_12_1665 (.fluid_in(k_12_1665), .fluid_out(k_11_832), .air_in(c_12_1));
valve v_12_1666 (.fluid_in(k_12_1666), .fluid_out(k_11_833), .air_in(c_12_0));
valve v_12_1667 (.fluid_in(k_12_1667), .fluid_out(k_11_833), .air_in(c_12_1));
valve v_12_1668 (.fluid_in(k_12_1668), .fluid_out(k_11_834), .air_in(c_12_0));
valve v_12_1669 (.fluid_in(k_12_1669), .fluid_out(k_11_834), .air_in(c_12_1));
valve v_12_1670 (.fluid_in(k_12_1670), .fluid_out(k_11_835), .air_in(c_12_0));
valve v_12_1671 (.fluid_in(k_12_1671), .fluid_out(k_11_835), .air_in(c_12_1));
valve v_12_1672 (.fluid_in(k_12_1672), .fluid_out(k_11_836), .air_in(c_12_0));
valve v_12_1673 (.fluid_in(k_12_1673), .fluid_out(k_11_836), .air_in(c_12_1));
valve v_12_1674 (.fluid_in(k_12_1674), .fluid_out(k_11_837), .air_in(c_12_0));
valve v_12_1675 (.fluid_in(k_12_1675), .fluid_out(k_11_837), .air_in(c_12_1));
valve v_12_1676 (.fluid_in(k_12_1676), .fluid_out(k_11_838), .air_in(c_12_0));
valve v_12_1677 (.fluid_in(k_12_1677), .fluid_out(k_11_838), .air_in(c_12_1));
valve v_12_1678 (.fluid_in(k_12_1678), .fluid_out(k_11_839), .air_in(c_12_0));
valve v_12_1679 (.fluid_in(k_12_1679), .fluid_out(k_11_839), .air_in(c_12_1));
valve v_12_1680 (.fluid_in(k_12_1680), .fluid_out(k_11_840), .air_in(c_12_0));
valve v_12_1681 (.fluid_in(k_12_1681), .fluid_out(k_11_840), .air_in(c_12_1));
valve v_12_1682 (.fluid_in(k_12_1682), .fluid_out(k_11_841), .air_in(c_12_0));
valve v_12_1683 (.fluid_in(k_12_1683), .fluid_out(k_11_841), .air_in(c_12_1));
valve v_12_1684 (.fluid_in(k_12_1684), .fluid_out(k_11_842), .air_in(c_12_0));
valve v_12_1685 (.fluid_in(k_12_1685), .fluid_out(k_11_842), .air_in(c_12_1));
valve v_12_1686 (.fluid_in(k_12_1686), .fluid_out(k_11_843), .air_in(c_12_0));
valve v_12_1687 (.fluid_in(k_12_1687), .fluid_out(k_11_843), .air_in(c_12_1));
valve v_12_1688 (.fluid_in(k_12_1688), .fluid_out(k_11_844), .air_in(c_12_0));
valve v_12_1689 (.fluid_in(k_12_1689), .fluid_out(k_11_844), .air_in(c_12_1));
valve v_12_1690 (.fluid_in(k_12_1690), .fluid_out(k_11_845), .air_in(c_12_0));
valve v_12_1691 (.fluid_in(k_12_1691), .fluid_out(k_11_845), .air_in(c_12_1));
valve v_12_1692 (.fluid_in(k_12_1692), .fluid_out(k_11_846), .air_in(c_12_0));
valve v_12_1693 (.fluid_in(k_12_1693), .fluid_out(k_11_846), .air_in(c_12_1));
valve v_12_1694 (.fluid_in(k_12_1694), .fluid_out(k_11_847), .air_in(c_12_0));
valve v_12_1695 (.fluid_in(k_12_1695), .fluid_out(k_11_847), .air_in(c_12_1));
valve v_12_1696 (.fluid_in(k_12_1696), .fluid_out(k_11_848), .air_in(c_12_0));
valve v_12_1697 (.fluid_in(k_12_1697), .fluid_out(k_11_848), .air_in(c_12_1));
valve v_12_1698 (.fluid_in(k_12_1698), .fluid_out(k_11_849), .air_in(c_12_0));
valve v_12_1699 (.fluid_in(k_12_1699), .fluid_out(k_11_849), .air_in(c_12_1));
valve v_12_1700 (.fluid_in(k_12_1700), .fluid_out(k_11_850), .air_in(c_12_0));
valve v_12_1701 (.fluid_in(k_12_1701), .fluid_out(k_11_850), .air_in(c_12_1));
valve v_12_1702 (.fluid_in(k_12_1702), .fluid_out(k_11_851), .air_in(c_12_0));
valve v_12_1703 (.fluid_in(k_12_1703), .fluid_out(k_11_851), .air_in(c_12_1));
valve v_12_1704 (.fluid_in(k_12_1704), .fluid_out(k_11_852), .air_in(c_12_0));
valve v_12_1705 (.fluid_in(k_12_1705), .fluid_out(k_11_852), .air_in(c_12_1));
valve v_12_1706 (.fluid_in(k_12_1706), .fluid_out(k_11_853), .air_in(c_12_0));
valve v_12_1707 (.fluid_in(k_12_1707), .fluid_out(k_11_853), .air_in(c_12_1));
valve v_12_1708 (.fluid_in(k_12_1708), .fluid_out(k_11_854), .air_in(c_12_0));
valve v_12_1709 (.fluid_in(k_12_1709), .fluid_out(k_11_854), .air_in(c_12_1));
valve v_12_1710 (.fluid_in(k_12_1710), .fluid_out(k_11_855), .air_in(c_12_0));
valve v_12_1711 (.fluid_in(k_12_1711), .fluid_out(k_11_855), .air_in(c_12_1));
valve v_12_1712 (.fluid_in(k_12_1712), .fluid_out(k_11_856), .air_in(c_12_0));
valve v_12_1713 (.fluid_in(k_12_1713), .fluid_out(k_11_856), .air_in(c_12_1));
valve v_12_1714 (.fluid_in(k_12_1714), .fluid_out(k_11_857), .air_in(c_12_0));
valve v_12_1715 (.fluid_in(k_12_1715), .fluid_out(k_11_857), .air_in(c_12_1));
valve v_12_1716 (.fluid_in(k_12_1716), .fluid_out(k_11_858), .air_in(c_12_0));
valve v_12_1717 (.fluid_in(k_12_1717), .fluid_out(k_11_858), .air_in(c_12_1));
valve v_12_1718 (.fluid_in(k_12_1718), .fluid_out(k_11_859), .air_in(c_12_0));
valve v_12_1719 (.fluid_in(k_12_1719), .fluid_out(k_11_859), .air_in(c_12_1));
valve v_12_1720 (.fluid_in(k_12_1720), .fluid_out(k_11_860), .air_in(c_12_0));
valve v_12_1721 (.fluid_in(k_12_1721), .fluid_out(k_11_860), .air_in(c_12_1));
valve v_12_1722 (.fluid_in(k_12_1722), .fluid_out(k_11_861), .air_in(c_12_0));
valve v_12_1723 (.fluid_in(k_12_1723), .fluid_out(k_11_861), .air_in(c_12_1));
valve v_12_1724 (.fluid_in(k_12_1724), .fluid_out(k_11_862), .air_in(c_12_0));
valve v_12_1725 (.fluid_in(k_12_1725), .fluid_out(k_11_862), .air_in(c_12_1));
valve v_12_1726 (.fluid_in(k_12_1726), .fluid_out(k_11_863), .air_in(c_12_0));
valve v_12_1727 (.fluid_in(k_12_1727), .fluid_out(k_11_863), .air_in(c_12_1));
valve v_12_1728 (.fluid_in(k_12_1728), .fluid_out(k_11_864), .air_in(c_12_0));
valve v_12_1729 (.fluid_in(k_12_1729), .fluid_out(k_11_864), .air_in(c_12_1));
valve v_12_1730 (.fluid_in(k_12_1730), .fluid_out(k_11_865), .air_in(c_12_0));
valve v_12_1731 (.fluid_in(k_12_1731), .fluid_out(k_11_865), .air_in(c_12_1));
valve v_12_1732 (.fluid_in(k_12_1732), .fluid_out(k_11_866), .air_in(c_12_0));
valve v_12_1733 (.fluid_in(k_12_1733), .fluid_out(k_11_866), .air_in(c_12_1));
valve v_12_1734 (.fluid_in(k_12_1734), .fluid_out(k_11_867), .air_in(c_12_0));
valve v_12_1735 (.fluid_in(k_12_1735), .fluid_out(k_11_867), .air_in(c_12_1));
valve v_12_1736 (.fluid_in(k_12_1736), .fluid_out(k_11_868), .air_in(c_12_0));
valve v_12_1737 (.fluid_in(k_12_1737), .fluid_out(k_11_868), .air_in(c_12_1));
valve v_12_1738 (.fluid_in(k_12_1738), .fluid_out(k_11_869), .air_in(c_12_0));
valve v_12_1739 (.fluid_in(k_12_1739), .fluid_out(k_11_869), .air_in(c_12_1));
valve v_12_1740 (.fluid_in(k_12_1740), .fluid_out(k_11_870), .air_in(c_12_0));
valve v_12_1741 (.fluid_in(k_12_1741), .fluid_out(k_11_870), .air_in(c_12_1));
valve v_12_1742 (.fluid_in(k_12_1742), .fluid_out(k_11_871), .air_in(c_12_0));
valve v_12_1743 (.fluid_in(k_12_1743), .fluid_out(k_11_871), .air_in(c_12_1));
valve v_12_1744 (.fluid_in(k_12_1744), .fluid_out(k_11_872), .air_in(c_12_0));
valve v_12_1745 (.fluid_in(k_12_1745), .fluid_out(k_11_872), .air_in(c_12_1));
valve v_12_1746 (.fluid_in(k_12_1746), .fluid_out(k_11_873), .air_in(c_12_0));
valve v_12_1747 (.fluid_in(k_12_1747), .fluid_out(k_11_873), .air_in(c_12_1));
valve v_12_1748 (.fluid_in(k_12_1748), .fluid_out(k_11_874), .air_in(c_12_0));
valve v_12_1749 (.fluid_in(k_12_1749), .fluid_out(k_11_874), .air_in(c_12_1));
valve v_12_1750 (.fluid_in(k_12_1750), .fluid_out(k_11_875), .air_in(c_12_0));
valve v_12_1751 (.fluid_in(k_12_1751), .fluid_out(k_11_875), .air_in(c_12_1));
valve v_12_1752 (.fluid_in(k_12_1752), .fluid_out(k_11_876), .air_in(c_12_0));
valve v_12_1753 (.fluid_in(k_12_1753), .fluid_out(k_11_876), .air_in(c_12_1));
valve v_12_1754 (.fluid_in(k_12_1754), .fluid_out(k_11_877), .air_in(c_12_0));
valve v_12_1755 (.fluid_in(k_12_1755), .fluid_out(k_11_877), .air_in(c_12_1));
valve v_12_1756 (.fluid_in(k_12_1756), .fluid_out(k_11_878), .air_in(c_12_0));
valve v_12_1757 (.fluid_in(k_12_1757), .fluid_out(k_11_878), .air_in(c_12_1));
valve v_12_1758 (.fluid_in(k_12_1758), .fluid_out(k_11_879), .air_in(c_12_0));
valve v_12_1759 (.fluid_in(k_12_1759), .fluid_out(k_11_879), .air_in(c_12_1));
valve v_12_1760 (.fluid_in(k_12_1760), .fluid_out(k_11_880), .air_in(c_12_0));
valve v_12_1761 (.fluid_in(k_12_1761), .fluid_out(k_11_880), .air_in(c_12_1));
valve v_12_1762 (.fluid_in(k_12_1762), .fluid_out(k_11_881), .air_in(c_12_0));
valve v_12_1763 (.fluid_in(k_12_1763), .fluid_out(k_11_881), .air_in(c_12_1));
valve v_12_1764 (.fluid_in(k_12_1764), .fluid_out(k_11_882), .air_in(c_12_0));
valve v_12_1765 (.fluid_in(k_12_1765), .fluid_out(k_11_882), .air_in(c_12_1));
valve v_12_1766 (.fluid_in(k_12_1766), .fluid_out(k_11_883), .air_in(c_12_0));
valve v_12_1767 (.fluid_in(k_12_1767), .fluid_out(k_11_883), .air_in(c_12_1));
valve v_12_1768 (.fluid_in(k_12_1768), .fluid_out(k_11_884), .air_in(c_12_0));
valve v_12_1769 (.fluid_in(k_12_1769), .fluid_out(k_11_884), .air_in(c_12_1));
valve v_12_1770 (.fluid_in(k_12_1770), .fluid_out(k_11_885), .air_in(c_12_0));
valve v_12_1771 (.fluid_in(k_12_1771), .fluid_out(k_11_885), .air_in(c_12_1));
valve v_12_1772 (.fluid_in(k_12_1772), .fluid_out(k_11_886), .air_in(c_12_0));
valve v_12_1773 (.fluid_in(k_12_1773), .fluid_out(k_11_886), .air_in(c_12_1));
valve v_12_1774 (.fluid_in(k_12_1774), .fluid_out(k_11_887), .air_in(c_12_0));
valve v_12_1775 (.fluid_in(k_12_1775), .fluid_out(k_11_887), .air_in(c_12_1));
valve v_12_1776 (.fluid_in(k_12_1776), .fluid_out(k_11_888), .air_in(c_12_0));
valve v_12_1777 (.fluid_in(k_12_1777), .fluid_out(k_11_888), .air_in(c_12_1));
valve v_12_1778 (.fluid_in(k_12_1778), .fluid_out(k_11_889), .air_in(c_12_0));
valve v_12_1779 (.fluid_in(k_12_1779), .fluid_out(k_11_889), .air_in(c_12_1));
valve v_12_1780 (.fluid_in(k_12_1780), .fluid_out(k_11_890), .air_in(c_12_0));
valve v_12_1781 (.fluid_in(k_12_1781), .fluid_out(k_11_890), .air_in(c_12_1));
valve v_12_1782 (.fluid_in(k_12_1782), .fluid_out(k_11_891), .air_in(c_12_0));
valve v_12_1783 (.fluid_in(k_12_1783), .fluid_out(k_11_891), .air_in(c_12_1));
valve v_12_1784 (.fluid_in(k_12_1784), .fluid_out(k_11_892), .air_in(c_12_0));
valve v_12_1785 (.fluid_in(k_12_1785), .fluid_out(k_11_892), .air_in(c_12_1));
valve v_12_1786 (.fluid_in(k_12_1786), .fluid_out(k_11_893), .air_in(c_12_0));
valve v_12_1787 (.fluid_in(k_12_1787), .fluid_out(k_11_893), .air_in(c_12_1));
valve v_12_1788 (.fluid_in(k_12_1788), .fluid_out(k_11_894), .air_in(c_12_0));
valve v_12_1789 (.fluid_in(k_12_1789), .fluid_out(k_11_894), .air_in(c_12_1));
valve v_12_1790 (.fluid_in(k_12_1790), .fluid_out(k_11_895), .air_in(c_12_0));
valve v_12_1791 (.fluid_in(k_12_1791), .fluid_out(k_11_895), .air_in(c_12_1));
valve v_12_1792 (.fluid_in(k_12_1792), .fluid_out(k_11_896), .air_in(c_12_0));
valve v_12_1793 (.fluid_in(k_12_1793), .fluid_out(k_11_896), .air_in(c_12_1));
valve v_12_1794 (.fluid_in(k_12_1794), .fluid_out(k_11_897), .air_in(c_12_0));
valve v_12_1795 (.fluid_in(k_12_1795), .fluid_out(k_11_897), .air_in(c_12_1));
valve v_12_1796 (.fluid_in(k_12_1796), .fluid_out(k_11_898), .air_in(c_12_0));
valve v_12_1797 (.fluid_in(k_12_1797), .fluid_out(k_11_898), .air_in(c_12_1));
valve v_12_1798 (.fluid_in(k_12_1798), .fluid_out(k_11_899), .air_in(c_12_0));
valve v_12_1799 (.fluid_in(k_12_1799), .fluid_out(k_11_899), .air_in(c_12_1));
valve v_12_1800 (.fluid_in(k_12_1800), .fluid_out(k_11_900), .air_in(c_12_0));
valve v_12_1801 (.fluid_in(k_12_1801), .fluid_out(k_11_900), .air_in(c_12_1));
valve v_12_1802 (.fluid_in(k_12_1802), .fluid_out(k_11_901), .air_in(c_12_0));
valve v_12_1803 (.fluid_in(k_12_1803), .fluid_out(k_11_901), .air_in(c_12_1));
valve v_12_1804 (.fluid_in(k_12_1804), .fluid_out(k_11_902), .air_in(c_12_0));
valve v_12_1805 (.fluid_in(k_12_1805), .fluid_out(k_11_902), .air_in(c_12_1));
valve v_12_1806 (.fluid_in(k_12_1806), .fluid_out(k_11_903), .air_in(c_12_0));
valve v_12_1807 (.fluid_in(k_12_1807), .fluid_out(k_11_903), .air_in(c_12_1));
valve v_12_1808 (.fluid_in(k_12_1808), .fluid_out(k_11_904), .air_in(c_12_0));
valve v_12_1809 (.fluid_in(k_12_1809), .fluid_out(k_11_904), .air_in(c_12_1));
valve v_12_1810 (.fluid_in(k_12_1810), .fluid_out(k_11_905), .air_in(c_12_0));
valve v_12_1811 (.fluid_in(k_12_1811), .fluid_out(k_11_905), .air_in(c_12_1));
valve v_12_1812 (.fluid_in(k_12_1812), .fluid_out(k_11_906), .air_in(c_12_0));
valve v_12_1813 (.fluid_in(k_12_1813), .fluid_out(k_11_906), .air_in(c_12_1));
valve v_12_1814 (.fluid_in(k_12_1814), .fluid_out(k_11_907), .air_in(c_12_0));
valve v_12_1815 (.fluid_in(k_12_1815), .fluid_out(k_11_907), .air_in(c_12_1));
valve v_12_1816 (.fluid_in(k_12_1816), .fluid_out(k_11_908), .air_in(c_12_0));
valve v_12_1817 (.fluid_in(k_12_1817), .fluid_out(k_11_908), .air_in(c_12_1));
valve v_12_1818 (.fluid_in(k_12_1818), .fluid_out(k_11_909), .air_in(c_12_0));
valve v_12_1819 (.fluid_in(k_12_1819), .fluid_out(k_11_909), .air_in(c_12_1));
valve v_12_1820 (.fluid_in(k_12_1820), .fluid_out(k_11_910), .air_in(c_12_0));
valve v_12_1821 (.fluid_in(k_12_1821), .fluid_out(k_11_910), .air_in(c_12_1));
valve v_12_1822 (.fluid_in(k_12_1822), .fluid_out(k_11_911), .air_in(c_12_0));
valve v_12_1823 (.fluid_in(k_12_1823), .fluid_out(k_11_911), .air_in(c_12_1));
valve v_12_1824 (.fluid_in(k_12_1824), .fluid_out(k_11_912), .air_in(c_12_0));
valve v_12_1825 (.fluid_in(k_12_1825), .fluid_out(k_11_912), .air_in(c_12_1));
valve v_12_1826 (.fluid_in(k_12_1826), .fluid_out(k_11_913), .air_in(c_12_0));
valve v_12_1827 (.fluid_in(k_12_1827), .fluid_out(k_11_913), .air_in(c_12_1));
valve v_12_1828 (.fluid_in(k_12_1828), .fluid_out(k_11_914), .air_in(c_12_0));
valve v_12_1829 (.fluid_in(k_12_1829), .fluid_out(k_11_914), .air_in(c_12_1));
valve v_12_1830 (.fluid_in(k_12_1830), .fluid_out(k_11_915), .air_in(c_12_0));
valve v_12_1831 (.fluid_in(k_12_1831), .fluid_out(k_11_915), .air_in(c_12_1));
valve v_12_1832 (.fluid_in(k_12_1832), .fluid_out(k_11_916), .air_in(c_12_0));
valve v_12_1833 (.fluid_in(k_12_1833), .fluid_out(k_11_916), .air_in(c_12_1));
valve v_12_1834 (.fluid_in(k_12_1834), .fluid_out(k_11_917), .air_in(c_12_0));
valve v_12_1835 (.fluid_in(k_12_1835), .fluid_out(k_11_917), .air_in(c_12_1));
valve v_12_1836 (.fluid_in(k_12_1836), .fluid_out(k_11_918), .air_in(c_12_0));
valve v_12_1837 (.fluid_in(k_12_1837), .fluid_out(k_11_918), .air_in(c_12_1));
valve v_12_1838 (.fluid_in(k_12_1838), .fluid_out(k_11_919), .air_in(c_12_0));
valve v_12_1839 (.fluid_in(k_12_1839), .fluid_out(k_11_919), .air_in(c_12_1));
valve v_12_1840 (.fluid_in(k_12_1840), .fluid_out(k_11_920), .air_in(c_12_0));
valve v_12_1841 (.fluid_in(k_12_1841), .fluid_out(k_11_920), .air_in(c_12_1));
valve v_12_1842 (.fluid_in(k_12_1842), .fluid_out(k_11_921), .air_in(c_12_0));
valve v_12_1843 (.fluid_in(k_12_1843), .fluid_out(k_11_921), .air_in(c_12_1));
valve v_12_1844 (.fluid_in(k_12_1844), .fluid_out(k_11_922), .air_in(c_12_0));
valve v_12_1845 (.fluid_in(k_12_1845), .fluid_out(k_11_922), .air_in(c_12_1));
valve v_12_1846 (.fluid_in(k_12_1846), .fluid_out(k_11_923), .air_in(c_12_0));
valve v_12_1847 (.fluid_in(k_12_1847), .fluid_out(k_11_923), .air_in(c_12_1));
valve v_12_1848 (.fluid_in(k_12_1848), .fluid_out(k_11_924), .air_in(c_12_0));
valve v_12_1849 (.fluid_in(k_12_1849), .fluid_out(k_11_924), .air_in(c_12_1));
valve v_12_1850 (.fluid_in(k_12_1850), .fluid_out(k_11_925), .air_in(c_12_0));
valve v_12_1851 (.fluid_in(k_12_1851), .fluid_out(k_11_925), .air_in(c_12_1));
valve v_12_1852 (.fluid_in(k_12_1852), .fluid_out(k_11_926), .air_in(c_12_0));
valve v_12_1853 (.fluid_in(k_12_1853), .fluid_out(k_11_926), .air_in(c_12_1));
valve v_12_1854 (.fluid_in(k_12_1854), .fluid_out(k_11_927), .air_in(c_12_0));
valve v_12_1855 (.fluid_in(k_12_1855), .fluid_out(k_11_927), .air_in(c_12_1));
valve v_12_1856 (.fluid_in(k_12_1856), .fluid_out(k_11_928), .air_in(c_12_0));
valve v_12_1857 (.fluid_in(k_12_1857), .fluid_out(k_11_928), .air_in(c_12_1));
valve v_12_1858 (.fluid_in(k_12_1858), .fluid_out(k_11_929), .air_in(c_12_0));
valve v_12_1859 (.fluid_in(k_12_1859), .fluid_out(k_11_929), .air_in(c_12_1));
valve v_12_1860 (.fluid_in(k_12_1860), .fluid_out(k_11_930), .air_in(c_12_0));
valve v_12_1861 (.fluid_in(k_12_1861), .fluid_out(k_11_930), .air_in(c_12_1));
valve v_12_1862 (.fluid_in(k_12_1862), .fluid_out(k_11_931), .air_in(c_12_0));
valve v_12_1863 (.fluid_in(k_12_1863), .fluid_out(k_11_931), .air_in(c_12_1));
valve v_12_1864 (.fluid_in(k_12_1864), .fluid_out(k_11_932), .air_in(c_12_0));
valve v_12_1865 (.fluid_in(k_12_1865), .fluid_out(k_11_932), .air_in(c_12_1));
valve v_12_1866 (.fluid_in(k_12_1866), .fluid_out(k_11_933), .air_in(c_12_0));
valve v_12_1867 (.fluid_in(k_12_1867), .fluid_out(k_11_933), .air_in(c_12_1));
valve v_12_1868 (.fluid_in(k_12_1868), .fluid_out(k_11_934), .air_in(c_12_0));
valve v_12_1869 (.fluid_in(k_12_1869), .fluid_out(k_11_934), .air_in(c_12_1));
valve v_12_1870 (.fluid_in(k_12_1870), .fluid_out(k_11_935), .air_in(c_12_0));
valve v_12_1871 (.fluid_in(k_12_1871), .fluid_out(k_11_935), .air_in(c_12_1));
valve v_12_1872 (.fluid_in(k_12_1872), .fluid_out(k_11_936), .air_in(c_12_0));
valve v_12_1873 (.fluid_in(k_12_1873), .fluid_out(k_11_936), .air_in(c_12_1));
valve v_12_1874 (.fluid_in(k_12_1874), .fluid_out(k_11_937), .air_in(c_12_0));
valve v_12_1875 (.fluid_in(k_12_1875), .fluid_out(k_11_937), .air_in(c_12_1));
valve v_12_1876 (.fluid_in(k_12_1876), .fluid_out(k_11_938), .air_in(c_12_0));
valve v_12_1877 (.fluid_in(k_12_1877), .fluid_out(k_11_938), .air_in(c_12_1));
valve v_12_1878 (.fluid_in(k_12_1878), .fluid_out(k_11_939), .air_in(c_12_0));
valve v_12_1879 (.fluid_in(k_12_1879), .fluid_out(k_11_939), .air_in(c_12_1));
valve v_12_1880 (.fluid_in(k_12_1880), .fluid_out(k_11_940), .air_in(c_12_0));
valve v_12_1881 (.fluid_in(k_12_1881), .fluid_out(k_11_940), .air_in(c_12_1));
valve v_12_1882 (.fluid_in(k_12_1882), .fluid_out(k_11_941), .air_in(c_12_0));
valve v_12_1883 (.fluid_in(k_12_1883), .fluid_out(k_11_941), .air_in(c_12_1));
valve v_12_1884 (.fluid_in(k_12_1884), .fluid_out(k_11_942), .air_in(c_12_0));
valve v_12_1885 (.fluid_in(k_12_1885), .fluid_out(k_11_942), .air_in(c_12_1));
valve v_12_1886 (.fluid_in(k_12_1886), .fluid_out(k_11_943), .air_in(c_12_0));
valve v_12_1887 (.fluid_in(k_12_1887), .fluid_out(k_11_943), .air_in(c_12_1));
valve v_12_1888 (.fluid_in(k_12_1888), .fluid_out(k_11_944), .air_in(c_12_0));
valve v_12_1889 (.fluid_in(k_12_1889), .fluid_out(k_11_944), .air_in(c_12_1));
valve v_12_1890 (.fluid_in(k_12_1890), .fluid_out(k_11_945), .air_in(c_12_0));
valve v_12_1891 (.fluid_in(k_12_1891), .fluid_out(k_11_945), .air_in(c_12_1));
valve v_12_1892 (.fluid_in(k_12_1892), .fluid_out(k_11_946), .air_in(c_12_0));
valve v_12_1893 (.fluid_in(k_12_1893), .fluid_out(k_11_946), .air_in(c_12_1));
valve v_12_1894 (.fluid_in(k_12_1894), .fluid_out(k_11_947), .air_in(c_12_0));
valve v_12_1895 (.fluid_in(k_12_1895), .fluid_out(k_11_947), .air_in(c_12_1));
valve v_12_1896 (.fluid_in(k_12_1896), .fluid_out(k_11_948), .air_in(c_12_0));
valve v_12_1897 (.fluid_in(k_12_1897), .fluid_out(k_11_948), .air_in(c_12_1));
valve v_12_1898 (.fluid_in(k_12_1898), .fluid_out(k_11_949), .air_in(c_12_0));
valve v_12_1899 (.fluid_in(k_12_1899), .fluid_out(k_11_949), .air_in(c_12_1));
valve v_12_1900 (.fluid_in(k_12_1900), .fluid_out(k_11_950), .air_in(c_12_0));
valve v_12_1901 (.fluid_in(k_12_1901), .fluid_out(k_11_950), .air_in(c_12_1));
valve v_12_1902 (.fluid_in(k_12_1902), .fluid_out(k_11_951), .air_in(c_12_0));
valve v_12_1903 (.fluid_in(k_12_1903), .fluid_out(k_11_951), .air_in(c_12_1));
valve v_12_1904 (.fluid_in(k_12_1904), .fluid_out(k_11_952), .air_in(c_12_0));
valve v_12_1905 (.fluid_in(k_12_1905), .fluid_out(k_11_952), .air_in(c_12_1));
valve v_12_1906 (.fluid_in(k_12_1906), .fluid_out(k_11_953), .air_in(c_12_0));
valve v_12_1907 (.fluid_in(k_12_1907), .fluid_out(k_11_953), .air_in(c_12_1));
valve v_12_1908 (.fluid_in(k_12_1908), .fluid_out(k_11_954), .air_in(c_12_0));
valve v_12_1909 (.fluid_in(k_12_1909), .fluid_out(k_11_954), .air_in(c_12_1));
valve v_12_1910 (.fluid_in(k_12_1910), .fluid_out(k_11_955), .air_in(c_12_0));
valve v_12_1911 (.fluid_in(k_12_1911), .fluid_out(k_11_955), .air_in(c_12_1));
valve v_12_1912 (.fluid_in(k_12_1912), .fluid_out(k_11_956), .air_in(c_12_0));
valve v_12_1913 (.fluid_in(k_12_1913), .fluid_out(k_11_956), .air_in(c_12_1));
valve v_12_1914 (.fluid_in(k_12_1914), .fluid_out(k_11_957), .air_in(c_12_0));
valve v_12_1915 (.fluid_in(k_12_1915), .fluid_out(k_11_957), .air_in(c_12_1));
valve v_12_1916 (.fluid_in(k_12_1916), .fluid_out(k_11_958), .air_in(c_12_0));
valve v_12_1917 (.fluid_in(k_12_1917), .fluid_out(k_11_958), .air_in(c_12_1));
valve v_12_1918 (.fluid_in(k_12_1918), .fluid_out(k_11_959), .air_in(c_12_0));
valve v_12_1919 (.fluid_in(k_12_1919), .fluid_out(k_11_959), .air_in(c_12_1));
valve v_12_1920 (.fluid_in(k_12_1920), .fluid_out(k_11_960), .air_in(c_12_0));
valve v_12_1921 (.fluid_in(k_12_1921), .fluid_out(k_11_960), .air_in(c_12_1));
valve v_12_1922 (.fluid_in(k_12_1922), .fluid_out(k_11_961), .air_in(c_12_0));
valve v_12_1923 (.fluid_in(k_12_1923), .fluid_out(k_11_961), .air_in(c_12_1));
valve v_12_1924 (.fluid_in(k_12_1924), .fluid_out(k_11_962), .air_in(c_12_0));
valve v_12_1925 (.fluid_in(k_12_1925), .fluid_out(k_11_962), .air_in(c_12_1));
valve v_12_1926 (.fluid_in(k_12_1926), .fluid_out(k_11_963), .air_in(c_12_0));
valve v_12_1927 (.fluid_in(k_12_1927), .fluid_out(k_11_963), .air_in(c_12_1));
valve v_12_1928 (.fluid_in(k_12_1928), .fluid_out(k_11_964), .air_in(c_12_0));
valve v_12_1929 (.fluid_in(k_12_1929), .fluid_out(k_11_964), .air_in(c_12_1));
valve v_12_1930 (.fluid_in(k_12_1930), .fluid_out(k_11_965), .air_in(c_12_0));
valve v_12_1931 (.fluid_in(k_12_1931), .fluid_out(k_11_965), .air_in(c_12_1));
valve v_12_1932 (.fluid_in(k_12_1932), .fluid_out(k_11_966), .air_in(c_12_0));
valve v_12_1933 (.fluid_in(k_12_1933), .fluid_out(k_11_966), .air_in(c_12_1));
valve v_12_1934 (.fluid_in(k_12_1934), .fluid_out(k_11_967), .air_in(c_12_0));
valve v_12_1935 (.fluid_in(k_12_1935), .fluid_out(k_11_967), .air_in(c_12_1));
valve v_12_1936 (.fluid_in(k_12_1936), .fluid_out(k_11_968), .air_in(c_12_0));
valve v_12_1937 (.fluid_in(k_12_1937), .fluid_out(k_11_968), .air_in(c_12_1));
valve v_12_1938 (.fluid_in(k_12_1938), .fluid_out(k_11_969), .air_in(c_12_0));
valve v_12_1939 (.fluid_in(k_12_1939), .fluid_out(k_11_969), .air_in(c_12_1));
valve v_12_1940 (.fluid_in(k_12_1940), .fluid_out(k_11_970), .air_in(c_12_0));
valve v_12_1941 (.fluid_in(k_12_1941), .fluid_out(k_11_970), .air_in(c_12_1));
valve v_12_1942 (.fluid_in(k_12_1942), .fluid_out(k_11_971), .air_in(c_12_0));
valve v_12_1943 (.fluid_in(k_12_1943), .fluid_out(k_11_971), .air_in(c_12_1));
valve v_12_1944 (.fluid_in(k_12_1944), .fluid_out(k_11_972), .air_in(c_12_0));
valve v_12_1945 (.fluid_in(k_12_1945), .fluid_out(k_11_972), .air_in(c_12_1));
valve v_12_1946 (.fluid_in(k_12_1946), .fluid_out(k_11_973), .air_in(c_12_0));
valve v_12_1947 (.fluid_in(k_12_1947), .fluid_out(k_11_973), .air_in(c_12_1));
valve v_12_1948 (.fluid_in(k_12_1948), .fluid_out(k_11_974), .air_in(c_12_0));
valve v_12_1949 (.fluid_in(k_12_1949), .fluid_out(k_11_974), .air_in(c_12_1));
valve v_12_1950 (.fluid_in(k_12_1950), .fluid_out(k_11_975), .air_in(c_12_0));
valve v_12_1951 (.fluid_in(k_12_1951), .fluid_out(k_11_975), .air_in(c_12_1));
valve v_12_1952 (.fluid_in(k_12_1952), .fluid_out(k_11_976), .air_in(c_12_0));
valve v_12_1953 (.fluid_in(k_12_1953), .fluid_out(k_11_976), .air_in(c_12_1));
valve v_12_1954 (.fluid_in(k_12_1954), .fluid_out(k_11_977), .air_in(c_12_0));
valve v_12_1955 (.fluid_in(k_12_1955), .fluid_out(k_11_977), .air_in(c_12_1));
valve v_12_1956 (.fluid_in(k_12_1956), .fluid_out(k_11_978), .air_in(c_12_0));
valve v_12_1957 (.fluid_in(k_12_1957), .fluid_out(k_11_978), .air_in(c_12_1));
valve v_12_1958 (.fluid_in(k_12_1958), .fluid_out(k_11_979), .air_in(c_12_0));
valve v_12_1959 (.fluid_in(k_12_1959), .fluid_out(k_11_979), .air_in(c_12_1));
valve v_12_1960 (.fluid_in(k_12_1960), .fluid_out(k_11_980), .air_in(c_12_0));
valve v_12_1961 (.fluid_in(k_12_1961), .fluid_out(k_11_980), .air_in(c_12_1));
valve v_12_1962 (.fluid_in(k_12_1962), .fluid_out(k_11_981), .air_in(c_12_0));
valve v_12_1963 (.fluid_in(k_12_1963), .fluid_out(k_11_981), .air_in(c_12_1));
valve v_12_1964 (.fluid_in(k_12_1964), .fluid_out(k_11_982), .air_in(c_12_0));
valve v_12_1965 (.fluid_in(k_12_1965), .fluid_out(k_11_982), .air_in(c_12_1));
valve v_12_1966 (.fluid_in(k_12_1966), .fluid_out(k_11_983), .air_in(c_12_0));
valve v_12_1967 (.fluid_in(k_12_1967), .fluid_out(k_11_983), .air_in(c_12_1));
valve v_12_1968 (.fluid_in(k_12_1968), .fluid_out(k_11_984), .air_in(c_12_0));
valve v_12_1969 (.fluid_in(k_12_1969), .fluid_out(k_11_984), .air_in(c_12_1));
valve v_12_1970 (.fluid_in(k_12_1970), .fluid_out(k_11_985), .air_in(c_12_0));
valve v_12_1971 (.fluid_in(k_12_1971), .fluid_out(k_11_985), .air_in(c_12_1));
valve v_12_1972 (.fluid_in(k_12_1972), .fluid_out(k_11_986), .air_in(c_12_0));
valve v_12_1973 (.fluid_in(k_12_1973), .fluid_out(k_11_986), .air_in(c_12_1));
valve v_12_1974 (.fluid_in(k_12_1974), .fluid_out(k_11_987), .air_in(c_12_0));
valve v_12_1975 (.fluid_in(k_12_1975), .fluid_out(k_11_987), .air_in(c_12_1));
valve v_12_1976 (.fluid_in(k_12_1976), .fluid_out(k_11_988), .air_in(c_12_0));
valve v_12_1977 (.fluid_in(k_12_1977), .fluid_out(k_11_988), .air_in(c_12_1));
valve v_12_1978 (.fluid_in(k_12_1978), .fluid_out(k_11_989), .air_in(c_12_0));
valve v_12_1979 (.fluid_in(k_12_1979), .fluid_out(k_11_989), .air_in(c_12_1));
valve v_12_1980 (.fluid_in(k_12_1980), .fluid_out(k_11_990), .air_in(c_12_0));
valve v_12_1981 (.fluid_in(k_12_1981), .fluid_out(k_11_990), .air_in(c_12_1));
valve v_12_1982 (.fluid_in(k_12_1982), .fluid_out(k_11_991), .air_in(c_12_0));
valve v_12_1983 (.fluid_in(k_12_1983), .fluid_out(k_11_991), .air_in(c_12_1));
valve v_12_1984 (.fluid_in(k_12_1984), .fluid_out(k_11_992), .air_in(c_12_0));
valve v_12_1985 (.fluid_in(k_12_1985), .fluid_out(k_11_992), .air_in(c_12_1));
valve v_12_1986 (.fluid_in(k_12_1986), .fluid_out(k_11_993), .air_in(c_12_0));
valve v_12_1987 (.fluid_in(k_12_1987), .fluid_out(k_11_993), .air_in(c_12_1));
valve v_12_1988 (.fluid_in(k_12_1988), .fluid_out(k_11_994), .air_in(c_12_0));
valve v_12_1989 (.fluid_in(k_12_1989), .fluid_out(k_11_994), .air_in(c_12_1));
valve v_12_1990 (.fluid_in(k_12_1990), .fluid_out(k_11_995), .air_in(c_12_0));
valve v_12_1991 (.fluid_in(k_12_1991), .fluid_out(k_11_995), .air_in(c_12_1));
valve v_12_1992 (.fluid_in(k_12_1992), .fluid_out(k_11_996), .air_in(c_12_0));
valve v_12_1993 (.fluid_in(k_12_1993), .fluid_out(k_11_996), .air_in(c_12_1));
valve v_12_1994 (.fluid_in(k_12_1994), .fluid_out(k_11_997), .air_in(c_12_0));
valve v_12_1995 (.fluid_in(k_12_1995), .fluid_out(k_11_997), .air_in(c_12_1));
valve v_12_1996 (.fluid_in(k_12_1996), .fluid_out(k_11_998), .air_in(c_12_0));
valve v_12_1997 (.fluid_in(k_12_1997), .fluid_out(k_11_998), .air_in(c_12_1));
valve v_12_1998 (.fluid_in(k_12_1998), .fluid_out(k_11_999), .air_in(c_12_0));
valve v_12_1999 (.fluid_in(k_12_1999), .fluid_out(k_11_999), .air_in(c_12_1));
valve v_12_2000 (.fluid_in(k_12_2000), .fluid_out(k_11_1000), .air_in(c_12_0));
valve v_12_2001 (.fluid_in(k_12_2001), .fluid_out(k_11_1000), .air_in(c_12_1));
valve v_12_2002 (.fluid_in(k_12_2002), .fluid_out(k_11_1001), .air_in(c_12_0));
valve v_12_2003 (.fluid_in(k_12_2003), .fluid_out(k_11_1001), .air_in(c_12_1));
valve v_12_2004 (.fluid_in(k_12_2004), .fluid_out(k_11_1002), .air_in(c_12_0));
valve v_12_2005 (.fluid_in(k_12_2005), .fluid_out(k_11_1002), .air_in(c_12_1));
valve v_12_2006 (.fluid_in(k_12_2006), .fluid_out(k_11_1003), .air_in(c_12_0));
valve v_12_2007 (.fluid_in(k_12_2007), .fluid_out(k_11_1003), .air_in(c_12_1));
valve v_12_2008 (.fluid_in(k_12_2008), .fluid_out(k_11_1004), .air_in(c_12_0));
valve v_12_2009 (.fluid_in(k_12_2009), .fluid_out(k_11_1004), .air_in(c_12_1));
valve v_12_2010 (.fluid_in(k_12_2010), .fluid_out(k_11_1005), .air_in(c_12_0));
valve v_12_2011 (.fluid_in(k_12_2011), .fluid_out(k_11_1005), .air_in(c_12_1));
valve v_12_2012 (.fluid_in(k_12_2012), .fluid_out(k_11_1006), .air_in(c_12_0));
valve v_12_2013 (.fluid_in(k_12_2013), .fluid_out(k_11_1006), .air_in(c_12_1));
valve v_12_2014 (.fluid_in(k_12_2014), .fluid_out(k_11_1007), .air_in(c_12_0));
valve v_12_2015 (.fluid_in(k_12_2015), .fluid_out(k_11_1007), .air_in(c_12_1));
valve v_12_2016 (.fluid_in(k_12_2016), .fluid_out(k_11_1008), .air_in(c_12_0));
valve v_12_2017 (.fluid_in(k_12_2017), .fluid_out(k_11_1008), .air_in(c_12_1));
valve v_12_2018 (.fluid_in(k_12_2018), .fluid_out(k_11_1009), .air_in(c_12_0));
valve v_12_2019 (.fluid_in(k_12_2019), .fluid_out(k_11_1009), .air_in(c_12_1));
valve v_12_2020 (.fluid_in(k_12_2020), .fluid_out(k_11_1010), .air_in(c_12_0));
valve v_12_2021 (.fluid_in(k_12_2021), .fluid_out(k_11_1010), .air_in(c_12_1));
valve v_12_2022 (.fluid_in(k_12_2022), .fluid_out(k_11_1011), .air_in(c_12_0));
valve v_12_2023 (.fluid_in(k_12_2023), .fluid_out(k_11_1011), .air_in(c_12_1));
valve v_12_2024 (.fluid_in(k_12_2024), .fluid_out(k_11_1012), .air_in(c_12_0));
valve v_12_2025 (.fluid_in(k_12_2025), .fluid_out(k_11_1012), .air_in(c_12_1));
valve v_12_2026 (.fluid_in(k_12_2026), .fluid_out(k_11_1013), .air_in(c_12_0));
valve v_12_2027 (.fluid_in(k_12_2027), .fluid_out(k_11_1013), .air_in(c_12_1));
valve v_12_2028 (.fluid_in(k_12_2028), .fluid_out(k_11_1014), .air_in(c_12_0));
valve v_12_2029 (.fluid_in(k_12_2029), .fluid_out(k_11_1014), .air_in(c_12_1));
valve v_12_2030 (.fluid_in(k_12_2030), .fluid_out(k_11_1015), .air_in(c_12_0));
valve v_12_2031 (.fluid_in(k_12_2031), .fluid_out(k_11_1015), .air_in(c_12_1));
valve v_12_2032 (.fluid_in(k_12_2032), .fluid_out(k_11_1016), .air_in(c_12_0));
valve v_12_2033 (.fluid_in(k_12_2033), .fluid_out(k_11_1016), .air_in(c_12_1));
valve v_12_2034 (.fluid_in(k_12_2034), .fluid_out(k_11_1017), .air_in(c_12_0));
valve v_12_2035 (.fluid_in(k_12_2035), .fluid_out(k_11_1017), .air_in(c_12_1));
valve v_12_2036 (.fluid_in(k_12_2036), .fluid_out(k_11_1018), .air_in(c_12_0));
valve v_12_2037 (.fluid_in(k_12_2037), .fluid_out(k_11_1018), .air_in(c_12_1));
valve v_12_2038 (.fluid_in(k_12_2038), .fluid_out(k_11_1019), .air_in(c_12_0));
valve v_12_2039 (.fluid_in(k_12_2039), .fluid_out(k_11_1019), .air_in(c_12_1));
valve v_12_2040 (.fluid_in(k_12_2040), .fluid_out(k_11_1020), .air_in(c_12_0));
valve v_12_2041 (.fluid_in(k_12_2041), .fluid_out(k_11_1020), .air_in(c_12_1));
valve v_12_2042 (.fluid_in(k_12_2042), .fluid_out(k_11_1021), .air_in(c_12_0));
valve v_12_2043 (.fluid_in(k_12_2043), .fluid_out(k_11_1021), .air_in(c_12_1));
valve v_12_2044 (.fluid_in(k_12_2044), .fluid_out(k_11_1022), .air_in(c_12_0));
valve v_12_2045 (.fluid_in(k_12_2045), .fluid_out(k_11_1022), .air_in(c_12_1));
valve v_12_2046 (.fluid_in(k_12_2046), .fluid_out(k_11_1023), .air_in(c_12_0));
valve v_12_2047 (.fluid_in(k_12_2047), .fluid_out(k_11_1023), .air_in(c_12_1));
valve v_12_2048 (.fluid_in(k_12_2048), .fluid_out(k_11_1024), .air_in(c_12_0));
valve v_12_2049 (.fluid_in(k_12_2049), .fluid_out(k_11_1024), .air_in(c_12_1));
valve v_12_2050 (.fluid_in(k_12_2050), .fluid_out(k_11_1025), .air_in(c_12_0));
valve v_12_2051 (.fluid_in(k_12_2051), .fluid_out(k_11_1025), .air_in(c_12_1));
valve v_12_2052 (.fluid_in(k_12_2052), .fluid_out(k_11_1026), .air_in(c_12_0));
valve v_12_2053 (.fluid_in(k_12_2053), .fluid_out(k_11_1026), .air_in(c_12_1));
valve v_12_2054 (.fluid_in(k_12_2054), .fluid_out(k_11_1027), .air_in(c_12_0));
valve v_12_2055 (.fluid_in(k_12_2055), .fluid_out(k_11_1027), .air_in(c_12_1));
valve v_12_2056 (.fluid_in(k_12_2056), .fluid_out(k_11_1028), .air_in(c_12_0));
valve v_12_2057 (.fluid_in(k_12_2057), .fluid_out(k_11_1028), .air_in(c_12_1));
valve v_12_2058 (.fluid_in(k_12_2058), .fluid_out(k_11_1029), .air_in(c_12_0));
valve v_12_2059 (.fluid_in(k_12_2059), .fluid_out(k_11_1029), .air_in(c_12_1));
valve v_12_2060 (.fluid_in(k_12_2060), .fluid_out(k_11_1030), .air_in(c_12_0));
valve v_12_2061 (.fluid_in(k_12_2061), .fluid_out(k_11_1030), .air_in(c_12_1));
valve v_12_2062 (.fluid_in(k_12_2062), .fluid_out(k_11_1031), .air_in(c_12_0));
valve v_12_2063 (.fluid_in(k_12_2063), .fluid_out(k_11_1031), .air_in(c_12_1));
valve v_12_2064 (.fluid_in(k_12_2064), .fluid_out(k_11_1032), .air_in(c_12_0));
valve v_12_2065 (.fluid_in(k_12_2065), .fluid_out(k_11_1032), .air_in(c_12_1));
valve v_12_2066 (.fluid_in(k_12_2066), .fluid_out(k_11_1033), .air_in(c_12_0));
valve v_12_2067 (.fluid_in(k_12_2067), .fluid_out(k_11_1033), .air_in(c_12_1));
valve v_12_2068 (.fluid_in(k_12_2068), .fluid_out(k_11_1034), .air_in(c_12_0));
valve v_12_2069 (.fluid_in(k_12_2069), .fluid_out(k_11_1034), .air_in(c_12_1));
valve v_12_2070 (.fluid_in(k_12_2070), .fluid_out(k_11_1035), .air_in(c_12_0));
valve v_12_2071 (.fluid_in(k_12_2071), .fluid_out(k_11_1035), .air_in(c_12_1));
valve v_12_2072 (.fluid_in(k_12_2072), .fluid_out(k_11_1036), .air_in(c_12_0));
valve v_12_2073 (.fluid_in(k_12_2073), .fluid_out(k_11_1036), .air_in(c_12_1));
valve v_12_2074 (.fluid_in(k_12_2074), .fluid_out(k_11_1037), .air_in(c_12_0));
valve v_12_2075 (.fluid_in(k_12_2075), .fluid_out(k_11_1037), .air_in(c_12_1));
valve v_12_2076 (.fluid_in(k_12_2076), .fluid_out(k_11_1038), .air_in(c_12_0));
valve v_12_2077 (.fluid_in(k_12_2077), .fluid_out(k_11_1038), .air_in(c_12_1));
valve v_12_2078 (.fluid_in(k_12_2078), .fluid_out(k_11_1039), .air_in(c_12_0));
valve v_12_2079 (.fluid_in(k_12_2079), .fluid_out(k_11_1039), .air_in(c_12_1));
valve v_12_2080 (.fluid_in(k_12_2080), .fluid_out(k_11_1040), .air_in(c_12_0));
valve v_12_2081 (.fluid_in(k_12_2081), .fluid_out(k_11_1040), .air_in(c_12_1));
valve v_12_2082 (.fluid_in(k_12_2082), .fluid_out(k_11_1041), .air_in(c_12_0));
valve v_12_2083 (.fluid_in(k_12_2083), .fluid_out(k_11_1041), .air_in(c_12_1));
valve v_12_2084 (.fluid_in(k_12_2084), .fluid_out(k_11_1042), .air_in(c_12_0));
valve v_12_2085 (.fluid_in(k_12_2085), .fluid_out(k_11_1042), .air_in(c_12_1));
valve v_12_2086 (.fluid_in(k_12_2086), .fluid_out(k_11_1043), .air_in(c_12_0));
valve v_12_2087 (.fluid_in(k_12_2087), .fluid_out(k_11_1043), .air_in(c_12_1));
valve v_12_2088 (.fluid_in(k_12_2088), .fluid_out(k_11_1044), .air_in(c_12_0));
valve v_12_2089 (.fluid_in(k_12_2089), .fluid_out(k_11_1044), .air_in(c_12_1));
valve v_12_2090 (.fluid_in(k_12_2090), .fluid_out(k_11_1045), .air_in(c_12_0));
valve v_12_2091 (.fluid_in(k_12_2091), .fluid_out(k_11_1045), .air_in(c_12_1));
valve v_12_2092 (.fluid_in(k_12_2092), .fluid_out(k_11_1046), .air_in(c_12_0));
valve v_12_2093 (.fluid_in(k_12_2093), .fluid_out(k_11_1046), .air_in(c_12_1));
valve v_12_2094 (.fluid_in(k_12_2094), .fluid_out(k_11_1047), .air_in(c_12_0));
valve v_12_2095 (.fluid_in(k_12_2095), .fluid_out(k_11_1047), .air_in(c_12_1));
valve v_12_2096 (.fluid_in(k_12_2096), .fluid_out(k_11_1048), .air_in(c_12_0));
valve v_12_2097 (.fluid_in(k_12_2097), .fluid_out(k_11_1048), .air_in(c_12_1));
valve v_12_2098 (.fluid_in(k_12_2098), .fluid_out(k_11_1049), .air_in(c_12_0));
valve v_12_2099 (.fluid_in(k_12_2099), .fluid_out(k_11_1049), .air_in(c_12_1));
valve v_12_2100 (.fluid_in(k_12_2100), .fluid_out(k_11_1050), .air_in(c_12_0));
valve v_12_2101 (.fluid_in(k_12_2101), .fluid_out(k_11_1050), .air_in(c_12_1));
valve v_12_2102 (.fluid_in(k_12_2102), .fluid_out(k_11_1051), .air_in(c_12_0));
valve v_12_2103 (.fluid_in(k_12_2103), .fluid_out(k_11_1051), .air_in(c_12_1));
valve v_12_2104 (.fluid_in(k_12_2104), .fluid_out(k_11_1052), .air_in(c_12_0));
valve v_12_2105 (.fluid_in(k_12_2105), .fluid_out(k_11_1052), .air_in(c_12_1));
valve v_12_2106 (.fluid_in(k_12_2106), .fluid_out(k_11_1053), .air_in(c_12_0));
valve v_12_2107 (.fluid_in(k_12_2107), .fluid_out(k_11_1053), .air_in(c_12_1));
valve v_12_2108 (.fluid_in(k_12_2108), .fluid_out(k_11_1054), .air_in(c_12_0));
valve v_12_2109 (.fluid_in(k_12_2109), .fluid_out(k_11_1054), .air_in(c_12_1));
valve v_12_2110 (.fluid_in(k_12_2110), .fluid_out(k_11_1055), .air_in(c_12_0));
valve v_12_2111 (.fluid_in(k_12_2111), .fluid_out(k_11_1055), .air_in(c_12_1));
valve v_12_2112 (.fluid_in(k_12_2112), .fluid_out(k_11_1056), .air_in(c_12_0));
valve v_12_2113 (.fluid_in(k_12_2113), .fluid_out(k_11_1056), .air_in(c_12_1));
valve v_12_2114 (.fluid_in(k_12_2114), .fluid_out(k_11_1057), .air_in(c_12_0));
valve v_12_2115 (.fluid_in(k_12_2115), .fluid_out(k_11_1057), .air_in(c_12_1));
valve v_12_2116 (.fluid_in(k_12_2116), .fluid_out(k_11_1058), .air_in(c_12_0));
valve v_12_2117 (.fluid_in(k_12_2117), .fluid_out(k_11_1058), .air_in(c_12_1));
valve v_12_2118 (.fluid_in(k_12_2118), .fluid_out(k_11_1059), .air_in(c_12_0));
valve v_12_2119 (.fluid_in(k_12_2119), .fluid_out(k_11_1059), .air_in(c_12_1));
valve v_12_2120 (.fluid_in(k_12_2120), .fluid_out(k_11_1060), .air_in(c_12_0));
valve v_12_2121 (.fluid_in(k_12_2121), .fluid_out(k_11_1060), .air_in(c_12_1));
valve v_12_2122 (.fluid_in(k_12_2122), .fluid_out(k_11_1061), .air_in(c_12_0));
valve v_12_2123 (.fluid_in(k_12_2123), .fluid_out(k_11_1061), .air_in(c_12_1));
valve v_12_2124 (.fluid_in(k_12_2124), .fluid_out(k_11_1062), .air_in(c_12_0));
valve v_12_2125 (.fluid_in(k_12_2125), .fluid_out(k_11_1062), .air_in(c_12_1));
valve v_12_2126 (.fluid_in(k_12_2126), .fluid_out(k_11_1063), .air_in(c_12_0));
valve v_12_2127 (.fluid_in(k_12_2127), .fluid_out(k_11_1063), .air_in(c_12_1));
valve v_12_2128 (.fluid_in(k_12_2128), .fluid_out(k_11_1064), .air_in(c_12_0));
valve v_12_2129 (.fluid_in(k_12_2129), .fluid_out(k_11_1064), .air_in(c_12_1));
valve v_12_2130 (.fluid_in(k_12_2130), .fluid_out(k_11_1065), .air_in(c_12_0));
valve v_12_2131 (.fluid_in(k_12_2131), .fluid_out(k_11_1065), .air_in(c_12_1));
valve v_12_2132 (.fluid_in(k_12_2132), .fluid_out(k_11_1066), .air_in(c_12_0));
valve v_12_2133 (.fluid_in(k_12_2133), .fluid_out(k_11_1066), .air_in(c_12_1));
valve v_12_2134 (.fluid_in(k_12_2134), .fluid_out(k_11_1067), .air_in(c_12_0));
valve v_12_2135 (.fluid_in(k_12_2135), .fluid_out(k_11_1067), .air_in(c_12_1));
valve v_12_2136 (.fluid_in(k_12_2136), .fluid_out(k_11_1068), .air_in(c_12_0));
valve v_12_2137 (.fluid_in(k_12_2137), .fluid_out(k_11_1068), .air_in(c_12_1));
valve v_12_2138 (.fluid_in(k_12_2138), .fluid_out(k_11_1069), .air_in(c_12_0));
valve v_12_2139 (.fluid_in(k_12_2139), .fluid_out(k_11_1069), .air_in(c_12_1));
valve v_12_2140 (.fluid_in(k_12_2140), .fluid_out(k_11_1070), .air_in(c_12_0));
valve v_12_2141 (.fluid_in(k_12_2141), .fluid_out(k_11_1070), .air_in(c_12_1));
valve v_12_2142 (.fluid_in(k_12_2142), .fluid_out(k_11_1071), .air_in(c_12_0));
valve v_12_2143 (.fluid_in(k_12_2143), .fluid_out(k_11_1071), .air_in(c_12_1));
valve v_12_2144 (.fluid_in(k_12_2144), .fluid_out(k_11_1072), .air_in(c_12_0));
valve v_12_2145 (.fluid_in(k_12_2145), .fluid_out(k_11_1072), .air_in(c_12_1));
valve v_12_2146 (.fluid_in(k_12_2146), .fluid_out(k_11_1073), .air_in(c_12_0));
valve v_12_2147 (.fluid_in(k_12_2147), .fluid_out(k_11_1073), .air_in(c_12_1));
valve v_12_2148 (.fluid_in(k_12_2148), .fluid_out(k_11_1074), .air_in(c_12_0));
valve v_12_2149 (.fluid_in(k_12_2149), .fluid_out(k_11_1074), .air_in(c_12_1));
valve v_12_2150 (.fluid_in(k_12_2150), .fluid_out(k_11_1075), .air_in(c_12_0));
valve v_12_2151 (.fluid_in(k_12_2151), .fluid_out(k_11_1075), .air_in(c_12_1));
valve v_12_2152 (.fluid_in(k_12_2152), .fluid_out(k_11_1076), .air_in(c_12_0));
valve v_12_2153 (.fluid_in(k_12_2153), .fluid_out(k_11_1076), .air_in(c_12_1));
valve v_12_2154 (.fluid_in(k_12_2154), .fluid_out(k_11_1077), .air_in(c_12_0));
valve v_12_2155 (.fluid_in(k_12_2155), .fluid_out(k_11_1077), .air_in(c_12_1));
valve v_12_2156 (.fluid_in(k_12_2156), .fluid_out(k_11_1078), .air_in(c_12_0));
valve v_12_2157 (.fluid_in(k_12_2157), .fluid_out(k_11_1078), .air_in(c_12_1));
valve v_12_2158 (.fluid_in(k_12_2158), .fluid_out(k_11_1079), .air_in(c_12_0));
valve v_12_2159 (.fluid_in(k_12_2159), .fluid_out(k_11_1079), .air_in(c_12_1));
valve v_12_2160 (.fluid_in(k_12_2160), .fluid_out(k_11_1080), .air_in(c_12_0));
valve v_12_2161 (.fluid_in(k_12_2161), .fluid_out(k_11_1080), .air_in(c_12_1));
valve v_12_2162 (.fluid_in(k_12_2162), .fluid_out(k_11_1081), .air_in(c_12_0));
valve v_12_2163 (.fluid_in(k_12_2163), .fluid_out(k_11_1081), .air_in(c_12_1));
valve v_12_2164 (.fluid_in(k_12_2164), .fluid_out(k_11_1082), .air_in(c_12_0));
valve v_12_2165 (.fluid_in(k_12_2165), .fluid_out(k_11_1082), .air_in(c_12_1));
valve v_12_2166 (.fluid_in(k_12_2166), .fluid_out(k_11_1083), .air_in(c_12_0));
valve v_12_2167 (.fluid_in(k_12_2167), .fluid_out(k_11_1083), .air_in(c_12_1));
valve v_12_2168 (.fluid_in(k_12_2168), .fluid_out(k_11_1084), .air_in(c_12_0));
valve v_12_2169 (.fluid_in(k_12_2169), .fluid_out(k_11_1084), .air_in(c_12_1));
valve v_12_2170 (.fluid_in(k_12_2170), .fluid_out(k_11_1085), .air_in(c_12_0));
valve v_12_2171 (.fluid_in(k_12_2171), .fluid_out(k_11_1085), .air_in(c_12_1));
valve v_12_2172 (.fluid_in(k_12_2172), .fluid_out(k_11_1086), .air_in(c_12_0));
valve v_12_2173 (.fluid_in(k_12_2173), .fluid_out(k_11_1086), .air_in(c_12_1));
valve v_12_2174 (.fluid_in(k_12_2174), .fluid_out(k_11_1087), .air_in(c_12_0));
valve v_12_2175 (.fluid_in(k_12_2175), .fluid_out(k_11_1087), .air_in(c_12_1));
valve v_12_2176 (.fluid_in(k_12_2176), .fluid_out(k_11_1088), .air_in(c_12_0));
valve v_12_2177 (.fluid_in(k_12_2177), .fluid_out(k_11_1088), .air_in(c_12_1));
valve v_12_2178 (.fluid_in(k_12_2178), .fluid_out(k_11_1089), .air_in(c_12_0));
valve v_12_2179 (.fluid_in(k_12_2179), .fluid_out(k_11_1089), .air_in(c_12_1));
valve v_12_2180 (.fluid_in(k_12_2180), .fluid_out(k_11_1090), .air_in(c_12_0));
valve v_12_2181 (.fluid_in(k_12_2181), .fluid_out(k_11_1090), .air_in(c_12_1));
valve v_12_2182 (.fluid_in(k_12_2182), .fluid_out(k_11_1091), .air_in(c_12_0));
valve v_12_2183 (.fluid_in(k_12_2183), .fluid_out(k_11_1091), .air_in(c_12_1));
valve v_12_2184 (.fluid_in(k_12_2184), .fluid_out(k_11_1092), .air_in(c_12_0));
valve v_12_2185 (.fluid_in(k_12_2185), .fluid_out(k_11_1092), .air_in(c_12_1));
valve v_12_2186 (.fluid_in(k_12_2186), .fluid_out(k_11_1093), .air_in(c_12_0));
valve v_12_2187 (.fluid_in(k_12_2187), .fluid_out(k_11_1093), .air_in(c_12_1));
valve v_12_2188 (.fluid_in(k_12_2188), .fluid_out(k_11_1094), .air_in(c_12_0));
valve v_12_2189 (.fluid_in(k_12_2189), .fluid_out(k_11_1094), .air_in(c_12_1));
valve v_12_2190 (.fluid_in(k_12_2190), .fluid_out(k_11_1095), .air_in(c_12_0));
valve v_12_2191 (.fluid_in(k_12_2191), .fluid_out(k_11_1095), .air_in(c_12_1));
valve v_12_2192 (.fluid_in(k_12_2192), .fluid_out(k_11_1096), .air_in(c_12_0));
valve v_12_2193 (.fluid_in(k_12_2193), .fluid_out(k_11_1096), .air_in(c_12_1));
valve v_12_2194 (.fluid_in(k_12_2194), .fluid_out(k_11_1097), .air_in(c_12_0));
valve v_12_2195 (.fluid_in(k_12_2195), .fluid_out(k_11_1097), .air_in(c_12_1));
valve v_12_2196 (.fluid_in(k_12_2196), .fluid_out(k_11_1098), .air_in(c_12_0));
valve v_12_2197 (.fluid_in(k_12_2197), .fluid_out(k_11_1098), .air_in(c_12_1));
valve v_12_2198 (.fluid_in(k_12_2198), .fluid_out(k_11_1099), .air_in(c_12_0));
valve v_12_2199 (.fluid_in(k_12_2199), .fluid_out(k_11_1099), .air_in(c_12_1));
valve v_12_2200 (.fluid_in(k_12_2200), .fluid_out(k_11_1100), .air_in(c_12_0));
valve v_12_2201 (.fluid_in(k_12_2201), .fluid_out(k_11_1100), .air_in(c_12_1));
valve v_12_2202 (.fluid_in(k_12_2202), .fluid_out(k_11_1101), .air_in(c_12_0));
valve v_12_2203 (.fluid_in(k_12_2203), .fluid_out(k_11_1101), .air_in(c_12_1));
valve v_12_2204 (.fluid_in(k_12_2204), .fluid_out(k_11_1102), .air_in(c_12_0));
valve v_12_2205 (.fluid_in(k_12_2205), .fluid_out(k_11_1102), .air_in(c_12_1));
valve v_12_2206 (.fluid_in(k_12_2206), .fluid_out(k_11_1103), .air_in(c_12_0));
valve v_12_2207 (.fluid_in(k_12_2207), .fluid_out(k_11_1103), .air_in(c_12_1));
valve v_12_2208 (.fluid_in(k_12_2208), .fluid_out(k_11_1104), .air_in(c_12_0));
valve v_12_2209 (.fluid_in(k_12_2209), .fluid_out(k_11_1104), .air_in(c_12_1));
valve v_12_2210 (.fluid_in(k_12_2210), .fluid_out(k_11_1105), .air_in(c_12_0));
valve v_12_2211 (.fluid_in(k_12_2211), .fluid_out(k_11_1105), .air_in(c_12_1));
valve v_12_2212 (.fluid_in(k_12_2212), .fluid_out(k_11_1106), .air_in(c_12_0));
valve v_12_2213 (.fluid_in(k_12_2213), .fluid_out(k_11_1106), .air_in(c_12_1));
valve v_12_2214 (.fluid_in(k_12_2214), .fluid_out(k_11_1107), .air_in(c_12_0));
valve v_12_2215 (.fluid_in(k_12_2215), .fluid_out(k_11_1107), .air_in(c_12_1));
valve v_12_2216 (.fluid_in(k_12_2216), .fluid_out(k_11_1108), .air_in(c_12_0));
valve v_12_2217 (.fluid_in(k_12_2217), .fluid_out(k_11_1108), .air_in(c_12_1));
valve v_12_2218 (.fluid_in(k_12_2218), .fluid_out(k_11_1109), .air_in(c_12_0));
valve v_12_2219 (.fluid_in(k_12_2219), .fluid_out(k_11_1109), .air_in(c_12_1));
valve v_12_2220 (.fluid_in(k_12_2220), .fluid_out(k_11_1110), .air_in(c_12_0));
valve v_12_2221 (.fluid_in(k_12_2221), .fluid_out(k_11_1110), .air_in(c_12_1));
valve v_12_2222 (.fluid_in(k_12_2222), .fluid_out(k_11_1111), .air_in(c_12_0));
valve v_12_2223 (.fluid_in(k_12_2223), .fluid_out(k_11_1111), .air_in(c_12_1));
valve v_12_2224 (.fluid_in(k_12_2224), .fluid_out(k_11_1112), .air_in(c_12_0));
valve v_12_2225 (.fluid_in(k_12_2225), .fluid_out(k_11_1112), .air_in(c_12_1));
valve v_12_2226 (.fluid_in(k_12_2226), .fluid_out(k_11_1113), .air_in(c_12_0));
valve v_12_2227 (.fluid_in(k_12_2227), .fluid_out(k_11_1113), .air_in(c_12_1));
valve v_12_2228 (.fluid_in(k_12_2228), .fluid_out(k_11_1114), .air_in(c_12_0));
valve v_12_2229 (.fluid_in(k_12_2229), .fluid_out(k_11_1114), .air_in(c_12_1));
valve v_12_2230 (.fluid_in(k_12_2230), .fluid_out(k_11_1115), .air_in(c_12_0));
valve v_12_2231 (.fluid_in(k_12_2231), .fluid_out(k_11_1115), .air_in(c_12_1));
valve v_12_2232 (.fluid_in(k_12_2232), .fluid_out(k_11_1116), .air_in(c_12_0));
valve v_12_2233 (.fluid_in(k_12_2233), .fluid_out(k_11_1116), .air_in(c_12_1));
valve v_12_2234 (.fluid_in(k_12_2234), .fluid_out(k_11_1117), .air_in(c_12_0));
valve v_12_2235 (.fluid_in(k_12_2235), .fluid_out(k_11_1117), .air_in(c_12_1));
valve v_12_2236 (.fluid_in(k_12_2236), .fluid_out(k_11_1118), .air_in(c_12_0));
valve v_12_2237 (.fluid_in(k_12_2237), .fluid_out(k_11_1118), .air_in(c_12_1));
valve v_12_2238 (.fluid_in(k_12_2238), .fluid_out(k_11_1119), .air_in(c_12_0));
valve v_12_2239 (.fluid_in(k_12_2239), .fluid_out(k_11_1119), .air_in(c_12_1));
valve v_12_2240 (.fluid_in(k_12_2240), .fluid_out(k_11_1120), .air_in(c_12_0));
valve v_12_2241 (.fluid_in(k_12_2241), .fluid_out(k_11_1120), .air_in(c_12_1));
valve v_12_2242 (.fluid_in(k_12_2242), .fluid_out(k_11_1121), .air_in(c_12_0));
valve v_12_2243 (.fluid_in(k_12_2243), .fluid_out(k_11_1121), .air_in(c_12_1));
valve v_12_2244 (.fluid_in(k_12_2244), .fluid_out(k_11_1122), .air_in(c_12_0));
valve v_12_2245 (.fluid_in(k_12_2245), .fluid_out(k_11_1122), .air_in(c_12_1));
valve v_12_2246 (.fluid_in(k_12_2246), .fluid_out(k_11_1123), .air_in(c_12_0));
valve v_12_2247 (.fluid_in(k_12_2247), .fluid_out(k_11_1123), .air_in(c_12_1));
valve v_12_2248 (.fluid_in(k_12_2248), .fluid_out(k_11_1124), .air_in(c_12_0));
valve v_12_2249 (.fluid_in(k_12_2249), .fluid_out(k_11_1124), .air_in(c_12_1));
valve v_12_2250 (.fluid_in(k_12_2250), .fluid_out(k_11_1125), .air_in(c_12_0));
valve v_12_2251 (.fluid_in(k_12_2251), .fluid_out(k_11_1125), .air_in(c_12_1));
valve v_12_2252 (.fluid_in(k_12_2252), .fluid_out(k_11_1126), .air_in(c_12_0));
valve v_12_2253 (.fluid_in(k_12_2253), .fluid_out(k_11_1126), .air_in(c_12_1));
valve v_12_2254 (.fluid_in(k_12_2254), .fluid_out(k_11_1127), .air_in(c_12_0));
valve v_12_2255 (.fluid_in(k_12_2255), .fluid_out(k_11_1127), .air_in(c_12_1));
valve v_12_2256 (.fluid_in(k_12_2256), .fluid_out(k_11_1128), .air_in(c_12_0));
valve v_12_2257 (.fluid_in(k_12_2257), .fluid_out(k_11_1128), .air_in(c_12_1));
valve v_12_2258 (.fluid_in(k_12_2258), .fluid_out(k_11_1129), .air_in(c_12_0));
valve v_12_2259 (.fluid_in(k_12_2259), .fluid_out(k_11_1129), .air_in(c_12_1));
valve v_12_2260 (.fluid_in(k_12_2260), .fluid_out(k_11_1130), .air_in(c_12_0));
valve v_12_2261 (.fluid_in(k_12_2261), .fluid_out(k_11_1130), .air_in(c_12_1));
valve v_12_2262 (.fluid_in(k_12_2262), .fluid_out(k_11_1131), .air_in(c_12_0));
valve v_12_2263 (.fluid_in(k_12_2263), .fluid_out(k_11_1131), .air_in(c_12_1));
valve v_12_2264 (.fluid_in(k_12_2264), .fluid_out(k_11_1132), .air_in(c_12_0));
valve v_12_2265 (.fluid_in(k_12_2265), .fluid_out(k_11_1132), .air_in(c_12_1));
valve v_12_2266 (.fluid_in(k_12_2266), .fluid_out(k_11_1133), .air_in(c_12_0));
valve v_12_2267 (.fluid_in(k_12_2267), .fluid_out(k_11_1133), .air_in(c_12_1));
valve v_12_2268 (.fluid_in(k_12_2268), .fluid_out(k_11_1134), .air_in(c_12_0));
valve v_12_2269 (.fluid_in(k_12_2269), .fluid_out(k_11_1134), .air_in(c_12_1));
valve v_12_2270 (.fluid_in(k_12_2270), .fluid_out(k_11_1135), .air_in(c_12_0));
valve v_12_2271 (.fluid_in(k_12_2271), .fluid_out(k_11_1135), .air_in(c_12_1));
valve v_12_2272 (.fluid_in(k_12_2272), .fluid_out(k_11_1136), .air_in(c_12_0));
valve v_12_2273 (.fluid_in(k_12_2273), .fluid_out(k_11_1136), .air_in(c_12_1));
valve v_12_2274 (.fluid_in(k_12_2274), .fluid_out(k_11_1137), .air_in(c_12_0));
valve v_12_2275 (.fluid_in(k_12_2275), .fluid_out(k_11_1137), .air_in(c_12_1));
valve v_12_2276 (.fluid_in(k_12_2276), .fluid_out(k_11_1138), .air_in(c_12_0));
valve v_12_2277 (.fluid_in(k_12_2277), .fluid_out(k_11_1138), .air_in(c_12_1));
valve v_12_2278 (.fluid_in(k_12_2278), .fluid_out(k_11_1139), .air_in(c_12_0));
valve v_12_2279 (.fluid_in(k_12_2279), .fluid_out(k_11_1139), .air_in(c_12_1));
valve v_12_2280 (.fluid_in(k_12_2280), .fluid_out(k_11_1140), .air_in(c_12_0));
valve v_12_2281 (.fluid_in(k_12_2281), .fluid_out(k_11_1140), .air_in(c_12_1));
valve v_12_2282 (.fluid_in(k_12_2282), .fluid_out(k_11_1141), .air_in(c_12_0));
valve v_12_2283 (.fluid_in(k_12_2283), .fluid_out(k_11_1141), .air_in(c_12_1));
valve v_12_2284 (.fluid_in(k_12_2284), .fluid_out(k_11_1142), .air_in(c_12_0));
valve v_12_2285 (.fluid_in(k_12_2285), .fluid_out(k_11_1142), .air_in(c_12_1));
valve v_12_2286 (.fluid_in(k_12_2286), .fluid_out(k_11_1143), .air_in(c_12_0));
valve v_12_2287 (.fluid_in(k_12_2287), .fluid_out(k_11_1143), .air_in(c_12_1));
valve v_12_2288 (.fluid_in(k_12_2288), .fluid_out(k_11_1144), .air_in(c_12_0));
valve v_12_2289 (.fluid_in(k_12_2289), .fluid_out(k_11_1144), .air_in(c_12_1));
valve v_12_2290 (.fluid_in(k_12_2290), .fluid_out(k_11_1145), .air_in(c_12_0));
valve v_12_2291 (.fluid_in(k_12_2291), .fluid_out(k_11_1145), .air_in(c_12_1));
valve v_12_2292 (.fluid_in(k_12_2292), .fluid_out(k_11_1146), .air_in(c_12_0));
valve v_12_2293 (.fluid_in(k_12_2293), .fluid_out(k_11_1146), .air_in(c_12_1));
valve v_12_2294 (.fluid_in(k_12_2294), .fluid_out(k_11_1147), .air_in(c_12_0));
valve v_12_2295 (.fluid_in(k_12_2295), .fluid_out(k_11_1147), .air_in(c_12_1));
valve v_12_2296 (.fluid_in(k_12_2296), .fluid_out(k_11_1148), .air_in(c_12_0));
valve v_12_2297 (.fluid_in(k_12_2297), .fluid_out(k_11_1148), .air_in(c_12_1));
valve v_12_2298 (.fluid_in(k_12_2298), .fluid_out(k_11_1149), .air_in(c_12_0));
valve v_12_2299 (.fluid_in(k_12_2299), .fluid_out(k_11_1149), .air_in(c_12_1));
valve v_12_2300 (.fluid_in(k_12_2300), .fluid_out(k_11_1150), .air_in(c_12_0));
valve v_12_2301 (.fluid_in(k_12_2301), .fluid_out(k_11_1150), .air_in(c_12_1));
valve v_12_2302 (.fluid_in(k_12_2302), .fluid_out(k_11_1151), .air_in(c_12_0));
valve v_12_2303 (.fluid_in(k_12_2303), .fluid_out(k_11_1151), .air_in(c_12_1));
valve v_12_2304 (.fluid_in(k_12_2304), .fluid_out(k_11_1152), .air_in(c_12_0));
valve v_12_2305 (.fluid_in(k_12_2305), .fluid_out(k_11_1152), .air_in(c_12_1));
valve v_12_2306 (.fluid_in(k_12_2306), .fluid_out(k_11_1153), .air_in(c_12_0));
valve v_12_2307 (.fluid_in(k_12_2307), .fluid_out(k_11_1153), .air_in(c_12_1));
valve v_12_2308 (.fluid_in(k_12_2308), .fluid_out(k_11_1154), .air_in(c_12_0));
valve v_12_2309 (.fluid_in(k_12_2309), .fluid_out(k_11_1154), .air_in(c_12_1));
valve v_12_2310 (.fluid_in(k_12_2310), .fluid_out(k_11_1155), .air_in(c_12_0));
valve v_12_2311 (.fluid_in(k_12_2311), .fluid_out(k_11_1155), .air_in(c_12_1));
valve v_12_2312 (.fluid_in(k_12_2312), .fluid_out(k_11_1156), .air_in(c_12_0));
valve v_12_2313 (.fluid_in(k_12_2313), .fluid_out(k_11_1156), .air_in(c_12_1));
valve v_12_2314 (.fluid_in(k_12_2314), .fluid_out(k_11_1157), .air_in(c_12_0));
valve v_12_2315 (.fluid_in(k_12_2315), .fluid_out(k_11_1157), .air_in(c_12_1));
valve v_12_2316 (.fluid_in(k_12_2316), .fluid_out(k_11_1158), .air_in(c_12_0));
valve v_12_2317 (.fluid_in(k_12_2317), .fluid_out(k_11_1158), .air_in(c_12_1));
valve v_12_2318 (.fluid_in(k_12_2318), .fluid_out(k_11_1159), .air_in(c_12_0));
valve v_12_2319 (.fluid_in(k_12_2319), .fluid_out(k_11_1159), .air_in(c_12_1));
valve v_12_2320 (.fluid_in(k_12_2320), .fluid_out(k_11_1160), .air_in(c_12_0));
valve v_12_2321 (.fluid_in(k_12_2321), .fluid_out(k_11_1160), .air_in(c_12_1));
valve v_12_2322 (.fluid_in(k_12_2322), .fluid_out(k_11_1161), .air_in(c_12_0));
valve v_12_2323 (.fluid_in(k_12_2323), .fluid_out(k_11_1161), .air_in(c_12_1));
valve v_12_2324 (.fluid_in(k_12_2324), .fluid_out(k_11_1162), .air_in(c_12_0));
valve v_12_2325 (.fluid_in(k_12_2325), .fluid_out(k_11_1162), .air_in(c_12_1));
valve v_12_2326 (.fluid_in(k_12_2326), .fluid_out(k_11_1163), .air_in(c_12_0));
valve v_12_2327 (.fluid_in(k_12_2327), .fluid_out(k_11_1163), .air_in(c_12_1));
valve v_12_2328 (.fluid_in(k_12_2328), .fluid_out(k_11_1164), .air_in(c_12_0));
valve v_12_2329 (.fluid_in(k_12_2329), .fluid_out(k_11_1164), .air_in(c_12_1));
valve v_12_2330 (.fluid_in(k_12_2330), .fluid_out(k_11_1165), .air_in(c_12_0));
valve v_12_2331 (.fluid_in(k_12_2331), .fluid_out(k_11_1165), .air_in(c_12_1));
valve v_12_2332 (.fluid_in(k_12_2332), .fluid_out(k_11_1166), .air_in(c_12_0));
valve v_12_2333 (.fluid_in(k_12_2333), .fluid_out(k_11_1166), .air_in(c_12_1));
valve v_12_2334 (.fluid_in(k_12_2334), .fluid_out(k_11_1167), .air_in(c_12_0));
valve v_12_2335 (.fluid_in(k_12_2335), .fluid_out(k_11_1167), .air_in(c_12_1));
valve v_12_2336 (.fluid_in(k_12_2336), .fluid_out(k_11_1168), .air_in(c_12_0));
valve v_12_2337 (.fluid_in(k_12_2337), .fluid_out(k_11_1168), .air_in(c_12_1));
valve v_12_2338 (.fluid_in(k_12_2338), .fluid_out(k_11_1169), .air_in(c_12_0));
valve v_12_2339 (.fluid_in(k_12_2339), .fluid_out(k_11_1169), .air_in(c_12_1));
valve v_12_2340 (.fluid_in(k_12_2340), .fluid_out(k_11_1170), .air_in(c_12_0));
valve v_12_2341 (.fluid_in(k_12_2341), .fluid_out(k_11_1170), .air_in(c_12_1));
valve v_12_2342 (.fluid_in(k_12_2342), .fluid_out(k_11_1171), .air_in(c_12_0));
valve v_12_2343 (.fluid_in(k_12_2343), .fluid_out(k_11_1171), .air_in(c_12_1));
valve v_12_2344 (.fluid_in(k_12_2344), .fluid_out(k_11_1172), .air_in(c_12_0));
valve v_12_2345 (.fluid_in(k_12_2345), .fluid_out(k_11_1172), .air_in(c_12_1));
valve v_12_2346 (.fluid_in(k_12_2346), .fluid_out(k_11_1173), .air_in(c_12_0));
valve v_12_2347 (.fluid_in(k_12_2347), .fluid_out(k_11_1173), .air_in(c_12_1));
valve v_12_2348 (.fluid_in(k_12_2348), .fluid_out(k_11_1174), .air_in(c_12_0));
valve v_12_2349 (.fluid_in(k_12_2349), .fluid_out(k_11_1174), .air_in(c_12_1));
valve v_12_2350 (.fluid_in(k_12_2350), .fluid_out(k_11_1175), .air_in(c_12_0));
valve v_12_2351 (.fluid_in(k_12_2351), .fluid_out(k_11_1175), .air_in(c_12_1));
valve v_12_2352 (.fluid_in(k_12_2352), .fluid_out(k_11_1176), .air_in(c_12_0));
valve v_12_2353 (.fluid_in(k_12_2353), .fluid_out(k_11_1176), .air_in(c_12_1));
valve v_12_2354 (.fluid_in(k_12_2354), .fluid_out(k_11_1177), .air_in(c_12_0));
valve v_12_2355 (.fluid_in(k_12_2355), .fluid_out(k_11_1177), .air_in(c_12_1));
valve v_12_2356 (.fluid_in(k_12_2356), .fluid_out(k_11_1178), .air_in(c_12_0));
valve v_12_2357 (.fluid_in(k_12_2357), .fluid_out(k_11_1178), .air_in(c_12_1));
valve v_12_2358 (.fluid_in(k_12_2358), .fluid_out(k_11_1179), .air_in(c_12_0));
valve v_12_2359 (.fluid_in(k_12_2359), .fluid_out(k_11_1179), .air_in(c_12_1));
valve v_12_2360 (.fluid_in(k_12_2360), .fluid_out(k_11_1180), .air_in(c_12_0));
valve v_12_2361 (.fluid_in(k_12_2361), .fluid_out(k_11_1180), .air_in(c_12_1));
valve v_12_2362 (.fluid_in(k_12_2362), .fluid_out(k_11_1181), .air_in(c_12_0));
valve v_12_2363 (.fluid_in(k_12_2363), .fluid_out(k_11_1181), .air_in(c_12_1));
valve v_12_2364 (.fluid_in(k_12_2364), .fluid_out(k_11_1182), .air_in(c_12_0));
valve v_12_2365 (.fluid_in(k_12_2365), .fluid_out(k_11_1182), .air_in(c_12_1));
valve v_12_2366 (.fluid_in(k_12_2366), .fluid_out(k_11_1183), .air_in(c_12_0));
valve v_12_2367 (.fluid_in(k_12_2367), .fluid_out(k_11_1183), .air_in(c_12_1));
valve v_12_2368 (.fluid_in(k_12_2368), .fluid_out(k_11_1184), .air_in(c_12_0));
valve v_12_2369 (.fluid_in(k_12_2369), .fluid_out(k_11_1184), .air_in(c_12_1));
valve v_12_2370 (.fluid_in(k_12_2370), .fluid_out(k_11_1185), .air_in(c_12_0));
valve v_12_2371 (.fluid_in(k_12_2371), .fluid_out(k_11_1185), .air_in(c_12_1));
valve v_12_2372 (.fluid_in(k_12_2372), .fluid_out(k_11_1186), .air_in(c_12_0));
valve v_12_2373 (.fluid_in(k_12_2373), .fluid_out(k_11_1186), .air_in(c_12_1));
valve v_12_2374 (.fluid_in(k_12_2374), .fluid_out(k_11_1187), .air_in(c_12_0));
valve v_12_2375 (.fluid_in(k_12_2375), .fluid_out(k_11_1187), .air_in(c_12_1));
valve v_12_2376 (.fluid_in(k_12_2376), .fluid_out(k_11_1188), .air_in(c_12_0));
valve v_12_2377 (.fluid_in(k_12_2377), .fluid_out(k_11_1188), .air_in(c_12_1));
valve v_12_2378 (.fluid_in(k_12_2378), .fluid_out(k_11_1189), .air_in(c_12_0));
valve v_12_2379 (.fluid_in(k_12_2379), .fluid_out(k_11_1189), .air_in(c_12_1));
valve v_12_2380 (.fluid_in(k_12_2380), .fluid_out(k_11_1190), .air_in(c_12_0));
valve v_12_2381 (.fluid_in(k_12_2381), .fluid_out(k_11_1190), .air_in(c_12_1));
valve v_12_2382 (.fluid_in(k_12_2382), .fluid_out(k_11_1191), .air_in(c_12_0));
valve v_12_2383 (.fluid_in(k_12_2383), .fluid_out(k_11_1191), .air_in(c_12_1));
valve v_12_2384 (.fluid_in(k_12_2384), .fluid_out(k_11_1192), .air_in(c_12_0));
valve v_12_2385 (.fluid_in(k_12_2385), .fluid_out(k_11_1192), .air_in(c_12_1));
valve v_12_2386 (.fluid_in(k_12_2386), .fluid_out(k_11_1193), .air_in(c_12_0));
valve v_12_2387 (.fluid_in(k_12_2387), .fluid_out(k_11_1193), .air_in(c_12_1));
valve v_12_2388 (.fluid_in(k_12_2388), .fluid_out(k_11_1194), .air_in(c_12_0));
valve v_12_2389 (.fluid_in(k_12_2389), .fluid_out(k_11_1194), .air_in(c_12_1));
valve v_12_2390 (.fluid_in(k_12_2390), .fluid_out(k_11_1195), .air_in(c_12_0));
valve v_12_2391 (.fluid_in(k_12_2391), .fluid_out(k_11_1195), .air_in(c_12_1));
valve v_12_2392 (.fluid_in(k_12_2392), .fluid_out(k_11_1196), .air_in(c_12_0));
valve v_12_2393 (.fluid_in(k_12_2393), .fluid_out(k_11_1196), .air_in(c_12_1));
valve v_12_2394 (.fluid_in(k_12_2394), .fluid_out(k_11_1197), .air_in(c_12_0));
valve v_12_2395 (.fluid_in(k_12_2395), .fluid_out(k_11_1197), .air_in(c_12_1));
valve v_12_2396 (.fluid_in(k_12_2396), .fluid_out(k_11_1198), .air_in(c_12_0));
valve v_12_2397 (.fluid_in(k_12_2397), .fluid_out(k_11_1198), .air_in(c_12_1));
valve v_12_2398 (.fluid_in(k_12_2398), .fluid_out(k_11_1199), .air_in(c_12_0));
valve v_12_2399 (.fluid_in(k_12_2399), .fluid_out(k_11_1199), .air_in(c_12_1));
valve v_12_2400 (.fluid_in(k_12_2400), .fluid_out(k_11_1200), .air_in(c_12_0));
valve v_12_2401 (.fluid_in(k_12_2401), .fluid_out(k_11_1200), .air_in(c_12_1));
valve v_12_2402 (.fluid_in(k_12_2402), .fluid_out(k_11_1201), .air_in(c_12_0));
valve v_12_2403 (.fluid_in(k_12_2403), .fluid_out(k_11_1201), .air_in(c_12_1));
valve v_12_2404 (.fluid_in(k_12_2404), .fluid_out(k_11_1202), .air_in(c_12_0));
valve v_12_2405 (.fluid_in(k_12_2405), .fluid_out(k_11_1202), .air_in(c_12_1));
valve v_12_2406 (.fluid_in(k_12_2406), .fluid_out(k_11_1203), .air_in(c_12_0));
valve v_12_2407 (.fluid_in(k_12_2407), .fluid_out(k_11_1203), .air_in(c_12_1));
valve v_12_2408 (.fluid_in(k_12_2408), .fluid_out(k_11_1204), .air_in(c_12_0));
valve v_12_2409 (.fluid_in(k_12_2409), .fluid_out(k_11_1204), .air_in(c_12_1));
valve v_12_2410 (.fluid_in(k_12_2410), .fluid_out(k_11_1205), .air_in(c_12_0));
valve v_12_2411 (.fluid_in(k_12_2411), .fluid_out(k_11_1205), .air_in(c_12_1));
valve v_12_2412 (.fluid_in(k_12_2412), .fluid_out(k_11_1206), .air_in(c_12_0));
valve v_12_2413 (.fluid_in(k_12_2413), .fluid_out(k_11_1206), .air_in(c_12_1));
valve v_12_2414 (.fluid_in(k_12_2414), .fluid_out(k_11_1207), .air_in(c_12_0));
valve v_12_2415 (.fluid_in(k_12_2415), .fluid_out(k_11_1207), .air_in(c_12_1));
valve v_12_2416 (.fluid_in(k_12_2416), .fluid_out(k_11_1208), .air_in(c_12_0));
valve v_12_2417 (.fluid_in(k_12_2417), .fluid_out(k_11_1208), .air_in(c_12_1));
valve v_12_2418 (.fluid_in(k_12_2418), .fluid_out(k_11_1209), .air_in(c_12_0));
valve v_12_2419 (.fluid_in(k_12_2419), .fluid_out(k_11_1209), .air_in(c_12_1));
valve v_12_2420 (.fluid_in(k_12_2420), .fluid_out(k_11_1210), .air_in(c_12_0));
valve v_12_2421 (.fluid_in(k_12_2421), .fluid_out(k_11_1210), .air_in(c_12_1));
valve v_12_2422 (.fluid_in(k_12_2422), .fluid_out(k_11_1211), .air_in(c_12_0));
valve v_12_2423 (.fluid_in(k_12_2423), .fluid_out(k_11_1211), .air_in(c_12_1));
valve v_12_2424 (.fluid_in(k_12_2424), .fluid_out(k_11_1212), .air_in(c_12_0));
valve v_12_2425 (.fluid_in(k_12_2425), .fluid_out(k_11_1212), .air_in(c_12_1));
valve v_12_2426 (.fluid_in(k_12_2426), .fluid_out(k_11_1213), .air_in(c_12_0));
valve v_12_2427 (.fluid_in(k_12_2427), .fluid_out(k_11_1213), .air_in(c_12_1));
valve v_12_2428 (.fluid_in(k_12_2428), .fluid_out(k_11_1214), .air_in(c_12_0));
valve v_12_2429 (.fluid_in(k_12_2429), .fluid_out(k_11_1214), .air_in(c_12_1));
valve v_12_2430 (.fluid_in(k_12_2430), .fluid_out(k_11_1215), .air_in(c_12_0));
valve v_12_2431 (.fluid_in(k_12_2431), .fluid_out(k_11_1215), .air_in(c_12_1));
valve v_12_2432 (.fluid_in(k_12_2432), .fluid_out(k_11_1216), .air_in(c_12_0));
valve v_12_2433 (.fluid_in(k_12_2433), .fluid_out(k_11_1216), .air_in(c_12_1));
valve v_12_2434 (.fluid_in(k_12_2434), .fluid_out(k_11_1217), .air_in(c_12_0));
valve v_12_2435 (.fluid_in(k_12_2435), .fluid_out(k_11_1217), .air_in(c_12_1));
valve v_12_2436 (.fluid_in(k_12_2436), .fluid_out(k_11_1218), .air_in(c_12_0));
valve v_12_2437 (.fluid_in(k_12_2437), .fluid_out(k_11_1218), .air_in(c_12_1));
valve v_12_2438 (.fluid_in(k_12_2438), .fluid_out(k_11_1219), .air_in(c_12_0));
valve v_12_2439 (.fluid_in(k_12_2439), .fluid_out(k_11_1219), .air_in(c_12_1));
valve v_12_2440 (.fluid_in(k_12_2440), .fluid_out(k_11_1220), .air_in(c_12_0));
valve v_12_2441 (.fluid_in(k_12_2441), .fluid_out(k_11_1220), .air_in(c_12_1));
valve v_12_2442 (.fluid_in(k_12_2442), .fluid_out(k_11_1221), .air_in(c_12_0));
valve v_12_2443 (.fluid_in(k_12_2443), .fluid_out(k_11_1221), .air_in(c_12_1));
valve v_12_2444 (.fluid_in(k_12_2444), .fluid_out(k_11_1222), .air_in(c_12_0));
valve v_12_2445 (.fluid_in(k_12_2445), .fluid_out(k_11_1222), .air_in(c_12_1));
valve v_12_2446 (.fluid_in(k_12_2446), .fluid_out(k_11_1223), .air_in(c_12_0));
valve v_12_2447 (.fluid_in(k_12_2447), .fluid_out(k_11_1223), .air_in(c_12_1));
valve v_12_2448 (.fluid_in(k_12_2448), .fluid_out(k_11_1224), .air_in(c_12_0));
valve v_12_2449 (.fluid_in(k_12_2449), .fluid_out(k_11_1224), .air_in(c_12_1));
valve v_12_2450 (.fluid_in(k_12_2450), .fluid_out(k_11_1225), .air_in(c_12_0));
valve v_12_2451 (.fluid_in(k_12_2451), .fluid_out(k_11_1225), .air_in(c_12_1));
valve v_12_2452 (.fluid_in(k_12_2452), .fluid_out(k_11_1226), .air_in(c_12_0));
valve v_12_2453 (.fluid_in(k_12_2453), .fluid_out(k_11_1226), .air_in(c_12_1));
valve v_12_2454 (.fluid_in(k_12_2454), .fluid_out(k_11_1227), .air_in(c_12_0));
valve v_12_2455 (.fluid_in(k_12_2455), .fluid_out(k_11_1227), .air_in(c_12_1));
valve v_12_2456 (.fluid_in(k_12_2456), .fluid_out(k_11_1228), .air_in(c_12_0));
valve v_12_2457 (.fluid_in(k_12_2457), .fluid_out(k_11_1228), .air_in(c_12_1));
valve v_12_2458 (.fluid_in(k_12_2458), .fluid_out(k_11_1229), .air_in(c_12_0));
valve v_12_2459 (.fluid_in(k_12_2459), .fluid_out(k_11_1229), .air_in(c_12_1));
valve v_12_2460 (.fluid_in(k_12_2460), .fluid_out(k_11_1230), .air_in(c_12_0));
valve v_12_2461 (.fluid_in(k_12_2461), .fluid_out(k_11_1230), .air_in(c_12_1));
valve v_12_2462 (.fluid_in(k_12_2462), .fluid_out(k_11_1231), .air_in(c_12_0));
valve v_12_2463 (.fluid_in(k_12_2463), .fluid_out(k_11_1231), .air_in(c_12_1));
valve v_12_2464 (.fluid_in(k_12_2464), .fluid_out(k_11_1232), .air_in(c_12_0));
valve v_12_2465 (.fluid_in(k_12_2465), .fluid_out(k_11_1232), .air_in(c_12_1));
valve v_12_2466 (.fluid_in(k_12_2466), .fluid_out(k_11_1233), .air_in(c_12_0));
valve v_12_2467 (.fluid_in(k_12_2467), .fluid_out(k_11_1233), .air_in(c_12_1));
valve v_12_2468 (.fluid_in(k_12_2468), .fluid_out(k_11_1234), .air_in(c_12_0));
valve v_12_2469 (.fluid_in(k_12_2469), .fluid_out(k_11_1234), .air_in(c_12_1));
valve v_12_2470 (.fluid_in(k_12_2470), .fluid_out(k_11_1235), .air_in(c_12_0));
valve v_12_2471 (.fluid_in(k_12_2471), .fluid_out(k_11_1235), .air_in(c_12_1));
valve v_12_2472 (.fluid_in(k_12_2472), .fluid_out(k_11_1236), .air_in(c_12_0));
valve v_12_2473 (.fluid_in(k_12_2473), .fluid_out(k_11_1236), .air_in(c_12_1));
valve v_12_2474 (.fluid_in(k_12_2474), .fluid_out(k_11_1237), .air_in(c_12_0));
valve v_12_2475 (.fluid_in(k_12_2475), .fluid_out(k_11_1237), .air_in(c_12_1));
valve v_12_2476 (.fluid_in(k_12_2476), .fluid_out(k_11_1238), .air_in(c_12_0));
valve v_12_2477 (.fluid_in(k_12_2477), .fluid_out(k_11_1238), .air_in(c_12_1));
valve v_12_2478 (.fluid_in(k_12_2478), .fluid_out(k_11_1239), .air_in(c_12_0));
valve v_12_2479 (.fluid_in(k_12_2479), .fluid_out(k_11_1239), .air_in(c_12_1));
valve v_12_2480 (.fluid_in(k_12_2480), .fluid_out(k_11_1240), .air_in(c_12_0));
valve v_12_2481 (.fluid_in(k_12_2481), .fluid_out(k_11_1240), .air_in(c_12_1));
valve v_12_2482 (.fluid_in(k_12_2482), .fluid_out(k_11_1241), .air_in(c_12_0));
valve v_12_2483 (.fluid_in(k_12_2483), .fluid_out(k_11_1241), .air_in(c_12_1));
valve v_12_2484 (.fluid_in(k_12_2484), .fluid_out(k_11_1242), .air_in(c_12_0));
valve v_12_2485 (.fluid_in(k_12_2485), .fluid_out(k_11_1242), .air_in(c_12_1));
valve v_12_2486 (.fluid_in(k_12_2486), .fluid_out(k_11_1243), .air_in(c_12_0));
valve v_12_2487 (.fluid_in(k_12_2487), .fluid_out(k_11_1243), .air_in(c_12_1));
valve v_12_2488 (.fluid_in(k_12_2488), .fluid_out(k_11_1244), .air_in(c_12_0));
valve v_12_2489 (.fluid_in(k_12_2489), .fluid_out(k_11_1244), .air_in(c_12_1));
valve v_12_2490 (.fluid_in(k_12_2490), .fluid_out(k_11_1245), .air_in(c_12_0));
valve v_12_2491 (.fluid_in(k_12_2491), .fluid_out(k_11_1245), .air_in(c_12_1));
valve v_12_2492 (.fluid_in(k_12_2492), .fluid_out(k_11_1246), .air_in(c_12_0));
valve v_12_2493 (.fluid_in(k_12_2493), .fluid_out(k_11_1246), .air_in(c_12_1));
valve v_12_2494 (.fluid_in(k_12_2494), .fluid_out(k_11_1247), .air_in(c_12_0));
valve v_12_2495 (.fluid_in(k_12_2495), .fluid_out(k_11_1247), .air_in(c_12_1));
valve v_12_2496 (.fluid_in(k_12_2496), .fluid_out(k_11_1248), .air_in(c_12_0));
valve v_12_2497 (.fluid_in(k_12_2497), .fluid_out(k_11_1248), .air_in(c_12_1));
valve v_12_2498 (.fluid_in(k_12_2498), .fluid_out(k_11_1249), .air_in(c_12_0));
valve v_12_2499 (.fluid_in(k_12_2499), .fluid_out(k_11_1249), .air_in(c_12_1));
valve v_12_2500 (.fluid_in(k_12_2500), .fluid_out(k_11_1250), .air_in(c_12_0));
valve v_12_2501 (.fluid_in(k_12_2501), .fluid_out(k_11_1250), .air_in(c_12_1));
valve v_12_2502 (.fluid_in(k_12_2502), .fluid_out(k_11_1251), .air_in(c_12_0));
valve v_12_2503 (.fluid_in(k_12_2503), .fluid_out(k_11_1251), .air_in(c_12_1));
valve v_12_2504 (.fluid_in(k_12_2504), .fluid_out(k_11_1252), .air_in(c_12_0));
valve v_12_2505 (.fluid_in(k_12_2505), .fluid_out(k_11_1252), .air_in(c_12_1));
valve v_12_2506 (.fluid_in(k_12_2506), .fluid_out(k_11_1253), .air_in(c_12_0));
valve v_12_2507 (.fluid_in(k_12_2507), .fluid_out(k_11_1253), .air_in(c_12_1));
valve v_12_2508 (.fluid_in(k_12_2508), .fluid_out(k_11_1254), .air_in(c_12_0));
valve v_12_2509 (.fluid_in(k_12_2509), .fluid_out(k_11_1254), .air_in(c_12_1));
valve v_12_2510 (.fluid_in(k_12_2510), .fluid_out(k_11_1255), .air_in(c_12_0));
valve v_12_2511 (.fluid_in(k_12_2511), .fluid_out(k_11_1255), .air_in(c_12_1));
valve v_12_2512 (.fluid_in(k_12_2512), .fluid_out(k_11_1256), .air_in(c_12_0));
valve v_12_2513 (.fluid_in(k_12_2513), .fluid_out(k_11_1256), .air_in(c_12_1));
valve v_12_2514 (.fluid_in(k_12_2514), .fluid_out(k_11_1257), .air_in(c_12_0));
valve v_12_2515 (.fluid_in(k_12_2515), .fluid_out(k_11_1257), .air_in(c_12_1));
valve v_12_2516 (.fluid_in(k_12_2516), .fluid_out(k_11_1258), .air_in(c_12_0));
valve v_12_2517 (.fluid_in(k_12_2517), .fluid_out(k_11_1258), .air_in(c_12_1));
valve v_12_2518 (.fluid_in(k_12_2518), .fluid_out(k_11_1259), .air_in(c_12_0));
valve v_12_2519 (.fluid_in(k_12_2519), .fluid_out(k_11_1259), .air_in(c_12_1));
valve v_12_2520 (.fluid_in(k_12_2520), .fluid_out(k_11_1260), .air_in(c_12_0));
valve v_12_2521 (.fluid_in(k_12_2521), .fluid_out(k_11_1260), .air_in(c_12_1));
valve v_12_2522 (.fluid_in(k_12_2522), .fluid_out(k_11_1261), .air_in(c_12_0));
valve v_12_2523 (.fluid_in(k_12_2523), .fluid_out(k_11_1261), .air_in(c_12_1));
valve v_12_2524 (.fluid_in(k_12_2524), .fluid_out(k_11_1262), .air_in(c_12_0));
valve v_12_2525 (.fluid_in(k_12_2525), .fluid_out(k_11_1262), .air_in(c_12_1));
valve v_12_2526 (.fluid_in(k_12_2526), .fluid_out(k_11_1263), .air_in(c_12_0));
valve v_12_2527 (.fluid_in(k_12_2527), .fluid_out(k_11_1263), .air_in(c_12_1));
valve v_12_2528 (.fluid_in(k_12_2528), .fluid_out(k_11_1264), .air_in(c_12_0));
valve v_12_2529 (.fluid_in(k_12_2529), .fluid_out(k_11_1264), .air_in(c_12_1));
valve v_12_2530 (.fluid_in(k_12_2530), .fluid_out(k_11_1265), .air_in(c_12_0));
valve v_12_2531 (.fluid_in(k_12_2531), .fluid_out(k_11_1265), .air_in(c_12_1));
valve v_12_2532 (.fluid_in(k_12_2532), .fluid_out(k_11_1266), .air_in(c_12_0));
valve v_12_2533 (.fluid_in(k_12_2533), .fluid_out(k_11_1266), .air_in(c_12_1));
valve v_12_2534 (.fluid_in(k_12_2534), .fluid_out(k_11_1267), .air_in(c_12_0));
valve v_12_2535 (.fluid_in(k_12_2535), .fluid_out(k_11_1267), .air_in(c_12_1));
valve v_12_2536 (.fluid_in(k_12_2536), .fluid_out(k_11_1268), .air_in(c_12_0));
valve v_12_2537 (.fluid_in(k_12_2537), .fluid_out(k_11_1268), .air_in(c_12_1));
valve v_12_2538 (.fluid_in(k_12_2538), .fluid_out(k_11_1269), .air_in(c_12_0));
valve v_12_2539 (.fluid_in(k_12_2539), .fluid_out(k_11_1269), .air_in(c_12_1));
valve v_12_2540 (.fluid_in(k_12_2540), .fluid_out(k_11_1270), .air_in(c_12_0));
valve v_12_2541 (.fluid_in(k_12_2541), .fluid_out(k_11_1270), .air_in(c_12_1));
valve v_12_2542 (.fluid_in(k_12_2542), .fluid_out(k_11_1271), .air_in(c_12_0));
valve v_12_2543 (.fluid_in(k_12_2543), .fluid_out(k_11_1271), .air_in(c_12_1));
valve v_12_2544 (.fluid_in(k_12_2544), .fluid_out(k_11_1272), .air_in(c_12_0));
valve v_12_2545 (.fluid_in(k_12_2545), .fluid_out(k_11_1272), .air_in(c_12_1));
valve v_12_2546 (.fluid_in(k_12_2546), .fluid_out(k_11_1273), .air_in(c_12_0));
valve v_12_2547 (.fluid_in(k_12_2547), .fluid_out(k_11_1273), .air_in(c_12_1));
valve v_12_2548 (.fluid_in(k_12_2548), .fluid_out(k_11_1274), .air_in(c_12_0));
valve v_12_2549 (.fluid_in(k_12_2549), .fluid_out(k_11_1274), .air_in(c_12_1));
valve v_12_2550 (.fluid_in(k_12_2550), .fluid_out(k_11_1275), .air_in(c_12_0));
valve v_12_2551 (.fluid_in(k_12_2551), .fluid_out(k_11_1275), .air_in(c_12_1));
valve v_12_2552 (.fluid_in(k_12_2552), .fluid_out(k_11_1276), .air_in(c_12_0));
valve v_12_2553 (.fluid_in(k_12_2553), .fluid_out(k_11_1276), .air_in(c_12_1));
valve v_12_2554 (.fluid_in(k_12_2554), .fluid_out(k_11_1277), .air_in(c_12_0));
valve v_12_2555 (.fluid_in(k_12_2555), .fluid_out(k_11_1277), .air_in(c_12_1));
valve v_12_2556 (.fluid_in(k_12_2556), .fluid_out(k_11_1278), .air_in(c_12_0));
valve v_12_2557 (.fluid_in(k_12_2557), .fluid_out(k_11_1278), .air_in(c_12_1));
valve v_12_2558 (.fluid_in(k_12_2558), .fluid_out(k_11_1279), .air_in(c_12_0));
valve v_12_2559 (.fluid_in(k_12_2559), .fluid_out(k_11_1279), .air_in(c_12_1));
valve v_12_2560 (.fluid_in(k_12_2560), .fluid_out(k_11_1280), .air_in(c_12_0));
valve v_12_2561 (.fluid_in(k_12_2561), .fluid_out(k_11_1280), .air_in(c_12_1));
valve v_12_2562 (.fluid_in(k_12_2562), .fluid_out(k_11_1281), .air_in(c_12_0));
valve v_12_2563 (.fluid_in(k_12_2563), .fluid_out(k_11_1281), .air_in(c_12_1));
valve v_12_2564 (.fluid_in(k_12_2564), .fluid_out(k_11_1282), .air_in(c_12_0));
valve v_12_2565 (.fluid_in(k_12_2565), .fluid_out(k_11_1282), .air_in(c_12_1));
valve v_12_2566 (.fluid_in(k_12_2566), .fluid_out(k_11_1283), .air_in(c_12_0));
valve v_12_2567 (.fluid_in(k_12_2567), .fluid_out(k_11_1283), .air_in(c_12_1));
valve v_12_2568 (.fluid_in(k_12_2568), .fluid_out(k_11_1284), .air_in(c_12_0));
valve v_12_2569 (.fluid_in(k_12_2569), .fluid_out(k_11_1284), .air_in(c_12_1));
valve v_12_2570 (.fluid_in(k_12_2570), .fluid_out(k_11_1285), .air_in(c_12_0));
valve v_12_2571 (.fluid_in(k_12_2571), .fluid_out(k_11_1285), .air_in(c_12_1));
valve v_12_2572 (.fluid_in(k_12_2572), .fluid_out(k_11_1286), .air_in(c_12_0));
valve v_12_2573 (.fluid_in(k_12_2573), .fluid_out(k_11_1286), .air_in(c_12_1));
valve v_12_2574 (.fluid_in(k_12_2574), .fluid_out(k_11_1287), .air_in(c_12_0));
valve v_12_2575 (.fluid_in(k_12_2575), .fluid_out(k_11_1287), .air_in(c_12_1));
valve v_12_2576 (.fluid_in(k_12_2576), .fluid_out(k_11_1288), .air_in(c_12_0));
valve v_12_2577 (.fluid_in(k_12_2577), .fluid_out(k_11_1288), .air_in(c_12_1));
valve v_12_2578 (.fluid_in(k_12_2578), .fluid_out(k_11_1289), .air_in(c_12_0));
valve v_12_2579 (.fluid_in(k_12_2579), .fluid_out(k_11_1289), .air_in(c_12_1));
valve v_12_2580 (.fluid_in(k_12_2580), .fluid_out(k_11_1290), .air_in(c_12_0));
valve v_12_2581 (.fluid_in(k_12_2581), .fluid_out(k_11_1290), .air_in(c_12_1));
valve v_12_2582 (.fluid_in(k_12_2582), .fluid_out(k_11_1291), .air_in(c_12_0));
valve v_12_2583 (.fluid_in(k_12_2583), .fluid_out(k_11_1291), .air_in(c_12_1));
valve v_12_2584 (.fluid_in(k_12_2584), .fluid_out(k_11_1292), .air_in(c_12_0));
valve v_12_2585 (.fluid_in(k_12_2585), .fluid_out(k_11_1292), .air_in(c_12_1));
valve v_12_2586 (.fluid_in(k_12_2586), .fluid_out(k_11_1293), .air_in(c_12_0));
valve v_12_2587 (.fluid_in(k_12_2587), .fluid_out(k_11_1293), .air_in(c_12_1));
valve v_12_2588 (.fluid_in(k_12_2588), .fluid_out(k_11_1294), .air_in(c_12_0));
valve v_12_2589 (.fluid_in(k_12_2589), .fluid_out(k_11_1294), .air_in(c_12_1));
valve v_12_2590 (.fluid_in(k_12_2590), .fluid_out(k_11_1295), .air_in(c_12_0));
valve v_12_2591 (.fluid_in(k_12_2591), .fluid_out(k_11_1295), .air_in(c_12_1));
valve v_12_2592 (.fluid_in(k_12_2592), .fluid_out(k_11_1296), .air_in(c_12_0));
valve v_12_2593 (.fluid_in(k_12_2593), .fluid_out(k_11_1296), .air_in(c_12_1));
valve v_12_2594 (.fluid_in(k_12_2594), .fluid_out(k_11_1297), .air_in(c_12_0));
valve v_12_2595 (.fluid_in(k_12_2595), .fluid_out(k_11_1297), .air_in(c_12_1));
valve v_12_2596 (.fluid_in(k_12_2596), .fluid_out(k_11_1298), .air_in(c_12_0));
valve v_12_2597 (.fluid_in(k_12_2597), .fluid_out(k_11_1298), .air_in(c_12_1));
valve v_12_2598 (.fluid_in(k_12_2598), .fluid_out(k_11_1299), .air_in(c_12_0));
valve v_12_2599 (.fluid_in(k_12_2599), .fluid_out(k_11_1299), .air_in(c_12_1));
valve v_12_2600 (.fluid_in(k_12_2600), .fluid_out(k_11_1300), .air_in(c_12_0));
valve v_12_2601 (.fluid_in(k_12_2601), .fluid_out(k_11_1300), .air_in(c_12_1));
valve v_12_2602 (.fluid_in(k_12_2602), .fluid_out(k_11_1301), .air_in(c_12_0));
valve v_12_2603 (.fluid_in(k_12_2603), .fluid_out(k_11_1301), .air_in(c_12_1));
valve v_12_2604 (.fluid_in(k_12_2604), .fluid_out(k_11_1302), .air_in(c_12_0));
valve v_12_2605 (.fluid_in(k_12_2605), .fluid_out(k_11_1302), .air_in(c_12_1));
valve v_12_2606 (.fluid_in(k_12_2606), .fluid_out(k_11_1303), .air_in(c_12_0));
valve v_12_2607 (.fluid_in(k_12_2607), .fluid_out(k_11_1303), .air_in(c_12_1));
valve v_12_2608 (.fluid_in(k_12_2608), .fluid_out(k_11_1304), .air_in(c_12_0));
valve v_12_2609 (.fluid_in(k_12_2609), .fluid_out(k_11_1304), .air_in(c_12_1));
valve v_12_2610 (.fluid_in(k_12_2610), .fluid_out(k_11_1305), .air_in(c_12_0));
valve v_12_2611 (.fluid_in(k_12_2611), .fluid_out(k_11_1305), .air_in(c_12_1));
valve v_12_2612 (.fluid_in(k_12_2612), .fluid_out(k_11_1306), .air_in(c_12_0));
valve v_12_2613 (.fluid_in(k_12_2613), .fluid_out(k_11_1306), .air_in(c_12_1));
valve v_12_2614 (.fluid_in(k_12_2614), .fluid_out(k_11_1307), .air_in(c_12_0));
valve v_12_2615 (.fluid_in(k_12_2615), .fluid_out(k_11_1307), .air_in(c_12_1));
valve v_12_2616 (.fluid_in(k_12_2616), .fluid_out(k_11_1308), .air_in(c_12_0));
valve v_12_2617 (.fluid_in(k_12_2617), .fluid_out(k_11_1308), .air_in(c_12_1));
valve v_12_2618 (.fluid_in(k_12_2618), .fluid_out(k_11_1309), .air_in(c_12_0));
valve v_12_2619 (.fluid_in(k_12_2619), .fluid_out(k_11_1309), .air_in(c_12_1));
valve v_12_2620 (.fluid_in(k_12_2620), .fluid_out(k_11_1310), .air_in(c_12_0));
valve v_12_2621 (.fluid_in(k_12_2621), .fluid_out(k_11_1310), .air_in(c_12_1));
valve v_12_2622 (.fluid_in(k_12_2622), .fluid_out(k_11_1311), .air_in(c_12_0));
valve v_12_2623 (.fluid_in(k_12_2623), .fluid_out(k_11_1311), .air_in(c_12_1));
valve v_12_2624 (.fluid_in(k_12_2624), .fluid_out(k_11_1312), .air_in(c_12_0));
valve v_12_2625 (.fluid_in(k_12_2625), .fluid_out(k_11_1312), .air_in(c_12_1));
valve v_12_2626 (.fluid_in(k_12_2626), .fluid_out(k_11_1313), .air_in(c_12_0));
valve v_12_2627 (.fluid_in(k_12_2627), .fluid_out(k_11_1313), .air_in(c_12_1));
valve v_12_2628 (.fluid_in(k_12_2628), .fluid_out(k_11_1314), .air_in(c_12_0));
valve v_12_2629 (.fluid_in(k_12_2629), .fluid_out(k_11_1314), .air_in(c_12_1));
valve v_12_2630 (.fluid_in(k_12_2630), .fluid_out(k_11_1315), .air_in(c_12_0));
valve v_12_2631 (.fluid_in(k_12_2631), .fluid_out(k_11_1315), .air_in(c_12_1));
valve v_12_2632 (.fluid_in(k_12_2632), .fluid_out(k_11_1316), .air_in(c_12_0));
valve v_12_2633 (.fluid_in(k_12_2633), .fluid_out(k_11_1316), .air_in(c_12_1));
valve v_12_2634 (.fluid_in(k_12_2634), .fluid_out(k_11_1317), .air_in(c_12_0));
valve v_12_2635 (.fluid_in(k_12_2635), .fluid_out(k_11_1317), .air_in(c_12_1));
valve v_12_2636 (.fluid_in(k_12_2636), .fluid_out(k_11_1318), .air_in(c_12_0));
valve v_12_2637 (.fluid_in(k_12_2637), .fluid_out(k_11_1318), .air_in(c_12_1));
valve v_12_2638 (.fluid_in(k_12_2638), .fluid_out(k_11_1319), .air_in(c_12_0));
valve v_12_2639 (.fluid_in(k_12_2639), .fluid_out(k_11_1319), .air_in(c_12_1));
valve v_12_2640 (.fluid_in(k_12_2640), .fluid_out(k_11_1320), .air_in(c_12_0));
valve v_12_2641 (.fluid_in(k_12_2641), .fluid_out(k_11_1320), .air_in(c_12_1));
valve v_12_2642 (.fluid_in(k_12_2642), .fluid_out(k_11_1321), .air_in(c_12_0));
valve v_12_2643 (.fluid_in(k_12_2643), .fluid_out(k_11_1321), .air_in(c_12_1));
valve v_12_2644 (.fluid_in(k_12_2644), .fluid_out(k_11_1322), .air_in(c_12_0));
valve v_12_2645 (.fluid_in(k_12_2645), .fluid_out(k_11_1322), .air_in(c_12_1));
valve v_12_2646 (.fluid_in(k_12_2646), .fluid_out(k_11_1323), .air_in(c_12_0));
valve v_12_2647 (.fluid_in(k_12_2647), .fluid_out(k_11_1323), .air_in(c_12_1));
valve v_12_2648 (.fluid_in(k_12_2648), .fluid_out(k_11_1324), .air_in(c_12_0));
valve v_12_2649 (.fluid_in(k_12_2649), .fluid_out(k_11_1324), .air_in(c_12_1));
valve v_12_2650 (.fluid_in(k_12_2650), .fluid_out(k_11_1325), .air_in(c_12_0));
valve v_12_2651 (.fluid_in(k_12_2651), .fluid_out(k_11_1325), .air_in(c_12_1));
valve v_12_2652 (.fluid_in(k_12_2652), .fluid_out(k_11_1326), .air_in(c_12_0));
valve v_12_2653 (.fluid_in(k_12_2653), .fluid_out(k_11_1326), .air_in(c_12_1));
valve v_12_2654 (.fluid_in(k_12_2654), .fluid_out(k_11_1327), .air_in(c_12_0));
valve v_12_2655 (.fluid_in(k_12_2655), .fluid_out(k_11_1327), .air_in(c_12_1));
valve v_12_2656 (.fluid_in(k_12_2656), .fluid_out(k_11_1328), .air_in(c_12_0));
valve v_12_2657 (.fluid_in(k_12_2657), .fluid_out(k_11_1328), .air_in(c_12_1));
valve v_12_2658 (.fluid_in(k_12_2658), .fluid_out(k_11_1329), .air_in(c_12_0));
valve v_12_2659 (.fluid_in(k_12_2659), .fluid_out(k_11_1329), .air_in(c_12_1));
valve v_12_2660 (.fluid_in(k_12_2660), .fluid_out(k_11_1330), .air_in(c_12_0));
valve v_12_2661 (.fluid_in(k_12_2661), .fluid_out(k_11_1330), .air_in(c_12_1));
valve v_12_2662 (.fluid_in(k_12_2662), .fluid_out(k_11_1331), .air_in(c_12_0));
valve v_12_2663 (.fluid_in(k_12_2663), .fluid_out(k_11_1331), .air_in(c_12_1));
valve v_12_2664 (.fluid_in(k_12_2664), .fluid_out(k_11_1332), .air_in(c_12_0));
valve v_12_2665 (.fluid_in(k_12_2665), .fluid_out(k_11_1332), .air_in(c_12_1));
valve v_12_2666 (.fluid_in(k_12_2666), .fluid_out(k_11_1333), .air_in(c_12_0));
valve v_12_2667 (.fluid_in(k_12_2667), .fluid_out(k_11_1333), .air_in(c_12_1));
valve v_12_2668 (.fluid_in(k_12_2668), .fluid_out(k_11_1334), .air_in(c_12_0));
valve v_12_2669 (.fluid_in(k_12_2669), .fluid_out(k_11_1334), .air_in(c_12_1));
valve v_12_2670 (.fluid_in(k_12_2670), .fluid_out(k_11_1335), .air_in(c_12_0));
valve v_12_2671 (.fluid_in(k_12_2671), .fluid_out(k_11_1335), .air_in(c_12_1));
valve v_12_2672 (.fluid_in(k_12_2672), .fluid_out(k_11_1336), .air_in(c_12_0));
valve v_12_2673 (.fluid_in(k_12_2673), .fluid_out(k_11_1336), .air_in(c_12_1));
valve v_12_2674 (.fluid_in(k_12_2674), .fluid_out(k_11_1337), .air_in(c_12_0));
valve v_12_2675 (.fluid_in(k_12_2675), .fluid_out(k_11_1337), .air_in(c_12_1));
valve v_12_2676 (.fluid_in(k_12_2676), .fluid_out(k_11_1338), .air_in(c_12_0));
valve v_12_2677 (.fluid_in(k_12_2677), .fluid_out(k_11_1338), .air_in(c_12_1));
valve v_12_2678 (.fluid_in(k_12_2678), .fluid_out(k_11_1339), .air_in(c_12_0));
valve v_12_2679 (.fluid_in(k_12_2679), .fluid_out(k_11_1339), .air_in(c_12_1));
valve v_12_2680 (.fluid_in(k_12_2680), .fluid_out(k_11_1340), .air_in(c_12_0));
valve v_12_2681 (.fluid_in(k_12_2681), .fluid_out(k_11_1340), .air_in(c_12_1));
valve v_12_2682 (.fluid_in(k_12_2682), .fluid_out(k_11_1341), .air_in(c_12_0));
valve v_12_2683 (.fluid_in(k_12_2683), .fluid_out(k_11_1341), .air_in(c_12_1));
valve v_12_2684 (.fluid_in(k_12_2684), .fluid_out(k_11_1342), .air_in(c_12_0));
valve v_12_2685 (.fluid_in(k_12_2685), .fluid_out(k_11_1342), .air_in(c_12_1));
valve v_12_2686 (.fluid_in(k_12_2686), .fluid_out(k_11_1343), .air_in(c_12_0));
valve v_12_2687 (.fluid_in(k_12_2687), .fluid_out(k_11_1343), .air_in(c_12_1));
valve v_12_2688 (.fluid_in(k_12_2688), .fluid_out(k_11_1344), .air_in(c_12_0));
valve v_12_2689 (.fluid_in(k_12_2689), .fluid_out(k_11_1344), .air_in(c_12_1));
valve v_12_2690 (.fluid_in(k_12_2690), .fluid_out(k_11_1345), .air_in(c_12_0));
valve v_12_2691 (.fluid_in(k_12_2691), .fluid_out(k_11_1345), .air_in(c_12_1));
valve v_12_2692 (.fluid_in(k_12_2692), .fluid_out(k_11_1346), .air_in(c_12_0));
valve v_12_2693 (.fluid_in(k_12_2693), .fluid_out(k_11_1346), .air_in(c_12_1));
valve v_12_2694 (.fluid_in(k_12_2694), .fluid_out(k_11_1347), .air_in(c_12_0));
valve v_12_2695 (.fluid_in(k_12_2695), .fluid_out(k_11_1347), .air_in(c_12_1));
valve v_12_2696 (.fluid_in(k_12_2696), .fluid_out(k_11_1348), .air_in(c_12_0));
valve v_12_2697 (.fluid_in(k_12_2697), .fluid_out(k_11_1348), .air_in(c_12_1));
valve v_12_2698 (.fluid_in(k_12_2698), .fluid_out(k_11_1349), .air_in(c_12_0));
valve v_12_2699 (.fluid_in(k_12_2699), .fluid_out(k_11_1349), .air_in(c_12_1));
valve v_12_2700 (.fluid_in(k_12_2700), .fluid_out(k_11_1350), .air_in(c_12_0));
valve v_12_2701 (.fluid_in(k_12_2701), .fluid_out(k_11_1350), .air_in(c_12_1));
valve v_12_2702 (.fluid_in(k_12_2702), .fluid_out(k_11_1351), .air_in(c_12_0));
valve v_12_2703 (.fluid_in(k_12_2703), .fluid_out(k_11_1351), .air_in(c_12_1));
valve v_12_2704 (.fluid_in(k_12_2704), .fluid_out(k_11_1352), .air_in(c_12_0));
valve v_12_2705 (.fluid_in(k_12_2705), .fluid_out(k_11_1352), .air_in(c_12_1));
valve v_12_2706 (.fluid_in(k_12_2706), .fluid_out(k_11_1353), .air_in(c_12_0));
valve v_12_2707 (.fluid_in(k_12_2707), .fluid_out(k_11_1353), .air_in(c_12_1));
valve v_12_2708 (.fluid_in(k_12_2708), .fluid_out(k_11_1354), .air_in(c_12_0));
valve v_12_2709 (.fluid_in(k_12_2709), .fluid_out(k_11_1354), .air_in(c_12_1));
valve v_12_2710 (.fluid_in(k_12_2710), .fluid_out(k_11_1355), .air_in(c_12_0));
valve v_12_2711 (.fluid_in(k_12_2711), .fluid_out(k_11_1355), .air_in(c_12_1));
valve v_12_2712 (.fluid_in(k_12_2712), .fluid_out(k_11_1356), .air_in(c_12_0));
valve v_12_2713 (.fluid_in(k_12_2713), .fluid_out(k_11_1356), .air_in(c_12_1));
valve v_12_2714 (.fluid_in(k_12_2714), .fluid_out(k_11_1357), .air_in(c_12_0));
valve v_12_2715 (.fluid_in(k_12_2715), .fluid_out(k_11_1357), .air_in(c_12_1));
valve v_12_2716 (.fluid_in(k_12_2716), .fluid_out(k_11_1358), .air_in(c_12_0));
valve v_12_2717 (.fluid_in(k_12_2717), .fluid_out(k_11_1358), .air_in(c_12_1));
valve v_12_2718 (.fluid_in(k_12_2718), .fluid_out(k_11_1359), .air_in(c_12_0));
valve v_12_2719 (.fluid_in(k_12_2719), .fluid_out(k_11_1359), .air_in(c_12_1));
valve v_12_2720 (.fluid_in(k_12_2720), .fluid_out(k_11_1360), .air_in(c_12_0));
valve v_12_2721 (.fluid_in(k_12_2721), .fluid_out(k_11_1360), .air_in(c_12_1));
valve v_12_2722 (.fluid_in(k_12_2722), .fluid_out(k_11_1361), .air_in(c_12_0));
valve v_12_2723 (.fluid_in(k_12_2723), .fluid_out(k_11_1361), .air_in(c_12_1));
valve v_12_2724 (.fluid_in(k_12_2724), .fluid_out(k_11_1362), .air_in(c_12_0));
valve v_12_2725 (.fluid_in(k_12_2725), .fluid_out(k_11_1362), .air_in(c_12_1));
valve v_12_2726 (.fluid_in(k_12_2726), .fluid_out(k_11_1363), .air_in(c_12_0));
valve v_12_2727 (.fluid_in(k_12_2727), .fluid_out(k_11_1363), .air_in(c_12_1));
valve v_12_2728 (.fluid_in(k_12_2728), .fluid_out(k_11_1364), .air_in(c_12_0));
valve v_12_2729 (.fluid_in(k_12_2729), .fluid_out(k_11_1364), .air_in(c_12_1));
valve v_12_2730 (.fluid_in(k_12_2730), .fluid_out(k_11_1365), .air_in(c_12_0));
valve v_12_2731 (.fluid_in(k_12_2731), .fluid_out(k_11_1365), .air_in(c_12_1));
valve v_12_2732 (.fluid_in(k_12_2732), .fluid_out(k_11_1366), .air_in(c_12_0));
valve v_12_2733 (.fluid_in(k_12_2733), .fluid_out(k_11_1366), .air_in(c_12_1));
valve v_12_2734 (.fluid_in(k_12_2734), .fluid_out(k_11_1367), .air_in(c_12_0));
valve v_12_2735 (.fluid_in(k_12_2735), .fluid_out(k_11_1367), .air_in(c_12_1));
valve v_12_2736 (.fluid_in(k_12_2736), .fluid_out(k_11_1368), .air_in(c_12_0));
valve v_12_2737 (.fluid_in(k_12_2737), .fluid_out(k_11_1368), .air_in(c_12_1));
valve v_12_2738 (.fluid_in(k_12_2738), .fluid_out(k_11_1369), .air_in(c_12_0));
valve v_12_2739 (.fluid_in(k_12_2739), .fluid_out(k_11_1369), .air_in(c_12_1));
valve v_12_2740 (.fluid_in(k_12_2740), .fluid_out(k_11_1370), .air_in(c_12_0));
valve v_12_2741 (.fluid_in(k_12_2741), .fluid_out(k_11_1370), .air_in(c_12_1));
valve v_12_2742 (.fluid_in(k_12_2742), .fluid_out(k_11_1371), .air_in(c_12_0));
valve v_12_2743 (.fluid_in(k_12_2743), .fluid_out(k_11_1371), .air_in(c_12_1));
valve v_12_2744 (.fluid_in(k_12_2744), .fluid_out(k_11_1372), .air_in(c_12_0));
valve v_12_2745 (.fluid_in(k_12_2745), .fluid_out(k_11_1372), .air_in(c_12_1));
valve v_12_2746 (.fluid_in(k_12_2746), .fluid_out(k_11_1373), .air_in(c_12_0));
valve v_12_2747 (.fluid_in(k_12_2747), .fluid_out(k_11_1373), .air_in(c_12_1));
valve v_12_2748 (.fluid_in(k_12_2748), .fluid_out(k_11_1374), .air_in(c_12_0));
valve v_12_2749 (.fluid_in(k_12_2749), .fluid_out(k_11_1374), .air_in(c_12_1));
valve v_12_2750 (.fluid_in(k_12_2750), .fluid_out(k_11_1375), .air_in(c_12_0));
valve v_12_2751 (.fluid_in(k_12_2751), .fluid_out(k_11_1375), .air_in(c_12_1));
valve v_12_2752 (.fluid_in(k_12_2752), .fluid_out(k_11_1376), .air_in(c_12_0));
valve v_12_2753 (.fluid_in(k_12_2753), .fluid_out(k_11_1376), .air_in(c_12_1));
valve v_12_2754 (.fluid_in(k_12_2754), .fluid_out(k_11_1377), .air_in(c_12_0));
valve v_12_2755 (.fluid_in(k_12_2755), .fluid_out(k_11_1377), .air_in(c_12_1));
valve v_12_2756 (.fluid_in(k_12_2756), .fluid_out(k_11_1378), .air_in(c_12_0));
valve v_12_2757 (.fluid_in(k_12_2757), .fluid_out(k_11_1378), .air_in(c_12_1));
valve v_12_2758 (.fluid_in(k_12_2758), .fluid_out(k_11_1379), .air_in(c_12_0));
valve v_12_2759 (.fluid_in(k_12_2759), .fluid_out(k_11_1379), .air_in(c_12_1));
valve v_12_2760 (.fluid_in(k_12_2760), .fluid_out(k_11_1380), .air_in(c_12_0));
valve v_12_2761 (.fluid_in(k_12_2761), .fluid_out(k_11_1380), .air_in(c_12_1));
valve v_12_2762 (.fluid_in(k_12_2762), .fluid_out(k_11_1381), .air_in(c_12_0));
valve v_12_2763 (.fluid_in(k_12_2763), .fluid_out(k_11_1381), .air_in(c_12_1));
valve v_12_2764 (.fluid_in(k_12_2764), .fluid_out(k_11_1382), .air_in(c_12_0));
valve v_12_2765 (.fluid_in(k_12_2765), .fluid_out(k_11_1382), .air_in(c_12_1));
valve v_12_2766 (.fluid_in(k_12_2766), .fluid_out(k_11_1383), .air_in(c_12_0));
valve v_12_2767 (.fluid_in(k_12_2767), .fluid_out(k_11_1383), .air_in(c_12_1));
valve v_12_2768 (.fluid_in(k_12_2768), .fluid_out(k_11_1384), .air_in(c_12_0));
valve v_12_2769 (.fluid_in(k_12_2769), .fluid_out(k_11_1384), .air_in(c_12_1));
valve v_12_2770 (.fluid_in(k_12_2770), .fluid_out(k_11_1385), .air_in(c_12_0));
valve v_12_2771 (.fluid_in(k_12_2771), .fluid_out(k_11_1385), .air_in(c_12_1));
valve v_12_2772 (.fluid_in(k_12_2772), .fluid_out(k_11_1386), .air_in(c_12_0));
valve v_12_2773 (.fluid_in(k_12_2773), .fluid_out(k_11_1386), .air_in(c_12_1));
valve v_12_2774 (.fluid_in(k_12_2774), .fluid_out(k_11_1387), .air_in(c_12_0));
valve v_12_2775 (.fluid_in(k_12_2775), .fluid_out(k_11_1387), .air_in(c_12_1));
valve v_12_2776 (.fluid_in(k_12_2776), .fluid_out(k_11_1388), .air_in(c_12_0));
valve v_12_2777 (.fluid_in(k_12_2777), .fluid_out(k_11_1388), .air_in(c_12_1));
valve v_12_2778 (.fluid_in(k_12_2778), .fluid_out(k_11_1389), .air_in(c_12_0));
valve v_12_2779 (.fluid_in(k_12_2779), .fluid_out(k_11_1389), .air_in(c_12_1));
valve v_12_2780 (.fluid_in(k_12_2780), .fluid_out(k_11_1390), .air_in(c_12_0));
valve v_12_2781 (.fluid_in(k_12_2781), .fluid_out(k_11_1390), .air_in(c_12_1));
valve v_12_2782 (.fluid_in(k_12_2782), .fluid_out(k_11_1391), .air_in(c_12_0));
valve v_12_2783 (.fluid_in(k_12_2783), .fluid_out(k_11_1391), .air_in(c_12_1));
valve v_12_2784 (.fluid_in(k_12_2784), .fluid_out(k_11_1392), .air_in(c_12_0));
valve v_12_2785 (.fluid_in(k_12_2785), .fluid_out(k_11_1392), .air_in(c_12_1));
valve v_12_2786 (.fluid_in(k_12_2786), .fluid_out(k_11_1393), .air_in(c_12_0));
valve v_12_2787 (.fluid_in(k_12_2787), .fluid_out(k_11_1393), .air_in(c_12_1));
valve v_12_2788 (.fluid_in(k_12_2788), .fluid_out(k_11_1394), .air_in(c_12_0));
valve v_12_2789 (.fluid_in(k_12_2789), .fluid_out(k_11_1394), .air_in(c_12_1));
valve v_12_2790 (.fluid_in(k_12_2790), .fluid_out(k_11_1395), .air_in(c_12_0));
valve v_12_2791 (.fluid_in(k_12_2791), .fluid_out(k_11_1395), .air_in(c_12_1));
valve v_12_2792 (.fluid_in(k_12_2792), .fluid_out(k_11_1396), .air_in(c_12_0));
valve v_12_2793 (.fluid_in(k_12_2793), .fluid_out(k_11_1396), .air_in(c_12_1));
valve v_12_2794 (.fluid_in(k_12_2794), .fluid_out(k_11_1397), .air_in(c_12_0));
valve v_12_2795 (.fluid_in(k_12_2795), .fluid_out(k_11_1397), .air_in(c_12_1));
valve v_12_2796 (.fluid_in(k_12_2796), .fluid_out(k_11_1398), .air_in(c_12_0));
valve v_12_2797 (.fluid_in(k_12_2797), .fluid_out(k_11_1398), .air_in(c_12_1));
valve v_12_2798 (.fluid_in(k_12_2798), .fluid_out(k_11_1399), .air_in(c_12_0));
valve v_12_2799 (.fluid_in(k_12_2799), .fluid_out(k_11_1399), .air_in(c_12_1));
valve v_12_2800 (.fluid_in(k_12_2800), .fluid_out(k_11_1400), .air_in(c_12_0));
valve v_12_2801 (.fluid_in(k_12_2801), .fluid_out(k_11_1400), .air_in(c_12_1));
valve v_12_2802 (.fluid_in(k_12_2802), .fluid_out(k_11_1401), .air_in(c_12_0));
valve v_12_2803 (.fluid_in(k_12_2803), .fluid_out(k_11_1401), .air_in(c_12_1));
valve v_12_2804 (.fluid_in(k_12_2804), .fluid_out(k_11_1402), .air_in(c_12_0));
valve v_12_2805 (.fluid_in(k_12_2805), .fluid_out(k_11_1402), .air_in(c_12_1));
valve v_12_2806 (.fluid_in(k_12_2806), .fluid_out(k_11_1403), .air_in(c_12_0));
valve v_12_2807 (.fluid_in(k_12_2807), .fluid_out(k_11_1403), .air_in(c_12_1));
valve v_12_2808 (.fluid_in(k_12_2808), .fluid_out(k_11_1404), .air_in(c_12_0));
valve v_12_2809 (.fluid_in(k_12_2809), .fluid_out(k_11_1404), .air_in(c_12_1));
valve v_12_2810 (.fluid_in(k_12_2810), .fluid_out(k_11_1405), .air_in(c_12_0));
valve v_12_2811 (.fluid_in(k_12_2811), .fluid_out(k_11_1405), .air_in(c_12_1));
valve v_12_2812 (.fluid_in(k_12_2812), .fluid_out(k_11_1406), .air_in(c_12_0));
valve v_12_2813 (.fluid_in(k_12_2813), .fluid_out(k_11_1406), .air_in(c_12_1));
valve v_12_2814 (.fluid_in(k_12_2814), .fluid_out(k_11_1407), .air_in(c_12_0));
valve v_12_2815 (.fluid_in(k_12_2815), .fluid_out(k_11_1407), .air_in(c_12_1));
valve v_12_2816 (.fluid_in(k_12_2816), .fluid_out(k_11_1408), .air_in(c_12_0));
valve v_12_2817 (.fluid_in(k_12_2817), .fluid_out(k_11_1408), .air_in(c_12_1));
valve v_12_2818 (.fluid_in(k_12_2818), .fluid_out(k_11_1409), .air_in(c_12_0));
valve v_12_2819 (.fluid_in(k_12_2819), .fluid_out(k_11_1409), .air_in(c_12_1));
valve v_12_2820 (.fluid_in(k_12_2820), .fluid_out(k_11_1410), .air_in(c_12_0));
valve v_12_2821 (.fluid_in(k_12_2821), .fluid_out(k_11_1410), .air_in(c_12_1));
valve v_12_2822 (.fluid_in(k_12_2822), .fluid_out(k_11_1411), .air_in(c_12_0));
valve v_12_2823 (.fluid_in(k_12_2823), .fluid_out(k_11_1411), .air_in(c_12_1));
valve v_12_2824 (.fluid_in(k_12_2824), .fluid_out(k_11_1412), .air_in(c_12_0));
valve v_12_2825 (.fluid_in(k_12_2825), .fluid_out(k_11_1412), .air_in(c_12_1));
valve v_12_2826 (.fluid_in(k_12_2826), .fluid_out(k_11_1413), .air_in(c_12_0));
valve v_12_2827 (.fluid_in(k_12_2827), .fluid_out(k_11_1413), .air_in(c_12_1));
valve v_12_2828 (.fluid_in(k_12_2828), .fluid_out(k_11_1414), .air_in(c_12_0));
valve v_12_2829 (.fluid_in(k_12_2829), .fluid_out(k_11_1414), .air_in(c_12_1));
valve v_12_2830 (.fluid_in(k_12_2830), .fluid_out(k_11_1415), .air_in(c_12_0));
valve v_12_2831 (.fluid_in(k_12_2831), .fluid_out(k_11_1415), .air_in(c_12_1));
valve v_12_2832 (.fluid_in(k_12_2832), .fluid_out(k_11_1416), .air_in(c_12_0));
valve v_12_2833 (.fluid_in(k_12_2833), .fluid_out(k_11_1416), .air_in(c_12_1));
valve v_12_2834 (.fluid_in(k_12_2834), .fluid_out(k_11_1417), .air_in(c_12_0));
valve v_12_2835 (.fluid_in(k_12_2835), .fluid_out(k_11_1417), .air_in(c_12_1));
valve v_12_2836 (.fluid_in(k_12_2836), .fluid_out(k_11_1418), .air_in(c_12_0));
valve v_12_2837 (.fluid_in(k_12_2837), .fluid_out(k_11_1418), .air_in(c_12_1));
valve v_12_2838 (.fluid_in(k_12_2838), .fluid_out(k_11_1419), .air_in(c_12_0));
valve v_12_2839 (.fluid_in(k_12_2839), .fluid_out(k_11_1419), .air_in(c_12_1));
valve v_12_2840 (.fluid_in(k_12_2840), .fluid_out(k_11_1420), .air_in(c_12_0));
valve v_12_2841 (.fluid_in(k_12_2841), .fluid_out(k_11_1420), .air_in(c_12_1));
valve v_12_2842 (.fluid_in(k_12_2842), .fluid_out(k_11_1421), .air_in(c_12_0));
valve v_12_2843 (.fluid_in(k_12_2843), .fluid_out(k_11_1421), .air_in(c_12_1));
valve v_12_2844 (.fluid_in(k_12_2844), .fluid_out(k_11_1422), .air_in(c_12_0));
valve v_12_2845 (.fluid_in(k_12_2845), .fluid_out(k_11_1422), .air_in(c_12_1));
valve v_12_2846 (.fluid_in(k_12_2846), .fluid_out(k_11_1423), .air_in(c_12_0));
valve v_12_2847 (.fluid_in(k_12_2847), .fluid_out(k_11_1423), .air_in(c_12_1));
valve v_12_2848 (.fluid_in(k_12_2848), .fluid_out(k_11_1424), .air_in(c_12_0));
valve v_12_2849 (.fluid_in(k_12_2849), .fluid_out(k_11_1424), .air_in(c_12_1));
valve v_12_2850 (.fluid_in(k_12_2850), .fluid_out(k_11_1425), .air_in(c_12_0));
valve v_12_2851 (.fluid_in(k_12_2851), .fluid_out(k_11_1425), .air_in(c_12_1));
valve v_12_2852 (.fluid_in(k_12_2852), .fluid_out(k_11_1426), .air_in(c_12_0));
valve v_12_2853 (.fluid_in(k_12_2853), .fluid_out(k_11_1426), .air_in(c_12_1));
valve v_12_2854 (.fluid_in(k_12_2854), .fluid_out(k_11_1427), .air_in(c_12_0));
valve v_12_2855 (.fluid_in(k_12_2855), .fluid_out(k_11_1427), .air_in(c_12_1));
valve v_12_2856 (.fluid_in(k_12_2856), .fluid_out(k_11_1428), .air_in(c_12_0));
valve v_12_2857 (.fluid_in(k_12_2857), .fluid_out(k_11_1428), .air_in(c_12_1));
valve v_12_2858 (.fluid_in(k_12_2858), .fluid_out(k_11_1429), .air_in(c_12_0));
valve v_12_2859 (.fluid_in(k_12_2859), .fluid_out(k_11_1429), .air_in(c_12_1));
valve v_12_2860 (.fluid_in(k_12_2860), .fluid_out(k_11_1430), .air_in(c_12_0));
valve v_12_2861 (.fluid_in(k_12_2861), .fluid_out(k_11_1430), .air_in(c_12_1));
valve v_12_2862 (.fluid_in(k_12_2862), .fluid_out(k_11_1431), .air_in(c_12_0));
valve v_12_2863 (.fluid_in(k_12_2863), .fluid_out(k_11_1431), .air_in(c_12_1));
valve v_12_2864 (.fluid_in(k_12_2864), .fluid_out(k_11_1432), .air_in(c_12_0));
valve v_12_2865 (.fluid_in(k_12_2865), .fluid_out(k_11_1432), .air_in(c_12_1));
valve v_12_2866 (.fluid_in(k_12_2866), .fluid_out(k_11_1433), .air_in(c_12_0));
valve v_12_2867 (.fluid_in(k_12_2867), .fluid_out(k_11_1433), .air_in(c_12_1));
valve v_12_2868 (.fluid_in(k_12_2868), .fluid_out(k_11_1434), .air_in(c_12_0));
valve v_12_2869 (.fluid_in(k_12_2869), .fluid_out(k_11_1434), .air_in(c_12_1));
valve v_12_2870 (.fluid_in(k_12_2870), .fluid_out(k_11_1435), .air_in(c_12_0));
valve v_12_2871 (.fluid_in(k_12_2871), .fluid_out(k_11_1435), .air_in(c_12_1));
valve v_12_2872 (.fluid_in(k_12_2872), .fluid_out(k_11_1436), .air_in(c_12_0));
valve v_12_2873 (.fluid_in(k_12_2873), .fluid_out(k_11_1436), .air_in(c_12_1));
valve v_12_2874 (.fluid_in(k_12_2874), .fluid_out(k_11_1437), .air_in(c_12_0));
valve v_12_2875 (.fluid_in(k_12_2875), .fluid_out(k_11_1437), .air_in(c_12_1));
valve v_12_2876 (.fluid_in(k_12_2876), .fluid_out(k_11_1438), .air_in(c_12_0));
valve v_12_2877 (.fluid_in(k_12_2877), .fluid_out(k_11_1438), .air_in(c_12_1));
valve v_12_2878 (.fluid_in(k_12_2878), .fluid_out(k_11_1439), .air_in(c_12_0));
valve v_12_2879 (.fluid_in(k_12_2879), .fluid_out(k_11_1439), .air_in(c_12_1));
valve v_12_2880 (.fluid_in(k_12_2880), .fluid_out(k_11_1440), .air_in(c_12_0));
valve v_12_2881 (.fluid_in(k_12_2881), .fluid_out(k_11_1440), .air_in(c_12_1));
valve v_12_2882 (.fluid_in(k_12_2882), .fluid_out(k_11_1441), .air_in(c_12_0));
valve v_12_2883 (.fluid_in(k_12_2883), .fluid_out(k_11_1441), .air_in(c_12_1));
valve v_12_2884 (.fluid_in(k_12_2884), .fluid_out(k_11_1442), .air_in(c_12_0));
valve v_12_2885 (.fluid_in(k_12_2885), .fluid_out(k_11_1442), .air_in(c_12_1));
valve v_12_2886 (.fluid_in(k_12_2886), .fluid_out(k_11_1443), .air_in(c_12_0));
valve v_12_2887 (.fluid_in(k_12_2887), .fluid_out(k_11_1443), .air_in(c_12_1));
valve v_12_2888 (.fluid_in(k_12_2888), .fluid_out(k_11_1444), .air_in(c_12_0));
valve v_12_2889 (.fluid_in(k_12_2889), .fluid_out(k_11_1444), .air_in(c_12_1));
valve v_12_2890 (.fluid_in(k_12_2890), .fluid_out(k_11_1445), .air_in(c_12_0));
valve v_12_2891 (.fluid_in(k_12_2891), .fluid_out(k_11_1445), .air_in(c_12_1));
valve v_12_2892 (.fluid_in(k_12_2892), .fluid_out(k_11_1446), .air_in(c_12_0));
valve v_12_2893 (.fluid_in(k_12_2893), .fluid_out(k_11_1446), .air_in(c_12_1));
valve v_12_2894 (.fluid_in(k_12_2894), .fluid_out(k_11_1447), .air_in(c_12_0));
valve v_12_2895 (.fluid_in(k_12_2895), .fluid_out(k_11_1447), .air_in(c_12_1));
valve v_12_2896 (.fluid_in(k_12_2896), .fluid_out(k_11_1448), .air_in(c_12_0));
valve v_12_2897 (.fluid_in(k_12_2897), .fluid_out(k_11_1448), .air_in(c_12_1));
valve v_12_2898 (.fluid_in(k_12_2898), .fluid_out(k_11_1449), .air_in(c_12_0));
valve v_12_2899 (.fluid_in(k_12_2899), .fluid_out(k_11_1449), .air_in(c_12_1));
valve v_12_2900 (.fluid_in(k_12_2900), .fluid_out(k_11_1450), .air_in(c_12_0));
valve v_12_2901 (.fluid_in(k_12_2901), .fluid_out(k_11_1450), .air_in(c_12_1));
valve v_12_2902 (.fluid_in(k_12_2902), .fluid_out(k_11_1451), .air_in(c_12_0));
valve v_12_2903 (.fluid_in(k_12_2903), .fluid_out(k_11_1451), .air_in(c_12_1));
valve v_12_2904 (.fluid_in(k_12_2904), .fluid_out(k_11_1452), .air_in(c_12_0));
valve v_12_2905 (.fluid_in(k_12_2905), .fluid_out(k_11_1452), .air_in(c_12_1));
valve v_12_2906 (.fluid_in(k_12_2906), .fluid_out(k_11_1453), .air_in(c_12_0));
valve v_12_2907 (.fluid_in(k_12_2907), .fluid_out(k_11_1453), .air_in(c_12_1));
valve v_12_2908 (.fluid_in(k_12_2908), .fluid_out(k_11_1454), .air_in(c_12_0));
valve v_12_2909 (.fluid_in(k_12_2909), .fluid_out(k_11_1454), .air_in(c_12_1));
valve v_12_2910 (.fluid_in(k_12_2910), .fluid_out(k_11_1455), .air_in(c_12_0));
valve v_12_2911 (.fluid_in(k_12_2911), .fluid_out(k_11_1455), .air_in(c_12_1));
valve v_12_2912 (.fluid_in(k_12_2912), .fluid_out(k_11_1456), .air_in(c_12_0));
valve v_12_2913 (.fluid_in(k_12_2913), .fluid_out(k_11_1456), .air_in(c_12_1));
valve v_12_2914 (.fluid_in(k_12_2914), .fluid_out(k_11_1457), .air_in(c_12_0));
valve v_12_2915 (.fluid_in(k_12_2915), .fluid_out(k_11_1457), .air_in(c_12_1));
valve v_12_2916 (.fluid_in(k_12_2916), .fluid_out(k_11_1458), .air_in(c_12_0));
valve v_12_2917 (.fluid_in(k_12_2917), .fluid_out(k_11_1458), .air_in(c_12_1));
valve v_12_2918 (.fluid_in(k_12_2918), .fluid_out(k_11_1459), .air_in(c_12_0));
valve v_12_2919 (.fluid_in(k_12_2919), .fluid_out(k_11_1459), .air_in(c_12_1));
valve v_12_2920 (.fluid_in(k_12_2920), .fluid_out(k_11_1460), .air_in(c_12_0));
valve v_12_2921 (.fluid_in(k_12_2921), .fluid_out(k_11_1460), .air_in(c_12_1));
valve v_12_2922 (.fluid_in(k_12_2922), .fluid_out(k_11_1461), .air_in(c_12_0));
valve v_12_2923 (.fluid_in(k_12_2923), .fluid_out(k_11_1461), .air_in(c_12_1));
valve v_12_2924 (.fluid_in(k_12_2924), .fluid_out(k_11_1462), .air_in(c_12_0));
valve v_12_2925 (.fluid_in(k_12_2925), .fluid_out(k_11_1462), .air_in(c_12_1));
valve v_12_2926 (.fluid_in(k_12_2926), .fluid_out(k_11_1463), .air_in(c_12_0));
valve v_12_2927 (.fluid_in(k_12_2927), .fluid_out(k_11_1463), .air_in(c_12_1));
valve v_12_2928 (.fluid_in(k_12_2928), .fluid_out(k_11_1464), .air_in(c_12_0));
valve v_12_2929 (.fluid_in(k_12_2929), .fluid_out(k_11_1464), .air_in(c_12_1));
valve v_12_2930 (.fluid_in(k_12_2930), .fluid_out(k_11_1465), .air_in(c_12_0));
valve v_12_2931 (.fluid_in(k_12_2931), .fluid_out(k_11_1465), .air_in(c_12_1));
valve v_12_2932 (.fluid_in(k_12_2932), .fluid_out(k_11_1466), .air_in(c_12_0));
valve v_12_2933 (.fluid_in(k_12_2933), .fluid_out(k_11_1466), .air_in(c_12_1));
valve v_12_2934 (.fluid_in(k_12_2934), .fluid_out(k_11_1467), .air_in(c_12_0));
valve v_12_2935 (.fluid_in(k_12_2935), .fluid_out(k_11_1467), .air_in(c_12_1));
valve v_12_2936 (.fluid_in(k_12_2936), .fluid_out(k_11_1468), .air_in(c_12_0));
valve v_12_2937 (.fluid_in(k_12_2937), .fluid_out(k_11_1468), .air_in(c_12_1));
valve v_12_2938 (.fluid_in(k_12_2938), .fluid_out(k_11_1469), .air_in(c_12_0));
valve v_12_2939 (.fluid_in(k_12_2939), .fluid_out(k_11_1469), .air_in(c_12_1));
valve v_12_2940 (.fluid_in(k_12_2940), .fluid_out(k_11_1470), .air_in(c_12_0));
valve v_12_2941 (.fluid_in(k_12_2941), .fluid_out(k_11_1470), .air_in(c_12_1));
valve v_12_2942 (.fluid_in(k_12_2942), .fluid_out(k_11_1471), .air_in(c_12_0));
valve v_12_2943 (.fluid_in(k_12_2943), .fluid_out(k_11_1471), .air_in(c_12_1));
valve v_12_2944 (.fluid_in(k_12_2944), .fluid_out(k_11_1472), .air_in(c_12_0));
valve v_12_2945 (.fluid_in(k_12_2945), .fluid_out(k_11_1472), .air_in(c_12_1));
valve v_12_2946 (.fluid_in(k_12_2946), .fluid_out(k_11_1473), .air_in(c_12_0));
valve v_12_2947 (.fluid_in(k_12_2947), .fluid_out(k_11_1473), .air_in(c_12_1));
valve v_12_2948 (.fluid_in(k_12_2948), .fluid_out(k_11_1474), .air_in(c_12_0));
valve v_12_2949 (.fluid_in(k_12_2949), .fluid_out(k_11_1474), .air_in(c_12_1));
valve v_12_2950 (.fluid_in(k_12_2950), .fluid_out(k_11_1475), .air_in(c_12_0));
valve v_12_2951 (.fluid_in(k_12_2951), .fluid_out(k_11_1475), .air_in(c_12_1));
valve v_12_2952 (.fluid_in(k_12_2952), .fluid_out(k_11_1476), .air_in(c_12_0));
valve v_12_2953 (.fluid_in(k_12_2953), .fluid_out(k_11_1476), .air_in(c_12_1));
valve v_12_2954 (.fluid_in(k_12_2954), .fluid_out(k_11_1477), .air_in(c_12_0));
valve v_12_2955 (.fluid_in(k_12_2955), .fluid_out(k_11_1477), .air_in(c_12_1));
valve v_12_2956 (.fluid_in(k_12_2956), .fluid_out(k_11_1478), .air_in(c_12_0));
valve v_12_2957 (.fluid_in(k_12_2957), .fluid_out(k_11_1478), .air_in(c_12_1));
valve v_12_2958 (.fluid_in(k_12_2958), .fluid_out(k_11_1479), .air_in(c_12_0));
valve v_12_2959 (.fluid_in(k_12_2959), .fluid_out(k_11_1479), .air_in(c_12_1));
valve v_12_2960 (.fluid_in(k_12_2960), .fluid_out(k_11_1480), .air_in(c_12_0));
valve v_12_2961 (.fluid_in(k_12_2961), .fluid_out(k_11_1480), .air_in(c_12_1));
valve v_12_2962 (.fluid_in(k_12_2962), .fluid_out(k_11_1481), .air_in(c_12_0));
valve v_12_2963 (.fluid_in(k_12_2963), .fluid_out(k_11_1481), .air_in(c_12_1));
valve v_12_2964 (.fluid_in(k_12_2964), .fluid_out(k_11_1482), .air_in(c_12_0));
valve v_12_2965 (.fluid_in(k_12_2965), .fluid_out(k_11_1482), .air_in(c_12_1));
valve v_12_2966 (.fluid_in(k_12_2966), .fluid_out(k_11_1483), .air_in(c_12_0));
valve v_12_2967 (.fluid_in(k_12_2967), .fluid_out(k_11_1483), .air_in(c_12_1));
valve v_12_2968 (.fluid_in(k_12_2968), .fluid_out(k_11_1484), .air_in(c_12_0));
valve v_12_2969 (.fluid_in(k_12_2969), .fluid_out(k_11_1484), .air_in(c_12_1));
valve v_12_2970 (.fluid_in(k_12_2970), .fluid_out(k_11_1485), .air_in(c_12_0));
valve v_12_2971 (.fluid_in(k_12_2971), .fluid_out(k_11_1485), .air_in(c_12_1));
valve v_12_2972 (.fluid_in(k_12_2972), .fluid_out(k_11_1486), .air_in(c_12_0));
valve v_12_2973 (.fluid_in(k_12_2973), .fluid_out(k_11_1486), .air_in(c_12_1));
valve v_12_2974 (.fluid_in(k_12_2974), .fluid_out(k_11_1487), .air_in(c_12_0));
valve v_12_2975 (.fluid_in(k_12_2975), .fluid_out(k_11_1487), .air_in(c_12_1));
valve v_12_2976 (.fluid_in(k_12_2976), .fluid_out(k_11_1488), .air_in(c_12_0));
valve v_12_2977 (.fluid_in(k_12_2977), .fluid_out(k_11_1488), .air_in(c_12_1));
valve v_12_2978 (.fluid_in(k_12_2978), .fluid_out(k_11_1489), .air_in(c_12_0));
valve v_12_2979 (.fluid_in(k_12_2979), .fluid_out(k_11_1489), .air_in(c_12_1));
valve v_12_2980 (.fluid_in(k_12_2980), .fluid_out(k_11_1490), .air_in(c_12_0));
valve v_12_2981 (.fluid_in(k_12_2981), .fluid_out(k_11_1490), .air_in(c_12_1));
valve v_12_2982 (.fluid_in(k_12_2982), .fluid_out(k_11_1491), .air_in(c_12_0));
valve v_12_2983 (.fluid_in(k_12_2983), .fluid_out(k_11_1491), .air_in(c_12_1));
valve v_12_2984 (.fluid_in(k_12_2984), .fluid_out(k_11_1492), .air_in(c_12_0));
valve v_12_2985 (.fluid_in(k_12_2985), .fluid_out(k_11_1492), .air_in(c_12_1));
valve v_12_2986 (.fluid_in(k_12_2986), .fluid_out(k_11_1493), .air_in(c_12_0));
valve v_12_2987 (.fluid_in(k_12_2987), .fluid_out(k_11_1493), .air_in(c_12_1));
valve v_12_2988 (.fluid_in(k_12_2988), .fluid_out(k_11_1494), .air_in(c_12_0));
valve v_12_2989 (.fluid_in(k_12_2989), .fluid_out(k_11_1494), .air_in(c_12_1));
valve v_12_2990 (.fluid_in(k_12_2990), .fluid_out(k_11_1495), .air_in(c_12_0));
valve v_12_2991 (.fluid_in(k_12_2991), .fluid_out(k_11_1495), .air_in(c_12_1));
valve v_12_2992 (.fluid_in(k_12_2992), .fluid_out(k_11_1496), .air_in(c_12_0));
valve v_12_2993 (.fluid_in(k_12_2993), .fluid_out(k_11_1496), .air_in(c_12_1));
valve v_12_2994 (.fluid_in(k_12_2994), .fluid_out(k_11_1497), .air_in(c_12_0));
valve v_12_2995 (.fluid_in(k_12_2995), .fluid_out(k_11_1497), .air_in(c_12_1));
valve v_12_2996 (.fluid_in(k_12_2996), .fluid_out(k_11_1498), .air_in(c_12_0));
valve v_12_2997 (.fluid_in(k_12_2997), .fluid_out(k_11_1498), .air_in(c_12_1));
valve v_12_2998 (.fluid_in(k_12_2998), .fluid_out(k_11_1499), .air_in(c_12_0));
valve v_12_2999 (.fluid_in(k_12_2999), .fluid_out(k_11_1499), .air_in(c_12_1));
valve v_12_3000 (.fluid_in(k_12_3000), .fluid_out(k_11_1500), .air_in(c_12_0));
valve v_12_3001 (.fluid_in(k_12_3001), .fluid_out(k_11_1500), .air_in(c_12_1));
valve v_12_3002 (.fluid_in(k_12_3002), .fluid_out(k_11_1501), .air_in(c_12_0));
valve v_12_3003 (.fluid_in(k_12_3003), .fluid_out(k_11_1501), .air_in(c_12_1));
valve v_12_3004 (.fluid_in(k_12_3004), .fluid_out(k_11_1502), .air_in(c_12_0));
valve v_12_3005 (.fluid_in(k_12_3005), .fluid_out(k_11_1502), .air_in(c_12_1));
valve v_12_3006 (.fluid_in(k_12_3006), .fluid_out(k_11_1503), .air_in(c_12_0));
valve v_12_3007 (.fluid_in(k_12_3007), .fluid_out(k_11_1503), .air_in(c_12_1));
valve v_12_3008 (.fluid_in(k_12_3008), .fluid_out(k_11_1504), .air_in(c_12_0));
valve v_12_3009 (.fluid_in(k_12_3009), .fluid_out(k_11_1504), .air_in(c_12_1));
valve v_12_3010 (.fluid_in(k_12_3010), .fluid_out(k_11_1505), .air_in(c_12_0));
valve v_12_3011 (.fluid_in(k_12_3011), .fluid_out(k_11_1505), .air_in(c_12_1));
valve v_12_3012 (.fluid_in(k_12_3012), .fluid_out(k_11_1506), .air_in(c_12_0));
valve v_12_3013 (.fluid_in(k_12_3013), .fluid_out(k_11_1506), .air_in(c_12_1));
valve v_12_3014 (.fluid_in(k_12_3014), .fluid_out(k_11_1507), .air_in(c_12_0));
valve v_12_3015 (.fluid_in(k_12_3015), .fluid_out(k_11_1507), .air_in(c_12_1));
valve v_12_3016 (.fluid_in(k_12_3016), .fluid_out(k_11_1508), .air_in(c_12_0));
valve v_12_3017 (.fluid_in(k_12_3017), .fluid_out(k_11_1508), .air_in(c_12_1));
valve v_12_3018 (.fluid_in(k_12_3018), .fluid_out(k_11_1509), .air_in(c_12_0));
valve v_12_3019 (.fluid_in(k_12_3019), .fluid_out(k_11_1509), .air_in(c_12_1));
valve v_12_3020 (.fluid_in(k_12_3020), .fluid_out(k_11_1510), .air_in(c_12_0));
valve v_12_3021 (.fluid_in(k_12_3021), .fluid_out(k_11_1510), .air_in(c_12_1));
valve v_12_3022 (.fluid_in(k_12_3022), .fluid_out(k_11_1511), .air_in(c_12_0));
valve v_12_3023 (.fluid_in(k_12_3023), .fluid_out(k_11_1511), .air_in(c_12_1));
valve v_12_3024 (.fluid_in(k_12_3024), .fluid_out(k_11_1512), .air_in(c_12_0));
valve v_12_3025 (.fluid_in(k_12_3025), .fluid_out(k_11_1512), .air_in(c_12_1));
valve v_12_3026 (.fluid_in(k_12_3026), .fluid_out(k_11_1513), .air_in(c_12_0));
valve v_12_3027 (.fluid_in(k_12_3027), .fluid_out(k_11_1513), .air_in(c_12_1));
valve v_12_3028 (.fluid_in(k_12_3028), .fluid_out(k_11_1514), .air_in(c_12_0));
valve v_12_3029 (.fluid_in(k_12_3029), .fluid_out(k_11_1514), .air_in(c_12_1));
valve v_12_3030 (.fluid_in(k_12_3030), .fluid_out(k_11_1515), .air_in(c_12_0));
valve v_12_3031 (.fluid_in(k_12_3031), .fluid_out(k_11_1515), .air_in(c_12_1));
valve v_12_3032 (.fluid_in(k_12_3032), .fluid_out(k_11_1516), .air_in(c_12_0));
valve v_12_3033 (.fluid_in(k_12_3033), .fluid_out(k_11_1516), .air_in(c_12_1));
valve v_12_3034 (.fluid_in(k_12_3034), .fluid_out(k_11_1517), .air_in(c_12_0));
valve v_12_3035 (.fluid_in(k_12_3035), .fluid_out(k_11_1517), .air_in(c_12_1));
valve v_12_3036 (.fluid_in(k_12_3036), .fluid_out(k_11_1518), .air_in(c_12_0));
valve v_12_3037 (.fluid_in(k_12_3037), .fluid_out(k_11_1518), .air_in(c_12_1));
valve v_12_3038 (.fluid_in(k_12_3038), .fluid_out(k_11_1519), .air_in(c_12_0));
valve v_12_3039 (.fluid_in(k_12_3039), .fluid_out(k_11_1519), .air_in(c_12_1));
valve v_12_3040 (.fluid_in(k_12_3040), .fluid_out(k_11_1520), .air_in(c_12_0));
valve v_12_3041 (.fluid_in(k_12_3041), .fluid_out(k_11_1520), .air_in(c_12_1));
valve v_12_3042 (.fluid_in(k_12_3042), .fluid_out(k_11_1521), .air_in(c_12_0));
valve v_12_3043 (.fluid_in(k_12_3043), .fluid_out(k_11_1521), .air_in(c_12_1));
valve v_12_3044 (.fluid_in(k_12_3044), .fluid_out(k_11_1522), .air_in(c_12_0));
valve v_12_3045 (.fluid_in(k_12_3045), .fluid_out(k_11_1522), .air_in(c_12_1));
valve v_12_3046 (.fluid_in(k_12_3046), .fluid_out(k_11_1523), .air_in(c_12_0));
valve v_12_3047 (.fluid_in(k_12_3047), .fluid_out(k_11_1523), .air_in(c_12_1));
valve v_12_3048 (.fluid_in(k_12_3048), .fluid_out(k_11_1524), .air_in(c_12_0));
valve v_12_3049 (.fluid_in(k_12_3049), .fluid_out(k_11_1524), .air_in(c_12_1));
valve v_12_3050 (.fluid_in(k_12_3050), .fluid_out(k_11_1525), .air_in(c_12_0));
valve v_12_3051 (.fluid_in(k_12_3051), .fluid_out(k_11_1525), .air_in(c_12_1));
valve v_12_3052 (.fluid_in(k_12_3052), .fluid_out(k_11_1526), .air_in(c_12_0));
valve v_12_3053 (.fluid_in(k_12_3053), .fluid_out(k_11_1526), .air_in(c_12_1));
valve v_12_3054 (.fluid_in(k_12_3054), .fluid_out(k_11_1527), .air_in(c_12_0));
valve v_12_3055 (.fluid_in(k_12_3055), .fluid_out(k_11_1527), .air_in(c_12_1));
valve v_12_3056 (.fluid_in(k_12_3056), .fluid_out(k_11_1528), .air_in(c_12_0));
valve v_12_3057 (.fluid_in(k_12_3057), .fluid_out(k_11_1528), .air_in(c_12_1));
valve v_12_3058 (.fluid_in(k_12_3058), .fluid_out(k_11_1529), .air_in(c_12_0));
valve v_12_3059 (.fluid_in(k_12_3059), .fluid_out(k_11_1529), .air_in(c_12_1));
valve v_12_3060 (.fluid_in(k_12_3060), .fluid_out(k_11_1530), .air_in(c_12_0));
valve v_12_3061 (.fluid_in(k_12_3061), .fluid_out(k_11_1530), .air_in(c_12_1));
valve v_12_3062 (.fluid_in(k_12_3062), .fluid_out(k_11_1531), .air_in(c_12_0));
valve v_12_3063 (.fluid_in(k_12_3063), .fluid_out(k_11_1531), .air_in(c_12_1));
valve v_12_3064 (.fluid_in(k_12_3064), .fluid_out(k_11_1532), .air_in(c_12_0));
valve v_12_3065 (.fluid_in(k_12_3065), .fluid_out(k_11_1532), .air_in(c_12_1));
valve v_12_3066 (.fluid_in(k_12_3066), .fluid_out(k_11_1533), .air_in(c_12_0));
valve v_12_3067 (.fluid_in(k_12_3067), .fluid_out(k_11_1533), .air_in(c_12_1));
valve v_12_3068 (.fluid_in(k_12_3068), .fluid_out(k_11_1534), .air_in(c_12_0));
valve v_12_3069 (.fluid_in(k_12_3069), .fluid_out(k_11_1534), .air_in(c_12_1));
valve v_12_3070 (.fluid_in(k_12_3070), .fluid_out(k_11_1535), .air_in(c_12_0));
valve v_12_3071 (.fluid_in(k_12_3071), .fluid_out(k_11_1535), .air_in(c_12_1));
valve v_12_3072 (.fluid_in(k_12_3072), .fluid_out(k_11_1536), .air_in(c_12_0));
valve v_12_3073 (.fluid_in(k_12_3073), .fluid_out(k_11_1536), .air_in(c_12_1));
valve v_12_3074 (.fluid_in(k_12_3074), .fluid_out(k_11_1537), .air_in(c_12_0));
valve v_12_3075 (.fluid_in(k_12_3075), .fluid_out(k_11_1537), .air_in(c_12_1));
valve v_12_3076 (.fluid_in(k_12_3076), .fluid_out(k_11_1538), .air_in(c_12_0));
valve v_12_3077 (.fluid_in(k_12_3077), .fluid_out(k_11_1538), .air_in(c_12_1));
valve v_12_3078 (.fluid_in(k_12_3078), .fluid_out(k_11_1539), .air_in(c_12_0));
valve v_12_3079 (.fluid_in(k_12_3079), .fluid_out(k_11_1539), .air_in(c_12_1));
valve v_12_3080 (.fluid_in(k_12_3080), .fluid_out(k_11_1540), .air_in(c_12_0));
valve v_12_3081 (.fluid_in(k_12_3081), .fluid_out(k_11_1540), .air_in(c_12_1));
valve v_12_3082 (.fluid_in(k_12_3082), .fluid_out(k_11_1541), .air_in(c_12_0));
valve v_12_3083 (.fluid_in(k_12_3083), .fluid_out(k_11_1541), .air_in(c_12_1));
valve v_12_3084 (.fluid_in(k_12_3084), .fluid_out(k_11_1542), .air_in(c_12_0));
valve v_12_3085 (.fluid_in(k_12_3085), .fluid_out(k_11_1542), .air_in(c_12_1));
valve v_12_3086 (.fluid_in(k_12_3086), .fluid_out(k_11_1543), .air_in(c_12_0));
valve v_12_3087 (.fluid_in(k_12_3087), .fluid_out(k_11_1543), .air_in(c_12_1));
valve v_12_3088 (.fluid_in(k_12_3088), .fluid_out(k_11_1544), .air_in(c_12_0));
valve v_12_3089 (.fluid_in(k_12_3089), .fluid_out(k_11_1544), .air_in(c_12_1));
valve v_12_3090 (.fluid_in(k_12_3090), .fluid_out(k_11_1545), .air_in(c_12_0));
valve v_12_3091 (.fluid_in(k_12_3091), .fluid_out(k_11_1545), .air_in(c_12_1));
valve v_12_3092 (.fluid_in(k_12_3092), .fluid_out(k_11_1546), .air_in(c_12_0));
valve v_12_3093 (.fluid_in(k_12_3093), .fluid_out(k_11_1546), .air_in(c_12_1));
valve v_12_3094 (.fluid_in(k_12_3094), .fluid_out(k_11_1547), .air_in(c_12_0));
valve v_12_3095 (.fluid_in(k_12_3095), .fluid_out(k_11_1547), .air_in(c_12_1));
valve v_12_3096 (.fluid_in(k_12_3096), .fluid_out(k_11_1548), .air_in(c_12_0));
valve v_12_3097 (.fluid_in(k_12_3097), .fluid_out(k_11_1548), .air_in(c_12_1));
valve v_12_3098 (.fluid_in(k_12_3098), .fluid_out(k_11_1549), .air_in(c_12_0));
valve v_12_3099 (.fluid_in(k_12_3099), .fluid_out(k_11_1549), .air_in(c_12_1));
valve v_12_3100 (.fluid_in(k_12_3100), .fluid_out(k_11_1550), .air_in(c_12_0));
valve v_12_3101 (.fluid_in(k_12_3101), .fluid_out(k_11_1550), .air_in(c_12_1));
valve v_12_3102 (.fluid_in(k_12_3102), .fluid_out(k_11_1551), .air_in(c_12_0));
valve v_12_3103 (.fluid_in(k_12_3103), .fluid_out(k_11_1551), .air_in(c_12_1));
valve v_12_3104 (.fluid_in(k_12_3104), .fluid_out(k_11_1552), .air_in(c_12_0));
valve v_12_3105 (.fluid_in(k_12_3105), .fluid_out(k_11_1552), .air_in(c_12_1));
valve v_12_3106 (.fluid_in(k_12_3106), .fluid_out(k_11_1553), .air_in(c_12_0));
valve v_12_3107 (.fluid_in(k_12_3107), .fluid_out(k_11_1553), .air_in(c_12_1));
valve v_12_3108 (.fluid_in(k_12_3108), .fluid_out(k_11_1554), .air_in(c_12_0));
valve v_12_3109 (.fluid_in(k_12_3109), .fluid_out(k_11_1554), .air_in(c_12_1));
valve v_12_3110 (.fluid_in(k_12_3110), .fluid_out(k_11_1555), .air_in(c_12_0));
valve v_12_3111 (.fluid_in(k_12_3111), .fluid_out(k_11_1555), .air_in(c_12_1));
valve v_12_3112 (.fluid_in(k_12_3112), .fluid_out(k_11_1556), .air_in(c_12_0));
valve v_12_3113 (.fluid_in(k_12_3113), .fluid_out(k_11_1556), .air_in(c_12_1));
valve v_12_3114 (.fluid_in(k_12_3114), .fluid_out(k_11_1557), .air_in(c_12_0));
valve v_12_3115 (.fluid_in(k_12_3115), .fluid_out(k_11_1557), .air_in(c_12_1));
valve v_12_3116 (.fluid_in(k_12_3116), .fluid_out(k_11_1558), .air_in(c_12_0));
valve v_12_3117 (.fluid_in(k_12_3117), .fluid_out(k_11_1558), .air_in(c_12_1));
valve v_12_3118 (.fluid_in(k_12_3118), .fluid_out(k_11_1559), .air_in(c_12_0));
valve v_12_3119 (.fluid_in(k_12_3119), .fluid_out(k_11_1559), .air_in(c_12_1));
valve v_12_3120 (.fluid_in(k_12_3120), .fluid_out(k_11_1560), .air_in(c_12_0));
valve v_12_3121 (.fluid_in(k_12_3121), .fluid_out(k_11_1560), .air_in(c_12_1));
valve v_12_3122 (.fluid_in(k_12_3122), .fluid_out(k_11_1561), .air_in(c_12_0));
valve v_12_3123 (.fluid_in(k_12_3123), .fluid_out(k_11_1561), .air_in(c_12_1));
valve v_12_3124 (.fluid_in(k_12_3124), .fluid_out(k_11_1562), .air_in(c_12_0));
valve v_12_3125 (.fluid_in(k_12_3125), .fluid_out(k_11_1562), .air_in(c_12_1));
valve v_12_3126 (.fluid_in(k_12_3126), .fluid_out(k_11_1563), .air_in(c_12_0));
valve v_12_3127 (.fluid_in(k_12_3127), .fluid_out(k_11_1563), .air_in(c_12_1));
valve v_12_3128 (.fluid_in(k_12_3128), .fluid_out(k_11_1564), .air_in(c_12_0));
valve v_12_3129 (.fluid_in(k_12_3129), .fluid_out(k_11_1564), .air_in(c_12_1));
valve v_12_3130 (.fluid_in(k_12_3130), .fluid_out(k_11_1565), .air_in(c_12_0));
valve v_12_3131 (.fluid_in(k_12_3131), .fluid_out(k_11_1565), .air_in(c_12_1));
valve v_12_3132 (.fluid_in(k_12_3132), .fluid_out(k_11_1566), .air_in(c_12_0));
valve v_12_3133 (.fluid_in(k_12_3133), .fluid_out(k_11_1566), .air_in(c_12_1));
valve v_12_3134 (.fluid_in(k_12_3134), .fluid_out(k_11_1567), .air_in(c_12_0));
valve v_12_3135 (.fluid_in(k_12_3135), .fluid_out(k_11_1567), .air_in(c_12_1));
valve v_12_3136 (.fluid_in(k_12_3136), .fluid_out(k_11_1568), .air_in(c_12_0));
valve v_12_3137 (.fluid_in(k_12_3137), .fluid_out(k_11_1568), .air_in(c_12_1));
valve v_12_3138 (.fluid_in(k_12_3138), .fluid_out(k_11_1569), .air_in(c_12_0));
valve v_12_3139 (.fluid_in(k_12_3139), .fluid_out(k_11_1569), .air_in(c_12_1));
valve v_12_3140 (.fluid_in(k_12_3140), .fluid_out(k_11_1570), .air_in(c_12_0));
valve v_12_3141 (.fluid_in(k_12_3141), .fluid_out(k_11_1570), .air_in(c_12_1));
valve v_12_3142 (.fluid_in(k_12_3142), .fluid_out(k_11_1571), .air_in(c_12_0));
valve v_12_3143 (.fluid_in(k_12_3143), .fluid_out(k_11_1571), .air_in(c_12_1));
valve v_12_3144 (.fluid_in(k_12_3144), .fluid_out(k_11_1572), .air_in(c_12_0));
valve v_12_3145 (.fluid_in(k_12_3145), .fluid_out(k_11_1572), .air_in(c_12_1));
valve v_12_3146 (.fluid_in(k_12_3146), .fluid_out(k_11_1573), .air_in(c_12_0));
valve v_12_3147 (.fluid_in(k_12_3147), .fluid_out(k_11_1573), .air_in(c_12_1));
valve v_12_3148 (.fluid_in(k_12_3148), .fluid_out(k_11_1574), .air_in(c_12_0));
valve v_12_3149 (.fluid_in(k_12_3149), .fluid_out(k_11_1574), .air_in(c_12_1));
valve v_12_3150 (.fluid_in(k_12_3150), .fluid_out(k_11_1575), .air_in(c_12_0));
valve v_12_3151 (.fluid_in(k_12_3151), .fluid_out(k_11_1575), .air_in(c_12_1));
valve v_12_3152 (.fluid_in(k_12_3152), .fluid_out(k_11_1576), .air_in(c_12_0));
valve v_12_3153 (.fluid_in(k_12_3153), .fluid_out(k_11_1576), .air_in(c_12_1));
valve v_12_3154 (.fluid_in(k_12_3154), .fluid_out(k_11_1577), .air_in(c_12_0));
valve v_12_3155 (.fluid_in(k_12_3155), .fluid_out(k_11_1577), .air_in(c_12_1));
valve v_12_3156 (.fluid_in(k_12_3156), .fluid_out(k_11_1578), .air_in(c_12_0));
valve v_12_3157 (.fluid_in(k_12_3157), .fluid_out(k_11_1578), .air_in(c_12_1));
valve v_12_3158 (.fluid_in(k_12_3158), .fluid_out(k_11_1579), .air_in(c_12_0));
valve v_12_3159 (.fluid_in(k_12_3159), .fluid_out(k_11_1579), .air_in(c_12_1));
valve v_12_3160 (.fluid_in(k_12_3160), .fluid_out(k_11_1580), .air_in(c_12_0));
valve v_12_3161 (.fluid_in(k_12_3161), .fluid_out(k_11_1580), .air_in(c_12_1));
valve v_12_3162 (.fluid_in(k_12_3162), .fluid_out(k_11_1581), .air_in(c_12_0));
valve v_12_3163 (.fluid_in(k_12_3163), .fluid_out(k_11_1581), .air_in(c_12_1));
valve v_12_3164 (.fluid_in(k_12_3164), .fluid_out(k_11_1582), .air_in(c_12_0));
valve v_12_3165 (.fluid_in(k_12_3165), .fluid_out(k_11_1582), .air_in(c_12_1));
valve v_12_3166 (.fluid_in(k_12_3166), .fluid_out(k_11_1583), .air_in(c_12_0));
valve v_12_3167 (.fluid_in(k_12_3167), .fluid_out(k_11_1583), .air_in(c_12_1));
valve v_12_3168 (.fluid_in(k_12_3168), .fluid_out(k_11_1584), .air_in(c_12_0));
valve v_12_3169 (.fluid_in(k_12_3169), .fluid_out(k_11_1584), .air_in(c_12_1));
valve v_12_3170 (.fluid_in(k_12_3170), .fluid_out(k_11_1585), .air_in(c_12_0));
valve v_12_3171 (.fluid_in(k_12_3171), .fluid_out(k_11_1585), .air_in(c_12_1));
valve v_12_3172 (.fluid_in(k_12_3172), .fluid_out(k_11_1586), .air_in(c_12_0));
valve v_12_3173 (.fluid_in(k_12_3173), .fluid_out(k_11_1586), .air_in(c_12_1));
valve v_12_3174 (.fluid_in(k_12_3174), .fluid_out(k_11_1587), .air_in(c_12_0));
valve v_12_3175 (.fluid_in(k_12_3175), .fluid_out(k_11_1587), .air_in(c_12_1));
valve v_12_3176 (.fluid_in(k_12_3176), .fluid_out(k_11_1588), .air_in(c_12_0));
valve v_12_3177 (.fluid_in(k_12_3177), .fluid_out(k_11_1588), .air_in(c_12_1));
valve v_12_3178 (.fluid_in(k_12_3178), .fluid_out(k_11_1589), .air_in(c_12_0));
valve v_12_3179 (.fluid_in(k_12_3179), .fluid_out(k_11_1589), .air_in(c_12_1));
valve v_12_3180 (.fluid_in(k_12_3180), .fluid_out(k_11_1590), .air_in(c_12_0));
valve v_12_3181 (.fluid_in(k_12_3181), .fluid_out(k_11_1590), .air_in(c_12_1));
valve v_12_3182 (.fluid_in(k_12_3182), .fluid_out(k_11_1591), .air_in(c_12_0));
valve v_12_3183 (.fluid_in(k_12_3183), .fluid_out(k_11_1591), .air_in(c_12_1));
valve v_12_3184 (.fluid_in(k_12_3184), .fluid_out(k_11_1592), .air_in(c_12_0));
valve v_12_3185 (.fluid_in(k_12_3185), .fluid_out(k_11_1592), .air_in(c_12_1));
valve v_12_3186 (.fluid_in(k_12_3186), .fluid_out(k_11_1593), .air_in(c_12_0));
valve v_12_3187 (.fluid_in(k_12_3187), .fluid_out(k_11_1593), .air_in(c_12_1));
valve v_12_3188 (.fluid_in(k_12_3188), .fluid_out(k_11_1594), .air_in(c_12_0));
valve v_12_3189 (.fluid_in(k_12_3189), .fluid_out(k_11_1594), .air_in(c_12_1));
valve v_12_3190 (.fluid_in(k_12_3190), .fluid_out(k_11_1595), .air_in(c_12_0));
valve v_12_3191 (.fluid_in(k_12_3191), .fluid_out(k_11_1595), .air_in(c_12_1));
valve v_12_3192 (.fluid_in(k_12_3192), .fluid_out(k_11_1596), .air_in(c_12_0));
valve v_12_3193 (.fluid_in(k_12_3193), .fluid_out(k_11_1596), .air_in(c_12_1));
valve v_12_3194 (.fluid_in(k_12_3194), .fluid_out(k_11_1597), .air_in(c_12_0));
valve v_12_3195 (.fluid_in(k_12_3195), .fluid_out(k_11_1597), .air_in(c_12_1));
valve v_12_3196 (.fluid_in(k_12_3196), .fluid_out(k_11_1598), .air_in(c_12_0));
valve v_12_3197 (.fluid_in(k_12_3197), .fluid_out(k_11_1598), .air_in(c_12_1));
valve v_12_3198 (.fluid_in(k_12_3198), .fluid_out(k_11_1599), .air_in(c_12_0));
valve v_12_3199 (.fluid_in(k_12_3199), .fluid_out(k_11_1599), .air_in(c_12_1));
valve v_12_3200 (.fluid_in(k_12_3200), .fluid_out(k_11_1600), .air_in(c_12_0));
valve v_12_3201 (.fluid_in(k_12_3201), .fluid_out(k_11_1600), .air_in(c_12_1));
valve v_12_3202 (.fluid_in(k_12_3202), .fluid_out(k_11_1601), .air_in(c_12_0));
valve v_12_3203 (.fluid_in(k_12_3203), .fluid_out(k_11_1601), .air_in(c_12_1));
valve v_12_3204 (.fluid_in(k_12_3204), .fluid_out(k_11_1602), .air_in(c_12_0));
valve v_12_3205 (.fluid_in(k_12_3205), .fluid_out(k_11_1602), .air_in(c_12_1));
valve v_12_3206 (.fluid_in(k_12_3206), .fluid_out(k_11_1603), .air_in(c_12_0));
valve v_12_3207 (.fluid_in(k_12_3207), .fluid_out(k_11_1603), .air_in(c_12_1));
valve v_12_3208 (.fluid_in(k_12_3208), .fluid_out(k_11_1604), .air_in(c_12_0));
valve v_12_3209 (.fluid_in(k_12_3209), .fluid_out(k_11_1604), .air_in(c_12_1));
valve v_12_3210 (.fluid_in(k_12_3210), .fluid_out(k_11_1605), .air_in(c_12_0));
valve v_12_3211 (.fluid_in(k_12_3211), .fluid_out(k_11_1605), .air_in(c_12_1));
valve v_12_3212 (.fluid_in(k_12_3212), .fluid_out(k_11_1606), .air_in(c_12_0));
valve v_12_3213 (.fluid_in(k_12_3213), .fluid_out(k_11_1606), .air_in(c_12_1));
valve v_12_3214 (.fluid_in(k_12_3214), .fluid_out(k_11_1607), .air_in(c_12_0));
valve v_12_3215 (.fluid_in(k_12_3215), .fluid_out(k_11_1607), .air_in(c_12_1));
valve v_12_3216 (.fluid_in(k_12_3216), .fluid_out(k_11_1608), .air_in(c_12_0));
valve v_12_3217 (.fluid_in(k_12_3217), .fluid_out(k_11_1608), .air_in(c_12_1));
valve v_12_3218 (.fluid_in(k_12_3218), .fluid_out(k_11_1609), .air_in(c_12_0));
valve v_12_3219 (.fluid_in(k_12_3219), .fluid_out(k_11_1609), .air_in(c_12_1));
valve v_12_3220 (.fluid_in(k_12_3220), .fluid_out(k_11_1610), .air_in(c_12_0));
valve v_12_3221 (.fluid_in(k_12_3221), .fluid_out(k_11_1610), .air_in(c_12_1));
valve v_12_3222 (.fluid_in(k_12_3222), .fluid_out(k_11_1611), .air_in(c_12_0));
valve v_12_3223 (.fluid_in(k_12_3223), .fluid_out(k_11_1611), .air_in(c_12_1));
valve v_12_3224 (.fluid_in(k_12_3224), .fluid_out(k_11_1612), .air_in(c_12_0));
valve v_12_3225 (.fluid_in(k_12_3225), .fluid_out(k_11_1612), .air_in(c_12_1));
valve v_12_3226 (.fluid_in(k_12_3226), .fluid_out(k_11_1613), .air_in(c_12_0));
valve v_12_3227 (.fluid_in(k_12_3227), .fluid_out(k_11_1613), .air_in(c_12_1));
valve v_12_3228 (.fluid_in(k_12_3228), .fluid_out(k_11_1614), .air_in(c_12_0));
valve v_12_3229 (.fluid_in(k_12_3229), .fluid_out(k_11_1614), .air_in(c_12_1));
valve v_12_3230 (.fluid_in(k_12_3230), .fluid_out(k_11_1615), .air_in(c_12_0));
valve v_12_3231 (.fluid_in(k_12_3231), .fluid_out(k_11_1615), .air_in(c_12_1));
valve v_12_3232 (.fluid_in(k_12_3232), .fluid_out(k_11_1616), .air_in(c_12_0));
valve v_12_3233 (.fluid_in(k_12_3233), .fluid_out(k_11_1616), .air_in(c_12_1));
valve v_12_3234 (.fluid_in(k_12_3234), .fluid_out(k_11_1617), .air_in(c_12_0));
valve v_12_3235 (.fluid_in(k_12_3235), .fluid_out(k_11_1617), .air_in(c_12_1));
valve v_12_3236 (.fluid_in(k_12_3236), .fluid_out(k_11_1618), .air_in(c_12_0));
valve v_12_3237 (.fluid_in(k_12_3237), .fluid_out(k_11_1618), .air_in(c_12_1));
valve v_12_3238 (.fluid_in(k_12_3238), .fluid_out(k_11_1619), .air_in(c_12_0));
valve v_12_3239 (.fluid_in(k_12_3239), .fluid_out(k_11_1619), .air_in(c_12_1));
valve v_12_3240 (.fluid_in(k_12_3240), .fluid_out(k_11_1620), .air_in(c_12_0));
valve v_12_3241 (.fluid_in(k_12_3241), .fluid_out(k_11_1620), .air_in(c_12_1));
valve v_12_3242 (.fluid_in(k_12_3242), .fluid_out(k_11_1621), .air_in(c_12_0));
valve v_12_3243 (.fluid_in(k_12_3243), .fluid_out(k_11_1621), .air_in(c_12_1));
valve v_12_3244 (.fluid_in(k_12_3244), .fluid_out(k_11_1622), .air_in(c_12_0));
valve v_12_3245 (.fluid_in(k_12_3245), .fluid_out(k_11_1622), .air_in(c_12_1));
valve v_12_3246 (.fluid_in(k_12_3246), .fluid_out(k_11_1623), .air_in(c_12_0));
valve v_12_3247 (.fluid_in(k_12_3247), .fluid_out(k_11_1623), .air_in(c_12_1));
valve v_12_3248 (.fluid_in(k_12_3248), .fluid_out(k_11_1624), .air_in(c_12_0));
valve v_12_3249 (.fluid_in(k_12_3249), .fluid_out(k_11_1624), .air_in(c_12_1));
valve v_12_3250 (.fluid_in(k_12_3250), .fluid_out(k_11_1625), .air_in(c_12_0));
valve v_12_3251 (.fluid_in(k_12_3251), .fluid_out(k_11_1625), .air_in(c_12_1));
valve v_12_3252 (.fluid_in(k_12_3252), .fluid_out(k_11_1626), .air_in(c_12_0));
valve v_12_3253 (.fluid_in(k_12_3253), .fluid_out(k_11_1626), .air_in(c_12_1));
valve v_12_3254 (.fluid_in(k_12_3254), .fluid_out(k_11_1627), .air_in(c_12_0));
valve v_12_3255 (.fluid_in(k_12_3255), .fluid_out(k_11_1627), .air_in(c_12_1));
valve v_12_3256 (.fluid_in(k_12_3256), .fluid_out(k_11_1628), .air_in(c_12_0));
valve v_12_3257 (.fluid_in(k_12_3257), .fluid_out(k_11_1628), .air_in(c_12_1));
valve v_12_3258 (.fluid_in(k_12_3258), .fluid_out(k_11_1629), .air_in(c_12_0));
valve v_12_3259 (.fluid_in(k_12_3259), .fluid_out(k_11_1629), .air_in(c_12_1));
valve v_12_3260 (.fluid_in(k_12_3260), .fluid_out(k_11_1630), .air_in(c_12_0));
valve v_12_3261 (.fluid_in(k_12_3261), .fluid_out(k_11_1630), .air_in(c_12_1));
valve v_12_3262 (.fluid_in(k_12_3262), .fluid_out(k_11_1631), .air_in(c_12_0));
valve v_12_3263 (.fluid_in(k_12_3263), .fluid_out(k_11_1631), .air_in(c_12_1));
valve v_12_3264 (.fluid_in(k_12_3264), .fluid_out(k_11_1632), .air_in(c_12_0));
valve v_12_3265 (.fluid_in(k_12_3265), .fluid_out(k_11_1632), .air_in(c_12_1));
valve v_12_3266 (.fluid_in(k_12_3266), .fluid_out(k_11_1633), .air_in(c_12_0));
valve v_12_3267 (.fluid_in(k_12_3267), .fluid_out(k_11_1633), .air_in(c_12_1));
valve v_12_3268 (.fluid_in(k_12_3268), .fluid_out(k_11_1634), .air_in(c_12_0));
valve v_12_3269 (.fluid_in(k_12_3269), .fluid_out(k_11_1634), .air_in(c_12_1));
valve v_12_3270 (.fluid_in(k_12_3270), .fluid_out(k_11_1635), .air_in(c_12_0));
valve v_12_3271 (.fluid_in(k_12_3271), .fluid_out(k_11_1635), .air_in(c_12_1));
valve v_12_3272 (.fluid_in(k_12_3272), .fluid_out(k_11_1636), .air_in(c_12_0));
valve v_12_3273 (.fluid_in(k_12_3273), .fluid_out(k_11_1636), .air_in(c_12_1));
valve v_12_3274 (.fluid_in(k_12_3274), .fluid_out(k_11_1637), .air_in(c_12_0));
valve v_12_3275 (.fluid_in(k_12_3275), .fluid_out(k_11_1637), .air_in(c_12_1));
valve v_12_3276 (.fluid_in(k_12_3276), .fluid_out(k_11_1638), .air_in(c_12_0));
valve v_12_3277 (.fluid_in(k_12_3277), .fluid_out(k_11_1638), .air_in(c_12_1));
valve v_12_3278 (.fluid_in(k_12_3278), .fluid_out(k_11_1639), .air_in(c_12_0));
valve v_12_3279 (.fluid_in(k_12_3279), .fluid_out(k_11_1639), .air_in(c_12_1));
valve v_12_3280 (.fluid_in(k_12_3280), .fluid_out(k_11_1640), .air_in(c_12_0));
valve v_12_3281 (.fluid_in(k_12_3281), .fluid_out(k_11_1640), .air_in(c_12_1));
valve v_12_3282 (.fluid_in(k_12_3282), .fluid_out(k_11_1641), .air_in(c_12_0));
valve v_12_3283 (.fluid_in(k_12_3283), .fluid_out(k_11_1641), .air_in(c_12_1));
valve v_12_3284 (.fluid_in(k_12_3284), .fluid_out(k_11_1642), .air_in(c_12_0));
valve v_12_3285 (.fluid_in(k_12_3285), .fluid_out(k_11_1642), .air_in(c_12_1));
valve v_12_3286 (.fluid_in(k_12_3286), .fluid_out(k_11_1643), .air_in(c_12_0));
valve v_12_3287 (.fluid_in(k_12_3287), .fluid_out(k_11_1643), .air_in(c_12_1));
valve v_12_3288 (.fluid_in(k_12_3288), .fluid_out(k_11_1644), .air_in(c_12_0));
valve v_12_3289 (.fluid_in(k_12_3289), .fluid_out(k_11_1644), .air_in(c_12_1));
valve v_12_3290 (.fluid_in(k_12_3290), .fluid_out(k_11_1645), .air_in(c_12_0));
valve v_12_3291 (.fluid_in(k_12_3291), .fluid_out(k_11_1645), .air_in(c_12_1));
valve v_12_3292 (.fluid_in(k_12_3292), .fluid_out(k_11_1646), .air_in(c_12_0));
valve v_12_3293 (.fluid_in(k_12_3293), .fluid_out(k_11_1646), .air_in(c_12_1));
valve v_12_3294 (.fluid_in(k_12_3294), .fluid_out(k_11_1647), .air_in(c_12_0));
valve v_12_3295 (.fluid_in(k_12_3295), .fluid_out(k_11_1647), .air_in(c_12_1));
valve v_12_3296 (.fluid_in(k_12_3296), .fluid_out(k_11_1648), .air_in(c_12_0));
valve v_12_3297 (.fluid_in(k_12_3297), .fluid_out(k_11_1648), .air_in(c_12_1));
valve v_12_3298 (.fluid_in(k_12_3298), .fluid_out(k_11_1649), .air_in(c_12_0));
valve v_12_3299 (.fluid_in(k_12_3299), .fluid_out(k_11_1649), .air_in(c_12_1));
valve v_12_3300 (.fluid_in(k_12_3300), .fluid_out(k_11_1650), .air_in(c_12_0));
valve v_12_3301 (.fluid_in(k_12_3301), .fluid_out(k_11_1650), .air_in(c_12_1));
valve v_12_3302 (.fluid_in(k_12_3302), .fluid_out(k_11_1651), .air_in(c_12_0));
valve v_12_3303 (.fluid_in(k_12_3303), .fluid_out(k_11_1651), .air_in(c_12_1));
valve v_12_3304 (.fluid_in(k_12_3304), .fluid_out(k_11_1652), .air_in(c_12_0));
valve v_12_3305 (.fluid_in(k_12_3305), .fluid_out(k_11_1652), .air_in(c_12_1));
valve v_12_3306 (.fluid_in(k_12_3306), .fluid_out(k_11_1653), .air_in(c_12_0));
valve v_12_3307 (.fluid_in(k_12_3307), .fluid_out(k_11_1653), .air_in(c_12_1));
valve v_12_3308 (.fluid_in(k_12_3308), .fluid_out(k_11_1654), .air_in(c_12_0));
valve v_12_3309 (.fluid_in(k_12_3309), .fluid_out(k_11_1654), .air_in(c_12_1));
valve v_12_3310 (.fluid_in(k_12_3310), .fluid_out(k_11_1655), .air_in(c_12_0));
valve v_12_3311 (.fluid_in(k_12_3311), .fluid_out(k_11_1655), .air_in(c_12_1));
valve v_12_3312 (.fluid_in(k_12_3312), .fluid_out(k_11_1656), .air_in(c_12_0));
valve v_12_3313 (.fluid_in(k_12_3313), .fluid_out(k_11_1656), .air_in(c_12_1));
valve v_12_3314 (.fluid_in(k_12_3314), .fluid_out(k_11_1657), .air_in(c_12_0));
valve v_12_3315 (.fluid_in(k_12_3315), .fluid_out(k_11_1657), .air_in(c_12_1));
valve v_12_3316 (.fluid_in(k_12_3316), .fluid_out(k_11_1658), .air_in(c_12_0));
valve v_12_3317 (.fluid_in(k_12_3317), .fluid_out(k_11_1658), .air_in(c_12_1));
valve v_12_3318 (.fluid_in(k_12_3318), .fluid_out(k_11_1659), .air_in(c_12_0));
valve v_12_3319 (.fluid_in(k_12_3319), .fluid_out(k_11_1659), .air_in(c_12_1));
valve v_12_3320 (.fluid_in(k_12_3320), .fluid_out(k_11_1660), .air_in(c_12_0));
valve v_12_3321 (.fluid_in(k_12_3321), .fluid_out(k_11_1660), .air_in(c_12_1));
valve v_12_3322 (.fluid_in(k_12_3322), .fluid_out(k_11_1661), .air_in(c_12_0));
valve v_12_3323 (.fluid_in(k_12_3323), .fluid_out(k_11_1661), .air_in(c_12_1));
valve v_12_3324 (.fluid_in(k_12_3324), .fluid_out(k_11_1662), .air_in(c_12_0));
valve v_12_3325 (.fluid_in(k_12_3325), .fluid_out(k_11_1662), .air_in(c_12_1));
valve v_12_3326 (.fluid_in(k_12_3326), .fluid_out(k_11_1663), .air_in(c_12_0));
valve v_12_3327 (.fluid_in(k_12_3327), .fluid_out(k_11_1663), .air_in(c_12_1));
valve v_12_3328 (.fluid_in(k_12_3328), .fluid_out(k_11_1664), .air_in(c_12_0));
valve v_12_3329 (.fluid_in(k_12_3329), .fluid_out(k_11_1664), .air_in(c_12_1));
valve v_12_3330 (.fluid_in(k_12_3330), .fluid_out(k_11_1665), .air_in(c_12_0));
valve v_12_3331 (.fluid_in(k_12_3331), .fluid_out(k_11_1665), .air_in(c_12_1));
valve v_12_3332 (.fluid_in(k_12_3332), .fluid_out(k_11_1666), .air_in(c_12_0));
valve v_12_3333 (.fluid_in(k_12_3333), .fluid_out(k_11_1666), .air_in(c_12_1));
valve v_12_3334 (.fluid_in(k_12_3334), .fluid_out(k_11_1667), .air_in(c_12_0));
valve v_12_3335 (.fluid_in(k_12_3335), .fluid_out(k_11_1667), .air_in(c_12_1));
valve v_12_3336 (.fluid_in(k_12_3336), .fluid_out(k_11_1668), .air_in(c_12_0));
valve v_12_3337 (.fluid_in(k_12_3337), .fluid_out(k_11_1668), .air_in(c_12_1));
valve v_12_3338 (.fluid_in(k_12_3338), .fluid_out(k_11_1669), .air_in(c_12_0));
valve v_12_3339 (.fluid_in(k_12_3339), .fluid_out(k_11_1669), .air_in(c_12_1));
valve v_12_3340 (.fluid_in(k_12_3340), .fluid_out(k_11_1670), .air_in(c_12_0));
valve v_12_3341 (.fluid_in(k_12_3341), .fluid_out(k_11_1670), .air_in(c_12_1));
valve v_12_3342 (.fluid_in(k_12_3342), .fluid_out(k_11_1671), .air_in(c_12_0));
valve v_12_3343 (.fluid_in(k_12_3343), .fluid_out(k_11_1671), .air_in(c_12_1));
valve v_12_3344 (.fluid_in(k_12_3344), .fluid_out(k_11_1672), .air_in(c_12_0));
valve v_12_3345 (.fluid_in(k_12_3345), .fluid_out(k_11_1672), .air_in(c_12_1));
valve v_12_3346 (.fluid_in(k_12_3346), .fluid_out(k_11_1673), .air_in(c_12_0));
valve v_12_3347 (.fluid_in(k_12_3347), .fluid_out(k_11_1673), .air_in(c_12_1));
valve v_12_3348 (.fluid_in(k_12_3348), .fluid_out(k_11_1674), .air_in(c_12_0));
valve v_12_3349 (.fluid_in(k_12_3349), .fluid_out(k_11_1674), .air_in(c_12_1));
valve v_12_3350 (.fluid_in(k_12_3350), .fluid_out(k_11_1675), .air_in(c_12_0));
valve v_12_3351 (.fluid_in(k_12_3351), .fluid_out(k_11_1675), .air_in(c_12_1));
valve v_12_3352 (.fluid_in(k_12_3352), .fluid_out(k_11_1676), .air_in(c_12_0));
valve v_12_3353 (.fluid_in(k_12_3353), .fluid_out(k_11_1676), .air_in(c_12_1));
valve v_12_3354 (.fluid_in(k_12_3354), .fluid_out(k_11_1677), .air_in(c_12_0));
valve v_12_3355 (.fluid_in(k_12_3355), .fluid_out(k_11_1677), .air_in(c_12_1));
valve v_12_3356 (.fluid_in(k_12_3356), .fluid_out(k_11_1678), .air_in(c_12_0));
valve v_12_3357 (.fluid_in(k_12_3357), .fluid_out(k_11_1678), .air_in(c_12_1));
valve v_12_3358 (.fluid_in(k_12_3358), .fluid_out(k_11_1679), .air_in(c_12_0));
valve v_12_3359 (.fluid_in(k_12_3359), .fluid_out(k_11_1679), .air_in(c_12_1));
valve v_12_3360 (.fluid_in(k_12_3360), .fluid_out(k_11_1680), .air_in(c_12_0));
valve v_12_3361 (.fluid_in(k_12_3361), .fluid_out(k_11_1680), .air_in(c_12_1));
valve v_12_3362 (.fluid_in(k_12_3362), .fluid_out(k_11_1681), .air_in(c_12_0));
valve v_12_3363 (.fluid_in(k_12_3363), .fluid_out(k_11_1681), .air_in(c_12_1));
valve v_12_3364 (.fluid_in(k_12_3364), .fluid_out(k_11_1682), .air_in(c_12_0));
valve v_12_3365 (.fluid_in(k_12_3365), .fluid_out(k_11_1682), .air_in(c_12_1));
valve v_12_3366 (.fluid_in(k_12_3366), .fluid_out(k_11_1683), .air_in(c_12_0));
valve v_12_3367 (.fluid_in(k_12_3367), .fluid_out(k_11_1683), .air_in(c_12_1));
valve v_12_3368 (.fluid_in(k_12_3368), .fluid_out(k_11_1684), .air_in(c_12_0));
valve v_12_3369 (.fluid_in(k_12_3369), .fluid_out(k_11_1684), .air_in(c_12_1));
valve v_12_3370 (.fluid_in(k_12_3370), .fluid_out(k_11_1685), .air_in(c_12_0));
valve v_12_3371 (.fluid_in(k_12_3371), .fluid_out(k_11_1685), .air_in(c_12_1));
valve v_12_3372 (.fluid_in(k_12_3372), .fluid_out(k_11_1686), .air_in(c_12_0));
valve v_12_3373 (.fluid_in(k_12_3373), .fluid_out(k_11_1686), .air_in(c_12_1));
valve v_12_3374 (.fluid_in(k_12_3374), .fluid_out(k_11_1687), .air_in(c_12_0));
valve v_12_3375 (.fluid_in(k_12_3375), .fluid_out(k_11_1687), .air_in(c_12_1));
valve v_12_3376 (.fluid_in(k_12_3376), .fluid_out(k_11_1688), .air_in(c_12_0));
valve v_12_3377 (.fluid_in(k_12_3377), .fluid_out(k_11_1688), .air_in(c_12_1));
valve v_12_3378 (.fluid_in(k_12_3378), .fluid_out(k_11_1689), .air_in(c_12_0));
valve v_12_3379 (.fluid_in(k_12_3379), .fluid_out(k_11_1689), .air_in(c_12_1));
valve v_12_3380 (.fluid_in(k_12_3380), .fluid_out(k_11_1690), .air_in(c_12_0));
valve v_12_3381 (.fluid_in(k_12_3381), .fluid_out(k_11_1690), .air_in(c_12_1));
valve v_12_3382 (.fluid_in(k_12_3382), .fluid_out(k_11_1691), .air_in(c_12_0));
valve v_12_3383 (.fluid_in(k_12_3383), .fluid_out(k_11_1691), .air_in(c_12_1));
valve v_12_3384 (.fluid_in(k_12_3384), .fluid_out(k_11_1692), .air_in(c_12_0));
valve v_12_3385 (.fluid_in(k_12_3385), .fluid_out(k_11_1692), .air_in(c_12_1));
valve v_12_3386 (.fluid_in(k_12_3386), .fluid_out(k_11_1693), .air_in(c_12_0));
valve v_12_3387 (.fluid_in(k_12_3387), .fluid_out(k_11_1693), .air_in(c_12_1));
valve v_12_3388 (.fluid_in(k_12_3388), .fluid_out(k_11_1694), .air_in(c_12_0));
valve v_12_3389 (.fluid_in(k_12_3389), .fluid_out(k_11_1694), .air_in(c_12_1));
valve v_12_3390 (.fluid_in(k_12_3390), .fluid_out(k_11_1695), .air_in(c_12_0));
valve v_12_3391 (.fluid_in(k_12_3391), .fluid_out(k_11_1695), .air_in(c_12_1));
valve v_12_3392 (.fluid_in(k_12_3392), .fluid_out(k_11_1696), .air_in(c_12_0));
valve v_12_3393 (.fluid_in(k_12_3393), .fluid_out(k_11_1696), .air_in(c_12_1));
valve v_12_3394 (.fluid_in(k_12_3394), .fluid_out(k_11_1697), .air_in(c_12_0));
valve v_12_3395 (.fluid_in(k_12_3395), .fluid_out(k_11_1697), .air_in(c_12_1));
valve v_12_3396 (.fluid_in(k_12_3396), .fluid_out(k_11_1698), .air_in(c_12_0));
valve v_12_3397 (.fluid_in(k_12_3397), .fluid_out(k_11_1698), .air_in(c_12_1));
valve v_12_3398 (.fluid_in(k_12_3398), .fluid_out(k_11_1699), .air_in(c_12_0));
valve v_12_3399 (.fluid_in(k_12_3399), .fluid_out(k_11_1699), .air_in(c_12_1));
valve v_12_3400 (.fluid_in(k_12_3400), .fluid_out(k_11_1700), .air_in(c_12_0));
valve v_12_3401 (.fluid_in(k_12_3401), .fluid_out(k_11_1700), .air_in(c_12_1));
valve v_12_3402 (.fluid_in(k_12_3402), .fluid_out(k_11_1701), .air_in(c_12_0));
valve v_12_3403 (.fluid_in(k_12_3403), .fluid_out(k_11_1701), .air_in(c_12_1));
valve v_12_3404 (.fluid_in(k_12_3404), .fluid_out(k_11_1702), .air_in(c_12_0));
valve v_12_3405 (.fluid_in(k_12_3405), .fluid_out(k_11_1702), .air_in(c_12_1));
valve v_12_3406 (.fluid_in(k_12_3406), .fluid_out(k_11_1703), .air_in(c_12_0));
valve v_12_3407 (.fluid_in(k_12_3407), .fluid_out(k_11_1703), .air_in(c_12_1));
valve v_12_3408 (.fluid_in(k_12_3408), .fluid_out(k_11_1704), .air_in(c_12_0));
valve v_12_3409 (.fluid_in(k_12_3409), .fluid_out(k_11_1704), .air_in(c_12_1));
valve v_12_3410 (.fluid_in(k_12_3410), .fluid_out(k_11_1705), .air_in(c_12_0));
valve v_12_3411 (.fluid_in(k_12_3411), .fluid_out(k_11_1705), .air_in(c_12_1));
valve v_12_3412 (.fluid_in(k_12_3412), .fluid_out(k_11_1706), .air_in(c_12_0));
valve v_12_3413 (.fluid_in(k_12_3413), .fluid_out(k_11_1706), .air_in(c_12_1));
valve v_12_3414 (.fluid_in(k_12_3414), .fluid_out(k_11_1707), .air_in(c_12_0));
valve v_12_3415 (.fluid_in(k_12_3415), .fluid_out(k_11_1707), .air_in(c_12_1));
valve v_12_3416 (.fluid_in(k_12_3416), .fluid_out(k_11_1708), .air_in(c_12_0));
valve v_12_3417 (.fluid_in(k_12_3417), .fluid_out(k_11_1708), .air_in(c_12_1));
valve v_12_3418 (.fluid_in(k_12_3418), .fluid_out(k_11_1709), .air_in(c_12_0));
valve v_12_3419 (.fluid_in(k_12_3419), .fluid_out(k_11_1709), .air_in(c_12_1));
valve v_12_3420 (.fluid_in(k_12_3420), .fluid_out(k_11_1710), .air_in(c_12_0));
valve v_12_3421 (.fluid_in(k_12_3421), .fluid_out(k_11_1710), .air_in(c_12_1));
valve v_12_3422 (.fluid_in(k_12_3422), .fluid_out(k_11_1711), .air_in(c_12_0));
valve v_12_3423 (.fluid_in(k_12_3423), .fluid_out(k_11_1711), .air_in(c_12_1));
valve v_12_3424 (.fluid_in(k_12_3424), .fluid_out(k_11_1712), .air_in(c_12_0));
valve v_12_3425 (.fluid_in(k_12_3425), .fluid_out(k_11_1712), .air_in(c_12_1));
valve v_12_3426 (.fluid_in(k_12_3426), .fluid_out(k_11_1713), .air_in(c_12_0));
valve v_12_3427 (.fluid_in(k_12_3427), .fluid_out(k_11_1713), .air_in(c_12_1));
valve v_12_3428 (.fluid_in(k_12_3428), .fluid_out(k_11_1714), .air_in(c_12_0));
valve v_12_3429 (.fluid_in(k_12_3429), .fluid_out(k_11_1714), .air_in(c_12_1));
valve v_12_3430 (.fluid_in(k_12_3430), .fluid_out(k_11_1715), .air_in(c_12_0));
valve v_12_3431 (.fluid_in(k_12_3431), .fluid_out(k_11_1715), .air_in(c_12_1));
valve v_12_3432 (.fluid_in(k_12_3432), .fluid_out(k_11_1716), .air_in(c_12_0));
valve v_12_3433 (.fluid_in(k_12_3433), .fluid_out(k_11_1716), .air_in(c_12_1));
valve v_12_3434 (.fluid_in(k_12_3434), .fluid_out(k_11_1717), .air_in(c_12_0));
valve v_12_3435 (.fluid_in(k_12_3435), .fluid_out(k_11_1717), .air_in(c_12_1));
valve v_12_3436 (.fluid_in(k_12_3436), .fluid_out(k_11_1718), .air_in(c_12_0));
valve v_12_3437 (.fluid_in(k_12_3437), .fluid_out(k_11_1718), .air_in(c_12_1));
valve v_12_3438 (.fluid_in(k_12_3438), .fluid_out(k_11_1719), .air_in(c_12_0));
valve v_12_3439 (.fluid_in(k_12_3439), .fluid_out(k_11_1719), .air_in(c_12_1));
valve v_12_3440 (.fluid_in(k_12_3440), .fluid_out(k_11_1720), .air_in(c_12_0));
valve v_12_3441 (.fluid_in(k_12_3441), .fluid_out(k_11_1720), .air_in(c_12_1));
valve v_12_3442 (.fluid_in(k_12_3442), .fluid_out(k_11_1721), .air_in(c_12_0));
valve v_12_3443 (.fluid_in(k_12_3443), .fluid_out(k_11_1721), .air_in(c_12_1));
valve v_12_3444 (.fluid_in(k_12_3444), .fluid_out(k_11_1722), .air_in(c_12_0));
valve v_12_3445 (.fluid_in(k_12_3445), .fluid_out(k_11_1722), .air_in(c_12_1));
valve v_12_3446 (.fluid_in(k_12_3446), .fluid_out(k_11_1723), .air_in(c_12_0));
valve v_12_3447 (.fluid_in(k_12_3447), .fluid_out(k_11_1723), .air_in(c_12_1));
valve v_12_3448 (.fluid_in(k_12_3448), .fluid_out(k_11_1724), .air_in(c_12_0));
valve v_12_3449 (.fluid_in(k_12_3449), .fluid_out(k_11_1724), .air_in(c_12_1));
valve v_12_3450 (.fluid_in(k_12_3450), .fluid_out(k_11_1725), .air_in(c_12_0));
valve v_12_3451 (.fluid_in(k_12_3451), .fluid_out(k_11_1725), .air_in(c_12_1));
valve v_12_3452 (.fluid_in(k_12_3452), .fluid_out(k_11_1726), .air_in(c_12_0));
valve v_12_3453 (.fluid_in(k_12_3453), .fluid_out(k_11_1726), .air_in(c_12_1));
valve v_12_3454 (.fluid_in(k_12_3454), .fluid_out(k_11_1727), .air_in(c_12_0));
valve v_12_3455 (.fluid_in(k_12_3455), .fluid_out(k_11_1727), .air_in(c_12_1));
valve v_12_3456 (.fluid_in(k_12_3456), .fluid_out(k_11_1728), .air_in(c_12_0));
valve v_12_3457 (.fluid_in(k_12_3457), .fluid_out(k_11_1728), .air_in(c_12_1));
valve v_12_3458 (.fluid_in(k_12_3458), .fluid_out(k_11_1729), .air_in(c_12_0));
valve v_12_3459 (.fluid_in(k_12_3459), .fluid_out(k_11_1729), .air_in(c_12_1));
valve v_12_3460 (.fluid_in(k_12_3460), .fluid_out(k_11_1730), .air_in(c_12_0));
valve v_12_3461 (.fluid_in(k_12_3461), .fluid_out(k_11_1730), .air_in(c_12_1));
valve v_12_3462 (.fluid_in(k_12_3462), .fluid_out(k_11_1731), .air_in(c_12_0));
valve v_12_3463 (.fluid_in(k_12_3463), .fluid_out(k_11_1731), .air_in(c_12_1));
valve v_12_3464 (.fluid_in(k_12_3464), .fluid_out(k_11_1732), .air_in(c_12_0));
valve v_12_3465 (.fluid_in(k_12_3465), .fluid_out(k_11_1732), .air_in(c_12_1));
valve v_12_3466 (.fluid_in(k_12_3466), .fluid_out(k_11_1733), .air_in(c_12_0));
valve v_12_3467 (.fluid_in(k_12_3467), .fluid_out(k_11_1733), .air_in(c_12_1));
valve v_12_3468 (.fluid_in(k_12_3468), .fluid_out(k_11_1734), .air_in(c_12_0));
valve v_12_3469 (.fluid_in(k_12_3469), .fluid_out(k_11_1734), .air_in(c_12_1));
valve v_12_3470 (.fluid_in(k_12_3470), .fluid_out(k_11_1735), .air_in(c_12_0));
valve v_12_3471 (.fluid_in(k_12_3471), .fluid_out(k_11_1735), .air_in(c_12_1));
valve v_12_3472 (.fluid_in(k_12_3472), .fluid_out(k_11_1736), .air_in(c_12_0));
valve v_12_3473 (.fluid_in(k_12_3473), .fluid_out(k_11_1736), .air_in(c_12_1));
valve v_12_3474 (.fluid_in(k_12_3474), .fluid_out(k_11_1737), .air_in(c_12_0));
valve v_12_3475 (.fluid_in(k_12_3475), .fluid_out(k_11_1737), .air_in(c_12_1));
valve v_12_3476 (.fluid_in(k_12_3476), .fluid_out(k_11_1738), .air_in(c_12_0));
valve v_12_3477 (.fluid_in(k_12_3477), .fluid_out(k_11_1738), .air_in(c_12_1));
valve v_12_3478 (.fluid_in(k_12_3478), .fluid_out(k_11_1739), .air_in(c_12_0));
valve v_12_3479 (.fluid_in(k_12_3479), .fluid_out(k_11_1739), .air_in(c_12_1));
valve v_12_3480 (.fluid_in(k_12_3480), .fluid_out(k_11_1740), .air_in(c_12_0));
valve v_12_3481 (.fluid_in(k_12_3481), .fluid_out(k_11_1740), .air_in(c_12_1));
valve v_12_3482 (.fluid_in(k_12_3482), .fluid_out(k_11_1741), .air_in(c_12_0));
valve v_12_3483 (.fluid_in(k_12_3483), .fluid_out(k_11_1741), .air_in(c_12_1));
valve v_12_3484 (.fluid_in(k_12_3484), .fluid_out(k_11_1742), .air_in(c_12_0));
valve v_12_3485 (.fluid_in(k_12_3485), .fluid_out(k_11_1742), .air_in(c_12_1));
valve v_12_3486 (.fluid_in(k_12_3486), .fluid_out(k_11_1743), .air_in(c_12_0));
valve v_12_3487 (.fluid_in(k_12_3487), .fluid_out(k_11_1743), .air_in(c_12_1));
valve v_12_3488 (.fluid_in(k_12_3488), .fluid_out(k_11_1744), .air_in(c_12_0));
valve v_12_3489 (.fluid_in(k_12_3489), .fluid_out(k_11_1744), .air_in(c_12_1));
valve v_12_3490 (.fluid_in(k_12_3490), .fluid_out(k_11_1745), .air_in(c_12_0));
valve v_12_3491 (.fluid_in(k_12_3491), .fluid_out(k_11_1745), .air_in(c_12_1));
valve v_12_3492 (.fluid_in(k_12_3492), .fluid_out(k_11_1746), .air_in(c_12_0));
valve v_12_3493 (.fluid_in(k_12_3493), .fluid_out(k_11_1746), .air_in(c_12_1));
valve v_12_3494 (.fluid_in(k_12_3494), .fluid_out(k_11_1747), .air_in(c_12_0));
valve v_12_3495 (.fluid_in(k_12_3495), .fluid_out(k_11_1747), .air_in(c_12_1));
valve v_12_3496 (.fluid_in(k_12_3496), .fluid_out(k_11_1748), .air_in(c_12_0));
valve v_12_3497 (.fluid_in(k_12_3497), .fluid_out(k_11_1748), .air_in(c_12_1));
valve v_12_3498 (.fluid_in(k_12_3498), .fluid_out(k_11_1749), .air_in(c_12_0));
valve v_12_3499 (.fluid_in(k_12_3499), .fluid_out(k_11_1749), .air_in(c_12_1));
valve v_12_3500 (.fluid_in(k_12_3500), .fluid_out(k_11_1750), .air_in(c_12_0));
valve v_12_3501 (.fluid_in(k_12_3501), .fluid_out(k_11_1750), .air_in(c_12_1));
valve v_12_3502 (.fluid_in(k_12_3502), .fluid_out(k_11_1751), .air_in(c_12_0));
valve v_12_3503 (.fluid_in(k_12_3503), .fluid_out(k_11_1751), .air_in(c_12_1));
valve v_12_3504 (.fluid_in(k_12_3504), .fluid_out(k_11_1752), .air_in(c_12_0));
valve v_12_3505 (.fluid_in(k_12_3505), .fluid_out(k_11_1752), .air_in(c_12_1));
valve v_12_3506 (.fluid_in(k_12_3506), .fluid_out(k_11_1753), .air_in(c_12_0));
valve v_12_3507 (.fluid_in(k_12_3507), .fluid_out(k_11_1753), .air_in(c_12_1));
valve v_12_3508 (.fluid_in(k_12_3508), .fluid_out(k_11_1754), .air_in(c_12_0));
valve v_12_3509 (.fluid_in(k_12_3509), .fluid_out(k_11_1754), .air_in(c_12_1));
valve v_12_3510 (.fluid_in(k_12_3510), .fluid_out(k_11_1755), .air_in(c_12_0));
valve v_12_3511 (.fluid_in(k_12_3511), .fluid_out(k_11_1755), .air_in(c_12_1));
valve v_12_3512 (.fluid_in(k_12_3512), .fluid_out(k_11_1756), .air_in(c_12_0));
valve v_12_3513 (.fluid_in(k_12_3513), .fluid_out(k_11_1756), .air_in(c_12_1));
valve v_12_3514 (.fluid_in(k_12_3514), .fluid_out(k_11_1757), .air_in(c_12_0));
valve v_12_3515 (.fluid_in(k_12_3515), .fluid_out(k_11_1757), .air_in(c_12_1));
valve v_12_3516 (.fluid_in(k_12_3516), .fluid_out(k_11_1758), .air_in(c_12_0));
valve v_12_3517 (.fluid_in(k_12_3517), .fluid_out(k_11_1758), .air_in(c_12_1));
valve v_12_3518 (.fluid_in(k_12_3518), .fluid_out(k_11_1759), .air_in(c_12_0));
valve v_12_3519 (.fluid_in(k_12_3519), .fluid_out(k_11_1759), .air_in(c_12_1));
valve v_12_3520 (.fluid_in(k_12_3520), .fluid_out(k_11_1760), .air_in(c_12_0));
valve v_12_3521 (.fluid_in(k_12_3521), .fluid_out(k_11_1760), .air_in(c_12_1));
valve v_12_3522 (.fluid_in(k_12_3522), .fluid_out(k_11_1761), .air_in(c_12_0));
valve v_12_3523 (.fluid_in(k_12_3523), .fluid_out(k_11_1761), .air_in(c_12_1));
valve v_12_3524 (.fluid_in(k_12_3524), .fluid_out(k_11_1762), .air_in(c_12_0));
valve v_12_3525 (.fluid_in(k_12_3525), .fluid_out(k_11_1762), .air_in(c_12_1));
valve v_12_3526 (.fluid_in(k_12_3526), .fluid_out(k_11_1763), .air_in(c_12_0));
valve v_12_3527 (.fluid_in(k_12_3527), .fluid_out(k_11_1763), .air_in(c_12_1));
valve v_12_3528 (.fluid_in(k_12_3528), .fluid_out(k_11_1764), .air_in(c_12_0));
valve v_12_3529 (.fluid_in(k_12_3529), .fluid_out(k_11_1764), .air_in(c_12_1));
valve v_12_3530 (.fluid_in(k_12_3530), .fluid_out(k_11_1765), .air_in(c_12_0));
valve v_12_3531 (.fluid_in(k_12_3531), .fluid_out(k_11_1765), .air_in(c_12_1));
valve v_12_3532 (.fluid_in(k_12_3532), .fluid_out(k_11_1766), .air_in(c_12_0));
valve v_12_3533 (.fluid_in(k_12_3533), .fluid_out(k_11_1766), .air_in(c_12_1));
valve v_12_3534 (.fluid_in(k_12_3534), .fluid_out(k_11_1767), .air_in(c_12_0));
valve v_12_3535 (.fluid_in(k_12_3535), .fluid_out(k_11_1767), .air_in(c_12_1));
valve v_12_3536 (.fluid_in(k_12_3536), .fluid_out(k_11_1768), .air_in(c_12_0));
valve v_12_3537 (.fluid_in(k_12_3537), .fluid_out(k_11_1768), .air_in(c_12_1));
valve v_12_3538 (.fluid_in(k_12_3538), .fluid_out(k_11_1769), .air_in(c_12_0));
valve v_12_3539 (.fluid_in(k_12_3539), .fluid_out(k_11_1769), .air_in(c_12_1));
valve v_12_3540 (.fluid_in(k_12_3540), .fluid_out(k_11_1770), .air_in(c_12_0));
valve v_12_3541 (.fluid_in(k_12_3541), .fluid_out(k_11_1770), .air_in(c_12_1));
valve v_12_3542 (.fluid_in(k_12_3542), .fluid_out(k_11_1771), .air_in(c_12_0));
valve v_12_3543 (.fluid_in(k_12_3543), .fluid_out(k_11_1771), .air_in(c_12_1));
valve v_12_3544 (.fluid_in(k_12_3544), .fluid_out(k_11_1772), .air_in(c_12_0));
valve v_12_3545 (.fluid_in(k_12_3545), .fluid_out(k_11_1772), .air_in(c_12_1));
valve v_12_3546 (.fluid_in(k_12_3546), .fluid_out(k_11_1773), .air_in(c_12_0));
valve v_12_3547 (.fluid_in(k_12_3547), .fluid_out(k_11_1773), .air_in(c_12_1));
valve v_12_3548 (.fluid_in(k_12_3548), .fluid_out(k_11_1774), .air_in(c_12_0));
valve v_12_3549 (.fluid_in(k_12_3549), .fluid_out(k_11_1774), .air_in(c_12_1));
valve v_12_3550 (.fluid_in(k_12_3550), .fluid_out(k_11_1775), .air_in(c_12_0));
valve v_12_3551 (.fluid_in(k_12_3551), .fluid_out(k_11_1775), .air_in(c_12_1));
valve v_12_3552 (.fluid_in(k_12_3552), .fluid_out(k_11_1776), .air_in(c_12_0));
valve v_12_3553 (.fluid_in(k_12_3553), .fluid_out(k_11_1776), .air_in(c_12_1));
valve v_12_3554 (.fluid_in(k_12_3554), .fluid_out(k_11_1777), .air_in(c_12_0));
valve v_12_3555 (.fluid_in(k_12_3555), .fluid_out(k_11_1777), .air_in(c_12_1));
valve v_12_3556 (.fluid_in(k_12_3556), .fluid_out(k_11_1778), .air_in(c_12_0));
valve v_12_3557 (.fluid_in(k_12_3557), .fluid_out(k_11_1778), .air_in(c_12_1));
valve v_12_3558 (.fluid_in(k_12_3558), .fluid_out(k_11_1779), .air_in(c_12_0));
valve v_12_3559 (.fluid_in(k_12_3559), .fluid_out(k_11_1779), .air_in(c_12_1));
valve v_12_3560 (.fluid_in(k_12_3560), .fluid_out(k_11_1780), .air_in(c_12_0));
valve v_12_3561 (.fluid_in(k_12_3561), .fluid_out(k_11_1780), .air_in(c_12_1));
valve v_12_3562 (.fluid_in(k_12_3562), .fluid_out(k_11_1781), .air_in(c_12_0));
valve v_12_3563 (.fluid_in(k_12_3563), .fluid_out(k_11_1781), .air_in(c_12_1));
valve v_12_3564 (.fluid_in(k_12_3564), .fluid_out(k_11_1782), .air_in(c_12_0));
valve v_12_3565 (.fluid_in(k_12_3565), .fluid_out(k_11_1782), .air_in(c_12_1));
valve v_12_3566 (.fluid_in(k_12_3566), .fluid_out(k_11_1783), .air_in(c_12_0));
valve v_12_3567 (.fluid_in(k_12_3567), .fluid_out(k_11_1783), .air_in(c_12_1));
valve v_12_3568 (.fluid_in(k_12_3568), .fluid_out(k_11_1784), .air_in(c_12_0));
valve v_12_3569 (.fluid_in(k_12_3569), .fluid_out(k_11_1784), .air_in(c_12_1));
valve v_12_3570 (.fluid_in(k_12_3570), .fluid_out(k_11_1785), .air_in(c_12_0));
valve v_12_3571 (.fluid_in(k_12_3571), .fluid_out(k_11_1785), .air_in(c_12_1));
valve v_12_3572 (.fluid_in(k_12_3572), .fluid_out(k_11_1786), .air_in(c_12_0));
valve v_12_3573 (.fluid_in(k_12_3573), .fluid_out(k_11_1786), .air_in(c_12_1));
valve v_12_3574 (.fluid_in(k_12_3574), .fluid_out(k_11_1787), .air_in(c_12_0));
valve v_12_3575 (.fluid_in(k_12_3575), .fluid_out(k_11_1787), .air_in(c_12_1));
valve v_12_3576 (.fluid_in(k_12_3576), .fluid_out(k_11_1788), .air_in(c_12_0));
valve v_12_3577 (.fluid_in(k_12_3577), .fluid_out(k_11_1788), .air_in(c_12_1));
valve v_12_3578 (.fluid_in(k_12_3578), .fluid_out(k_11_1789), .air_in(c_12_0));
valve v_12_3579 (.fluid_in(k_12_3579), .fluid_out(k_11_1789), .air_in(c_12_1));
valve v_12_3580 (.fluid_in(k_12_3580), .fluid_out(k_11_1790), .air_in(c_12_0));
valve v_12_3581 (.fluid_in(k_12_3581), .fluid_out(k_11_1790), .air_in(c_12_1));
valve v_12_3582 (.fluid_in(k_12_3582), .fluid_out(k_11_1791), .air_in(c_12_0));
valve v_12_3583 (.fluid_in(k_12_3583), .fluid_out(k_11_1791), .air_in(c_12_1));
valve v_12_3584 (.fluid_in(k_12_3584), .fluid_out(k_11_1792), .air_in(c_12_0));
valve v_12_3585 (.fluid_in(k_12_3585), .fluid_out(k_11_1792), .air_in(c_12_1));
valve v_12_3586 (.fluid_in(k_12_3586), .fluid_out(k_11_1793), .air_in(c_12_0));
valve v_12_3587 (.fluid_in(k_12_3587), .fluid_out(k_11_1793), .air_in(c_12_1));
valve v_12_3588 (.fluid_in(k_12_3588), .fluid_out(k_11_1794), .air_in(c_12_0));
valve v_12_3589 (.fluid_in(k_12_3589), .fluid_out(k_11_1794), .air_in(c_12_1));
valve v_12_3590 (.fluid_in(k_12_3590), .fluid_out(k_11_1795), .air_in(c_12_0));
valve v_12_3591 (.fluid_in(k_12_3591), .fluid_out(k_11_1795), .air_in(c_12_1));
valve v_12_3592 (.fluid_in(k_12_3592), .fluid_out(k_11_1796), .air_in(c_12_0));
valve v_12_3593 (.fluid_in(k_12_3593), .fluid_out(k_11_1796), .air_in(c_12_1));
valve v_12_3594 (.fluid_in(k_12_3594), .fluid_out(k_11_1797), .air_in(c_12_0));
valve v_12_3595 (.fluid_in(k_12_3595), .fluid_out(k_11_1797), .air_in(c_12_1));
valve v_12_3596 (.fluid_in(k_12_3596), .fluid_out(k_11_1798), .air_in(c_12_0));
valve v_12_3597 (.fluid_in(k_12_3597), .fluid_out(k_11_1798), .air_in(c_12_1));
valve v_12_3598 (.fluid_in(k_12_3598), .fluid_out(k_11_1799), .air_in(c_12_0));
valve v_12_3599 (.fluid_in(k_12_3599), .fluid_out(k_11_1799), .air_in(c_12_1));
valve v_12_3600 (.fluid_in(k_12_3600), .fluid_out(k_11_1800), .air_in(c_12_0));
valve v_12_3601 (.fluid_in(k_12_3601), .fluid_out(k_11_1800), .air_in(c_12_1));
valve v_12_3602 (.fluid_in(k_12_3602), .fluid_out(k_11_1801), .air_in(c_12_0));
valve v_12_3603 (.fluid_in(k_12_3603), .fluid_out(k_11_1801), .air_in(c_12_1));
valve v_12_3604 (.fluid_in(k_12_3604), .fluid_out(k_11_1802), .air_in(c_12_0));
valve v_12_3605 (.fluid_in(k_12_3605), .fluid_out(k_11_1802), .air_in(c_12_1));
valve v_12_3606 (.fluid_in(k_12_3606), .fluid_out(k_11_1803), .air_in(c_12_0));
valve v_12_3607 (.fluid_in(k_12_3607), .fluid_out(k_11_1803), .air_in(c_12_1));
valve v_12_3608 (.fluid_in(k_12_3608), .fluid_out(k_11_1804), .air_in(c_12_0));
valve v_12_3609 (.fluid_in(k_12_3609), .fluid_out(k_11_1804), .air_in(c_12_1));
valve v_12_3610 (.fluid_in(k_12_3610), .fluid_out(k_11_1805), .air_in(c_12_0));
valve v_12_3611 (.fluid_in(k_12_3611), .fluid_out(k_11_1805), .air_in(c_12_1));
valve v_12_3612 (.fluid_in(k_12_3612), .fluid_out(k_11_1806), .air_in(c_12_0));
valve v_12_3613 (.fluid_in(k_12_3613), .fluid_out(k_11_1806), .air_in(c_12_1));
valve v_12_3614 (.fluid_in(k_12_3614), .fluid_out(k_11_1807), .air_in(c_12_0));
valve v_12_3615 (.fluid_in(k_12_3615), .fluid_out(k_11_1807), .air_in(c_12_1));
valve v_12_3616 (.fluid_in(k_12_3616), .fluid_out(k_11_1808), .air_in(c_12_0));
valve v_12_3617 (.fluid_in(k_12_3617), .fluid_out(k_11_1808), .air_in(c_12_1));
valve v_12_3618 (.fluid_in(k_12_3618), .fluid_out(k_11_1809), .air_in(c_12_0));
valve v_12_3619 (.fluid_in(k_12_3619), .fluid_out(k_11_1809), .air_in(c_12_1));
valve v_12_3620 (.fluid_in(k_12_3620), .fluid_out(k_11_1810), .air_in(c_12_0));
valve v_12_3621 (.fluid_in(k_12_3621), .fluid_out(k_11_1810), .air_in(c_12_1));
valve v_12_3622 (.fluid_in(k_12_3622), .fluid_out(k_11_1811), .air_in(c_12_0));
valve v_12_3623 (.fluid_in(k_12_3623), .fluid_out(k_11_1811), .air_in(c_12_1));
valve v_12_3624 (.fluid_in(k_12_3624), .fluid_out(k_11_1812), .air_in(c_12_0));
valve v_12_3625 (.fluid_in(k_12_3625), .fluid_out(k_11_1812), .air_in(c_12_1));
valve v_12_3626 (.fluid_in(k_12_3626), .fluid_out(k_11_1813), .air_in(c_12_0));
valve v_12_3627 (.fluid_in(k_12_3627), .fluid_out(k_11_1813), .air_in(c_12_1));
valve v_12_3628 (.fluid_in(k_12_3628), .fluid_out(k_11_1814), .air_in(c_12_0));
valve v_12_3629 (.fluid_in(k_12_3629), .fluid_out(k_11_1814), .air_in(c_12_1));
valve v_12_3630 (.fluid_in(k_12_3630), .fluid_out(k_11_1815), .air_in(c_12_0));
valve v_12_3631 (.fluid_in(k_12_3631), .fluid_out(k_11_1815), .air_in(c_12_1));
valve v_12_3632 (.fluid_in(k_12_3632), .fluid_out(k_11_1816), .air_in(c_12_0));
valve v_12_3633 (.fluid_in(k_12_3633), .fluid_out(k_11_1816), .air_in(c_12_1));
valve v_12_3634 (.fluid_in(k_12_3634), .fluid_out(k_11_1817), .air_in(c_12_0));
valve v_12_3635 (.fluid_in(k_12_3635), .fluid_out(k_11_1817), .air_in(c_12_1));
valve v_12_3636 (.fluid_in(k_12_3636), .fluid_out(k_11_1818), .air_in(c_12_0));
valve v_12_3637 (.fluid_in(k_12_3637), .fluid_out(k_11_1818), .air_in(c_12_1));
valve v_12_3638 (.fluid_in(k_12_3638), .fluid_out(k_11_1819), .air_in(c_12_0));
valve v_12_3639 (.fluid_in(k_12_3639), .fluid_out(k_11_1819), .air_in(c_12_1));
valve v_12_3640 (.fluid_in(k_12_3640), .fluid_out(k_11_1820), .air_in(c_12_0));
valve v_12_3641 (.fluid_in(k_12_3641), .fluid_out(k_11_1820), .air_in(c_12_1));
valve v_12_3642 (.fluid_in(k_12_3642), .fluid_out(k_11_1821), .air_in(c_12_0));
valve v_12_3643 (.fluid_in(k_12_3643), .fluid_out(k_11_1821), .air_in(c_12_1));
valve v_12_3644 (.fluid_in(k_12_3644), .fluid_out(k_11_1822), .air_in(c_12_0));
valve v_12_3645 (.fluid_in(k_12_3645), .fluid_out(k_11_1822), .air_in(c_12_1));
valve v_12_3646 (.fluid_in(k_12_3646), .fluid_out(k_11_1823), .air_in(c_12_0));
valve v_12_3647 (.fluid_in(k_12_3647), .fluid_out(k_11_1823), .air_in(c_12_1));
valve v_12_3648 (.fluid_in(k_12_3648), .fluid_out(k_11_1824), .air_in(c_12_0));
valve v_12_3649 (.fluid_in(k_12_3649), .fluid_out(k_11_1824), .air_in(c_12_1));
valve v_12_3650 (.fluid_in(k_12_3650), .fluid_out(k_11_1825), .air_in(c_12_0));
valve v_12_3651 (.fluid_in(k_12_3651), .fluid_out(k_11_1825), .air_in(c_12_1));
valve v_12_3652 (.fluid_in(k_12_3652), .fluid_out(k_11_1826), .air_in(c_12_0));
valve v_12_3653 (.fluid_in(k_12_3653), .fluid_out(k_11_1826), .air_in(c_12_1));
valve v_12_3654 (.fluid_in(k_12_3654), .fluid_out(k_11_1827), .air_in(c_12_0));
valve v_12_3655 (.fluid_in(k_12_3655), .fluid_out(k_11_1827), .air_in(c_12_1));
valve v_12_3656 (.fluid_in(k_12_3656), .fluid_out(k_11_1828), .air_in(c_12_0));
valve v_12_3657 (.fluid_in(k_12_3657), .fluid_out(k_11_1828), .air_in(c_12_1));
valve v_12_3658 (.fluid_in(k_12_3658), .fluid_out(k_11_1829), .air_in(c_12_0));
valve v_12_3659 (.fluid_in(k_12_3659), .fluid_out(k_11_1829), .air_in(c_12_1));
valve v_12_3660 (.fluid_in(k_12_3660), .fluid_out(k_11_1830), .air_in(c_12_0));
valve v_12_3661 (.fluid_in(k_12_3661), .fluid_out(k_11_1830), .air_in(c_12_1));
valve v_12_3662 (.fluid_in(k_12_3662), .fluid_out(k_11_1831), .air_in(c_12_0));
valve v_12_3663 (.fluid_in(k_12_3663), .fluid_out(k_11_1831), .air_in(c_12_1));
valve v_12_3664 (.fluid_in(k_12_3664), .fluid_out(k_11_1832), .air_in(c_12_0));
valve v_12_3665 (.fluid_in(k_12_3665), .fluid_out(k_11_1832), .air_in(c_12_1));
valve v_12_3666 (.fluid_in(k_12_3666), .fluid_out(k_11_1833), .air_in(c_12_0));
valve v_12_3667 (.fluid_in(k_12_3667), .fluid_out(k_11_1833), .air_in(c_12_1));
valve v_12_3668 (.fluid_in(k_12_3668), .fluid_out(k_11_1834), .air_in(c_12_0));
valve v_12_3669 (.fluid_in(k_12_3669), .fluid_out(k_11_1834), .air_in(c_12_1));
valve v_12_3670 (.fluid_in(k_12_3670), .fluid_out(k_11_1835), .air_in(c_12_0));
valve v_12_3671 (.fluid_in(k_12_3671), .fluid_out(k_11_1835), .air_in(c_12_1));
valve v_12_3672 (.fluid_in(k_12_3672), .fluid_out(k_11_1836), .air_in(c_12_0));
valve v_12_3673 (.fluid_in(k_12_3673), .fluid_out(k_11_1836), .air_in(c_12_1));
valve v_12_3674 (.fluid_in(k_12_3674), .fluid_out(k_11_1837), .air_in(c_12_0));
valve v_12_3675 (.fluid_in(k_12_3675), .fluid_out(k_11_1837), .air_in(c_12_1));
valve v_12_3676 (.fluid_in(k_12_3676), .fluid_out(k_11_1838), .air_in(c_12_0));
valve v_12_3677 (.fluid_in(k_12_3677), .fluid_out(k_11_1838), .air_in(c_12_1));
valve v_12_3678 (.fluid_in(k_12_3678), .fluid_out(k_11_1839), .air_in(c_12_0));
valve v_12_3679 (.fluid_in(k_12_3679), .fluid_out(k_11_1839), .air_in(c_12_1));
valve v_12_3680 (.fluid_in(k_12_3680), .fluid_out(k_11_1840), .air_in(c_12_0));
valve v_12_3681 (.fluid_in(k_12_3681), .fluid_out(k_11_1840), .air_in(c_12_1));
valve v_12_3682 (.fluid_in(k_12_3682), .fluid_out(k_11_1841), .air_in(c_12_0));
valve v_12_3683 (.fluid_in(k_12_3683), .fluid_out(k_11_1841), .air_in(c_12_1));
valve v_12_3684 (.fluid_in(k_12_3684), .fluid_out(k_11_1842), .air_in(c_12_0));
valve v_12_3685 (.fluid_in(k_12_3685), .fluid_out(k_11_1842), .air_in(c_12_1));
valve v_12_3686 (.fluid_in(k_12_3686), .fluid_out(k_11_1843), .air_in(c_12_0));
valve v_12_3687 (.fluid_in(k_12_3687), .fluid_out(k_11_1843), .air_in(c_12_1));
valve v_12_3688 (.fluid_in(k_12_3688), .fluid_out(k_11_1844), .air_in(c_12_0));
valve v_12_3689 (.fluid_in(k_12_3689), .fluid_out(k_11_1844), .air_in(c_12_1));
valve v_12_3690 (.fluid_in(k_12_3690), .fluid_out(k_11_1845), .air_in(c_12_0));
valve v_12_3691 (.fluid_in(k_12_3691), .fluid_out(k_11_1845), .air_in(c_12_1));
valve v_12_3692 (.fluid_in(k_12_3692), .fluid_out(k_11_1846), .air_in(c_12_0));
valve v_12_3693 (.fluid_in(k_12_3693), .fluid_out(k_11_1846), .air_in(c_12_1));
valve v_12_3694 (.fluid_in(k_12_3694), .fluid_out(k_11_1847), .air_in(c_12_0));
valve v_12_3695 (.fluid_in(k_12_3695), .fluid_out(k_11_1847), .air_in(c_12_1));
valve v_12_3696 (.fluid_in(k_12_3696), .fluid_out(k_11_1848), .air_in(c_12_0));
valve v_12_3697 (.fluid_in(k_12_3697), .fluid_out(k_11_1848), .air_in(c_12_1));
valve v_12_3698 (.fluid_in(k_12_3698), .fluid_out(k_11_1849), .air_in(c_12_0));
valve v_12_3699 (.fluid_in(k_12_3699), .fluid_out(k_11_1849), .air_in(c_12_1));
valve v_12_3700 (.fluid_in(k_12_3700), .fluid_out(k_11_1850), .air_in(c_12_0));
valve v_12_3701 (.fluid_in(k_12_3701), .fluid_out(k_11_1850), .air_in(c_12_1));
valve v_12_3702 (.fluid_in(k_12_3702), .fluid_out(k_11_1851), .air_in(c_12_0));
valve v_12_3703 (.fluid_in(k_12_3703), .fluid_out(k_11_1851), .air_in(c_12_1));
valve v_12_3704 (.fluid_in(k_12_3704), .fluid_out(k_11_1852), .air_in(c_12_0));
valve v_12_3705 (.fluid_in(k_12_3705), .fluid_out(k_11_1852), .air_in(c_12_1));
valve v_12_3706 (.fluid_in(k_12_3706), .fluid_out(k_11_1853), .air_in(c_12_0));
valve v_12_3707 (.fluid_in(k_12_3707), .fluid_out(k_11_1853), .air_in(c_12_1));
valve v_12_3708 (.fluid_in(k_12_3708), .fluid_out(k_11_1854), .air_in(c_12_0));
valve v_12_3709 (.fluid_in(k_12_3709), .fluid_out(k_11_1854), .air_in(c_12_1));
valve v_12_3710 (.fluid_in(k_12_3710), .fluid_out(k_11_1855), .air_in(c_12_0));
valve v_12_3711 (.fluid_in(k_12_3711), .fluid_out(k_11_1855), .air_in(c_12_1));
valve v_12_3712 (.fluid_in(k_12_3712), .fluid_out(k_11_1856), .air_in(c_12_0));
valve v_12_3713 (.fluid_in(k_12_3713), .fluid_out(k_11_1856), .air_in(c_12_1));
valve v_12_3714 (.fluid_in(k_12_3714), .fluid_out(k_11_1857), .air_in(c_12_0));
valve v_12_3715 (.fluid_in(k_12_3715), .fluid_out(k_11_1857), .air_in(c_12_1));
valve v_12_3716 (.fluid_in(k_12_3716), .fluid_out(k_11_1858), .air_in(c_12_0));
valve v_12_3717 (.fluid_in(k_12_3717), .fluid_out(k_11_1858), .air_in(c_12_1));
valve v_12_3718 (.fluid_in(k_12_3718), .fluid_out(k_11_1859), .air_in(c_12_0));
valve v_12_3719 (.fluid_in(k_12_3719), .fluid_out(k_11_1859), .air_in(c_12_1));
valve v_12_3720 (.fluid_in(k_12_3720), .fluid_out(k_11_1860), .air_in(c_12_0));
valve v_12_3721 (.fluid_in(k_12_3721), .fluid_out(k_11_1860), .air_in(c_12_1));
valve v_12_3722 (.fluid_in(k_12_3722), .fluid_out(k_11_1861), .air_in(c_12_0));
valve v_12_3723 (.fluid_in(k_12_3723), .fluid_out(k_11_1861), .air_in(c_12_1));
valve v_12_3724 (.fluid_in(k_12_3724), .fluid_out(k_11_1862), .air_in(c_12_0));
valve v_12_3725 (.fluid_in(k_12_3725), .fluid_out(k_11_1862), .air_in(c_12_1));
valve v_12_3726 (.fluid_in(k_12_3726), .fluid_out(k_11_1863), .air_in(c_12_0));
valve v_12_3727 (.fluid_in(k_12_3727), .fluid_out(k_11_1863), .air_in(c_12_1));
valve v_12_3728 (.fluid_in(k_12_3728), .fluid_out(k_11_1864), .air_in(c_12_0));
valve v_12_3729 (.fluid_in(k_12_3729), .fluid_out(k_11_1864), .air_in(c_12_1));
valve v_12_3730 (.fluid_in(k_12_3730), .fluid_out(k_11_1865), .air_in(c_12_0));
valve v_12_3731 (.fluid_in(k_12_3731), .fluid_out(k_11_1865), .air_in(c_12_1));
valve v_12_3732 (.fluid_in(k_12_3732), .fluid_out(k_11_1866), .air_in(c_12_0));
valve v_12_3733 (.fluid_in(k_12_3733), .fluid_out(k_11_1866), .air_in(c_12_1));
valve v_12_3734 (.fluid_in(k_12_3734), .fluid_out(k_11_1867), .air_in(c_12_0));
valve v_12_3735 (.fluid_in(k_12_3735), .fluid_out(k_11_1867), .air_in(c_12_1));
valve v_12_3736 (.fluid_in(k_12_3736), .fluid_out(k_11_1868), .air_in(c_12_0));
valve v_12_3737 (.fluid_in(k_12_3737), .fluid_out(k_11_1868), .air_in(c_12_1));
valve v_12_3738 (.fluid_in(k_12_3738), .fluid_out(k_11_1869), .air_in(c_12_0));
valve v_12_3739 (.fluid_in(k_12_3739), .fluid_out(k_11_1869), .air_in(c_12_1));
valve v_12_3740 (.fluid_in(k_12_3740), .fluid_out(k_11_1870), .air_in(c_12_0));
valve v_12_3741 (.fluid_in(k_12_3741), .fluid_out(k_11_1870), .air_in(c_12_1));
valve v_12_3742 (.fluid_in(k_12_3742), .fluid_out(k_11_1871), .air_in(c_12_0));
valve v_12_3743 (.fluid_in(k_12_3743), .fluid_out(k_11_1871), .air_in(c_12_1));
valve v_12_3744 (.fluid_in(k_12_3744), .fluid_out(k_11_1872), .air_in(c_12_0));
valve v_12_3745 (.fluid_in(k_12_3745), .fluid_out(k_11_1872), .air_in(c_12_1));
valve v_12_3746 (.fluid_in(k_12_3746), .fluid_out(k_11_1873), .air_in(c_12_0));
valve v_12_3747 (.fluid_in(k_12_3747), .fluid_out(k_11_1873), .air_in(c_12_1));
valve v_12_3748 (.fluid_in(k_12_3748), .fluid_out(k_11_1874), .air_in(c_12_0));
valve v_12_3749 (.fluid_in(k_12_3749), .fluid_out(k_11_1874), .air_in(c_12_1));
valve v_12_3750 (.fluid_in(k_12_3750), .fluid_out(k_11_1875), .air_in(c_12_0));
valve v_12_3751 (.fluid_in(k_12_3751), .fluid_out(k_11_1875), .air_in(c_12_1));
valve v_12_3752 (.fluid_in(k_12_3752), .fluid_out(k_11_1876), .air_in(c_12_0));
valve v_12_3753 (.fluid_in(k_12_3753), .fluid_out(k_11_1876), .air_in(c_12_1));
valve v_12_3754 (.fluid_in(k_12_3754), .fluid_out(k_11_1877), .air_in(c_12_0));
valve v_12_3755 (.fluid_in(k_12_3755), .fluid_out(k_11_1877), .air_in(c_12_1));
valve v_12_3756 (.fluid_in(k_12_3756), .fluid_out(k_11_1878), .air_in(c_12_0));
valve v_12_3757 (.fluid_in(k_12_3757), .fluid_out(k_11_1878), .air_in(c_12_1));
valve v_12_3758 (.fluid_in(k_12_3758), .fluid_out(k_11_1879), .air_in(c_12_0));
valve v_12_3759 (.fluid_in(k_12_3759), .fluid_out(k_11_1879), .air_in(c_12_1));
valve v_12_3760 (.fluid_in(k_12_3760), .fluid_out(k_11_1880), .air_in(c_12_0));
valve v_12_3761 (.fluid_in(k_12_3761), .fluid_out(k_11_1880), .air_in(c_12_1));
valve v_12_3762 (.fluid_in(k_12_3762), .fluid_out(k_11_1881), .air_in(c_12_0));
valve v_12_3763 (.fluid_in(k_12_3763), .fluid_out(k_11_1881), .air_in(c_12_1));
valve v_12_3764 (.fluid_in(k_12_3764), .fluid_out(k_11_1882), .air_in(c_12_0));
valve v_12_3765 (.fluid_in(k_12_3765), .fluid_out(k_11_1882), .air_in(c_12_1));
valve v_12_3766 (.fluid_in(k_12_3766), .fluid_out(k_11_1883), .air_in(c_12_0));
valve v_12_3767 (.fluid_in(k_12_3767), .fluid_out(k_11_1883), .air_in(c_12_1));
valve v_12_3768 (.fluid_in(k_12_3768), .fluid_out(k_11_1884), .air_in(c_12_0));
valve v_12_3769 (.fluid_in(k_12_3769), .fluid_out(k_11_1884), .air_in(c_12_1));
valve v_12_3770 (.fluid_in(k_12_3770), .fluid_out(k_11_1885), .air_in(c_12_0));
valve v_12_3771 (.fluid_in(k_12_3771), .fluid_out(k_11_1885), .air_in(c_12_1));
valve v_12_3772 (.fluid_in(k_12_3772), .fluid_out(k_11_1886), .air_in(c_12_0));
valve v_12_3773 (.fluid_in(k_12_3773), .fluid_out(k_11_1886), .air_in(c_12_1));
valve v_12_3774 (.fluid_in(k_12_3774), .fluid_out(k_11_1887), .air_in(c_12_0));
valve v_12_3775 (.fluid_in(k_12_3775), .fluid_out(k_11_1887), .air_in(c_12_1));
valve v_12_3776 (.fluid_in(k_12_3776), .fluid_out(k_11_1888), .air_in(c_12_0));
valve v_12_3777 (.fluid_in(k_12_3777), .fluid_out(k_11_1888), .air_in(c_12_1));
valve v_12_3778 (.fluid_in(k_12_3778), .fluid_out(k_11_1889), .air_in(c_12_0));
valve v_12_3779 (.fluid_in(k_12_3779), .fluid_out(k_11_1889), .air_in(c_12_1));
valve v_12_3780 (.fluid_in(k_12_3780), .fluid_out(k_11_1890), .air_in(c_12_0));
valve v_12_3781 (.fluid_in(k_12_3781), .fluid_out(k_11_1890), .air_in(c_12_1));
valve v_12_3782 (.fluid_in(k_12_3782), .fluid_out(k_11_1891), .air_in(c_12_0));
valve v_12_3783 (.fluid_in(k_12_3783), .fluid_out(k_11_1891), .air_in(c_12_1));
valve v_12_3784 (.fluid_in(k_12_3784), .fluid_out(k_11_1892), .air_in(c_12_0));
valve v_12_3785 (.fluid_in(k_12_3785), .fluid_out(k_11_1892), .air_in(c_12_1));
valve v_12_3786 (.fluid_in(k_12_3786), .fluid_out(k_11_1893), .air_in(c_12_0));
valve v_12_3787 (.fluid_in(k_12_3787), .fluid_out(k_11_1893), .air_in(c_12_1));
valve v_12_3788 (.fluid_in(k_12_3788), .fluid_out(k_11_1894), .air_in(c_12_0));
valve v_12_3789 (.fluid_in(k_12_3789), .fluid_out(k_11_1894), .air_in(c_12_1));
valve v_12_3790 (.fluid_in(k_12_3790), .fluid_out(k_11_1895), .air_in(c_12_0));
valve v_12_3791 (.fluid_in(k_12_3791), .fluid_out(k_11_1895), .air_in(c_12_1));
valve v_12_3792 (.fluid_in(k_12_3792), .fluid_out(k_11_1896), .air_in(c_12_0));
valve v_12_3793 (.fluid_in(k_12_3793), .fluid_out(k_11_1896), .air_in(c_12_1));
valve v_12_3794 (.fluid_in(k_12_3794), .fluid_out(k_11_1897), .air_in(c_12_0));
valve v_12_3795 (.fluid_in(k_12_3795), .fluid_out(k_11_1897), .air_in(c_12_1));
valve v_12_3796 (.fluid_in(k_12_3796), .fluid_out(k_11_1898), .air_in(c_12_0));
valve v_12_3797 (.fluid_in(k_12_3797), .fluid_out(k_11_1898), .air_in(c_12_1));
valve v_12_3798 (.fluid_in(k_12_3798), .fluid_out(k_11_1899), .air_in(c_12_0));
valve v_12_3799 (.fluid_in(k_12_3799), .fluid_out(k_11_1899), .air_in(c_12_1));
valve v_12_3800 (.fluid_in(k_12_3800), .fluid_out(k_11_1900), .air_in(c_12_0));
valve v_12_3801 (.fluid_in(k_12_3801), .fluid_out(k_11_1900), .air_in(c_12_1));
valve v_12_3802 (.fluid_in(k_12_3802), .fluid_out(k_11_1901), .air_in(c_12_0));
valve v_12_3803 (.fluid_in(k_12_3803), .fluid_out(k_11_1901), .air_in(c_12_1));
valve v_12_3804 (.fluid_in(k_12_3804), .fluid_out(k_11_1902), .air_in(c_12_0));
valve v_12_3805 (.fluid_in(k_12_3805), .fluid_out(k_11_1902), .air_in(c_12_1));
valve v_12_3806 (.fluid_in(k_12_3806), .fluid_out(k_11_1903), .air_in(c_12_0));
valve v_12_3807 (.fluid_in(k_12_3807), .fluid_out(k_11_1903), .air_in(c_12_1));
valve v_12_3808 (.fluid_in(k_12_3808), .fluid_out(k_11_1904), .air_in(c_12_0));
valve v_12_3809 (.fluid_in(k_12_3809), .fluid_out(k_11_1904), .air_in(c_12_1));
valve v_12_3810 (.fluid_in(k_12_3810), .fluid_out(k_11_1905), .air_in(c_12_0));
valve v_12_3811 (.fluid_in(k_12_3811), .fluid_out(k_11_1905), .air_in(c_12_1));
valve v_12_3812 (.fluid_in(k_12_3812), .fluid_out(k_11_1906), .air_in(c_12_0));
valve v_12_3813 (.fluid_in(k_12_3813), .fluid_out(k_11_1906), .air_in(c_12_1));
valve v_12_3814 (.fluid_in(k_12_3814), .fluid_out(k_11_1907), .air_in(c_12_0));
valve v_12_3815 (.fluid_in(k_12_3815), .fluid_out(k_11_1907), .air_in(c_12_1));
valve v_12_3816 (.fluid_in(k_12_3816), .fluid_out(k_11_1908), .air_in(c_12_0));
valve v_12_3817 (.fluid_in(k_12_3817), .fluid_out(k_11_1908), .air_in(c_12_1));
valve v_12_3818 (.fluid_in(k_12_3818), .fluid_out(k_11_1909), .air_in(c_12_0));
valve v_12_3819 (.fluid_in(k_12_3819), .fluid_out(k_11_1909), .air_in(c_12_1));
valve v_12_3820 (.fluid_in(k_12_3820), .fluid_out(k_11_1910), .air_in(c_12_0));
valve v_12_3821 (.fluid_in(k_12_3821), .fluid_out(k_11_1910), .air_in(c_12_1));
valve v_12_3822 (.fluid_in(k_12_3822), .fluid_out(k_11_1911), .air_in(c_12_0));
valve v_12_3823 (.fluid_in(k_12_3823), .fluid_out(k_11_1911), .air_in(c_12_1));
valve v_12_3824 (.fluid_in(k_12_3824), .fluid_out(k_11_1912), .air_in(c_12_0));
valve v_12_3825 (.fluid_in(k_12_3825), .fluid_out(k_11_1912), .air_in(c_12_1));
valve v_12_3826 (.fluid_in(k_12_3826), .fluid_out(k_11_1913), .air_in(c_12_0));
valve v_12_3827 (.fluid_in(k_12_3827), .fluid_out(k_11_1913), .air_in(c_12_1));
valve v_12_3828 (.fluid_in(k_12_3828), .fluid_out(k_11_1914), .air_in(c_12_0));
valve v_12_3829 (.fluid_in(k_12_3829), .fluid_out(k_11_1914), .air_in(c_12_1));
valve v_12_3830 (.fluid_in(k_12_3830), .fluid_out(k_11_1915), .air_in(c_12_0));
valve v_12_3831 (.fluid_in(k_12_3831), .fluid_out(k_11_1915), .air_in(c_12_1));
valve v_12_3832 (.fluid_in(k_12_3832), .fluid_out(k_11_1916), .air_in(c_12_0));
valve v_12_3833 (.fluid_in(k_12_3833), .fluid_out(k_11_1916), .air_in(c_12_1));
valve v_12_3834 (.fluid_in(k_12_3834), .fluid_out(k_11_1917), .air_in(c_12_0));
valve v_12_3835 (.fluid_in(k_12_3835), .fluid_out(k_11_1917), .air_in(c_12_1));
valve v_12_3836 (.fluid_in(k_12_3836), .fluid_out(k_11_1918), .air_in(c_12_0));
valve v_12_3837 (.fluid_in(k_12_3837), .fluid_out(k_11_1918), .air_in(c_12_1));
valve v_12_3838 (.fluid_in(k_12_3838), .fluid_out(k_11_1919), .air_in(c_12_0));
valve v_12_3839 (.fluid_in(k_12_3839), .fluid_out(k_11_1919), .air_in(c_12_1));
valve v_12_3840 (.fluid_in(k_12_3840), .fluid_out(k_11_1920), .air_in(c_12_0));
valve v_12_3841 (.fluid_in(k_12_3841), .fluid_out(k_11_1920), .air_in(c_12_1));
valve v_12_3842 (.fluid_in(k_12_3842), .fluid_out(k_11_1921), .air_in(c_12_0));
valve v_12_3843 (.fluid_in(k_12_3843), .fluid_out(k_11_1921), .air_in(c_12_1));
valve v_12_3844 (.fluid_in(k_12_3844), .fluid_out(k_11_1922), .air_in(c_12_0));
valve v_12_3845 (.fluid_in(k_12_3845), .fluid_out(k_11_1922), .air_in(c_12_1));
valve v_12_3846 (.fluid_in(k_12_3846), .fluid_out(k_11_1923), .air_in(c_12_0));
valve v_12_3847 (.fluid_in(k_12_3847), .fluid_out(k_11_1923), .air_in(c_12_1));
valve v_12_3848 (.fluid_in(k_12_3848), .fluid_out(k_11_1924), .air_in(c_12_0));
valve v_12_3849 (.fluid_in(k_12_3849), .fluid_out(k_11_1924), .air_in(c_12_1));
valve v_12_3850 (.fluid_in(k_12_3850), .fluid_out(k_11_1925), .air_in(c_12_0));
valve v_12_3851 (.fluid_in(k_12_3851), .fluid_out(k_11_1925), .air_in(c_12_1));
valve v_12_3852 (.fluid_in(k_12_3852), .fluid_out(k_11_1926), .air_in(c_12_0));
valve v_12_3853 (.fluid_in(k_12_3853), .fluid_out(k_11_1926), .air_in(c_12_1));
valve v_12_3854 (.fluid_in(k_12_3854), .fluid_out(k_11_1927), .air_in(c_12_0));
valve v_12_3855 (.fluid_in(k_12_3855), .fluid_out(k_11_1927), .air_in(c_12_1));
valve v_12_3856 (.fluid_in(k_12_3856), .fluid_out(k_11_1928), .air_in(c_12_0));
valve v_12_3857 (.fluid_in(k_12_3857), .fluid_out(k_11_1928), .air_in(c_12_1));
valve v_12_3858 (.fluid_in(k_12_3858), .fluid_out(k_11_1929), .air_in(c_12_0));
valve v_12_3859 (.fluid_in(k_12_3859), .fluid_out(k_11_1929), .air_in(c_12_1));
valve v_12_3860 (.fluid_in(k_12_3860), .fluid_out(k_11_1930), .air_in(c_12_0));
valve v_12_3861 (.fluid_in(k_12_3861), .fluid_out(k_11_1930), .air_in(c_12_1));
valve v_12_3862 (.fluid_in(k_12_3862), .fluid_out(k_11_1931), .air_in(c_12_0));
valve v_12_3863 (.fluid_in(k_12_3863), .fluid_out(k_11_1931), .air_in(c_12_1));
valve v_12_3864 (.fluid_in(k_12_3864), .fluid_out(k_11_1932), .air_in(c_12_0));
valve v_12_3865 (.fluid_in(k_12_3865), .fluid_out(k_11_1932), .air_in(c_12_1));
valve v_12_3866 (.fluid_in(k_12_3866), .fluid_out(k_11_1933), .air_in(c_12_0));
valve v_12_3867 (.fluid_in(k_12_3867), .fluid_out(k_11_1933), .air_in(c_12_1));
valve v_12_3868 (.fluid_in(k_12_3868), .fluid_out(k_11_1934), .air_in(c_12_0));
valve v_12_3869 (.fluid_in(k_12_3869), .fluid_out(k_11_1934), .air_in(c_12_1));
valve v_12_3870 (.fluid_in(k_12_3870), .fluid_out(k_11_1935), .air_in(c_12_0));
valve v_12_3871 (.fluid_in(k_12_3871), .fluid_out(k_11_1935), .air_in(c_12_1));
valve v_12_3872 (.fluid_in(k_12_3872), .fluid_out(k_11_1936), .air_in(c_12_0));
valve v_12_3873 (.fluid_in(k_12_3873), .fluid_out(k_11_1936), .air_in(c_12_1));
valve v_12_3874 (.fluid_in(k_12_3874), .fluid_out(k_11_1937), .air_in(c_12_0));
valve v_12_3875 (.fluid_in(k_12_3875), .fluid_out(k_11_1937), .air_in(c_12_1));
valve v_12_3876 (.fluid_in(k_12_3876), .fluid_out(k_11_1938), .air_in(c_12_0));
valve v_12_3877 (.fluid_in(k_12_3877), .fluid_out(k_11_1938), .air_in(c_12_1));
valve v_12_3878 (.fluid_in(k_12_3878), .fluid_out(k_11_1939), .air_in(c_12_0));
valve v_12_3879 (.fluid_in(k_12_3879), .fluid_out(k_11_1939), .air_in(c_12_1));
valve v_12_3880 (.fluid_in(k_12_3880), .fluid_out(k_11_1940), .air_in(c_12_0));
valve v_12_3881 (.fluid_in(k_12_3881), .fluid_out(k_11_1940), .air_in(c_12_1));
valve v_12_3882 (.fluid_in(k_12_3882), .fluid_out(k_11_1941), .air_in(c_12_0));
valve v_12_3883 (.fluid_in(k_12_3883), .fluid_out(k_11_1941), .air_in(c_12_1));
valve v_12_3884 (.fluid_in(k_12_3884), .fluid_out(k_11_1942), .air_in(c_12_0));
valve v_12_3885 (.fluid_in(k_12_3885), .fluid_out(k_11_1942), .air_in(c_12_1));
valve v_12_3886 (.fluid_in(k_12_3886), .fluid_out(k_11_1943), .air_in(c_12_0));
valve v_12_3887 (.fluid_in(k_12_3887), .fluid_out(k_11_1943), .air_in(c_12_1));
valve v_12_3888 (.fluid_in(k_12_3888), .fluid_out(k_11_1944), .air_in(c_12_0));
valve v_12_3889 (.fluid_in(k_12_3889), .fluid_out(k_11_1944), .air_in(c_12_1));
valve v_12_3890 (.fluid_in(k_12_3890), .fluid_out(k_11_1945), .air_in(c_12_0));
valve v_12_3891 (.fluid_in(k_12_3891), .fluid_out(k_11_1945), .air_in(c_12_1));
valve v_12_3892 (.fluid_in(k_12_3892), .fluid_out(k_11_1946), .air_in(c_12_0));
valve v_12_3893 (.fluid_in(k_12_3893), .fluid_out(k_11_1946), .air_in(c_12_1));
valve v_12_3894 (.fluid_in(k_12_3894), .fluid_out(k_11_1947), .air_in(c_12_0));
valve v_12_3895 (.fluid_in(k_12_3895), .fluid_out(k_11_1947), .air_in(c_12_1));
valve v_12_3896 (.fluid_in(k_12_3896), .fluid_out(k_11_1948), .air_in(c_12_0));
valve v_12_3897 (.fluid_in(k_12_3897), .fluid_out(k_11_1948), .air_in(c_12_1));
valve v_12_3898 (.fluid_in(k_12_3898), .fluid_out(k_11_1949), .air_in(c_12_0));
valve v_12_3899 (.fluid_in(k_12_3899), .fluid_out(k_11_1949), .air_in(c_12_1));
valve v_12_3900 (.fluid_in(k_12_3900), .fluid_out(k_11_1950), .air_in(c_12_0));
valve v_12_3901 (.fluid_in(k_12_3901), .fluid_out(k_11_1950), .air_in(c_12_1));
valve v_12_3902 (.fluid_in(k_12_3902), .fluid_out(k_11_1951), .air_in(c_12_0));
valve v_12_3903 (.fluid_in(k_12_3903), .fluid_out(k_11_1951), .air_in(c_12_1));
valve v_12_3904 (.fluid_in(k_12_3904), .fluid_out(k_11_1952), .air_in(c_12_0));
valve v_12_3905 (.fluid_in(k_12_3905), .fluid_out(k_11_1952), .air_in(c_12_1));
valve v_12_3906 (.fluid_in(k_12_3906), .fluid_out(k_11_1953), .air_in(c_12_0));
valve v_12_3907 (.fluid_in(k_12_3907), .fluid_out(k_11_1953), .air_in(c_12_1));
valve v_12_3908 (.fluid_in(k_12_3908), .fluid_out(k_11_1954), .air_in(c_12_0));
valve v_12_3909 (.fluid_in(k_12_3909), .fluid_out(k_11_1954), .air_in(c_12_1));
valve v_12_3910 (.fluid_in(k_12_3910), .fluid_out(k_11_1955), .air_in(c_12_0));
valve v_12_3911 (.fluid_in(k_12_3911), .fluid_out(k_11_1955), .air_in(c_12_1));
valve v_12_3912 (.fluid_in(k_12_3912), .fluid_out(k_11_1956), .air_in(c_12_0));
valve v_12_3913 (.fluid_in(k_12_3913), .fluid_out(k_11_1956), .air_in(c_12_1));
valve v_12_3914 (.fluid_in(k_12_3914), .fluid_out(k_11_1957), .air_in(c_12_0));
valve v_12_3915 (.fluid_in(k_12_3915), .fluid_out(k_11_1957), .air_in(c_12_1));
valve v_12_3916 (.fluid_in(k_12_3916), .fluid_out(k_11_1958), .air_in(c_12_0));
valve v_12_3917 (.fluid_in(k_12_3917), .fluid_out(k_11_1958), .air_in(c_12_1));
valve v_12_3918 (.fluid_in(k_12_3918), .fluid_out(k_11_1959), .air_in(c_12_0));
valve v_12_3919 (.fluid_in(k_12_3919), .fluid_out(k_11_1959), .air_in(c_12_1));
valve v_12_3920 (.fluid_in(k_12_3920), .fluid_out(k_11_1960), .air_in(c_12_0));
valve v_12_3921 (.fluid_in(k_12_3921), .fluid_out(k_11_1960), .air_in(c_12_1));
valve v_12_3922 (.fluid_in(k_12_3922), .fluid_out(k_11_1961), .air_in(c_12_0));
valve v_12_3923 (.fluid_in(k_12_3923), .fluid_out(k_11_1961), .air_in(c_12_1));
valve v_12_3924 (.fluid_in(k_12_3924), .fluid_out(k_11_1962), .air_in(c_12_0));
valve v_12_3925 (.fluid_in(k_12_3925), .fluid_out(k_11_1962), .air_in(c_12_1));
valve v_12_3926 (.fluid_in(k_12_3926), .fluid_out(k_11_1963), .air_in(c_12_0));
valve v_12_3927 (.fluid_in(k_12_3927), .fluid_out(k_11_1963), .air_in(c_12_1));
valve v_12_3928 (.fluid_in(k_12_3928), .fluid_out(k_11_1964), .air_in(c_12_0));
valve v_12_3929 (.fluid_in(k_12_3929), .fluid_out(k_11_1964), .air_in(c_12_1));
valve v_12_3930 (.fluid_in(k_12_3930), .fluid_out(k_11_1965), .air_in(c_12_0));
valve v_12_3931 (.fluid_in(k_12_3931), .fluid_out(k_11_1965), .air_in(c_12_1));
valve v_12_3932 (.fluid_in(k_12_3932), .fluid_out(k_11_1966), .air_in(c_12_0));
valve v_12_3933 (.fluid_in(k_12_3933), .fluid_out(k_11_1966), .air_in(c_12_1));
valve v_12_3934 (.fluid_in(k_12_3934), .fluid_out(k_11_1967), .air_in(c_12_0));
valve v_12_3935 (.fluid_in(k_12_3935), .fluid_out(k_11_1967), .air_in(c_12_1));
valve v_12_3936 (.fluid_in(k_12_3936), .fluid_out(k_11_1968), .air_in(c_12_0));
valve v_12_3937 (.fluid_in(k_12_3937), .fluid_out(k_11_1968), .air_in(c_12_1));
valve v_12_3938 (.fluid_in(k_12_3938), .fluid_out(k_11_1969), .air_in(c_12_0));
valve v_12_3939 (.fluid_in(k_12_3939), .fluid_out(k_11_1969), .air_in(c_12_1));
valve v_12_3940 (.fluid_in(k_12_3940), .fluid_out(k_11_1970), .air_in(c_12_0));
valve v_12_3941 (.fluid_in(k_12_3941), .fluid_out(k_11_1970), .air_in(c_12_1));
valve v_12_3942 (.fluid_in(k_12_3942), .fluid_out(k_11_1971), .air_in(c_12_0));
valve v_12_3943 (.fluid_in(k_12_3943), .fluid_out(k_11_1971), .air_in(c_12_1));
valve v_12_3944 (.fluid_in(k_12_3944), .fluid_out(k_11_1972), .air_in(c_12_0));
valve v_12_3945 (.fluid_in(k_12_3945), .fluid_out(k_11_1972), .air_in(c_12_1));
valve v_12_3946 (.fluid_in(k_12_3946), .fluid_out(k_11_1973), .air_in(c_12_0));
valve v_12_3947 (.fluid_in(k_12_3947), .fluid_out(k_11_1973), .air_in(c_12_1));
valve v_12_3948 (.fluid_in(k_12_3948), .fluid_out(k_11_1974), .air_in(c_12_0));
valve v_12_3949 (.fluid_in(k_12_3949), .fluid_out(k_11_1974), .air_in(c_12_1));
valve v_12_3950 (.fluid_in(k_12_3950), .fluid_out(k_11_1975), .air_in(c_12_0));
valve v_12_3951 (.fluid_in(k_12_3951), .fluid_out(k_11_1975), .air_in(c_12_1));
valve v_12_3952 (.fluid_in(k_12_3952), .fluid_out(k_11_1976), .air_in(c_12_0));
valve v_12_3953 (.fluid_in(k_12_3953), .fluid_out(k_11_1976), .air_in(c_12_1));
valve v_12_3954 (.fluid_in(k_12_3954), .fluid_out(k_11_1977), .air_in(c_12_0));
valve v_12_3955 (.fluid_in(k_12_3955), .fluid_out(k_11_1977), .air_in(c_12_1));
valve v_12_3956 (.fluid_in(k_12_3956), .fluid_out(k_11_1978), .air_in(c_12_0));
valve v_12_3957 (.fluid_in(k_12_3957), .fluid_out(k_11_1978), .air_in(c_12_1));
valve v_12_3958 (.fluid_in(k_12_3958), .fluid_out(k_11_1979), .air_in(c_12_0));
valve v_12_3959 (.fluid_in(k_12_3959), .fluid_out(k_11_1979), .air_in(c_12_1));
valve v_12_3960 (.fluid_in(k_12_3960), .fluid_out(k_11_1980), .air_in(c_12_0));
valve v_12_3961 (.fluid_in(k_12_3961), .fluid_out(k_11_1980), .air_in(c_12_1));
valve v_12_3962 (.fluid_in(k_12_3962), .fluid_out(k_11_1981), .air_in(c_12_0));
valve v_12_3963 (.fluid_in(k_12_3963), .fluid_out(k_11_1981), .air_in(c_12_1));
valve v_12_3964 (.fluid_in(k_12_3964), .fluid_out(k_11_1982), .air_in(c_12_0));
valve v_12_3965 (.fluid_in(k_12_3965), .fluid_out(k_11_1982), .air_in(c_12_1));
valve v_12_3966 (.fluid_in(k_12_3966), .fluid_out(k_11_1983), .air_in(c_12_0));
valve v_12_3967 (.fluid_in(k_12_3967), .fluid_out(k_11_1983), .air_in(c_12_1));
valve v_12_3968 (.fluid_in(k_12_3968), .fluid_out(k_11_1984), .air_in(c_12_0));
valve v_12_3969 (.fluid_in(k_12_3969), .fluid_out(k_11_1984), .air_in(c_12_1));
valve v_12_3970 (.fluid_in(k_12_3970), .fluid_out(k_11_1985), .air_in(c_12_0));
valve v_12_3971 (.fluid_in(k_12_3971), .fluid_out(k_11_1985), .air_in(c_12_1));
valve v_12_3972 (.fluid_in(k_12_3972), .fluid_out(k_11_1986), .air_in(c_12_0));
valve v_12_3973 (.fluid_in(k_12_3973), .fluid_out(k_11_1986), .air_in(c_12_1));
valve v_12_3974 (.fluid_in(k_12_3974), .fluid_out(k_11_1987), .air_in(c_12_0));
valve v_12_3975 (.fluid_in(k_12_3975), .fluid_out(k_11_1987), .air_in(c_12_1));
valve v_12_3976 (.fluid_in(k_12_3976), .fluid_out(k_11_1988), .air_in(c_12_0));
valve v_12_3977 (.fluid_in(k_12_3977), .fluid_out(k_11_1988), .air_in(c_12_1));
valve v_12_3978 (.fluid_in(k_12_3978), .fluid_out(k_11_1989), .air_in(c_12_0));
valve v_12_3979 (.fluid_in(k_12_3979), .fluid_out(k_11_1989), .air_in(c_12_1));
valve v_12_3980 (.fluid_in(k_12_3980), .fluid_out(k_11_1990), .air_in(c_12_0));
valve v_12_3981 (.fluid_in(k_12_3981), .fluid_out(k_11_1990), .air_in(c_12_1));
valve v_12_3982 (.fluid_in(k_12_3982), .fluid_out(k_11_1991), .air_in(c_12_0));
valve v_12_3983 (.fluid_in(k_12_3983), .fluid_out(k_11_1991), .air_in(c_12_1));
valve v_12_3984 (.fluid_in(k_12_3984), .fluid_out(k_11_1992), .air_in(c_12_0));
valve v_12_3985 (.fluid_in(k_12_3985), .fluid_out(k_11_1992), .air_in(c_12_1));
valve v_12_3986 (.fluid_in(k_12_3986), .fluid_out(k_11_1993), .air_in(c_12_0));
valve v_12_3987 (.fluid_in(k_12_3987), .fluid_out(k_11_1993), .air_in(c_12_1));
valve v_12_3988 (.fluid_in(k_12_3988), .fluid_out(k_11_1994), .air_in(c_12_0));
valve v_12_3989 (.fluid_in(k_12_3989), .fluid_out(k_11_1994), .air_in(c_12_1));
valve v_12_3990 (.fluid_in(k_12_3990), .fluid_out(k_11_1995), .air_in(c_12_0));
valve v_12_3991 (.fluid_in(k_12_3991), .fluid_out(k_11_1995), .air_in(c_12_1));
valve v_12_3992 (.fluid_in(k_12_3992), .fluid_out(k_11_1996), .air_in(c_12_0));
valve v_12_3993 (.fluid_in(k_12_3993), .fluid_out(k_11_1996), .air_in(c_12_1));
valve v_12_3994 (.fluid_in(k_12_3994), .fluid_out(k_11_1997), .air_in(c_12_0));
valve v_12_3995 (.fluid_in(k_12_3995), .fluid_out(k_11_1997), .air_in(c_12_1));
valve v_12_3996 (.fluid_in(k_12_3996), .fluid_out(k_11_1998), .air_in(c_12_0));
valve v_12_3997 (.fluid_in(k_12_3997), .fluid_out(k_11_1998), .air_in(c_12_1));
valve v_12_3998 (.fluid_in(k_12_3998), .fluid_out(k_11_1999), .air_in(c_12_0));
valve v_12_3999 (.fluid_in(k_12_3999), .fluid_out(k_11_1999), .air_in(c_12_1));
valve v_12_4000 (.fluid_in(k_12_4000), .fluid_out(k_11_2000), .air_in(c_12_0));
valve v_12_4001 (.fluid_in(k_12_4001), .fluid_out(k_11_2000), .air_in(c_12_1));
valve v_12_4002 (.fluid_in(k_12_4002), .fluid_out(k_11_2001), .air_in(c_12_0));
valve v_12_4003 (.fluid_in(k_12_4003), .fluid_out(k_11_2001), .air_in(c_12_1));
valve v_12_4004 (.fluid_in(k_12_4004), .fluid_out(k_11_2002), .air_in(c_12_0));
valve v_12_4005 (.fluid_in(k_12_4005), .fluid_out(k_11_2002), .air_in(c_12_1));
valve v_12_4006 (.fluid_in(k_12_4006), .fluid_out(k_11_2003), .air_in(c_12_0));
valve v_12_4007 (.fluid_in(k_12_4007), .fluid_out(k_11_2003), .air_in(c_12_1));
valve v_12_4008 (.fluid_in(k_12_4008), .fluid_out(k_11_2004), .air_in(c_12_0));
valve v_12_4009 (.fluid_in(k_12_4009), .fluid_out(k_11_2004), .air_in(c_12_1));
valve v_12_4010 (.fluid_in(k_12_4010), .fluid_out(k_11_2005), .air_in(c_12_0));
valve v_12_4011 (.fluid_in(k_12_4011), .fluid_out(k_11_2005), .air_in(c_12_1));
valve v_12_4012 (.fluid_in(k_12_4012), .fluid_out(k_11_2006), .air_in(c_12_0));
valve v_12_4013 (.fluid_in(k_12_4013), .fluid_out(k_11_2006), .air_in(c_12_1));
valve v_12_4014 (.fluid_in(k_12_4014), .fluid_out(k_11_2007), .air_in(c_12_0));
valve v_12_4015 (.fluid_in(k_12_4015), .fluid_out(k_11_2007), .air_in(c_12_1));
valve v_12_4016 (.fluid_in(k_12_4016), .fluid_out(k_11_2008), .air_in(c_12_0));
valve v_12_4017 (.fluid_in(k_12_4017), .fluid_out(k_11_2008), .air_in(c_12_1));
valve v_12_4018 (.fluid_in(k_12_4018), .fluid_out(k_11_2009), .air_in(c_12_0));
valve v_12_4019 (.fluid_in(k_12_4019), .fluid_out(k_11_2009), .air_in(c_12_1));
valve v_12_4020 (.fluid_in(k_12_4020), .fluid_out(k_11_2010), .air_in(c_12_0));
valve v_12_4021 (.fluid_in(k_12_4021), .fluid_out(k_11_2010), .air_in(c_12_1));
valve v_12_4022 (.fluid_in(k_12_4022), .fluid_out(k_11_2011), .air_in(c_12_0));
valve v_12_4023 (.fluid_in(k_12_4023), .fluid_out(k_11_2011), .air_in(c_12_1));
valve v_12_4024 (.fluid_in(k_12_4024), .fluid_out(k_11_2012), .air_in(c_12_0));
valve v_12_4025 (.fluid_in(k_12_4025), .fluid_out(k_11_2012), .air_in(c_12_1));
valve v_12_4026 (.fluid_in(k_12_4026), .fluid_out(k_11_2013), .air_in(c_12_0));
valve v_12_4027 (.fluid_in(k_12_4027), .fluid_out(k_11_2013), .air_in(c_12_1));
valve v_12_4028 (.fluid_in(k_12_4028), .fluid_out(k_11_2014), .air_in(c_12_0));
valve v_12_4029 (.fluid_in(k_12_4029), .fluid_out(k_11_2014), .air_in(c_12_1));
valve v_12_4030 (.fluid_in(k_12_4030), .fluid_out(k_11_2015), .air_in(c_12_0));
valve v_12_4031 (.fluid_in(k_12_4031), .fluid_out(k_11_2015), .air_in(c_12_1));
valve v_12_4032 (.fluid_in(k_12_4032), .fluid_out(k_11_2016), .air_in(c_12_0));
valve v_12_4033 (.fluid_in(k_12_4033), .fluid_out(k_11_2016), .air_in(c_12_1));
valve v_12_4034 (.fluid_in(k_12_4034), .fluid_out(k_11_2017), .air_in(c_12_0));
valve v_12_4035 (.fluid_in(k_12_4035), .fluid_out(k_11_2017), .air_in(c_12_1));
valve v_12_4036 (.fluid_in(k_12_4036), .fluid_out(k_11_2018), .air_in(c_12_0));
valve v_12_4037 (.fluid_in(k_12_4037), .fluid_out(k_11_2018), .air_in(c_12_1));
valve v_12_4038 (.fluid_in(k_12_4038), .fluid_out(k_11_2019), .air_in(c_12_0));
valve v_12_4039 (.fluid_in(k_12_4039), .fluid_out(k_11_2019), .air_in(c_12_1));
valve v_12_4040 (.fluid_in(k_12_4040), .fluid_out(k_11_2020), .air_in(c_12_0));
valve v_12_4041 (.fluid_in(k_12_4041), .fluid_out(k_11_2020), .air_in(c_12_1));
valve v_12_4042 (.fluid_in(k_12_4042), .fluid_out(k_11_2021), .air_in(c_12_0));
valve v_12_4043 (.fluid_in(k_12_4043), .fluid_out(k_11_2021), .air_in(c_12_1));
valve v_12_4044 (.fluid_in(k_12_4044), .fluid_out(k_11_2022), .air_in(c_12_0));
valve v_12_4045 (.fluid_in(k_12_4045), .fluid_out(k_11_2022), .air_in(c_12_1));
valve v_12_4046 (.fluid_in(k_12_4046), .fluid_out(k_11_2023), .air_in(c_12_0));
valve v_12_4047 (.fluid_in(k_12_4047), .fluid_out(k_11_2023), .air_in(c_12_1));
valve v_12_4048 (.fluid_in(k_12_4048), .fluid_out(k_11_2024), .air_in(c_12_0));
valve v_12_4049 (.fluid_in(k_12_4049), .fluid_out(k_11_2024), .air_in(c_12_1));
valve v_12_4050 (.fluid_in(k_12_4050), .fluid_out(k_11_2025), .air_in(c_12_0));
valve v_12_4051 (.fluid_in(k_12_4051), .fluid_out(k_11_2025), .air_in(c_12_1));
valve v_12_4052 (.fluid_in(k_12_4052), .fluid_out(k_11_2026), .air_in(c_12_0));
valve v_12_4053 (.fluid_in(k_12_4053), .fluid_out(k_11_2026), .air_in(c_12_1));
valve v_12_4054 (.fluid_in(k_12_4054), .fluid_out(k_11_2027), .air_in(c_12_0));
valve v_12_4055 (.fluid_in(k_12_4055), .fluid_out(k_11_2027), .air_in(c_12_1));
valve v_12_4056 (.fluid_in(k_12_4056), .fluid_out(k_11_2028), .air_in(c_12_0));
valve v_12_4057 (.fluid_in(k_12_4057), .fluid_out(k_11_2028), .air_in(c_12_1));
valve v_12_4058 (.fluid_in(k_12_4058), .fluid_out(k_11_2029), .air_in(c_12_0));
valve v_12_4059 (.fluid_in(k_12_4059), .fluid_out(k_11_2029), .air_in(c_12_1));
valve v_12_4060 (.fluid_in(k_12_4060), .fluid_out(k_11_2030), .air_in(c_12_0));
valve v_12_4061 (.fluid_in(k_12_4061), .fluid_out(k_11_2030), .air_in(c_12_1));
valve v_12_4062 (.fluid_in(k_12_4062), .fluid_out(k_11_2031), .air_in(c_12_0));
valve v_12_4063 (.fluid_in(k_12_4063), .fluid_out(k_11_2031), .air_in(c_12_1));
valve v_12_4064 (.fluid_in(k_12_4064), .fluid_out(k_11_2032), .air_in(c_12_0));
valve v_12_4065 (.fluid_in(k_12_4065), .fluid_out(k_11_2032), .air_in(c_12_1));
valve v_12_4066 (.fluid_in(k_12_4066), .fluid_out(k_11_2033), .air_in(c_12_0));
valve v_12_4067 (.fluid_in(k_12_4067), .fluid_out(k_11_2033), .air_in(c_12_1));
valve v_12_4068 (.fluid_in(k_12_4068), .fluid_out(k_11_2034), .air_in(c_12_0));
valve v_12_4069 (.fluid_in(k_12_4069), .fluid_out(k_11_2034), .air_in(c_12_1));
valve v_12_4070 (.fluid_in(k_12_4070), .fluid_out(k_11_2035), .air_in(c_12_0));
valve v_12_4071 (.fluid_in(k_12_4071), .fluid_out(k_11_2035), .air_in(c_12_1));
valve v_12_4072 (.fluid_in(k_12_4072), .fluid_out(k_11_2036), .air_in(c_12_0));
valve v_12_4073 (.fluid_in(k_12_4073), .fluid_out(k_11_2036), .air_in(c_12_1));
valve v_12_4074 (.fluid_in(k_12_4074), .fluid_out(k_11_2037), .air_in(c_12_0));
valve v_12_4075 (.fluid_in(k_12_4075), .fluid_out(k_11_2037), .air_in(c_12_1));
valve v_12_4076 (.fluid_in(k_12_4076), .fluid_out(k_11_2038), .air_in(c_12_0));
valve v_12_4077 (.fluid_in(k_12_4077), .fluid_out(k_11_2038), .air_in(c_12_1));
valve v_12_4078 (.fluid_in(k_12_4078), .fluid_out(k_11_2039), .air_in(c_12_0));
valve v_12_4079 (.fluid_in(k_12_4079), .fluid_out(k_11_2039), .air_in(c_12_1));
valve v_12_4080 (.fluid_in(k_12_4080), .fluid_out(k_11_2040), .air_in(c_12_0));
valve v_12_4081 (.fluid_in(k_12_4081), .fluid_out(k_11_2040), .air_in(c_12_1));
valve v_12_4082 (.fluid_in(k_12_4082), .fluid_out(k_11_2041), .air_in(c_12_0));
valve v_12_4083 (.fluid_in(k_12_4083), .fluid_out(k_11_2041), .air_in(c_12_1));
valve v_12_4084 (.fluid_in(k_12_4084), .fluid_out(k_11_2042), .air_in(c_12_0));
valve v_12_4085 (.fluid_in(k_12_4085), .fluid_out(k_11_2042), .air_in(c_12_1));
valve v_12_4086 (.fluid_in(k_12_4086), .fluid_out(k_11_2043), .air_in(c_12_0));
valve v_12_4087 (.fluid_in(k_12_4087), .fluid_out(k_11_2043), .air_in(c_12_1));
valve v_12_4088 (.fluid_in(k_12_4088), .fluid_out(k_11_2044), .air_in(c_12_0));
valve v_12_4089 (.fluid_in(k_12_4089), .fluid_out(k_11_2044), .air_in(c_12_1));
valve v_12_4090 (.fluid_in(k_12_4090), .fluid_out(k_11_2045), .air_in(c_12_0));
valve v_12_4091 (.fluid_in(k_12_4091), .fluid_out(k_11_2045), .air_in(c_12_1));
valve v_12_4092 (.fluid_in(k_12_4092), .fluid_out(k_11_2046), .air_in(c_12_0));
valve v_12_4093 (.fluid_in(k_12_4093), .fluid_out(k_11_2046), .air_in(c_12_1));
valve v_12_4094 (.fluid_in(k_12_4094), .fluid_out(k_11_2047), .air_in(c_12_0));
valve v_12_4095 (.fluid_in(k_12_4095), .fluid_out(k_11_2047), .air_in(c_12_1));
endmodule
