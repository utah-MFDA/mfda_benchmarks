module fanout2_braid_16_96 (
output output_0,output output_1,output output_2,output output_3,output output_4,output output_5,output output_6,output output_7,output output_8,output output_9,output output_10,output output_11,output output_12,output output_13,output output_14,output output_15,input input_0,input input_1,input input_2,input input_3,input input_4,input input_5,input input_6,input input_7,input input_8,input input_9,input input_10,input input_11,input input_12,input input_13,input input_14,input input_15
);
wire output_1_0, output_1_1, output_0_0;
mixer gate_output_0_0(.a(output_1_0), .b(output_1_1), .y(output_0_0));
wire output_2_0, output_2_1, output_1_0;
mixer gate_output_1_0(.a(output_2_0), .b(output_2_1), .y(output_1_0));
wire output_3_0, output_3_1, output_2_0;
mixer gate_output_2_0(.a(output_3_0), .b(output_3_1), .y(output_2_0));
wire output_4_0, output_4_1, output_3_0;
mixer gate_output_3_0(.a(output_4_0), .b(output_4_1), .y(output_3_0));
wire output_5_0, output_5_1, output_4_0;
mixer gate_output_4_0(.a(output_5_0), .b(output_5_1), .y(output_4_0));
wire output_6_0, output_6_1, output_5_0;
mixer gate_output_5_0(.a(output_6_0), .b(output_6_1), .y(output_5_0));
wire output_7_0, output_7_1, output_6_0;
mixer gate_output_6_0(.a(output_7_0), .b(output_7_1), .y(output_6_0));
wire output_8_0, output_8_1, output_7_0;
mixer gate_output_7_0(.a(output_8_0), .b(output_8_1), .y(output_7_0));
wire output_9_0, output_9_1, output_8_0;
mixer gate_output_8_0(.a(output_9_0), .b(output_9_1), .y(output_8_0));
wire output_10_0, output_10_1, output_9_0;
mixer gate_output_9_0(.a(output_10_0), .b(output_10_1), .y(output_9_0));
wire output_11_0, output_11_1, output_10_0;
mixer gate_output_10_0(.a(output_11_0), .b(output_11_1), .y(output_10_0));
wire output_12_0, output_12_1, output_11_0;
mixer gate_output_11_0(.a(output_12_0), .b(output_12_1), .y(output_11_0));
wire output_13_0, output_13_1, output_12_0;
mixer gate_output_12_0(.a(output_13_0), .b(output_13_1), .y(output_12_0));
wire output_14_0, output_14_1, output_13_0;
mixer gate_output_13_0(.a(output_14_0), .b(output_14_1), .y(output_13_0));
wire output_15_0, output_15_1, output_14_0;
mixer gate_output_14_0(.a(output_15_0), .b(output_15_1), .y(output_14_0));
wire output_16_0, output_16_1, output_15_0;
mixer gate_output_15_0(.a(output_16_0), .b(output_16_1), .y(output_15_0));
wire output_1_1, output_1_2, output_0_1;
mixer gate_output_0_1(.a(output_1_1), .b(output_1_2), .y(output_0_1));
wire output_2_1, output_2_2, output_1_1;
mixer gate_output_1_1(.a(output_2_1), .b(output_2_2), .y(output_1_1));
wire output_3_1, output_3_2, output_2_1;
mixer gate_output_2_1(.a(output_3_1), .b(output_3_2), .y(output_2_1));
wire output_4_1, output_4_2, output_3_1;
mixer gate_output_3_1(.a(output_4_1), .b(output_4_2), .y(output_3_1));
wire output_5_1, output_5_2, output_4_1;
mixer gate_output_4_1(.a(output_5_1), .b(output_5_2), .y(output_4_1));
wire output_6_1, output_6_2, output_5_1;
mixer gate_output_5_1(.a(output_6_1), .b(output_6_2), .y(output_5_1));
wire output_7_1, output_7_2, output_6_1;
mixer gate_output_6_1(.a(output_7_1), .b(output_7_2), .y(output_6_1));
wire output_8_1, output_8_2, output_7_1;
mixer gate_output_7_1(.a(output_8_1), .b(output_8_2), .y(output_7_1));
wire output_9_1, output_9_2, output_8_1;
mixer gate_output_8_1(.a(output_9_1), .b(output_9_2), .y(output_8_1));
wire output_10_1, output_10_2, output_9_1;
mixer gate_output_9_1(.a(output_10_1), .b(output_10_2), .y(output_9_1));
wire output_11_1, output_11_2, output_10_1;
mixer gate_output_10_1(.a(output_11_1), .b(output_11_2), .y(output_10_1));
wire output_12_1, output_12_2, output_11_1;
mixer gate_output_11_1(.a(output_12_1), .b(output_12_2), .y(output_11_1));
wire output_13_1, output_13_2, output_12_1;
mixer gate_output_12_1(.a(output_13_1), .b(output_13_2), .y(output_12_1));
wire output_14_1, output_14_2, output_13_1;
mixer gate_output_13_1(.a(output_14_1), .b(output_14_2), .y(output_13_1));
wire output_15_1, output_15_2, output_14_1;
mixer gate_output_14_1(.a(output_15_1), .b(output_15_2), .y(output_14_1));
wire output_16_1, output_16_2, output_15_1;
mixer gate_output_15_1(.a(output_16_1), .b(output_16_2), .y(output_15_1));
wire output_1_2, output_1_3, output_0_2;
mixer gate_output_0_2(.a(output_1_2), .b(output_1_3), .y(output_0_2));
wire output_2_2, output_2_3, output_1_2;
mixer gate_output_1_2(.a(output_2_2), .b(output_2_3), .y(output_1_2));
wire output_3_2, output_3_3, output_2_2;
mixer gate_output_2_2(.a(output_3_2), .b(output_3_3), .y(output_2_2));
wire output_4_2, output_4_3, output_3_2;
mixer gate_output_3_2(.a(output_4_2), .b(output_4_3), .y(output_3_2));
wire output_5_2, output_5_3, output_4_2;
mixer gate_output_4_2(.a(output_5_2), .b(output_5_3), .y(output_4_2));
wire output_6_2, output_6_3, output_5_2;
mixer gate_output_5_2(.a(output_6_2), .b(output_6_3), .y(output_5_2));
wire output_7_2, output_7_3, output_6_2;
mixer gate_output_6_2(.a(output_7_2), .b(output_7_3), .y(output_6_2));
wire output_8_2, output_8_3, output_7_2;
mixer gate_output_7_2(.a(output_8_2), .b(output_8_3), .y(output_7_2));
wire output_9_2, output_9_3, output_8_2;
mixer gate_output_8_2(.a(output_9_2), .b(output_9_3), .y(output_8_2));
wire output_10_2, output_10_3, output_9_2;
mixer gate_output_9_2(.a(output_10_2), .b(output_10_3), .y(output_9_2));
wire output_11_2, output_11_3, output_10_2;
mixer gate_output_10_2(.a(output_11_2), .b(output_11_3), .y(output_10_2));
wire output_12_2, output_12_3, output_11_2;
mixer gate_output_11_2(.a(output_12_2), .b(output_12_3), .y(output_11_2));
wire output_13_2, output_13_3, output_12_2;
mixer gate_output_12_2(.a(output_13_2), .b(output_13_3), .y(output_12_2));
wire output_14_2, output_14_3, output_13_2;
mixer gate_output_13_2(.a(output_14_2), .b(output_14_3), .y(output_13_2));
wire output_15_2, output_15_3, output_14_2;
mixer gate_output_14_2(.a(output_15_2), .b(output_15_3), .y(output_14_2));
wire output_16_2, output_16_3, output_15_2;
mixer gate_output_15_2(.a(output_16_2), .b(output_16_3), .y(output_15_2));
wire output_1_3, output_1_4, output_0_3;
mixer gate_output_0_3(.a(output_1_3), .b(output_1_4), .y(output_0_3));
wire output_2_3, output_2_4, output_1_3;
mixer gate_output_1_3(.a(output_2_3), .b(output_2_4), .y(output_1_3));
wire output_3_3, output_3_4, output_2_3;
mixer gate_output_2_3(.a(output_3_3), .b(output_3_4), .y(output_2_3));
wire output_4_3, output_4_4, output_3_3;
mixer gate_output_3_3(.a(output_4_3), .b(output_4_4), .y(output_3_3));
wire output_5_3, output_5_4, output_4_3;
mixer gate_output_4_3(.a(output_5_3), .b(output_5_4), .y(output_4_3));
wire output_6_3, output_6_4, output_5_3;
mixer gate_output_5_3(.a(output_6_3), .b(output_6_4), .y(output_5_3));
wire output_7_3, output_7_4, output_6_3;
mixer gate_output_6_3(.a(output_7_3), .b(output_7_4), .y(output_6_3));
wire output_8_3, output_8_4, output_7_3;
mixer gate_output_7_3(.a(output_8_3), .b(output_8_4), .y(output_7_3));
wire output_9_3, output_9_4, output_8_3;
mixer gate_output_8_3(.a(output_9_3), .b(output_9_4), .y(output_8_3));
wire output_10_3, output_10_4, output_9_3;
mixer gate_output_9_3(.a(output_10_3), .b(output_10_4), .y(output_9_3));
wire output_11_3, output_11_4, output_10_3;
mixer gate_output_10_3(.a(output_11_3), .b(output_11_4), .y(output_10_3));
wire output_12_3, output_12_4, output_11_3;
mixer gate_output_11_3(.a(output_12_3), .b(output_12_4), .y(output_11_3));
wire output_13_3, output_13_4, output_12_3;
mixer gate_output_12_3(.a(output_13_3), .b(output_13_4), .y(output_12_3));
wire output_14_3, output_14_4, output_13_3;
mixer gate_output_13_3(.a(output_14_3), .b(output_14_4), .y(output_13_3));
wire output_15_3, output_15_4, output_14_3;
mixer gate_output_14_3(.a(output_15_3), .b(output_15_4), .y(output_14_3));
wire output_16_3, output_16_4, output_15_3;
mixer gate_output_15_3(.a(output_16_3), .b(output_16_4), .y(output_15_3));
wire output_1_4, output_1_5, output_0_4;
mixer gate_output_0_4(.a(output_1_4), .b(output_1_5), .y(output_0_4));
wire output_2_4, output_2_5, output_1_4;
mixer gate_output_1_4(.a(output_2_4), .b(output_2_5), .y(output_1_4));
wire output_3_4, output_3_5, output_2_4;
mixer gate_output_2_4(.a(output_3_4), .b(output_3_5), .y(output_2_4));
wire output_4_4, output_4_5, output_3_4;
mixer gate_output_3_4(.a(output_4_4), .b(output_4_5), .y(output_3_4));
wire output_5_4, output_5_5, output_4_4;
mixer gate_output_4_4(.a(output_5_4), .b(output_5_5), .y(output_4_4));
wire output_6_4, output_6_5, output_5_4;
mixer gate_output_5_4(.a(output_6_4), .b(output_6_5), .y(output_5_4));
wire output_7_4, output_7_5, output_6_4;
mixer gate_output_6_4(.a(output_7_4), .b(output_7_5), .y(output_6_4));
wire output_8_4, output_8_5, output_7_4;
mixer gate_output_7_4(.a(output_8_4), .b(output_8_5), .y(output_7_4));
wire output_9_4, output_9_5, output_8_4;
mixer gate_output_8_4(.a(output_9_4), .b(output_9_5), .y(output_8_4));
wire output_10_4, output_10_5, output_9_4;
mixer gate_output_9_4(.a(output_10_4), .b(output_10_5), .y(output_9_4));
wire output_11_4, output_11_5, output_10_4;
mixer gate_output_10_4(.a(output_11_4), .b(output_11_5), .y(output_10_4));
wire output_12_4, output_12_5, output_11_4;
mixer gate_output_11_4(.a(output_12_4), .b(output_12_5), .y(output_11_4));
wire output_13_4, output_13_5, output_12_4;
mixer gate_output_12_4(.a(output_13_4), .b(output_13_5), .y(output_12_4));
wire output_14_4, output_14_5, output_13_4;
mixer gate_output_13_4(.a(output_14_4), .b(output_14_5), .y(output_13_4));
wire output_15_4, output_15_5, output_14_4;
mixer gate_output_14_4(.a(output_15_4), .b(output_15_5), .y(output_14_4));
wire output_16_4, output_16_5, output_15_4;
mixer gate_output_15_4(.a(output_16_4), .b(output_16_5), .y(output_15_4));
wire output_1_5, output_1_6, output_0_5;
mixer gate_output_0_5(.a(output_1_5), .b(output_1_6), .y(output_0_5));
wire output_2_5, output_2_6, output_1_5;
mixer gate_output_1_5(.a(output_2_5), .b(output_2_6), .y(output_1_5));
wire output_3_5, output_3_6, output_2_5;
mixer gate_output_2_5(.a(output_3_5), .b(output_3_6), .y(output_2_5));
wire output_4_5, output_4_6, output_3_5;
mixer gate_output_3_5(.a(output_4_5), .b(output_4_6), .y(output_3_5));
wire output_5_5, output_5_6, output_4_5;
mixer gate_output_4_5(.a(output_5_5), .b(output_5_6), .y(output_4_5));
wire output_6_5, output_6_6, output_5_5;
mixer gate_output_5_5(.a(output_6_5), .b(output_6_6), .y(output_5_5));
wire output_7_5, output_7_6, output_6_5;
mixer gate_output_6_5(.a(output_7_5), .b(output_7_6), .y(output_6_5));
wire output_8_5, output_8_6, output_7_5;
mixer gate_output_7_5(.a(output_8_5), .b(output_8_6), .y(output_7_5));
wire output_9_5, output_9_6, output_8_5;
mixer gate_output_8_5(.a(output_9_5), .b(output_9_6), .y(output_8_5));
wire output_10_5, output_10_6, output_9_5;
mixer gate_output_9_5(.a(output_10_5), .b(output_10_6), .y(output_9_5));
wire output_11_5, output_11_6, output_10_5;
mixer gate_output_10_5(.a(output_11_5), .b(output_11_6), .y(output_10_5));
wire output_12_5, output_12_6, output_11_5;
mixer gate_output_11_5(.a(output_12_5), .b(output_12_6), .y(output_11_5));
wire output_13_5, output_13_6, output_12_5;
mixer gate_output_12_5(.a(output_13_5), .b(output_13_6), .y(output_12_5));
wire output_14_5, output_14_6, output_13_5;
mixer gate_output_13_5(.a(output_14_5), .b(output_14_6), .y(output_13_5));
wire output_15_5, output_15_6, output_14_5;
mixer gate_output_14_5(.a(output_15_5), .b(output_15_6), .y(output_14_5));
wire output_16_5, output_16_6, output_15_5;
mixer gate_output_15_5(.a(output_16_5), .b(output_16_6), .y(output_15_5));
wire output_1_6, output_1_7, output_0_6;
mixer gate_output_0_6(.a(output_1_6), .b(output_1_7), .y(output_0_6));
wire output_2_6, output_2_7, output_1_6;
mixer gate_output_1_6(.a(output_2_6), .b(output_2_7), .y(output_1_6));
wire output_3_6, output_3_7, output_2_6;
mixer gate_output_2_6(.a(output_3_6), .b(output_3_7), .y(output_2_6));
wire output_4_6, output_4_7, output_3_6;
mixer gate_output_3_6(.a(output_4_6), .b(output_4_7), .y(output_3_6));
wire output_5_6, output_5_7, output_4_6;
mixer gate_output_4_6(.a(output_5_6), .b(output_5_7), .y(output_4_6));
wire output_6_6, output_6_7, output_5_6;
mixer gate_output_5_6(.a(output_6_6), .b(output_6_7), .y(output_5_6));
wire output_7_6, output_7_7, output_6_6;
mixer gate_output_6_6(.a(output_7_6), .b(output_7_7), .y(output_6_6));
wire output_8_6, output_8_7, output_7_6;
mixer gate_output_7_6(.a(output_8_6), .b(output_8_7), .y(output_7_6));
wire output_9_6, output_9_7, output_8_6;
mixer gate_output_8_6(.a(output_9_6), .b(output_9_7), .y(output_8_6));
wire output_10_6, output_10_7, output_9_6;
mixer gate_output_9_6(.a(output_10_6), .b(output_10_7), .y(output_9_6));
wire output_11_6, output_11_7, output_10_6;
mixer gate_output_10_6(.a(output_11_6), .b(output_11_7), .y(output_10_6));
wire output_12_6, output_12_7, output_11_6;
mixer gate_output_11_6(.a(output_12_6), .b(output_12_7), .y(output_11_6));
wire output_13_6, output_13_7, output_12_6;
mixer gate_output_12_6(.a(output_13_6), .b(output_13_7), .y(output_12_6));
wire output_14_6, output_14_7, output_13_6;
mixer gate_output_13_6(.a(output_14_6), .b(output_14_7), .y(output_13_6));
wire output_15_6, output_15_7, output_14_6;
mixer gate_output_14_6(.a(output_15_6), .b(output_15_7), .y(output_14_6));
wire output_16_6, output_16_7, output_15_6;
mixer gate_output_15_6(.a(output_16_6), .b(output_16_7), .y(output_15_6));
wire output_1_7, output_1_8, output_0_7;
mixer gate_output_0_7(.a(output_1_7), .b(output_1_8), .y(output_0_7));
wire output_2_7, output_2_8, output_1_7;
mixer gate_output_1_7(.a(output_2_7), .b(output_2_8), .y(output_1_7));
wire output_3_7, output_3_8, output_2_7;
mixer gate_output_2_7(.a(output_3_7), .b(output_3_8), .y(output_2_7));
wire output_4_7, output_4_8, output_3_7;
mixer gate_output_3_7(.a(output_4_7), .b(output_4_8), .y(output_3_7));
wire output_5_7, output_5_8, output_4_7;
mixer gate_output_4_7(.a(output_5_7), .b(output_5_8), .y(output_4_7));
wire output_6_7, output_6_8, output_5_7;
mixer gate_output_5_7(.a(output_6_7), .b(output_6_8), .y(output_5_7));
wire output_7_7, output_7_8, output_6_7;
mixer gate_output_6_7(.a(output_7_7), .b(output_7_8), .y(output_6_7));
wire output_8_7, output_8_8, output_7_7;
mixer gate_output_7_7(.a(output_8_7), .b(output_8_8), .y(output_7_7));
wire output_9_7, output_9_8, output_8_7;
mixer gate_output_8_7(.a(output_9_7), .b(output_9_8), .y(output_8_7));
wire output_10_7, output_10_8, output_9_7;
mixer gate_output_9_7(.a(output_10_7), .b(output_10_8), .y(output_9_7));
wire output_11_7, output_11_8, output_10_7;
mixer gate_output_10_7(.a(output_11_7), .b(output_11_8), .y(output_10_7));
wire output_12_7, output_12_8, output_11_7;
mixer gate_output_11_7(.a(output_12_7), .b(output_12_8), .y(output_11_7));
wire output_13_7, output_13_8, output_12_7;
mixer gate_output_12_7(.a(output_13_7), .b(output_13_8), .y(output_12_7));
wire output_14_7, output_14_8, output_13_7;
mixer gate_output_13_7(.a(output_14_7), .b(output_14_8), .y(output_13_7));
wire output_15_7, output_15_8, output_14_7;
mixer gate_output_14_7(.a(output_15_7), .b(output_15_8), .y(output_14_7));
wire output_16_7, output_16_8, output_15_7;
mixer gate_output_15_7(.a(output_16_7), .b(output_16_8), .y(output_15_7));
wire output_1_8, output_1_9, output_0_8;
mixer gate_output_0_8(.a(output_1_8), .b(output_1_9), .y(output_0_8));
wire output_2_8, output_2_9, output_1_8;
mixer gate_output_1_8(.a(output_2_8), .b(output_2_9), .y(output_1_8));
wire output_3_8, output_3_9, output_2_8;
mixer gate_output_2_8(.a(output_3_8), .b(output_3_9), .y(output_2_8));
wire output_4_8, output_4_9, output_3_8;
mixer gate_output_3_8(.a(output_4_8), .b(output_4_9), .y(output_3_8));
wire output_5_8, output_5_9, output_4_8;
mixer gate_output_4_8(.a(output_5_8), .b(output_5_9), .y(output_4_8));
wire output_6_8, output_6_9, output_5_8;
mixer gate_output_5_8(.a(output_6_8), .b(output_6_9), .y(output_5_8));
wire output_7_8, output_7_9, output_6_8;
mixer gate_output_6_8(.a(output_7_8), .b(output_7_9), .y(output_6_8));
wire output_8_8, output_8_9, output_7_8;
mixer gate_output_7_8(.a(output_8_8), .b(output_8_9), .y(output_7_8));
wire output_9_8, output_9_9, output_8_8;
mixer gate_output_8_8(.a(output_9_8), .b(output_9_9), .y(output_8_8));
wire output_10_8, output_10_9, output_9_8;
mixer gate_output_9_8(.a(output_10_8), .b(output_10_9), .y(output_9_8));
wire output_11_8, output_11_9, output_10_8;
mixer gate_output_10_8(.a(output_11_8), .b(output_11_9), .y(output_10_8));
wire output_12_8, output_12_9, output_11_8;
mixer gate_output_11_8(.a(output_12_8), .b(output_12_9), .y(output_11_8));
wire output_13_8, output_13_9, output_12_8;
mixer gate_output_12_8(.a(output_13_8), .b(output_13_9), .y(output_12_8));
wire output_14_8, output_14_9, output_13_8;
mixer gate_output_13_8(.a(output_14_8), .b(output_14_9), .y(output_13_8));
wire output_15_8, output_15_9, output_14_8;
mixer gate_output_14_8(.a(output_15_8), .b(output_15_9), .y(output_14_8));
wire output_16_8, output_16_9, output_15_8;
mixer gate_output_15_8(.a(output_16_8), .b(output_16_9), .y(output_15_8));
wire output_1_9, output_1_10, output_0_9;
mixer gate_output_0_9(.a(output_1_9), .b(output_1_10), .y(output_0_9));
wire output_2_9, output_2_10, output_1_9;
mixer gate_output_1_9(.a(output_2_9), .b(output_2_10), .y(output_1_9));
wire output_3_9, output_3_10, output_2_9;
mixer gate_output_2_9(.a(output_3_9), .b(output_3_10), .y(output_2_9));
wire output_4_9, output_4_10, output_3_9;
mixer gate_output_3_9(.a(output_4_9), .b(output_4_10), .y(output_3_9));
wire output_5_9, output_5_10, output_4_9;
mixer gate_output_4_9(.a(output_5_9), .b(output_5_10), .y(output_4_9));
wire output_6_9, output_6_10, output_5_9;
mixer gate_output_5_9(.a(output_6_9), .b(output_6_10), .y(output_5_9));
wire output_7_9, output_7_10, output_6_9;
mixer gate_output_6_9(.a(output_7_9), .b(output_7_10), .y(output_6_9));
wire output_8_9, output_8_10, output_7_9;
mixer gate_output_7_9(.a(output_8_9), .b(output_8_10), .y(output_7_9));
wire output_9_9, output_9_10, output_8_9;
mixer gate_output_8_9(.a(output_9_9), .b(output_9_10), .y(output_8_9));
wire output_10_9, output_10_10, output_9_9;
mixer gate_output_9_9(.a(output_10_9), .b(output_10_10), .y(output_9_9));
wire output_11_9, output_11_10, output_10_9;
mixer gate_output_10_9(.a(output_11_9), .b(output_11_10), .y(output_10_9));
wire output_12_9, output_12_10, output_11_9;
mixer gate_output_11_9(.a(output_12_9), .b(output_12_10), .y(output_11_9));
wire output_13_9, output_13_10, output_12_9;
mixer gate_output_12_9(.a(output_13_9), .b(output_13_10), .y(output_12_9));
wire output_14_9, output_14_10, output_13_9;
mixer gate_output_13_9(.a(output_14_9), .b(output_14_10), .y(output_13_9));
wire output_15_9, output_15_10, output_14_9;
mixer gate_output_14_9(.a(output_15_9), .b(output_15_10), .y(output_14_9));
wire output_16_9, output_16_10, output_15_9;
mixer gate_output_15_9(.a(output_16_9), .b(output_16_10), .y(output_15_9));
wire output_1_10, output_1_11, output_0_10;
mixer gate_output_0_10(.a(output_1_10), .b(output_1_11), .y(output_0_10));
wire output_2_10, output_2_11, output_1_10;
mixer gate_output_1_10(.a(output_2_10), .b(output_2_11), .y(output_1_10));
wire output_3_10, output_3_11, output_2_10;
mixer gate_output_2_10(.a(output_3_10), .b(output_3_11), .y(output_2_10));
wire output_4_10, output_4_11, output_3_10;
mixer gate_output_3_10(.a(output_4_10), .b(output_4_11), .y(output_3_10));
wire output_5_10, output_5_11, output_4_10;
mixer gate_output_4_10(.a(output_5_10), .b(output_5_11), .y(output_4_10));
wire output_6_10, output_6_11, output_5_10;
mixer gate_output_5_10(.a(output_6_10), .b(output_6_11), .y(output_5_10));
wire output_7_10, output_7_11, output_6_10;
mixer gate_output_6_10(.a(output_7_10), .b(output_7_11), .y(output_6_10));
wire output_8_10, output_8_11, output_7_10;
mixer gate_output_7_10(.a(output_8_10), .b(output_8_11), .y(output_7_10));
wire output_9_10, output_9_11, output_8_10;
mixer gate_output_8_10(.a(output_9_10), .b(output_9_11), .y(output_8_10));
wire output_10_10, output_10_11, output_9_10;
mixer gate_output_9_10(.a(output_10_10), .b(output_10_11), .y(output_9_10));
wire output_11_10, output_11_11, output_10_10;
mixer gate_output_10_10(.a(output_11_10), .b(output_11_11), .y(output_10_10));
wire output_12_10, output_12_11, output_11_10;
mixer gate_output_11_10(.a(output_12_10), .b(output_12_11), .y(output_11_10));
wire output_13_10, output_13_11, output_12_10;
mixer gate_output_12_10(.a(output_13_10), .b(output_13_11), .y(output_12_10));
wire output_14_10, output_14_11, output_13_10;
mixer gate_output_13_10(.a(output_14_10), .b(output_14_11), .y(output_13_10));
wire output_15_10, output_15_11, output_14_10;
mixer gate_output_14_10(.a(output_15_10), .b(output_15_11), .y(output_14_10));
wire output_16_10, output_16_11, output_15_10;
mixer gate_output_15_10(.a(output_16_10), .b(output_16_11), .y(output_15_10));
wire output_1_11, output_1_12, output_0_11;
mixer gate_output_0_11(.a(output_1_11), .b(output_1_12), .y(output_0_11));
wire output_2_11, output_2_12, output_1_11;
mixer gate_output_1_11(.a(output_2_11), .b(output_2_12), .y(output_1_11));
wire output_3_11, output_3_12, output_2_11;
mixer gate_output_2_11(.a(output_3_11), .b(output_3_12), .y(output_2_11));
wire output_4_11, output_4_12, output_3_11;
mixer gate_output_3_11(.a(output_4_11), .b(output_4_12), .y(output_3_11));
wire output_5_11, output_5_12, output_4_11;
mixer gate_output_4_11(.a(output_5_11), .b(output_5_12), .y(output_4_11));
wire output_6_11, output_6_12, output_5_11;
mixer gate_output_5_11(.a(output_6_11), .b(output_6_12), .y(output_5_11));
wire output_7_11, output_7_12, output_6_11;
mixer gate_output_6_11(.a(output_7_11), .b(output_7_12), .y(output_6_11));
wire output_8_11, output_8_12, output_7_11;
mixer gate_output_7_11(.a(output_8_11), .b(output_8_12), .y(output_7_11));
wire output_9_11, output_9_12, output_8_11;
mixer gate_output_8_11(.a(output_9_11), .b(output_9_12), .y(output_8_11));
wire output_10_11, output_10_12, output_9_11;
mixer gate_output_9_11(.a(output_10_11), .b(output_10_12), .y(output_9_11));
wire output_11_11, output_11_12, output_10_11;
mixer gate_output_10_11(.a(output_11_11), .b(output_11_12), .y(output_10_11));
wire output_12_11, output_12_12, output_11_11;
mixer gate_output_11_11(.a(output_12_11), .b(output_12_12), .y(output_11_11));
wire output_13_11, output_13_12, output_12_11;
mixer gate_output_12_11(.a(output_13_11), .b(output_13_12), .y(output_12_11));
wire output_14_11, output_14_12, output_13_11;
mixer gate_output_13_11(.a(output_14_11), .b(output_14_12), .y(output_13_11));
wire output_15_11, output_15_12, output_14_11;
mixer gate_output_14_11(.a(output_15_11), .b(output_15_12), .y(output_14_11));
wire output_16_11, output_16_12, output_15_11;
mixer gate_output_15_11(.a(output_16_11), .b(output_16_12), .y(output_15_11));
wire output_1_12, output_1_13, output_0_12;
mixer gate_output_0_12(.a(output_1_12), .b(output_1_13), .y(output_0_12));
wire output_2_12, output_2_13, output_1_12;
mixer gate_output_1_12(.a(output_2_12), .b(output_2_13), .y(output_1_12));
wire output_3_12, output_3_13, output_2_12;
mixer gate_output_2_12(.a(output_3_12), .b(output_3_13), .y(output_2_12));
wire output_4_12, output_4_13, output_3_12;
mixer gate_output_3_12(.a(output_4_12), .b(output_4_13), .y(output_3_12));
wire output_5_12, output_5_13, output_4_12;
mixer gate_output_4_12(.a(output_5_12), .b(output_5_13), .y(output_4_12));
wire output_6_12, output_6_13, output_5_12;
mixer gate_output_5_12(.a(output_6_12), .b(output_6_13), .y(output_5_12));
wire output_7_12, output_7_13, output_6_12;
mixer gate_output_6_12(.a(output_7_12), .b(output_7_13), .y(output_6_12));
wire output_8_12, output_8_13, output_7_12;
mixer gate_output_7_12(.a(output_8_12), .b(output_8_13), .y(output_7_12));
wire output_9_12, output_9_13, output_8_12;
mixer gate_output_8_12(.a(output_9_12), .b(output_9_13), .y(output_8_12));
wire output_10_12, output_10_13, output_9_12;
mixer gate_output_9_12(.a(output_10_12), .b(output_10_13), .y(output_9_12));
wire output_11_12, output_11_13, output_10_12;
mixer gate_output_10_12(.a(output_11_12), .b(output_11_13), .y(output_10_12));
wire output_12_12, output_12_13, output_11_12;
mixer gate_output_11_12(.a(output_12_12), .b(output_12_13), .y(output_11_12));
wire output_13_12, output_13_13, output_12_12;
mixer gate_output_12_12(.a(output_13_12), .b(output_13_13), .y(output_12_12));
wire output_14_12, output_14_13, output_13_12;
mixer gate_output_13_12(.a(output_14_12), .b(output_14_13), .y(output_13_12));
wire output_15_12, output_15_13, output_14_12;
mixer gate_output_14_12(.a(output_15_12), .b(output_15_13), .y(output_14_12));
wire output_16_12, output_16_13, output_15_12;
mixer gate_output_15_12(.a(output_16_12), .b(output_16_13), .y(output_15_12));
wire output_1_13, output_1_14, output_0_13;
mixer gate_output_0_13(.a(output_1_13), .b(output_1_14), .y(output_0_13));
wire output_2_13, output_2_14, output_1_13;
mixer gate_output_1_13(.a(output_2_13), .b(output_2_14), .y(output_1_13));
wire output_3_13, output_3_14, output_2_13;
mixer gate_output_2_13(.a(output_3_13), .b(output_3_14), .y(output_2_13));
wire output_4_13, output_4_14, output_3_13;
mixer gate_output_3_13(.a(output_4_13), .b(output_4_14), .y(output_3_13));
wire output_5_13, output_5_14, output_4_13;
mixer gate_output_4_13(.a(output_5_13), .b(output_5_14), .y(output_4_13));
wire output_6_13, output_6_14, output_5_13;
mixer gate_output_5_13(.a(output_6_13), .b(output_6_14), .y(output_5_13));
wire output_7_13, output_7_14, output_6_13;
mixer gate_output_6_13(.a(output_7_13), .b(output_7_14), .y(output_6_13));
wire output_8_13, output_8_14, output_7_13;
mixer gate_output_7_13(.a(output_8_13), .b(output_8_14), .y(output_7_13));
wire output_9_13, output_9_14, output_8_13;
mixer gate_output_8_13(.a(output_9_13), .b(output_9_14), .y(output_8_13));
wire output_10_13, output_10_14, output_9_13;
mixer gate_output_9_13(.a(output_10_13), .b(output_10_14), .y(output_9_13));
wire output_11_13, output_11_14, output_10_13;
mixer gate_output_10_13(.a(output_11_13), .b(output_11_14), .y(output_10_13));
wire output_12_13, output_12_14, output_11_13;
mixer gate_output_11_13(.a(output_12_13), .b(output_12_14), .y(output_11_13));
wire output_13_13, output_13_14, output_12_13;
mixer gate_output_12_13(.a(output_13_13), .b(output_13_14), .y(output_12_13));
wire output_14_13, output_14_14, output_13_13;
mixer gate_output_13_13(.a(output_14_13), .b(output_14_14), .y(output_13_13));
wire output_15_13, output_15_14, output_14_13;
mixer gate_output_14_13(.a(output_15_13), .b(output_15_14), .y(output_14_13));
wire output_16_13, output_16_14, output_15_13;
mixer gate_output_15_13(.a(output_16_13), .b(output_16_14), .y(output_15_13));
wire output_1_14, output_1_15, output_0_14;
mixer gate_output_0_14(.a(output_1_14), .b(output_1_15), .y(output_0_14));
wire output_2_14, output_2_15, output_1_14;
mixer gate_output_1_14(.a(output_2_14), .b(output_2_15), .y(output_1_14));
wire output_3_14, output_3_15, output_2_14;
mixer gate_output_2_14(.a(output_3_14), .b(output_3_15), .y(output_2_14));
wire output_4_14, output_4_15, output_3_14;
mixer gate_output_3_14(.a(output_4_14), .b(output_4_15), .y(output_3_14));
wire output_5_14, output_5_15, output_4_14;
mixer gate_output_4_14(.a(output_5_14), .b(output_5_15), .y(output_4_14));
wire output_6_14, output_6_15, output_5_14;
mixer gate_output_5_14(.a(output_6_14), .b(output_6_15), .y(output_5_14));
wire output_7_14, output_7_15, output_6_14;
mixer gate_output_6_14(.a(output_7_14), .b(output_7_15), .y(output_6_14));
wire output_8_14, output_8_15, output_7_14;
mixer gate_output_7_14(.a(output_8_14), .b(output_8_15), .y(output_7_14));
wire output_9_14, output_9_15, output_8_14;
mixer gate_output_8_14(.a(output_9_14), .b(output_9_15), .y(output_8_14));
wire output_10_14, output_10_15, output_9_14;
mixer gate_output_9_14(.a(output_10_14), .b(output_10_15), .y(output_9_14));
wire output_11_14, output_11_15, output_10_14;
mixer gate_output_10_14(.a(output_11_14), .b(output_11_15), .y(output_10_14));
wire output_12_14, output_12_15, output_11_14;
mixer gate_output_11_14(.a(output_12_14), .b(output_12_15), .y(output_11_14));
wire output_13_14, output_13_15, output_12_14;
mixer gate_output_12_14(.a(output_13_14), .b(output_13_15), .y(output_12_14));
wire output_14_14, output_14_15, output_13_14;
mixer gate_output_13_14(.a(output_14_14), .b(output_14_15), .y(output_13_14));
wire output_15_14, output_15_15, output_14_14;
mixer gate_output_14_14(.a(output_15_14), .b(output_15_15), .y(output_14_14));
wire output_16_14, output_16_15, output_15_14;
mixer gate_output_15_14(.a(output_16_14), .b(output_16_15), .y(output_15_14));
wire output_1_15, output_1_0, output_0_15;
mixer gate_output_0_15(.a(output_1_15), .b(output_1_0), .y(output_0_15));
wire output_2_15, output_2_0, output_1_15;
mixer gate_output_1_15(.a(output_2_15), .b(output_2_0), .y(output_1_15));
wire output_3_15, output_3_0, output_2_15;
mixer gate_output_2_15(.a(output_3_15), .b(output_3_0), .y(output_2_15));
wire output_4_15, output_4_0, output_3_15;
mixer gate_output_3_15(.a(output_4_15), .b(output_4_0), .y(output_3_15));
wire output_5_15, output_5_0, output_4_15;
mixer gate_output_4_15(.a(output_5_15), .b(output_5_0), .y(output_4_15));
wire output_6_15, output_6_0, output_5_15;
mixer gate_output_5_15(.a(output_6_15), .b(output_6_0), .y(output_5_15));
wire output_7_15, output_7_0, output_6_15;
mixer gate_output_6_15(.a(output_7_15), .b(output_7_0), .y(output_6_15));
wire output_8_15, output_8_0, output_7_15;
mixer gate_output_7_15(.a(output_8_15), .b(output_8_0), .y(output_7_15));
wire output_9_15, output_9_0, output_8_15;
mixer gate_output_8_15(.a(output_9_15), .b(output_9_0), .y(output_8_15));
wire output_10_15, output_10_0, output_9_15;
mixer gate_output_9_15(.a(output_10_15), .b(output_10_0), .y(output_9_15));
wire output_11_15, output_11_0, output_10_15;
mixer gate_output_10_15(.a(output_11_15), .b(output_11_0), .y(output_10_15));
wire output_12_15, output_12_0, output_11_15;
mixer gate_output_11_15(.a(output_12_15), .b(output_12_0), .y(output_11_15));
wire output_13_15, output_13_0, output_12_15;
mixer gate_output_12_15(.a(output_13_15), .b(output_13_0), .y(output_12_15));
wire output_14_15, output_14_0, output_13_15;
mixer gate_output_13_15(.a(output_14_15), .b(output_14_0), .y(output_13_15));
wire output_15_15, output_15_0, output_14_15;
mixer gate_output_14_15(.a(output_15_15), .b(output_15_0), .y(output_14_15));
wire output_16_15, output_16_0, output_15_15;
mixer gate_output_15_15(.a(output_16_15), .b(output_16_0), .y(output_15_15));
wire output_1_16, output_1_1, output_0_16;
mixer gate_output_0_16(.a(output_1_16), .b(output_1_1), .y(output_0_16));
wire output_2_16, output_2_1, output_1_16;
mixer gate_output_1_16(.a(output_2_16), .b(output_2_1), .y(output_1_16));
wire output_3_16, output_3_1, output_2_16;
mixer gate_output_2_16(.a(output_3_16), .b(output_3_1), .y(output_2_16));
wire output_4_16, output_4_1, output_3_16;
mixer gate_output_3_16(.a(output_4_16), .b(output_4_1), .y(output_3_16));
wire output_5_16, output_5_1, output_4_16;
mixer gate_output_4_16(.a(output_5_16), .b(output_5_1), .y(output_4_16));
wire output_6_16, output_6_1, output_5_16;
mixer gate_output_5_16(.a(output_6_16), .b(output_6_1), .y(output_5_16));
wire output_7_16, output_7_1, output_6_16;
mixer gate_output_6_16(.a(output_7_16), .b(output_7_1), .y(output_6_16));
wire output_8_16, output_8_1, output_7_16;
mixer gate_output_7_16(.a(output_8_16), .b(output_8_1), .y(output_7_16));
wire output_9_16, output_9_1, output_8_16;
mixer gate_output_8_16(.a(output_9_16), .b(output_9_1), .y(output_8_16));
wire output_10_16, output_10_1, output_9_16;
mixer gate_output_9_16(.a(output_10_16), .b(output_10_1), .y(output_9_16));
wire output_11_16, output_11_1, output_10_16;
mixer gate_output_10_16(.a(output_11_16), .b(output_11_1), .y(output_10_16));
wire output_12_16, output_12_1, output_11_16;
mixer gate_output_11_16(.a(output_12_16), .b(output_12_1), .y(output_11_16));
wire output_13_16, output_13_1, output_12_16;
mixer gate_output_12_16(.a(output_13_16), .b(output_13_1), .y(output_12_16));
wire output_14_16, output_14_1, output_13_16;
mixer gate_output_13_16(.a(output_14_16), .b(output_14_1), .y(output_13_16));
wire output_15_16, output_15_1, output_14_16;
mixer gate_output_14_16(.a(output_15_16), .b(output_15_1), .y(output_14_16));
wire output_16_16, output_16_1, output_15_16;
mixer gate_output_15_16(.a(output_16_16), .b(output_16_1), .y(output_15_16));
wire output_1_17, output_1_2, output_0_17;
mixer gate_output_0_17(.a(output_1_17), .b(output_1_2), .y(output_0_17));
wire output_2_17, output_2_2, output_1_17;
mixer gate_output_1_17(.a(output_2_17), .b(output_2_2), .y(output_1_17));
wire output_3_17, output_3_2, output_2_17;
mixer gate_output_2_17(.a(output_3_17), .b(output_3_2), .y(output_2_17));
wire output_4_17, output_4_2, output_3_17;
mixer gate_output_3_17(.a(output_4_17), .b(output_4_2), .y(output_3_17));
wire output_5_17, output_5_2, output_4_17;
mixer gate_output_4_17(.a(output_5_17), .b(output_5_2), .y(output_4_17));
wire output_6_17, output_6_2, output_5_17;
mixer gate_output_5_17(.a(output_6_17), .b(output_6_2), .y(output_5_17));
wire output_7_17, output_7_2, output_6_17;
mixer gate_output_6_17(.a(output_7_17), .b(output_7_2), .y(output_6_17));
wire output_8_17, output_8_2, output_7_17;
mixer gate_output_7_17(.a(output_8_17), .b(output_8_2), .y(output_7_17));
wire output_9_17, output_9_2, output_8_17;
mixer gate_output_8_17(.a(output_9_17), .b(output_9_2), .y(output_8_17));
wire output_10_17, output_10_2, output_9_17;
mixer gate_output_9_17(.a(output_10_17), .b(output_10_2), .y(output_9_17));
wire output_11_17, output_11_2, output_10_17;
mixer gate_output_10_17(.a(output_11_17), .b(output_11_2), .y(output_10_17));
wire output_12_17, output_12_2, output_11_17;
mixer gate_output_11_17(.a(output_12_17), .b(output_12_2), .y(output_11_17));
wire output_13_17, output_13_2, output_12_17;
mixer gate_output_12_17(.a(output_13_17), .b(output_13_2), .y(output_12_17));
wire output_14_17, output_14_2, output_13_17;
mixer gate_output_13_17(.a(output_14_17), .b(output_14_2), .y(output_13_17));
wire output_15_17, output_15_2, output_14_17;
mixer gate_output_14_17(.a(output_15_17), .b(output_15_2), .y(output_14_17));
wire output_16_17, output_16_2, output_15_17;
mixer gate_output_15_17(.a(output_16_17), .b(output_16_2), .y(output_15_17));
wire output_1_18, output_1_3, output_0_18;
mixer gate_output_0_18(.a(output_1_18), .b(output_1_3), .y(output_0_18));
wire output_2_18, output_2_3, output_1_18;
mixer gate_output_1_18(.a(output_2_18), .b(output_2_3), .y(output_1_18));
wire output_3_18, output_3_3, output_2_18;
mixer gate_output_2_18(.a(output_3_18), .b(output_3_3), .y(output_2_18));
wire output_4_18, output_4_3, output_3_18;
mixer gate_output_3_18(.a(output_4_18), .b(output_4_3), .y(output_3_18));
wire output_5_18, output_5_3, output_4_18;
mixer gate_output_4_18(.a(output_5_18), .b(output_5_3), .y(output_4_18));
wire output_6_18, output_6_3, output_5_18;
mixer gate_output_5_18(.a(output_6_18), .b(output_6_3), .y(output_5_18));
wire output_7_18, output_7_3, output_6_18;
mixer gate_output_6_18(.a(output_7_18), .b(output_7_3), .y(output_6_18));
wire output_8_18, output_8_3, output_7_18;
mixer gate_output_7_18(.a(output_8_18), .b(output_8_3), .y(output_7_18));
wire output_9_18, output_9_3, output_8_18;
mixer gate_output_8_18(.a(output_9_18), .b(output_9_3), .y(output_8_18));
wire output_10_18, output_10_3, output_9_18;
mixer gate_output_9_18(.a(output_10_18), .b(output_10_3), .y(output_9_18));
wire output_11_18, output_11_3, output_10_18;
mixer gate_output_10_18(.a(output_11_18), .b(output_11_3), .y(output_10_18));
wire output_12_18, output_12_3, output_11_18;
mixer gate_output_11_18(.a(output_12_18), .b(output_12_3), .y(output_11_18));
wire output_13_18, output_13_3, output_12_18;
mixer gate_output_12_18(.a(output_13_18), .b(output_13_3), .y(output_12_18));
wire output_14_18, output_14_3, output_13_18;
mixer gate_output_13_18(.a(output_14_18), .b(output_14_3), .y(output_13_18));
wire output_15_18, output_15_3, output_14_18;
mixer gate_output_14_18(.a(output_15_18), .b(output_15_3), .y(output_14_18));
wire output_16_18, output_16_3, output_15_18;
mixer gate_output_15_18(.a(output_16_18), .b(output_16_3), .y(output_15_18));
wire output_1_19, output_1_4, output_0_19;
mixer gate_output_0_19(.a(output_1_19), .b(output_1_4), .y(output_0_19));
wire output_2_19, output_2_4, output_1_19;
mixer gate_output_1_19(.a(output_2_19), .b(output_2_4), .y(output_1_19));
wire output_3_19, output_3_4, output_2_19;
mixer gate_output_2_19(.a(output_3_19), .b(output_3_4), .y(output_2_19));
wire output_4_19, output_4_4, output_3_19;
mixer gate_output_3_19(.a(output_4_19), .b(output_4_4), .y(output_3_19));
wire output_5_19, output_5_4, output_4_19;
mixer gate_output_4_19(.a(output_5_19), .b(output_5_4), .y(output_4_19));
wire output_6_19, output_6_4, output_5_19;
mixer gate_output_5_19(.a(output_6_19), .b(output_6_4), .y(output_5_19));
wire output_7_19, output_7_4, output_6_19;
mixer gate_output_6_19(.a(output_7_19), .b(output_7_4), .y(output_6_19));
wire output_8_19, output_8_4, output_7_19;
mixer gate_output_7_19(.a(output_8_19), .b(output_8_4), .y(output_7_19));
wire output_9_19, output_9_4, output_8_19;
mixer gate_output_8_19(.a(output_9_19), .b(output_9_4), .y(output_8_19));
wire output_10_19, output_10_4, output_9_19;
mixer gate_output_9_19(.a(output_10_19), .b(output_10_4), .y(output_9_19));
wire output_11_19, output_11_4, output_10_19;
mixer gate_output_10_19(.a(output_11_19), .b(output_11_4), .y(output_10_19));
wire output_12_19, output_12_4, output_11_19;
mixer gate_output_11_19(.a(output_12_19), .b(output_12_4), .y(output_11_19));
wire output_13_19, output_13_4, output_12_19;
mixer gate_output_12_19(.a(output_13_19), .b(output_13_4), .y(output_12_19));
wire output_14_19, output_14_4, output_13_19;
mixer gate_output_13_19(.a(output_14_19), .b(output_14_4), .y(output_13_19));
wire output_15_19, output_15_4, output_14_19;
mixer gate_output_14_19(.a(output_15_19), .b(output_15_4), .y(output_14_19));
wire output_16_19, output_16_4, output_15_19;
mixer gate_output_15_19(.a(output_16_19), .b(output_16_4), .y(output_15_19));
wire output_1_20, output_1_5, output_0_20;
mixer gate_output_0_20(.a(output_1_20), .b(output_1_5), .y(output_0_20));
wire output_2_20, output_2_5, output_1_20;
mixer gate_output_1_20(.a(output_2_20), .b(output_2_5), .y(output_1_20));
wire output_3_20, output_3_5, output_2_20;
mixer gate_output_2_20(.a(output_3_20), .b(output_3_5), .y(output_2_20));
wire output_4_20, output_4_5, output_3_20;
mixer gate_output_3_20(.a(output_4_20), .b(output_4_5), .y(output_3_20));
wire output_5_20, output_5_5, output_4_20;
mixer gate_output_4_20(.a(output_5_20), .b(output_5_5), .y(output_4_20));
wire output_6_20, output_6_5, output_5_20;
mixer gate_output_5_20(.a(output_6_20), .b(output_6_5), .y(output_5_20));
wire output_7_20, output_7_5, output_6_20;
mixer gate_output_6_20(.a(output_7_20), .b(output_7_5), .y(output_6_20));
wire output_8_20, output_8_5, output_7_20;
mixer gate_output_7_20(.a(output_8_20), .b(output_8_5), .y(output_7_20));
wire output_9_20, output_9_5, output_8_20;
mixer gate_output_8_20(.a(output_9_20), .b(output_9_5), .y(output_8_20));
wire output_10_20, output_10_5, output_9_20;
mixer gate_output_9_20(.a(output_10_20), .b(output_10_5), .y(output_9_20));
wire output_11_20, output_11_5, output_10_20;
mixer gate_output_10_20(.a(output_11_20), .b(output_11_5), .y(output_10_20));
wire output_12_20, output_12_5, output_11_20;
mixer gate_output_11_20(.a(output_12_20), .b(output_12_5), .y(output_11_20));
wire output_13_20, output_13_5, output_12_20;
mixer gate_output_12_20(.a(output_13_20), .b(output_13_5), .y(output_12_20));
wire output_14_20, output_14_5, output_13_20;
mixer gate_output_13_20(.a(output_14_20), .b(output_14_5), .y(output_13_20));
wire output_15_20, output_15_5, output_14_20;
mixer gate_output_14_20(.a(output_15_20), .b(output_15_5), .y(output_14_20));
wire output_16_20, output_16_5, output_15_20;
mixer gate_output_15_20(.a(output_16_20), .b(output_16_5), .y(output_15_20));
wire output_1_21, output_1_6, output_0_21;
mixer gate_output_0_21(.a(output_1_21), .b(output_1_6), .y(output_0_21));
wire output_2_21, output_2_6, output_1_21;
mixer gate_output_1_21(.a(output_2_21), .b(output_2_6), .y(output_1_21));
wire output_3_21, output_3_6, output_2_21;
mixer gate_output_2_21(.a(output_3_21), .b(output_3_6), .y(output_2_21));
wire output_4_21, output_4_6, output_3_21;
mixer gate_output_3_21(.a(output_4_21), .b(output_4_6), .y(output_3_21));
wire output_5_21, output_5_6, output_4_21;
mixer gate_output_4_21(.a(output_5_21), .b(output_5_6), .y(output_4_21));
wire output_6_21, output_6_6, output_5_21;
mixer gate_output_5_21(.a(output_6_21), .b(output_6_6), .y(output_5_21));
wire output_7_21, output_7_6, output_6_21;
mixer gate_output_6_21(.a(output_7_21), .b(output_7_6), .y(output_6_21));
wire output_8_21, output_8_6, output_7_21;
mixer gate_output_7_21(.a(output_8_21), .b(output_8_6), .y(output_7_21));
wire output_9_21, output_9_6, output_8_21;
mixer gate_output_8_21(.a(output_9_21), .b(output_9_6), .y(output_8_21));
wire output_10_21, output_10_6, output_9_21;
mixer gate_output_9_21(.a(output_10_21), .b(output_10_6), .y(output_9_21));
wire output_11_21, output_11_6, output_10_21;
mixer gate_output_10_21(.a(output_11_21), .b(output_11_6), .y(output_10_21));
wire output_12_21, output_12_6, output_11_21;
mixer gate_output_11_21(.a(output_12_21), .b(output_12_6), .y(output_11_21));
wire output_13_21, output_13_6, output_12_21;
mixer gate_output_12_21(.a(output_13_21), .b(output_13_6), .y(output_12_21));
wire output_14_21, output_14_6, output_13_21;
mixer gate_output_13_21(.a(output_14_21), .b(output_14_6), .y(output_13_21));
wire output_15_21, output_15_6, output_14_21;
mixer gate_output_14_21(.a(output_15_21), .b(output_15_6), .y(output_14_21));
wire output_16_21, output_16_6, output_15_21;
mixer gate_output_15_21(.a(output_16_21), .b(output_16_6), .y(output_15_21));
wire output_1_22, output_1_7, output_0_22;
mixer gate_output_0_22(.a(output_1_22), .b(output_1_7), .y(output_0_22));
wire output_2_22, output_2_7, output_1_22;
mixer gate_output_1_22(.a(output_2_22), .b(output_2_7), .y(output_1_22));
wire output_3_22, output_3_7, output_2_22;
mixer gate_output_2_22(.a(output_3_22), .b(output_3_7), .y(output_2_22));
wire output_4_22, output_4_7, output_3_22;
mixer gate_output_3_22(.a(output_4_22), .b(output_4_7), .y(output_3_22));
wire output_5_22, output_5_7, output_4_22;
mixer gate_output_4_22(.a(output_5_22), .b(output_5_7), .y(output_4_22));
wire output_6_22, output_6_7, output_5_22;
mixer gate_output_5_22(.a(output_6_22), .b(output_6_7), .y(output_5_22));
wire output_7_22, output_7_7, output_6_22;
mixer gate_output_6_22(.a(output_7_22), .b(output_7_7), .y(output_6_22));
wire output_8_22, output_8_7, output_7_22;
mixer gate_output_7_22(.a(output_8_22), .b(output_8_7), .y(output_7_22));
wire output_9_22, output_9_7, output_8_22;
mixer gate_output_8_22(.a(output_9_22), .b(output_9_7), .y(output_8_22));
wire output_10_22, output_10_7, output_9_22;
mixer gate_output_9_22(.a(output_10_22), .b(output_10_7), .y(output_9_22));
wire output_11_22, output_11_7, output_10_22;
mixer gate_output_10_22(.a(output_11_22), .b(output_11_7), .y(output_10_22));
wire output_12_22, output_12_7, output_11_22;
mixer gate_output_11_22(.a(output_12_22), .b(output_12_7), .y(output_11_22));
wire output_13_22, output_13_7, output_12_22;
mixer gate_output_12_22(.a(output_13_22), .b(output_13_7), .y(output_12_22));
wire output_14_22, output_14_7, output_13_22;
mixer gate_output_13_22(.a(output_14_22), .b(output_14_7), .y(output_13_22));
wire output_15_22, output_15_7, output_14_22;
mixer gate_output_14_22(.a(output_15_22), .b(output_15_7), .y(output_14_22));
wire output_16_22, output_16_7, output_15_22;
mixer gate_output_15_22(.a(output_16_22), .b(output_16_7), .y(output_15_22));
wire output_1_23, output_1_8, output_0_23;
mixer gate_output_0_23(.a(output_1_23), .b(output_1_8), .y(output_0_23));
wire output_2_23, output_2_8, output_1_23;
mixer gate_output_1_23(.a(output_2_23), .b(output_2_8), .y(output_1_23));
wire output_3_23, output_3_8, output_2_23;
mixer gate_output_2_23(.a(output_3_23), .b(output_3_8), .y(output_2_23));
wire output_4_23, output_4_8, output_3_23;
mixer gate_output_3_23(.a(output_4_23), .b(output_4_8), .y(output_3_23));
wire output_5_23, output_5_8, output_4_23;
mixer gate_output_4_23(.a(output_5_23), .b(output_5_8), .y(output_4_23));
wire output_6_23, output_6_8, output_5_23;
mixer gate_output_5_23(.a(output_6_23), .b(output_6_8), .y(output_5_23));
wire output_7_23, output_7_8, output_6_23;
mixer gate_output_6_23(.a(output_7_23), .b(output_7_8), .y(output_6_23));
wire output_8_23, output_8_8, output_7_23;
mixer gate_output_7_23(.a(output_8_23), .b(output_8_8), .y(output_7_23));
wire output_9_23, output_9_8, output_8_23;
mixer gate_output_8_23(.a(output_9_23), .b(output_9_8), .y(output_8_23));
wire output_10_23, output_10_8, output_9_23;
mixer gate_output_9_23(.a(output_10_23), .b(output_10_8), .y(output_9_23));
wire output_11_23, output_11_8, output_10_23;
mixer gate_output_10_23(.a(output_11_23), .b(output_11_8), .y(output_10_23));
wire output_12_23, output_12_8, output_11_23;
mixer gate_output_11_23(.a(output_12_23), .b(output_12_8), .y(output_11_23));
wire output_13_23, output_13_8, output_12_23;
mixer gate_output_12_23(.a(output_13_23), .b(output_13_8), .y(output_12_23));
wire output_14_23, output_14_8, output_13_23;
mixer gate_output_13_23(.a(output_14_23), .b(output_14_8), .y(output_13_23));
wire output_15_23, output_15_8, output_14_23;
mixer gate_output_14_23(.a(output_15_23), .b(output_15_8), .y(output_14_23));
wire output_16_23, output_16_8, output_15_23;
mixer gate_output_15_23(.a(output_16_23), .b(output_16_8), .y(output_15_23));
wire output_1_24, output_1_9, output_0_24;
mixer gate_output_0_24(.a(output_1_24), .b(output_1_9), .y(output_0_24));
wire output_2_24, output_2_9, output_1_24;
mixer gate_output_1_24(.a(output_2_24), .b(output_2_9), .y(output_1_24));
wire output_3_24, output_3_9, output_2_24;
mixer gate_output_2_24(.a(output_3_24), .b(output_3_9), .y(output_2_24));
wire output_4_24, output_4_9, output_3_24;
mixer gate_output_3_24(.a(output_4_24), .b(output_4_9), .y(output_3_24));
wire output_5_24, output_5_9, output_4_24;
mixer gate_output_4_24(.a(output_5_24), .b(output_5_9), .y(output_4_24));
wire output_6_24, output_6_9, output_5_24;
mixer gate_output_5_24(.a(output_6_24), .b(output_6_9), .y(output_5_24));
wire output_7_24, output_7_9, output_6_24;
mixer gate_output_6_24(.a(output_7_24), .b(output_7_9), .y(output_6_24));
wire output_8_24, output_8_9, output_7_24;
mixer gate_output_7_24(.a(output_8_24), .b(output_8_9), .y(output_7_24));
wire output_9_24, output_9_9, output_8_24;
mixer gate_output_8_24(.a(output_9_24), .b(output_9_9), .y(output_8_24));
wire output_10_24, output_10_9, output_9_24;
mixer gate_output_9_24(.a(output_10_24), .b(output_10_9), .y(output_9_24));
wire output_11_24, output_11_9, output_10_24;
mixer gate_output_10_24(.a(output_11_24), .b(output_11_9), .y(output_10_24));
wire output_12_24, output_12_9, output_11_24;
mixer gate_output_11_24(.a(output_12_24), .b(output_12_9), .y(output_11_24));
wire output_13_24, output_13_9, output_12_24;
mixer gate_output_12_24(.a(output_13_24), .b(output_13_9), .y(output_12_24));
wire output_14_24, output_14_9, output_13_24;
mixer gate_output_13_24(.a(output_14_24), .b(output_14_9), .y(output_13_24));
wire output_15_24, output_15_9, output_14_24;
mixer gate_output_14_24(.a(output_15_24), .b(output_15_9), .y(output_14_24));
wire output_16_24, output_16_9, output_15_24;
mixer gate_output_15_24(.a(output_16_24), .b(output_16_9), .y(output_15_24));
wire output_1_25, output_1_10, output_0_25;
mixer gate_output_0_25(.a(output_1_25), .b(output_1_10), .y(output_0_25));
wire output_2_25, output_2_10, output_1_25;
mixer gate_output_1_25(.a(output_2_25), .b(output_2_10), .y(output_1_25));
wire output_3_25, output_3_10, output_2_25;
mixer gate_output_2_25(.a(output_3_25), .b(output_3_10), .y(output_2_25));
wire output_4_25, output_4_10, output_3_25;
mixer gate_output_3_25(.a(output_4_25), .b(output_4_10), .y(output_3_25));
wire output_5_25, output_5_10, output_4_25;
mixer gate_output_4_25(.a(output_5_25), .b(output_5_10), .y(output_4_25));
wire output_6_25, output_6_10, output_5_25;
mixer gate_output_5_25(.a(output_6_25), .b(output_6_10), .y(output_5_25));
wire output_7_25, output_7_10, output_6_25;
mixer gate_output_6_25(.a(output_7_25), .b(output_7_10), .y(output_6_25));
wire output_8_25, output_8_10, output_7_25;
mixer gate_output_7_25(.a(output_8_25), .b(output_8_10), .y(output_7_25));
wire output_9_25, output_9_10, output_8_25;
mixer gate_output_8_25(.a(output_9_25), .b(output_9_10), .y(output_8_25));
wire output_10_25, output_10_10, output_9_25;
mixer gate_output_9_25(.a(output_10_25), .b(output_10_10), .y(output_9_25));
wire output_11_25, output_11_10, output_10_25;
mixer gate_output_10_25(.a(output_11_25), .b(output_11_10), .y(output_10_25));
wire output_12_25, output_12_10, output_11_25;
mixer gate_output_11_25(.a(output_12_25), .b(output_12_10), .y(output_11_25));
wire output_13_25, output_13_10, output_12_25;
mixer gate_output_12_25(.a(output_13_25), .b(output_13_10), .y(output_12_25));
wire output_14_25, output_14_10, output_13_25;
mixer gate_output_13_25(.a(output_14_25), .b(output_14_10), .y(output_13_25));
wire output_15_25, output_15_10, output_14_25;
mixer gate_output_14_25(.a(output_15_25), .b(output_15_10), .y(output_14_25));
wire output_16_25, output_16_10, output_15_25;
mixer gate_output_15_25(.a(output_16_25), .b(output_16_10), .y(output_15_25));
wire output_1_26, output_1_11, output_0_26;
mixer gate_output_0_26(.a(output_1_26), .b(output_1_11), .y(output_0_26));
wire output_2_26, output_2_11, output_1_26;
mixer gate_output_1_26(.a(output_2_26), .b(output_2_11), .y(output_1_26));
wire output_3_26, output_3_11, output_2_26;
mixer gate_output_2_26(.a(output_3_26), .b(output_3_11), .y(output_2_26));
wire output_4_26, output_4_11, output_3_26;
mixer gate_output_3_26(.a(output_4_26), .b(output_4_11), .y(output_3_26));
wire output_5_26, output_5_11, output_4_26;
mixer gate_output_4_26(.a(output_5_26), .b(output_5_11), .y(output_4_26));
wire output_6_26, output_6_11, output_5_26;
mixer gate_output_5_26(.a(output_6_26), .b(output_6_11), .y(output_5_26));
wire output_7_26, output_7_11, output_6_26;
mixer gate_output_6_26(.a(output_7_26), .b(output_7_11), .y(output_6_26));
wire output_8_26, output_8_11, output_7_26;
mixer gate_output_7_26(.a(output_8_26), .b(output_8_11), .y(output_7_26));
wire output_9_26, output_9_11, output_8_26;
mixer gate_output_8_26(.a(output_9_26), .b(output_9_11), .y(output_8_26));
wire output_10_26, output_10_11, output_9_26;
mixer gate_output_9_26(.a(output_10_26), .b(output_10_11), .y(output_9_26));
wire output_11_26, output_11_11, output_10_26;
mixer gate_output_10_26(.a(output_11_26), .b(output_11_11), .y(output_10_26));
wire output_12_26, output_12_11, output_11_26;
mixer gate_output_11_26(.a(output_12_26), .b(output_12_11), .y(output_11_26));
wire output_13_26, output_13_11, output_12_26;
mixer gate_output_12_26(.a(output_13_26), .b(output_13_11), .y(output_12_26));
wire output_14_26, output_14_11, output_13_26;
mixer gate_output_13_26(.a(output_14_26), .b(output_14_11), .y(output_13_26));
wire output_15_26, output_15_11, output_14_26;
mixer gate_output_14_26(.a(output_15_26), .b(output_15_11), .y(output_14_26));
wire output_16_26, output_16_11, output_15_26;
mixer gate_output_15_26(.a(output_16_26), .b(output_16_11), .y(output_15_26));
wire output_1_27, output_1_12, output_0_27;
mixer gate_output_0_27(.a(output_1_27), .b(output_1_12), .y(output_0_27));
wire output_2_27, output_2_12, output_1_27;
mixer gate_output_1_27(.a(output_2_27), .b(output_2_12), .y(output_1_27));
wire output_3_27, output_3_12, output_2_27;
mixer gate_output_2_27(.a(output_3_27), .b(output_3_12), .y(output_2_27));
wire output_4_27, output_4_12, output_3_27;
mixer gate_output_3_27(.a(output_4_27), .b(output_4_12), .y(output_3_27));
wire output_5_27, output_5_12, output_4_27;
mixer gate_output_4_27(.a(output_5_27), .b(output_5_12), .y(output_4_27));
wire output_6_27, output_6_12, output_5_27;
mixer gate_output_5_27(.a(output_6_27), .b(output_6_12), .y(output_5_27));
wire output_7_27, output_7_12, output_6_27;
mixer gate_output_6_27(.a(output_7_27), .b(output_7_12), .y(output_6_27));
wire output_8_27, output_8_12, output_7_27;
mixer gate_output_7_27(.a(output_8_27), .b(output_8_12), .y(output_7_27));
wire output_9_27, output_9_12, output_8_27;
mixer gate_output_8_27(.a(output_9_27), .b(output_9_12), .y(output_8_27));
wire output_10_27, output_10_12, output_9_27;
mixer gate_output_9_27(.a(output_10_27), .b(output_10_12), .y(output_9_27));
wire output_11_27, output_11_12, output_10_27;
mixer gate_output_10_27(.a(output_11_27), .b(output_11_12), .y(output_10_27));
wire output_12_27, output_12_12, output_11_27;
mixer gate_output_11_27(.a(output_12_27), .b(output_12_12), .y(output_11_27));
wire output_13_27, output_13_12, output_12_27;
mixer gate_output_12_27(.a(output_13_27), .b(output_13_12), .y(output_12_27));
wire output_14_27, output_14_12, output_13_27;
mixer gate_output_13_27(.a(output_14_27), .b(output_14_12), .y(output_13_27));
wire output_15_27, output_15_12, output_14_27;
mixer gate_output_14_27(.a(output_15_27), .b(output_15_12), .y(output_14_27));
wire output_16_27, output_16_12, output_15_27;
mixer gate_output_15_27(.a(output_16_27), .b(output_16_12), .y(output_15_27));
wire output_1_28, output_1_13, output_0_28;
mixer gate_output_0_28(.a(output_1_28), .b(output_1_13), .y(output_0_28));
wire output_2_28, output_2_13, output_1_28;
mixer gate_output_1_28(.a(output_2_28), .b(output_2_13), .y(output_1_28));
wire output_3_28, output_3_13, output_2_28;
mixer gate_output_2_28(.a(output_3_28), .b(output_3_13), .y(output_2_28));
wire output_4_28, output_4_13, output_3_28;
mixer gate_output_3_28(.a(output_4_28), .b(output_4_13), .y(output_3_28));
wire output_5_28, output_5_13, output_4_28;
mixer gate_output_4_28(.a(output_5_28), .b(output_5_13), .y(output_4_28));
wire output_6_28, output_6_13, output_5_28;
mixer gate_output_5_28(.a(output_6_28), .b(output_6_13), .y(output_5_28));
wire output_7_28, output_7_13, output_6_28;
mixer gate_output_6_28(.a(output_7_28), .b(output_7_13), .y(output_6_28));
wire output_8_28, output_8_13, output_7_28;
mixer gate_output_7_28(.a(output_8_28), .b(output_8_13), .y(output_7_28));
wire output_9_28, output_9_13, output_8_28;
mixer gate_output_8_28(.a(output_9_28), .b(output_9_13), .y(output_8_28));
wire output_10_28, output_10_13, output_9_28;
mixer gate_output_9_28(.a(output_10_28), .b(output_10_13), .y(output_9_28));
wire output_11_28, output_11_13, output_10_28;
mixer gate_output_10_28(.a(output_11_28), .b(output_11_13), .y(output_10_28));
wire output_12_28, output_12_13, output_11_28;
mixer gate_output_11_28(.a(output_12_28), .b(output_12_13), .y(output_11_28));
wire output_13_28, output_13_13, output_12_28;
mixer gate_output_12_28(.a(output_13_28), .b(output_13_13), .y(output_12_28));
wire output_14_28, output_14_13, output_13_28;
mixer gate_output_13_28(.a(output_14_28), .b(output_14_13), .y(output_13_28));
wire output_15_28, output_15_13, output_14_28;
mixer gate_output_14_28(.a(output_15_28), .b(output_15_13), .y(output_14_28));
wire output_16_28, output_16_13, output_15_28;
mixer gate_output_15_28(.a(output_16_28), .b(output_16_13), .y(output_15_28));
wire output_1_29, output_1_14, output_0_29;
mixer gate_output_0_29(.a(output_1_29), .b(output_1_14), .y(output_0_29));
wire output_2_29, output_2_14, output_1_29;
mixer gate_output_1_29(.a(output_2_29), .b(output_2_14), .y(output_1_29));
wire output_3_29, output_3_14, output_2_29;
mixer gate_output_2_29(.a(output_3_29), .b(output_3_14), .y(output_2_29));
wire output_4_29, output_4_14, output_3_29;
mixer gate_output_3_29(.a(output_4_29), .b(output_4_14), .y(output_3_29));
wire output_5_29, output_5_14, output_4_29;
mixer gate_output_4_29(.a(output_5_29), .b(output_5_14), .y(output_4_29));
wire output_6_29, output_6_14, output_5_29;
mixer gate_output_5_29(.a(output_6_29), .b(output_6_14), .y(output_5_29));
wire output_7_29, output_7_14, output_6_29;
mixer gate_output_6_29(.a(output_7_29), .b(output_7_14), .y(output_6_29));
wire output_8_29, output_8_14, output_7_29;
mixer gate_output_7_29(.a(output_8_29), .b(output_8_14), .y(output_7_29));
wire output_9_29, output_9_14, output_8_29;
mixer gate_output_8_29(.a(output_9_29), .b(output_9_14), .y(output_8_29));
wire output_10_29, output_10_14, output_9_29;
mixer gate_output_9_29(.a(output_10_29), .b(output_10_14), .y(output_9_29));
wire output_11_29, output_11_14, output_10_29;
mixer gate_output_10_29(.a(output_11_29), .b(output_11_14), .y(output_10_29));
wire output_12_29, output_12_14, output_11_29;
mixer gate_output_11_29(.a(output_12_29), .b(output_12_14), .y(output_11_29));
wire output_13_29, output_13_14, output_12_29;
mixer gate_output_12_29(.a(output_13_29), .b(output_13_14), .y(output_12_29));
wire output_14_29, output_14_14, output_13_29;
mixer gate_output_13_29(.a(output_14_29), .b(output_14_14), .y(output_13_29));
wire output_15_29, output_15_14, output_14_29;
mixer gate_output_14_29(.a(output_15_29), .b(output_15_14), .y(output_14_29));
wire output_16_29, output_16_14, output_15_29;
mixer gate_output_15_29(.a(output_16_29), .b(output_16_14), .y(output_15_29));
wire output_1_30, output_1_15, output_0_30;
mixer gate_output_0_30(.a(output_1_30), .b(output_1_15), .y(output_0_30));
wire output_2_30, output_2_15, output_1_30;
mixer gate_output_1_30(.a(output_2_30), .b(output_2_15), .y(output_1_30));
wire output_3_30, output_3_15, output_2_30;
mixer gate_output_2_30(.a(output_3_30), .b(output_3_15), .y(output_2_30));
wire output_4_30, output_4_15, output_3_30;
mixer gate_output_3_30(.a(output_4_30), .b(output_4_15), .y(output_3_30));
wire output_5_30, output_5_15, output_4_30;
mixer gate_output_4_30(.a(output_5_30), .b(output_5_15), .y(output_4_30));
wire output_6_30, output_6_15, output_5_30;
mixer gate_output_5_30(.a(output_6_30), .b(output_6_15), .y(output_5_30));
wire output_7_30, output_7_15, output_6_30;
mixer gate_output_6_30(.a(output_7_30), .b(output_7_15), .y(output_6_30));
wire output_8_30, output_8_15, output_7_30;
mixer gate_output_7_30(.a(output_8_30), .b(output_8_15), .y(output_7_30));
wire output_9_30, output_9_15, output_8_30;
mixer gate_output_8_30(.a(output_9_30), .b(output_9_15), .y(output_8_30));
wire output_10_30, output_10_15, output_9_30;
mixer gate_output_9_30(.a(output_10_30), .b(output_10_15), .y(output_9_30));
wire output_11_30, output_11_15, output_10_30;
mixer gate_output_10_30(.a(output_11_30), .b(output_11_15), .y(output_10_30));
wire output_12_30, output_12_15, output_11_30;
mixer gate_output_11_30(.a(output_12_30), .b(output_12_15), .y(output_11_30));
wire output_13_30, output_13_15, output_12_30;
mixer gate_output_12_30(.a(output_13_30), .b(output_13_15), .y(output_12_30));
wire output_14_30, output_14_15, output_13_30;
mixer gate_output_13_30(.a(output_14_30), .b(output_14_15), .y(output_13_30));
wire output_15_30, output_15_15, output_14_30;
mixer gate_output_14_30(.a(output_15_30), .b(output_15_15), .y(output_14_30));
wire output_16_30, output_16_15, output_15_30;
mixer gate_output_15_30(.a(output_16_30), .b(output_16_15), .y(output_15_30));
wire output_1_31, output_1_0, output_0_31;
mixer gate_output_0_31(.a(output_1_31), .b(output_1_0), .y(output_0_31));
wire output_2_31, output_2_0, output_1_31;
mixer gate_output_1_31(.a(output_2_31), .b(output_2_0), .y(output_1_31));
wire output_3_31, output_3_0, output_2_31;
mixer gate_output_2_31(.a(output_3_31), .b(output_3_0), .y(output_2_31));
wire output_4_31, output_4_0, output_3_31;
mixer gate_output_3_31(.a(output_4_31), .b(output_4_0), .y(output_3_31));
wire output_5_31, output_5_0, output_4_31;
mixer gate_output_4_31(.a(output_5_31), .b(output_5_0), .y(output_4_31));
wire output_6_31, output_6_0, output_5_31;
mixer gate_output_5_31(.a(output_6_31), .b(output_6_0), .y(output_5_31));
wire output_7_31, output_7_0, output_6_31;
mixer gate_output_6_31(.a(output_7_31), .b(output_7_0), .y(output_6_31));
wire output_8_31, output_8_0, output_7_31;
mixer gate_output_7_31(.a(output_8_31), .b(output_8_0), .y(output_7_31));
wire output_9_31, output_9_0, output_8_31;
mixer gate_output_8_31(.a(output_9_31), .b(output_9_0), .y(output_8_31));
wire output_10_31, output_10_0, output_9_31;
mixer gate_output_9_31(.a(output_10_31), .b(output_10_0), .y(output_9_31));
wire output_11_31, output_11_0, output_10_31;
mixer gate_output_10_31(.a(output_11_31), .b(output_11_0), .y(output_10_31));
wire output_12_31, output_12_0, output_11_31;
mixer gate_output_11_31(.a(output_12_31), .b(output_12_0), .y(output_11_31));
wire output_13_31, output_13_0, output_12_31;
mixer gate_output_12_31(.a(output_13_31), .b(output_13_0), .y(output_12_31));
wire output_14_31, output_14_0, output_13_31;
mixer gate_output_13_31(.a(output_14_31), .b(output_14_0), .y(output_13_31));
wire output_15_31, output_15_0, output_14_31;
mixer gate_output_14_31(.a(output_15_31), .b(output_15_0), .y(output_14_31));
wire output_16_31, output_16_0, output_15_31;
mixer gate_output_15_31(.a(output_16_31), .b(output_16_0), .y(output_15_31));
wire output_1_32, output_1_1, output_0_32;
mixer gate_output_0_32(.a(output_1_32), .b(output_1_1), .y(output_0_32));
wire output_2_32, output_2_1, output_1_32;
mixer gate_output_1_32(.a(output_2_32), .b(output_2_1), .y(output_1_32));
wire output_3_32, output_3_1, output_2_32;
mixer gate_output_2_32(.a(output_3_32), .b(output_3_1), .y(output_2_32));
wire output_4_32, output_4_1, output_3_32;
mixer gate_output_3_32(.a(output_4_32), .b(output_4_1), .y(output_3_32));
wire output_5_32, output_5_1, output_4_32;
mixer gate_output_4_32(.a(output_5_32), .b(output_5_1), .y(output_4_32));
wire output_6_32, output_6_1, output_5_32;
mixer gate_output_5_32(.a(output_6_32), .b(output_6_1), .y(output_5_32));
wire output_7_32, output_7_1, output_6_32;
mixer gate_output_6_32(.a(output_7_32), .b(output_7_1), .y(output_6_32));
wire output_8_32, output_8_1, output_7_32;
mixer gate_output_7_32(.a(output_8_32), .b(output_8_1), .y(output_7_32));
wire output_9_32, output_9_1, output_8_32;
mixer gate_output_8_32(.a(output_9_32), .b(output_9_1), .y(output_8_32));
wire output_10_32, output_10_1, output_9_32;
mixer gate_output_9_32(.a(output_10_32), .b(output_10_1), .y(output_9_32));
wire output_11_32, output_11_1, output_10_32;
mixer gate_output_10_32(.a(output_11_32), .b(output_11_1), .y(output_10_32));
wire output_12_32, output_12_1, output_11_32;
mixer gate_output_11_32(.a(output_12_32), .b(output_12_1), .y(output_11_32));
wire output_13_32, output_13_1, output_12_32;
mixer gate_output_12_32(.a(output_13_32), .b(output_13_1), .y(output_12_32));
wire output_14_32, output_14_1, output_13_32;
mixer gate_output_13_32(.a(output_14_32), .b(output_14_1), .y(output_13_32));
wire output_15_32, output_15_1, output_14_32;
mixer gate_output_14_32(.a(output_15_32), .b(output_15_1), .y(output_14_32));
wire output_16_32, output_16_1, output_15_32;
mixer gate_output_15_32(.a(output_16_32), .b(output_16_1), .y(output_15_32));
wire output_1_33, output_1_2, output_0_33;
mixer gate_output_0_33(.a(output_1_33), .b(output_1_2), .y(output_0_33));
wire output_2_33, output_2_2, output_1_33;
mixer gate_output_1_33(.a(output_2_33), .b(output_2_2), .y(output_1_33));
wire output_3_33, output_3_2, output_2_33;
mixer gate_output_2_33(.a(output_3_33), .b(output_3_2), .y(output_2_33));
wire output_4_33, output_4_2, output_3_33;
mixer gate_output_3_33(.a(output_4_33), .b(output_4_2), .y(output_3_33));
wire output_5_33, output_5_2, output_4_33;
mixer gate_output_4_33(.a(output_5_33), .b(output_5_2), .y(output_4_33));
wire output_6_33, output_6_2, output_5_33;
mixer gate_output_5_33(.a(output_6_33), .b(output_6_2), .y(output_5_33));
wire output_7_33, output_7_2, output_6_33;
mixer gate_output_6_33(.a(output_7_33), .b(output_7_2), .y(output_6_33));
wire output_8_33, output_8_2, output_7_33;
mixer gate_output_7_33(.a(output_8_33), .b(output_8_2), .y(output_7_33));
wire output_9_33, output_9_2, output_8_33;
mixer gate_output_8_33(.a(output_9_33), .b(output_9_2), .y(output_8_33));
wire output_10_33, output_10_2, output_9_33;
mixer gate_output_9_33(.a(output_10_33), .b(output_10_2), .y(output_9_33));
wire output_11_33, output_11_2, output_10_33;
mixer gate_output_10_33(.a(output_11_33), .b(output_11_2), .y(output_10_33));
wire output_12_33, output_12_2, output_11_33;
mixer gate_output_11_33(.a(output_12_33), .b(output_12_2), .y(output_11_33));
wire output_13_33, output_13_2, output_12_33;
mixer gate_output_12_33(.a(output_13_33), .b(output_13_2), .y(output_12_33));
wire output_14_33, output_14_2, output_13_33;
mixer gate_output_13_33(.a(output_14_33), .b(output_14_2), .y(output_13_33));
wire output_15_33, output_15_2, output_14_33;
mixer gate_output_14_33(.a(output_15_33), .b(output_15_2), .y(output_14_33));
wire output_16_33, output_16_2, output_15_33;
mixer gate_output_15_33(.a(output_16_33), .b(output_16_2), .y(output_15_33));
wire output_1_34, output_1_3, output_0_34;
mixer gate_output_0_34(.a(output_1_34), .b(output_1_3), .y(output_0_34));
wire output_2_34, output_2_3, output_1_34;
mixer gate_output_1_34(.a(output_2_34), .b(output_2_3), .y(output_1_34));
wire output_3_34, output_3_3, output_2_34;
mixer gate_output_2_34(.a(output_3_34), .b(output_3_3), .y(output_2_34));
wire output_4_34, output_4_3, output_3_34;
mixer gate_output_3_34(.a(output_4_34), .b(output_4_3), .y(output_3_34));
wire output_5_34, output_5_3, output_4_34;
mixer gate_output_4_34(.a(output_5_34), .b(output_5_3), .y(output_4_34));
wire output_6_34, output_6_3, output_5_34;
mixer gate_output_5_34(.a(output_6_34), .b(output_6_3), .y(output_5_34));
wire output_7_34, output_7_3, output_6_34;
mixer gate_output_6_34(.a(output_7_34), .b(output_7_3), .y(output_6_34));
wire output_8_34, output_8_3, output_7_34;
mixer gate_output_7_34(.a(output_8_34), .b(output_8_3), .y(output_7_34));
wire output_9_34, output_9_3, output_8_34;
mixer gate_output_8_34(.a(output_9_34), .b(output_9_3), .y(output_8_34));
wire output_10_34, output_10_3, output_9_34;
mixer gate_output_9_34(.a(output_10_34), .b(output_10_3), .y(output_9_34));
wire output_11_34, output_11_3, output_10_34;
mixer gate_output_10_34(.a(output_11_34), .b(output_11_3), .y(output_10_34));
wire output_12_34, output_12_3, output_11_34;
mixer gate_output_11_34(.a(output_12_34), .b(output_12_3), .y(output_11_34));
wire output_13_34, output_13_3, output_12_34;
mixer gate_output_12_34(.a(output_13_34), .b(output_13_3), .y(output_12_34));
wire output_14_34, output_14_3, output_13_34;
mixer gate_output_13_34(.a(output_14_34), .b(output_14_3), .y(output_13_34));
wire output_15_34, output_15_3, output_14_34;
mixer gate_output_14_34(.a(output_15_34), .b(output_15_3), .y(output_14_34));
wire output_16_34, output_16_3, output_15_34;
mixer gate_output_15_34(.a(output_16_34), .b(output_16_3), .y(output_15_34));
wire output_1_35, output_1_4, output_0_35;
mixer gate_output_0_35(.a(output_1_35), .b(output_1_4), .y(output_0_35));
wire output_2_35, output_2_4, output_1_35;
mixer gate_output_1_35(.a(output_2_35), .b(output_2_4), .y(output_1_35));
wire output_3_35, output_3_4, output_2_35;
mixer gate_output_2_35(.a(output_3_35), .b(output_3_4), .y(output_2_35));
wire output_4_35, output_4_4, output_3_35;
mixer gate_output_3_35(.a(output_4_35), .b(output_4_4), .y(output_3_35));
wire output_5_35, output_5_4, output_4_35;
mixer gate_output_4_35(.a(output_5_35), .b(output_5_4), .y(output_4_35));
wire output_6_35, output_6_4, output_5_35;
mixer gate_output_5_35(.a(output_6_35), .b(output_6_4), .y(output_5_35));
wire output_7_35, output_7_4, output_6_35;
mixer gate_output_6_35(.a(output_7_35), .b(output_7_4), .y(output_6_35));
wire output_8_35, output_8_4, output_7_35;
mixer gate_output_7_35(.a(output_8_35), .b(output_8_4), .y(output_7_35));
wire output_9_35, output_9_4, output_8_35;
mixer gate_output_8_35(.a(output_9_35), .b(output_9_4), .y(output_8_35));
wire output_10_35, output_10_4, output_9_35;
mixer gate_output_9_35(.a(output_10_35), .b(output_10_4), .y(output_9_35));
wire output_11_35, output_11_4, output_10_35;
mixer gate_output_10_35(.a(output_11_35), .b(output_11_4), .y(output_10_35));
wire output_12_35, output_12_4, output_11_35;
mixer gate_output_11_35(.a(output_12_35), .b(output_12_4), .y(output_11_35));
wire output_13_35, output_13_4, output_12_35;
mixer gate_output_12_35(.a(output_13_35), .b(output_13_4), .y(output_12_35));
wire output_14_35, output_14_4, output_13_35;
mixer gate_output_13_35(.a(output_14_35), .b(output_14_4), .y(output_13_35));
wire output_15_35, output_15_4, output_14_35;
mixer gate_output_14_35(.a(output_15_35), .b(output_15_4), .y(output_14_35));
wire output_16_35, output_16_4, output_15_35;
mixer gate_output_15_35(.a(output_16_35), .b(output_16_4), .y(output_15_35));
wire output_1_36, output_1_5, output_0_36;
mixer gate_output_0_36(.a(output_1_36), .b(output_1_5), .y(output_0_36));
wire output_2_36, output_2_5, output_1_36;
mixer gate_output_1_36(.a(output_2_36), .b(output_2_5), .y(output_1_36));
wire output_3_36, output_3_5, output_2_36;
mixer gate_output_2_36(.a(output_3_36), .b(output_3_5), .y(output_2_36));
wire output_4_36, output_4_5, output_3_36;
mixer gate_output_3_36(.a(output_4_36), .b(output_4_5), .y(output_3_36));
wire output_5_36, output_5_5, output_4_36;
mixer gate_output_4_36(.a(output_5_36), .b(output_5_5), .y(output_4_36));
wire output_6_36, output_6_5, output_5_36;
mixer gate_output_5_36(.a(output_6_36), .b(output_6_5), .y(output_5_36));
wire output_7_36, output_7_5, output_6_36;
mixer gate_output_6_36(.a(output_7_36), .b(output_7_5), .y(output_6_36));
wire output_8_36, output_8_5, output_7_36;
mixer gate_output_7_36(.a(output_8_36), .b(output_8_5), .y(output_7_36));
wire output_9_36, output_9_5, output_8_36;
mixer gate_output_8_36(.a(output_9_36), .b(output_9_5), .y(output_8_36));
wire output_10_36, output_10_5, output_9_36;
mixer gate_output_9_36(.a(output_10_36), .b(output_10_5), .y(output_9_36));
wire output_11_36, output_11_5, output_10_36;
mixer gate_output_10_36(.a(output_11_36), .b(output_11_5), .y(output_10_36));
wire output_12_36, output_12_5, output_11_36;
mixer gate_output_11_36(.a(output_12_36), .b(output_12_5), .y(output_11_36));
wire output_13_36, output_13_5, output_12_36;
mixer gate_output_12_36(.a(output_13_36), .b(output_13_5), .y(output_12_36));
wire output_14_36, output_14_5, output_13_36;
mixer gate_output_13_36(.a(output_14_36), .b(output_14_5), .y(output_13_36));
wire output_15_36, output_15_5, output_14_36;
mixer gate_output_14_36(.a(output_15_36), .b(output_15_5), .y(output_14_36));
wire output_16_36, output_16_5, output_15_36;
mixer gate_output_15_36(.a(output_16_36), .b(output_16_5), .y(output_15_36));
wire output_1_37, output_1_6, output_0_37;
mixer gate_output_0_37(.a(output_1_37), .b(output_1_6), .y(output_0_37));
wire output_2_37, output_2_6, output_1_37;
mixer gate_output_1_37(.a(output_2_37), .b(output_2_6), .y(output_1_37));
wire output_3_37, output_3_6, output_2_37;
mixer gate_output_2_37(.a(output_3_37), .b(output_3_6), .y(output_2_37));
wire output_4_37, output_4_6, output_3_37;
mixer gate_output_3_37(.a(output_4_37), .b(output_4_6), .y(output_3_37));
wire output_5_37, output_5_6, output_4_37;
mixer gate_output_4_37(.a(output_5_37), .b(output_5_6), .y(output_4_37));
wire output_6_37, output_6_6, output_5_37;
mixer gate_output_5_37(.a(output_6_37), .b(output_6_6), .y(output_5_37));
wire output_7_37, output_7_6, output_6_37;
mixer gate_output_6_37(.a(output_7_37), .b(output_7_6), .y(output_6_37));
wire output_8_37, output_8_6, output_7_37;
mixer gate_output_7_37(.a(output_8_37), .b(output_8_6), .y(output_7_37));
wire output_9_37, output_9_6, output_8_37;
mixer gate_output_8_37(.a(output_9_37), .b(output_9_6), .y(output_8_37));
wire output_10_37, output_10_6, output_9_37;
mixer gate_output_9_37(.a(output_10_37), .b(output_10_6), .y(output_9_37));
wire output_11_37, output_11_6, output_10_37;
mixer gate_output_10_37(.a(output_11_37), .b(output_11_6), .y(output_10_37));
wire output_12_37, output_12_6, output_11_37;
mixer gate_output_11_37(.a(output_12_37), .b(output_12_6), .y(output_11_37));
wire output_13_37, output_13_6, output_12_37;
mixer gate_output_12_37(.a(output_13_37), .b(output_13_6), .y(output_12_37));
wire output_14_37, output_14_6, output_13_37;
mixer gate_output_13_37(.a(output_14_37), .b(output_14_6), .y(output_13_37));
wire output_15_37, output_15_6, output_14_37;
mixer gate_output_14_37(.a(output_15_37), .b(output_15_6), .y(output_14_37));
wire output_16_37, output_16_6, output_15_37;
mixer gate_output_15_37(.a(output_16_37), .b(output_16_6), .y(output_15_37));
wire output_1_38, output_1_7, output_0_38;
mixer gate_output_0_38(.a(output_1_38), .b(output_1_7), .y(output_0_38));
wire output_2_38, output_2_7, output_1_38;
mixer gate_output_1_38(.a(output_2_38), .b(output_2_7), .y(output_1_38));
wire output_3_38, output_3_7, output_2_38;
mixer gate_output_2_38(.a(output_3_38), .b(output_3_7), .y(output_2_38));
wire output_4_38, output_4_7, output_3_38;
mixer gate_output_3_38(.a(output_4_38), .b(output_4_7), .y(output_3_38));
wire output_5_38, output_5_7, output_4_38;
mixer gate_output_4_38(.a(output_5_38), .b(output_5_7), .y(output_4_38));
wire output_6_38, output_6_7, output_5_38;
mixer gate_output_5_38(.a(output_6_38), .b(output_6_7), .y(output_5_38));
wire output_7_38, output_7_7, output_6_38;
mixer gate_output_6_38(.a(output_7_38), .b(output_7_7), .y(output_6_38));
wire output_8_38, output_8_7, output_7_38;
mixer gate_output_7_38(.a(output_8_38), .b(output_8_7), .y(output_7_38));
wire output_9_38, output_9_7, output_8_38;
mixer gate_output_8_38(.a(output_9_38), .b(output_9_7), .y(output_8_38));
wire output_10_38, output_10_7, output_9_38;
mixer gate_output_9_38(.a(output_10_38), .b(output_10_7), .y(output_9_38));
wire output_11_38, output_11_7, output_10_38;
mixer gate_output_10_38(.a(output_11_38), .b(output_11_7), .y(output_10_38));
wire output_12_38, output_12_7, output_11_38;
mixer gate_output_11_38(.a(output_12_38), .b(output_12_7), .y(output_11_38));
wire output_13_38, output_13_7, output_12_38;
mixer gate_output_12_38(.a(output_13_38), .b(output_13_7), .y(output_12_38));
wire output_14_38, output_14_7, output_13_38;
mixer gate_output_13_38(.a(output_14_38), .b(output_14_7), .y(output_13_38));
wire output_15_38, output_15_7, output_14_38;
mixer gate_output_14_38(.a(output_15_38), .b(output_15_7), .y(output_14_38));
wire output_16_38, output_16_7, output_15_38;
mixer gate_output_15_38(.a(output_16_38), .b(output_16_7), .y(output_15_38));
wire output_1_39, output_1_8, output_0_39;
mixer gate_output_0_39(.a(output_1_39), .b(output_1_8), .y(output_0_39));
wire output_2_39, output_2_8, output_1_39;
mixer gate_output_1_39(.a(output_2_39), .b(output_2_8), .y(output_1_39));
wire output_3_39, output_3_8, output_2_39;
mixer gate_output_2_39(.a(output_3_39), .b(output_3_8), .y(output_2_39));
wire output_4_39, output_4_8, output_3_39;
mixer gate_output_3_39(.a(output_4_39), .b(output_4_8), .y(output_3_39));
wire output_5_39, output_5_8, output_4_39;
mixer gate_output_4_39(.a(output_5_39), .b(output_5_8), .y(output_4_39));
wire output_6_39, output_6_8, output_5_39;
mixer gate_output_5_39(.a(output_6_39), .b(output_6_8), .y(output_5_39));
wire output_7_39, output_7_8, output_6_39;
mixer gate_output_6_39(.a(output_7_39), .b(output_7_8), .y(output_6_39));
wire output_8_39, output_8_8, output_7_39;
mixer gate_output_7_39(.a(output_8_39), .b(output_8_8), .y(output_7_39));
wire output_9_39, output_9_8, output_8_39;
mixer gate_output_8_39(.a(output_9_39), .b(output_9_8), .y(output_8_39));
wire output_10_39, output_10_8, output_9_39;
mixer gate_output_9_39(.a(output_10_39), .b(output_10_8), .y(output_9_39));
wire output_11_39, output_11_8, output_10_39;
mixer gate_output_10_39(.a(output_11_39), .b(output_11_8), .y(output_10_39));
wire output_12_39, output_12_8, output_11_39;
mixer gate_output_11_39(.a(output_12_39), .b(output_12_8), .y(output_11_39));
wire output_13_39, output_13_8, output_12_39;
mixer gate_output_12_39(.a(output_13_39), .b(output_13_8), .y(output_12_39));
wire output_14_39, output_14_8, output_13_39;
mixer gate_output_13_39(.a(output_14_39), .b(output_14_8), .y(output_13_39));
wire output_15_39, output_15_8, output_14_39;
mixer gate_output_14_39(.a(output_15_39), .b(output_15_8), .y(output_14_39));
wire output_16_39, output_16_8, output_15_39;
mixer gate_output_15_39(.a(output_16_39), .b(output_16_8), .y(output_15_39));
wire output_1_40, output_1_9, output_0_40;
mixer gate_output_0_40(.a(output_1_40), .b(output_1_9), .y(output_0_40));
wire output_2_40, output_2_9, output_1_40;
mixer gate_output_1_40(.a(output_2_40), .b(output_2_9), .y(output_1_40));
wire output_3_40, output_3_9, output_2_40;
mixer gate_output_2_40(.a(output_3_40), .b(output_3_9), .y(output_2_40));
wire output_4_40, output_4_9, output_3_40;
mixer gate_output_3_40(.a(output_4_40), .b(output_4_9), .y(output_3_40));
wire output_5_40, output_5_9, output_4_40;
mixer gate_output_4_40(.a(output_5_40), .b(output_5_9), .y(output_4_40));
wire output_6_40, output_6_9, output_5_40;
mixer gate_output_5_40(.a(output_6_40), .b(output_6_9), .y(output_5_40));
wire output_7_40, output_7_9, output_6_40;
mixer gate_output_6_40(.a(output_7_40), .b(output_7_9), .y(output_6_40));
wire output_8_40, output_8_9, output_7_40;
mixer gate_output_7_40(.a(output_8_40), .b(output_8_9), .y(output_7_40));
wire output_9_40, output_9_9, output_8_40;
mixer gate_output_8_40(.a(output_9_40), .b(output_9_9), .y(output_8_40));
wire output_10_40, output_10_9, output_9_40;
mixer gate_output_9_40(.a(output_10_40), .b(output_10_9), .y(output_9_40));
wire output_11_40, output_11_9, output_10_40;
mixer gate_output_10_40(.a(output_11_40), .b(output_11_9), .y(output_10_40));
wire output_12_40, output_12_9, output_11_40;
mixer gate_output_11_40(.a(output_12_40), .b(output_12_9), .y(output_11_40));
wire output_13_40, output_13_9, output_12_40;
mixer gate_output_12_40(.a(output_13_40), .b(output_13_9), .y(output_12_40));
wire output_14_40, output_14_9, output_13_40;
mixer gate_output_13_40(.a(output_14_40), .b(output_14_9), .y(output_13_40));
wire output_15_40, output_15_9, output_14_40;
mixer gate_output_14_40(.a(output_15_40), .b(output_15_9), .y(output_14_40));
wire output_16_40, output_16_9, output_15_40;
mixer gate_output_15_40(.a(output_16_40), .b(output_16_9), .y(output_15_40));
wire output_1_41, output_1_10, output_0_41;
mixer gate_output_0_41(.a(output_1_41), .b(output_1_10), .y(output_0_41));
wire output_2_41, output_2_10, output_1_41;
mixer gate_output_1_41(.a(output_2_41), .b(output_2_10), .y(output_1_41));
wire output_3_41, output_3_10, output_2_41;
mixer gate_output_2_41(.a(output_3_41), .b(output_3_10), .y(output_2_41));
wire output_4_41, output_4_10, output_3_41;
mixer gate_output_3_41(.a(output_4_41), .b(output_4_10), .y(output_3_41));
wire output_5_41, output_5_10, output_4_41;
mixer gate_output_4_41(.a(output_5_41), .b(output_5_10), .y(output_4_41));
wire output_6_41, output_6_10, output_5_41;
mixer gate_output_5_41(.a(output_6_41), .b(output_6_10), .y(output_5_41));
wire output_7_41, output_7_10, output_6_41;
mixer gate_output_6_41(.a(output_7_41), .b(output_7_10), .y(output_6_41));
wire output_8_41, output_8_10, output_7_41;
mixer gate_output_7_41(.a(output_8_41), .b(output_8_10), .y(output_7_41));
wire output_9_41, output_9_10, output_8_41;
mixer gate_output_8_41(.a(output_9_41), .b(output_9_10), .y(output_8_41));
wire output_10_41, output_10_10, output_9_41;
mixer gate_output_9_41(.a(output_10_41), .b(output_10_10), .y(output_9_41));
wire output_11_41, output_11_10, output_10_41;
mixer gate_output_10_41(.a(output_11_41), .b(output_11_10), .y(output_10_41));
wire output_12_41, output_12_10, output_11_41;
mixer gate_output_11_41(.a(output_12_41), .b(output_12_10), .y(output_11_41));
wire output_13_41, output_13_10, output_12_41;
mixer gate_output_12_41(.a(output_13_41), .b(output_13_10), .y(output_12_41));
wire output_14_41, output_14_10, output_13_41;
mixer gate_output_13_41(.a(output_14_41), .b(output_14_10), .y(output_13_41));
wire output_15_41, output_15_10, output_14_41;
mixer gate_output_14_41(.a(output_15_41), .b(output_15_10), .y(output_14_41));
wire output_16_41, output_16_10, output_15_41;
mixer gate_output_15_41(.a(output_16_41), .b(output_16_10), .y(output_15_41));
wire output_1_42, output_1_11, output_0_42;
mixer gate_output_0_42(.a(output_1_42), .b(output_1_11), .y(output_0_42));
wire output_2_42, output_2_11, output_1_42;
mixer gate_output_1_42(.a(output_2_42), .b(output_2_11), .y(output_1_42));
wire output_3_42, output_3_11, output_2_42;
mixer gate_output_2_42(.a(output_3_42), .b(output_3_11), .y(output_2_42));
wire output_4_42, output_4_11, output_3_42;
mixer gate_output_3_42(.a(output_4_42), .b(output_4_11), .y(output_3_42));
wire output_5_42, output_5_11, output_4_42;
mixer gate_output_4_42(.a(output_5_42), .b(output_5_11), .y(output_4_42));
wire output_6_42, output_6_11, output_5_42;
mixer gate_output_5_42(.a(output_6_42), .b(output_6_11), .y(output_5_42));
wire output_7_42, output_7_11, output_6_42;
mixer gate_output_6_42(.a(output_7_42), .b(output_7_11), .y(output_6_42));
wire output_8_42, output_8_11, output_7_42;
mixer gate_output_7_42(.a(output_8_42), .b(output_8_11), .y(output_7_42));
wire output_9_42, output_9_11, output_8_42;
mixer gate_output_8_42(.a(output_9_42), .b(output_9_11), .y(output_8_42));
wire output_10_42, output_10_11, output_9_42;
mixer gate_output_9_42(.a(output_10_42), .b(output_10_11), .y(output_9_42));
wire output_11_42, output_11_11, output_10_42;
mixer gate_output_10_42(.a(output_11_42), .b(output_11_11), .y(output_10_42));
wire output_12_42, output_12_11, output_11_42;
mixer gate_output_11_42(.a(output_12_42), .b(output_12_11), .y(output_11_42));
wire output_13_42, output_13_11, output_12_42;
mixer gate_output_12_42(.a(output_13_42), .b(output_13_11), .y(output_12_42));
wire output_14_42, output_14_11, output_13_42;
mixer gate_output_13_42(.a(output_14_42), .b(output_14_11), .y(output_13_42));
wire output_15_42, output_15_11, output_14_42;
mixer gate_output_14_42(.a(output_15_42), .b(output_15_11), .y(output_14_42));
wire output_16_42, output_16_11, output_15_42;
mixer gate_output_15_42(.a(output_16_42), .b(output_16_11), .y(output_15_42));
wire output_1_43, output_1_12, output_0_43;
mixer gate_output_0_43(.a(output_1_43), .b(output_1_12), .y(output_0_43));
wire output_2_43, output_2_12, output_1_43;
mixer gate_output_1_43(.a(output_2_43), .b(output_2_12), .y(output_1_43));
wire output_3_43, output_3_12, output_2_43;
mixer gate_output_2_43(.a(output_3_43), .b(output_3_12), .y(output_2_43));
wire output_4_43, output_4_12, output_3_43;
mixer gate_output_3_43(.a(output_4_43), .b(output_4_12), .y(output_3_43));
wire output_5_43, output_5_12, output_4_43;
mixer gate_output_4_43(.a(output_5_43), .b(output_5_12), .y(output_4_43));
wire output_6_43, output_6_12, output_5_43;
mixer gate_output_5_43(.a(output_6_43), .b(output_6_12), .y(output_5_43));
wire output_7_43, output_7_12, output_6_43;
mixer gate_output_6_43(.a(output_7_43), .b(output_7_12), .y(output_6_43));
wire output_8_43, output_8_12, output_7_43;
mixer gate_output_7_43(.a(output_8_43), .b(output_8_12), .y(output_7_43));
wire output_9_43, output_9_12, output_8_43;
mixer gate_output_8_43(.a(output_9_43), .b(output_9_12), .y(output_8_43));
wire output_10_43, output_10_12, output_9_43;
mixer gate_output_9_43(.a(output_10_43), .b(output_10_12), .y(output_9_43));
wire output_11_43, output_11_12, output_10_43;
mixer gate_output_10_43(.a(output_11_43), .b(output_11_12), .y(output_10_43));
wire output_12_43, output_12_12, output_11_43;
mixer gate_output_11_43(.a(output_12_43), .b(output_12_12), .y(output_11_43));
wire output_13_43, output_13_12, output_12_43;
mixer gate_output_12_43(.a(output_13_43), .b(output_13_12), .y(output_12_43));
wire output_14_43, output_14_12, output_13_43;
mixer gate_output_13_43(.a(output_14_43), .b(output_14_12), .y(output_13_43));
wire output_15_43, output_15_12, output_14_43;
mixer gate_output_14_43(.a(output_15_43), .b(output_15_12), .y(output_14_43));
wire output_16_43, output_16_12, output_15_43;
mixer gate_output_15_43(.a(output_16_43), .b(output_16_12), .y(output_15_43));
wire output_1_44, output_1_13, output_0_44;
mixer gate_output_0_44(.a(output_1_44), .b(output_1_13), .y(output_0_44));
wire output_2_44, output_2_13, output_1_44;
mixer gate_output_1_44(.a(output_2_44), .b(output_2_13), .y(output_1_44));
wire output_3_44, output_3_13, output_2_44;
mixer gate_output_2_44(.a(output_3_44), .b(output_3_13), .y(output_2_44));
wire output_4_44, output_4_13, output_3_44;
mixer gate_output_3_44(.a(output_4_44), .b(output_4_13), .y(output_3_44));
wire output_5_44, output_5_13, output_4_44;
mixer gate_output_4_44(.a(output_5_44), .b(output_5_13), .y(output_4_44));
wire output_6_44, output_6_13, output_5_44;
mixer gate_output_5_44(.a(output_6_44), .b(output_6_13), .y(output_5_44));
wire output_7_44, output_7_13, output_6_44;
mixer gate_output_6_44(.a(output_7_44), .b(output_7_13), .y(output_6_44));
wire output_8_44, output_8_13, output_7_44;
mixer gate_output_7_44(.a(output_8_44), .b(output_8_13), .y(output_7_44));
wire output_9_44, output_9_13, output_8_44;
mixer gate_output_8_44(.a(output_9_44), .b(output_9_13), .y(output_8_44));
wire output_10_44, output_10_13, output_9_44;
mixer gate_output_9_44(.a(output_10_44), .b(output_10_13), .y(output_9_44));
wire output_11_44, output_11_13, output_10_44;
mixer gate_output_10_44(.a(output_11_44), .b(output_11_13), .y(output_10_44));
wire output_12_44, output_12_13, output_11_44;
mixer gate_output_11_44(.a(output_12_44), .b(output_12_13), .y(output_11_44));
wire output_13_44, output_13_13, output_12_44;
mixer gate_output_12_44(.a(output_13_44), .b(output_13_13), .y(output_12_44));
wire output_14_44, output_14_13, output_13_44;
mixer gate_output_13_44(.a(output_14_44), .b(output_14_13), .y(output_13_44));
wire output_15_44, output_15_13, output_14_44;
mixer gate_output_14_44(.a(output_15_44), .b(output_15_13), .y(output_14_44));
wire output_16_44, output_16_13, output_15_44;
mixer gate_output_15_44(.a(output_16_44), .b(output_16_13), .y(output_15_44));
wire output_1_45, output_1_14, output_0_45;
mixer gate_output_0_45(.a(output_1_45), .b(output_1_14), .y(output_0_45));
wire output_2_45, output_2_14, output_1_45;
mixer gate_output_1_45(.a(output_2_45), .b(output_2_14), .y(output_1_45));
wire output_3_45, output_3_14, output_2_45;
mixer gate_output_2_45(.a(output_3_45), .b(output_3_14), .y(output_2_45));
wire output_4_45, output_4_14, output_3_45;
mixer gate_output_3_45(.a(output_4_45), .b(output_4_14), .y(output_3_45));
wire output_5_45, output_5_14, output_4_45;
mixer gate_output_4_45(.a(output_5_45), .b(output_5_14), .y(output_4_45));
wire output_6_45, output_6_14, output_5_45;
mixer gate_output_5_45(.a(output_6_45), .b(output_6_14), .y(output_5_45));
wire output_7_45, output_7_14, output_6_45;
mixer gate_output_6_45(.a(output_7_45), .b(output_7_14), .y(output_6_45));
wire output_8_45, output_8_14, output_7_45;
mixer gate_output_7_45(.a(output_8_45), .b(output_8_14), .y(output_7_45));
wire output_9_45, output_9_14, output_8_45;
mixer gate_output_8_45(.a(output_9_45), .b(output_9_14), .y(output_8_45));
wire output_10_45, output_10_14, output_9_45;
mixer gate_output_9_45(.a(output_10_45), .b(output_10_14), .y(output_9_45));
wire output_11_45, output_11_14, output_10_45;
mixer gate_output_10_45(.a(output_11_45), .b(output_11_14), .y(output_10_45));
wire output_12_45, output_12_14, output_11_45;
mixer gate_output_11_45(.a(output_12_45), .b(output_12_14), .y(output_11_45));
wire output_13_45, output_13_14, output_12_45;
mixer gate_output_12_45(.a(output_13_45), .b(output_13_14), .y(output_12_45));
wire output_14_45, output_14_14, output_13_45;
mixer gate_output_13_45(.a(output_14_45), .b(output_14_14), .y(output_13_45));
wire output_15_45, output_15_14, output_14_45;
mixer gate_output_14_45(.a(output_15_45), .b(output_15_14), .y(output_14_45));
wire output_16_45, output_16_14, output_15_45;
mixer gate_output_15_45(.a(output_16_45), .b(output_16_14), .y(output_15_45));
wire output_1_46, output_1_15, output_0_46;
mixer gate_output_0_46(.a(output_1_46), .b(output_1_15), .y(output_0_46));
wire output_2_46, output_2_15, output_1_46;
mixer gate_output_1_46(.a(output_2_46), .b(output_2_15), .y(output_1_46));
wire output_3_46, output_3_15, output_2_46;
mixer gate_output_2_46(.a(output_3_46), .b(output_3_15), .y(output_2_46));
wire output_4_46, output_4_15, output_3_46;
mixer gate_output_3_46(.a(output_4_46), .b(output_4_15), .y(output_3_46));
wire output_5_46, output_5_15, output_4_46;
mixer gate_output_4_46(.a(output_5_46), .b(output_5_15), .y(output_4_46));
wire output_6_46, output_6_15, output_5_46;
mixer gate_output_5_46(.a(output_6_46), .b(output_6_15), .y(output_5_46));
wire output_7_46, output_7_15, output_6_46;
mixer gate_output_6_46(.a(output_7_46), .b(output_7_15), .y(output_6_46));
wire output_8_46, output_8_15, output_7_46;
mixer gate_output_7_46(.a(output_8_46), .b(output_8_15), .y(output_7_46));
wire output_9_46, output_9_15, output_8_46;
mixer gate_output_8_46(.a(output_9_46), .b(output_9_15), .y(output_8_46));
wire output_10_46, output_10_15, output_9_46;
mixer gate_output_9_46(.a(output_10_46), .b(output_10_15), .y(output_9_46));
wire output_11_46, output_11_15, output_10_46;
mixer gate_output_10_46(.a(output_11_46), .b(output_11_15), .y(output_10_46));
wire output_12_46, output_12_15, output_11_46;
mixer gate_output_11_46(.a(output_12_46), .b(output_12_15), .y(output_11_46));
wire output_13_46, output_13_15, output_12_46;
mixer gate_output_12_46(.a(output_13_46), .b(output_13_15), .y(output_12_46));
wire output_14_46, output_14_15, output_13_46;
mixer gate_output_13_46(.a(output_14_46), .b(output_14_15), .y(output_13_46));
wire output_15_46, output_15_15, output_14_46;
mixer gate_output_14_46(.a(output_15_46), .b(output_15_15), .y(output_14_46));
wire output_16_46, output_16_15, output_15_46;
mixer gate_output_15_46(.a(output_16_46), .b(output_16_15), .y(output_15_46));
wire output_1_47, output_1_0, output_0_47;
mixer gate_output_0_47(.a(output_1_47), .b(output_1_0), .y(output_0_47));
wire output_2_47, output_2_0, output_1_47;
mixer gate_output_1_47(.a(output_2_47), .b(output_2_0), .y(output_1_47));
wire output_3_47, output_3_0, output_2_47;
mixer gate_output_2_47(.a(output_3_47), .b(output_3_0), .y(output_2_47));
wire output_4_47, output_4_0, output_3_47;
mixer gate_output_3_47(.a(output_4_47), .b(output_4_0), .y(output_3_47));
wire output_5_47, output_5_0, output_4_47;
mixer gate_output_4_47(.a(output_5_47), .b(output_5_0), .y(output_4_47));
wire output_6_47, output_6_0, output_5_47;
mixer gate_output_5_47(.a(output_6_47), .b(output_6_0), .y(output_5_47));
wire output_7_47, output_7_0, output_6_47;
mixer gate_output_6_47(.a(output_7_47), .b(output_7_0), .y(output_6_47));
wire output_8_47, output_8_0, output_7_47;
mixer gate_output_7_47(.a(output_8_47), .b(output_8_0), .y(output_7_47));
wire output_9_47, output_9_0, output_8_47;
mixer gate_output_8_47(.a(output_9_47), .b(output_9_0), .y(output_8_47));
wire output_10_47, output_10_0, output_9_47;
mixer gate_output_9_47(.a(output_10_47), .b(output_10_0), .y(output_9_47));
wire output_11_47, output_11_0, output_10_47;
mixer gate_output_10_47(.a(output_11_47), .b(output_11_0), .y(output_10_47));
wire output_12_47, output_12_0, output_11_47;
mixer gate_output_11_47(.a(output_12_47), .b(output_12_0), .y(output_11_47));
wire output_13_47, output_13_0, output_12_47;
mixer gate_output_12_47(.a(output_13_47), .b(output_13_0), .y(output_12_47));
wire output_14_47, output_14_0, output_13_47;
mixer gate_output_13_47(.a(output_14_47), .b(output_14_0), .y(output_13_47));
wire output_15_47, output_15_0, output_14_47;
mixer gate_output_14_47(.a(output_15_47), .b(output_15_0), .y(output_14_47));
wire output_16_47, output_16_0, output_15_47;
mixer gate_output_15_47(.a(output_16_47), .b(output_16_0), .y(output_15_47));
wire output_1_48, output_1_1, output_0_48;
mixer gate_output_0_48(.a(output_1_48), .b(output_1_1), .y(output_0_48));
wire output_2_48, output_2_1, output_1_48;
mixer gate_output_1_48(.a(output_2_48), .b(output_2_1), .y(output_1_48));
wire output_3_48, output_3_1, output_2_48;
mixer gate_output_2_48(.a(output_3_48), .b(output_3_1), .y(output_2_48));
wire output_4_48, output_4_1, output_3_48;
mixer gate_output_3_48(.a(output_4_48), .b(output_4_1), .y(output_3_48));
wire output_5_48, output_5_1, output_4_48;
mixer gate_output_4_48(.a(output_5_48), .b(output_5_1), .y(output_4_48));
wire output_6_48, output_6_1, output_5_48;
mixer gate_output_5_48(.a(output_6_48), .b(output_6_1), .y(output_5_48));
wire output_7_48, output_7_1, output_6_48;
mixer gate_output_6_48(.a(output_7_48), .b(output_7_1), .y(output_6_48));
wire output_8_48, output_8_1, output_7_48;
mixer gate_output_7_48(.a(output_8_48), .b(output_8_1), .y(output_7_48));
wire output_9_48, output_9_1, output_8_48;
mixer gate_output_8_48(.a(output_9_48), .b(output_9_1), .y(output_8_48));
wire output_10_48, output_10_1, output_9_48;
mixer gate_output_9_48(.a(output_10_48), .b(output_10_1), .y(output_9_48));
wire output_11_48, output_11_1, output_10_48;
mixer gate_output_10_48(.a(output_11_48), .b(output_11_1), .y(output_10_48));
wire output_12_48, output_12_1, output_11_48;
mixer gate_output_11_48(.a(output_12_48), .b(output_12_1), .y(output_11_48));
wire output_13_48, output_13_1, output_12_48;
mixer gate_output_12_48(.a(output_13_48), .b(output_13_1), .y(output_12_48));
wire output_14_48, output_14_1, output_13_48;
mixer gate_output_13_48(.a(output_14_48), .b(output_14_1), .y(output_13_48));
wire output_15_48, output_15_1, output_14_48;
mixer gate_output_14_48(.a(output_15_48), .b(output_15_1), .y(output_14_48));
wire output_16_48, output_16_1, output_15_48;
mixer gate_output_15_48(.a(output_16_48), .b(output_16_1), .y(output_15_48));
wire output_1_49, output_1_2, output_0_49;
mixer gate_output_0_49(.a(output_1_49), .b(output_1_2), .y(output_0_49));
wire output_2_49, output_2_2, output_1_49;
mixer gate_output_1_49(.a(output_2_49), .b(output_2_2), .y(output_1_49));
wire output_3_49, output_3_2, output_2_49;
mixer gate_output_2_49(.a(output_3_49), .b(output_3_2), .y(output_2_49));
wire output_4_49, output_4_2, output_3_49;
mixer gate_output_3_49(.a(output_4_49), .b(output_4_2), .y(output_3_49));
wire output_5_49, output_5_2, output_4_49;
mixer gate_output_4_49(.a(output_5_49), .b(output_5_2), .y(output_4_49));
wire output_6_49, output_6_2, output_5_49;
mixer gate_output_5_49(.a(output_6_49), .b(output_6_2), .y(output_5_49));
wire output_7_49, output_7_2, output_6_49;
mixer gate_output_6_49(.a(output_7_49), .b(output_7_2), .y(output_6_49));
wire output_8_49, output_8_2, output_7_49;
mixer gate_output_7_49(.a(output_8_49), .b(output_8_2), .y(output_7_49));
wire output_9_49, output_9_2, output_8_49;
mixer gate_output_8_49(.a(output_9_49), .b(output_9_2), .y(output_8_49));
wire output_10_49, output_10_2, output_9_49;
mixer gate_output_9_49(.a(output_10_49), .b(output_10_2), .y(output_9_49));
wire output_11_49, output_11_2, output_10_49;
mixer gate_output_10_49(.a(output_11_49), .b(output_11_2), .y(output_10_49));
wire output_12_49, output_12_2, output_11_49;
mixer gate_output_11_49(.a(output_12_49), .b(output_12_2), .y(output_11_49));
wire output_13_49, output_13_2, output_12_49;
mixer gate_output_12_49(.a(output_13_49), .b(output_13_2), .y(output_12_49));
wire output_14_49, output_14_2, output_13_49;
mixer gate_output_13_49(.a(output_14_49), .b(output_14_2), .y(output_13_49));
wire output_15_49, output_15_2, output_14_49;
mixer gate_output_14_49(.a(output_15_49), .b(output_15_2), .y(output_14_49));
wire output_16_49, output_16_2, output_15_49;
mixer gate_output_15_49(.a(output_16_49), .b(output_16_2), .y(output_15_49));
wire output_1_50, output_1_3, output_0_50;
mixer gate_output_0_50(.a(output_1_50), .b(output_1_3), .y(output_0_50));
wire output_2_50, output_2_3, output_1_50;
mixer gate_output_1_50(.a(output_2_50), .b(output_2_3), .y(output_1_50));
wire output_3_50, output_3_3, output_2_50;
mixer gate_output_2_50(.a(output_3_50), .b(output_3_3), .y(output_2_50));
wire output_4_50, output_4_3, output_3_50;
mixer gate_output_3_50(.a(output_4_50), .b(output_4_3), .y(output_3_50));
wire output_5_50, output_5_3, output_4_50;
mixer gate_output_4_50(.a(output_5_50), .b(output_5_3), .y(output_4_50));
wire output_6_50, output_6_3, output_5_50;
mixer gate_output_5_50(.a(output_6_50), .b(output_6_3), .y(output_5_50));
wire output_7_50, output_7_3, output_6_50;
mixer gate_output_6_50(.a(output_7_50), .b(output_7_3), .y(output_6_50));
wire output_8_50, output_8_3, output_7_50;
mixer gate_output_7_50(.a(output_8_50), .b(output_8_3), .y(output_7_50));
wire output_9_50, output_9_3, output_8_50;
mixer gate_output_8_50(.a(output_9_50), .b(output_9_3), .y(output_8_50));
wire output_10_50, output_10_3, output_9_50;
mixer gate_output_9_50(.a(output_10_50), .b(output_10_3), .y(output_9_50));
wire output_11_50, output_11_3, output_10_50;
mixer gate_output_10_50(.a(output_11_50), .b(output_11_3), .y(output_10_50));
wire output_12_50, output_12_3, output_11_50;
mixer gate_output_11_50(.a(output_12_50), .b(output_12_3), .y(output_11_50));
wire output_13_50, output_13_3, output_12_50;
mixer gate_output_12_50(.a(output_13_50), .b(output_13_3), .y(output_12_50));
wire output_14_50, output_14_3, output_13_50;
mixer gate_output_13_50(.a(output_14_50), .b(output_14_3), .y(output_13_50));
wire output_15_50, output_15_3, output_14_50;
mixer gate_output_14_50(.a(output_15_50), .b(output_15_3), .y(output_14_50));
wire output_16_50, output_16_3, output_15_50;
mixer gate_output_15_50(.a(output_16_50), .b(output_16_3), .y(output_15_50));
wire output_1_51, output_1_4, output_0_51;
mixer gate_output_0_51(.a(output_1_51), .b(output_1_4), .y(output_0_51));
wire output_2_51, output_2_4, output_1_51;
mixer gate_output_1_51(.a(output_2_51), .b(output_2_4), .y(output_1_51));
wire output_3_51, output_3_4, output_2_51;
mixer gate_output_2_51(.a(output_3_51), .b(output_3_4), .y(output_2_51));
wire output_4_51, output_4_4, output_3_51;
mixer gate_output_3_51(.a(output_4_51), .b(output_4_4), .y(output_3_51));
wire output_5_51, output_5_4, output_4_51;
mixer gate_output_4_51(.a(output_5_51), .b(output_5_4), .y(output_4_51));
wire output_6_51, output_6_4, output_5_51;
mixer gate_output_5_51(.a(output_6_51), .b(output_6_4), .y(output_5_51));
wire output_7_51, output_7_4, output_6_51;
mixer gate_output_6_51(.a(output_7_51), .b(output_7_4), .y(output_6_51));
wire output_8_51, output_8_4, output_7_51;
mixer gate_output_7_51(.a(output_8_51), .b(output_8_4), .y(output_7_51));
wire output_9_51, output_9_4, output_8_51;
mixer gate_output_8_51(.a(output_9_51), .b(output_9_4), .y(output_8_51));
wire output_10_51, output_10_4, output_9_51;
mixer gate_output_9_51(.a(output_10_51), .b(output_10_4), .y(output_9_51));
wire output_11_51, output_11_4, output_10_51;
mixer gate_output_10_51(.a(output_11_51), .b(output_11_4), .y(output_10_51));
wire output_12_51, output_12_4, output_11_51;
mixer gate_output_11_51(.a(output_12_51), .b(output_12_4), .y(output_11_51));
wire output_13_51, output_13_4, output_12_51;
mixer gate_output_12_51(.a(output_13_51), .b(output_13_4), .y(output_12_51));
wire output_14_51, output_14_4, output_13_51;
mixer gate_output_13_51(.a(output_14_51), .b(output_14_4), .y(output_13_51));
wire output_15_51, output_15_4, output_14_51;
mixer gate_output_14_51(.a(output_15_51), .b(output_15_4), .y(output_14_51));
wire output_16_51, output_16_4, output_15_51;
mixer gate_output_15_51(.a(output_16_51), .b(output_16_4), .y(output_15_51));
wire output_1_52, output_1_5, output_0_52;
mixer gate_output_0_52(.a(output_1_52), .b(output_1_5), .y(output_0_52));
wire output_2_52, output_2_5, output_1_52;
mixer gate_output_1_52(.a(output_2_52), .b(output_2_5), .y(output_1_52));
wire output_3_52, output_3_5, output_2_52;
mixer gate_output_2_52(.a(output_3_52), .b(output_3_5), .y(output_2_52));
wire output_4_52, output_4_5, output_3_52;
mixer gate_output_3_52(.a(output_4_52), .b(output_4_5), .y(output_3_52));
wire output_5_52, output_5_5, output_4_52;
mixer gate_output_4_52(.a(output_5_52), .b(output_5_5), .y(output_4_52));
wire output_6_52, output_6_5, output_5_52;
mixer gate_output_5_52(.a(output_6_52), .b(output_6_5), .y(output_5_52));
wire output_7_52, output_7_5, output_6_52;
mixer gate_output_6_52(.a(output_7_52), .b(output_7_5), .y(output_6_52));
wire output_8_52, output_8_5, output_7_52;
mixer gate_output_7_52(.a(output_8_52), .b(output_8_5), .y(output_7_52));
wire output_9_52, output_9_5, output_8_52;
mixer gate_output_8_52(.a(output_9_52), .b(output_9_5), .y(output_8_52));
wire output_10_52, output_10_5, output_9_52;
mixer gate_output_9_52(.a(output_10_52), .b(output_10_5), .y(output_9_52));
wire output_11_52, output_11_5, output_10_52;
mixer gate_output_10_52(.a(output_11_52), .b(output_11_5), .y(output_10_52));
wire output_12_52, output_12_5, output_11_52;
mixer gate_output_11_52(.a(output_12_52), .b(output_12_5), .y(output_11_52));
wire output_13_52, output_13_5, output_12_52;
mixer gate_output_12_52(.a(output_13_52), .b(output_13_5), .y(output_12_52));
wire output_14_52, output_14_5, output_13_52;
mixer gate_output_13_52(.a(output_14_52), .b(output_14_5), .y(output_13_52));
wire output_15_52, output_15_5, output_14_52;
mixer gate_output_14_52(.a(output_15_52), .b(output_15_5), .y(output_14_52));
wire output_16_52, output_16_5, output_15_52;
mixer gate_output_15_52(.a(output_16_52), .b(output_16_5), .y(output_15_52));
wire output_1_53, output_1_6, output_0_53;
mixer gate_output_0_53(.a(output_1_53), .b(output_1_6), .y(output_0_53));
wire output_2_53, output_2_6, output_1_53;
mixer gate_output_1_53(.a(output_2_53), .b(output_2_6), .y(output_1_53));
wire output_3_53, output_3_6, output_2_53;
mixer gate_output_2_53(.a(output_3_53), .b(output_3_6), .y(output_2_53));
wire output_4_53, output_4_6, output_3_53;
mixer gate_output_3_53(.a(output_4_53), .b(output_4_6), .y(output_3_53));
wire output_5_53, output_5_6, output_4_53;
mixer gate_output_4_53(.a(output_5_53), .b(output_5_6), .y(output_4_53));
wire output_6_53, output_6_6, output_5_53;
mixer gate_output_5_53(.a(output_6_53), .b(output_6_6), .y(output_5_53));
wire output_7_53, output_7_6, output_6_53;
mixer gate_output_6_53(.a(output_7_53), .b(output_7_6), .y(output_6_53));
wire output_8_53, output_8_6, output_7_53;
mixer gate_output_7_53(.a(output_8_53), .b(output_8_6), .y(output_7_53));
wire output_9_53, output_9_6, output_8_53;
mixer gate_output_8_53(.a(output_9_53), .b(output_9_6), .y(output_8_53));
wire output_10_53, output_10_6, output_9_53;
mixer gate_output_9_53(.a(output_10_53), .b(output_10_6), .y(output_9_53));
wire output_11_53, output_11_6, output_10_53;
mixer gate_output_10_53(.a(output_11_53), .b(output_11_6), .y(output_10_53));
wire output_12_53, output_12_6, output_11_53;
mixer gate_output_11_53(.a(output_12_53), .b(output_12_6), .y(output_11_53));
wire output_13_53, output_13_6, output_12_53;
mixer gate_output_12_53(.a(output_13_53), .b(output_13_6), .y(output_12_53));
wire output_14_53, output_14_6, output_13_53;
mixer gate_output_13_53(.a(output_14_53), .b(output_14_6), .y(output_13_53));
wire output_15_53, output_15_6, output_14_53;
mixer gate_output_14_53(.a(output_15_53), .b(output_15_6), .y(output_14_53));
wire output_16_53, output_16_6, output_15_53;
mixer gate_output_15_53(.a(output_16_53), .b(output_16_6), .y(output_15_53));
wire output_1_54, output_1_7, output_0_54;
mixer gate_output_0_54(.a(output_1_54), .b(output_1_7), .y(output_0_54));
wire output_2_54, output_2_7, output_1_54;
mixer gate_output_1_54(.a(output_2_54), .b(output_2_7), .y(output_1_54));
wire output_3_54, output_3_7, output_2_54;
mixer gate_output_2_54(.a(output_3_54), .b(output_3_7), .y(output_2_54));
wire output_4_54, output_4_7, output_3_54;
mixer gate_output_3_54(.a(output_4_54), .b(output_4_7), .y(output_3_54));
wire output_5_54, output_5_7, output_4_54;
mixer gate_output_4_54(.a(output_5_54), .b(output_5_7), .y(output_4_54));
wire output_6_54, output_6_7, output_5_54;
mixer gate_output_5_54(.a(output_6_54), .b(output_6_7), .y(output_5_54));
wire output_7_54, output_7_7, output_6_54;
mixer gate_output_6_54(.a(output_7_54), .b(output_7_7), .y(output_6_54));
wire output_8_54, output_8_7, output_7_54;
mixer gate_output_7_54(.a(output_8_54), .b(output_8_7), .y(output_7_54));
wire output_9_54, output_9_7, output_8_54;
mixer gate_output_8_54(.a(output_9_54), .b(output_9_7), .y(output_8_54));
wire output_10_54, output_10_7, output_9_54;
mixer gate_output_9_54(.a(output_10_54), .b(output_10_7), .y(output_9_54));
wire output_11_54, output_11_7, output_10_54;
mixer gate_output_10_54(.a(output_11_54), .b(output_11_7), .y(output_10_54));
wire output_12_54, output_12_7, output_11_54;
mixer gate_output_11_54(.a(output_12_54), .b(output_12_7), .y(output_11_54));
wire output_13_54, output_13_7, output_12_54;
mixer gate_output_12_54(.a(output_13_54), .b(output_13_7), .y(output_12_54));
wire output_14_54, output_14_7, output_13_54;
mixer gate_output_13_54(.a(output_14_54), .b(output_14_7), .y(output_13_54));
wire output_15_54, output_15_7, output_14_54;
mixer gate_output_14_54(.a(output_15_54), .b(output_15_7), .y(output_14_54));
wire output_16_54, output_16_7, output_15_54;
mixer gate_output_15_54(.a(output_16_54), .b(output_16_7), .y(output_15_54));
wire output_1_55, output_1_8, output_0_55;
mixer gate_output_0_55(.a(output_1_55), .b(output_1_8), .y(output_0_55));
wire output_2_55, output_2_8, output_1_55;
mixer gate_output_1_55(.a(output_2_55), .b(output_2_8), .y(output_1_55));
wire output_3_55, output_3_8, output_2_55;
mixer gate_output_2_55(.a(output_3_55), .b(output_3_8), .y(output_2_55));
wire output_4_55, output_4_8, output_3_55;
mixer gate_output_3_55(.a(output_4_55), .b(output_4_8), .y(output_3_55));
wire output_5_55, output_5_8, output_4_55;
mixer gate_output_4_55(.a(output_5_55), .b(output_5_8), .y(output_4_55));
wire output_6_55, output_6_8, output_5_55;
mixer gate_output_5_55(.a(output_6_55), .b(output_6_8), .y(output_5_55));
wire output_7_55, output_7_8, output_6_55;
mixer gate_output_6_55(.a(output_7_55), .b(output_7_8), .y(output_6_55));
wire output_8_55, output_8_8, output_7_55;
mixer gate_output_7_55(.a(output_8_55), .b(output_8_8), .y(output_7_55));
wire output_9_55, output_9_8, output_8_55;
mixer gate_output_8_55(.a(output_9_55), .b(output_9_8), .y(output_8_55));
wire output_10_55, output_10_8, output_9_55;
mixer gate_output_9_55(.a(output_10_55), .b(output_10_8), .y(output_9_55));
wire output_11_55, output_11_8, output_10_55;
mixer gate_output_10_55(.a(output_11_55), .b(output_11_8), .y(output_10_55));
wire output_12_55, output_12_8, output_11_55;
mixer gate_output_11_55(.a(output_12_55), .b(output_12_8), .y(output_11_55));
wire output_13_55, output_13_8, output_12_55;
mixer gate_output_12_55(.a(output_13_55), .b(output_13_8), .y(output_12_55));
wire output_14_55, output_14_8, output_13_55;
mixer gate_output_13_55(.a(output_14_55), .b(output_14_8), .y(output_13_55));
wire output_15_55, output_15_8, output_14_55;
mixer gate_output_14_55(.a(output_15_55), .b(output_15_8), .y(output_14_55));
wire output_16_55, output_16_8, output_15_55;
mixer gate_output_15_55(.a(output_16_55), .b(output_16_8), .y(output_15_55));
wire output_1_56, output_1_9, output_0_56;
mixer gate_output_0_56(.a(output_1_56), .b(output_1_9), .y(output_0_56));
wire output_2_56, output_2_9, output_1_56;
mixer gate_output_1_56(.a(output_2_56), .b(output_2_9), .y(output_1_56));
wire output_3_56, output_3_9, output_2_56;
mixer gate_output_2_56(.a(output_3_56), .b(output_3_9), .y(output_2_56));
wire output_4_56, output_4_9, output_3_56;
mixer gate_output_3_56(.a(output_4_56), .b(output_4_9), .y(output_3_56));
wire output_5_56, output_5_9, output_4_56;
mixer gate_output_4_56(.a(output_5_56), .b(output_5_9), .y(output_4_56));
wire output_6_56, output_6_9, output_5_56;
mixer gate_output_5_56(.a(output_6_56), .b(output_6_9), .y(output_5_56));
wire output_7_56, output_7_9, output_6_56;
mixer gate_output_6_56(.a(output_7_56), .b(output_7_9), .y(output_6_56));
wire output_8_56, output_8_9, output_7_56;
mixer gate_output_7_56(.a(output_8_56), .b(output_8_9), .y(output_7_56));
wire output_9_56, output_9_9, output_8_56;
mixer gate_output_8_56(.a(output_9_56), .b(output_9_9), .y(output_8_56));
wire output_10_56, output_10_9, output_9_56;
mixer gate_output_9_56(.a(output_10_56), .b(output_10_9), .y(output_9_56));
wire output_11_56, output_11_9, output_10_56;
mixer gate_output_10_56(.a(output_11_56), .b(output_11_9), .y(output_10_56));
wire output_12_56, output_12_9, output_11_56;
mixer gate_output_11_56(.a(output_12_56), .b(output_12_9), .y(output_11_56));
wire output_13_56, output_13_9, output_12_56;
mixer gate_output_12_56(.a(output_13_56), .b(output_13_9), .y(output_12_56));
wire output_14_56, output_14_9, output_13_56;
mixer gate_output_13_56(.a(output_14_56), .b(output_14_9), .y(output_13_56));
wire output_15_56, output_15_9, output_14_56;
mixer gate_output_14_56(.a(output_15_56), .b(output_15_9), .y(output_14_56));
wire output_16_56, output_16_9, output_15_56;
mixer gate_output_15_56(.a(output_16_56), .b(output_16_9), .y(output_15_56));
wire output_1_57, output_1_10, output_0_57;
mixer gate_output_0_57(.a(output_1_57), .b(output_1_10), .y(output_0_57));
wire output_2_57, output_2_10, output_1_57;
mixer gate_output_1_57(.a(output_2_57), .b(output_2_10), .y(output_1_57));
wire output_3_57, output_3_10, output_2_57;
mixer gate_output_2_57(.a(output_3_57), .b(output_3_10), .y(output_2_57));
wire output_4_57, output_4_10, output_3_57;
mixer gate_output_3_57(.a(output_4_57), .b(output_4_10), .y(output_3_57));
wire output_5_57, output_5_10, output_4_57;
mixer gate_output_4_57(.a(output_5_57), .b(output_5_10), .y(output_4_57));
wire output_6_57, output_6_10, output_5_57;
mixer gate_output_5_57(.a(output_6_57), .b(output_6_10), .y(output_5_57));
wire output_7_57, output_7_10, output_6_57;
mixer gate_output_6_57(.a(output_7_57), .b(output_7_10), .y(output_6_57));
wire output_8_57, output_8_10, output_7_57;
mixer gate_output_7_57(.a(output_8_57), .b(output_8_10), .y(output_7_57));
wire output_9_57, output_9_10, output_8_57;
mixer gate_output_8_57(.a(output_9_57), .b(output_9_10), .y(output_8_57));
wire output_10_57, output_10_10, output_9_57;
mixer gate_output_9_57(.a(output_10_57), .b(output_10_10), .y(output_9_57));
wire output_11_57, output_11_10, output_10_57;
mixer gate_output_10_57(.a(output_11_57), .b(output_11_10), .y(output_10_57));
wire output_12_57, output_12_10, output_11_57;
mixer gate_output_11_57(.a(output_12_57), .b(output_12_10), .y(output_11_57));
wire output_13_57, output_13_10, output_12_57;
mixer gate_output_12_57(.a(output_13_57), .b(output_13_10), .y(output_12_57));
wire output_14_57, output_14_10, output_13_57;
mixer gate_output_13_57(.a(output_14_57), .b(output_14_10), .y(output_13_57));
wire output_15_57, output_15_10, output_14_57;
mixer gate_output_14_57(.a(output_15_57), .b(output_15_10), .y(output_14_57));
wire output_16_57, output_16_10, output_15_57;
mixer gate_output_15_57(.a(output_16_57), .b(output_16_10), .y(output_15_57));
wire output_1_58, output_1_11, output_0_58;
mixer gate_output_0_58(.a(output_1_58), .b(output_1_11), .y(output_0_58));
wire output_2_58, output_2_11, output_1_58;
mixer gate_output_1_58(.a(output_2_58), .b(output_2_11), .y(output_1_58));
wire output_3_58, output_3_11, output_2_58;
mixer gate_output_2_58(.a(output_3_58), .b(output_3_11), .y(output_2_58));
wire output_4_58, output_4_11, output_3_58;
mixer gate_output_3_58(.a(output_4_58), .b(output_4_11), .y(output_3_58));
wire output_5_58, output_5_11, output_4_58;
mixer gate_output_4_58(.a(output_5_58), .b(output_5_11), .y(output_4_58));
wire output_6_58, output_6_11, output_5_58;
mixer gate_output_5_58(.a(output_6_58), .b(output_6_11), .y(output_5_58));
wire output_7_58, output_7_11, output_6_58;
mixer gate_output_6_58(.a(output_7_58), .b(output_7_11), .y(output_6_58));
wire output_8_58, output_8_11, output_7_58;
mixer gate_output_7_58(.a(output_8_58), .b(output_8_11), .y(output_7_58));
wire output_9_58, output_9_11, output_8_58;
mixer gate_output_8_58(.a(output_9_58), .b(output_9_11), .y(output_8_58));
wire output_10_58, output_10_11, output_9_58;
mixer gate_output_9_58(.a(output_10_58), .b(output_10_11), .y(output_9_58));
wire output_11_58, output_11_11, output_10_58;
mixer gate_output_10_58(.a(output_11_58), .b(output_11_11), .y(output_10_58));
wire output_12_58, output_12_11, output_11_58;
mixer gate_output_11_58(.a(output_12_58), .b(output_12_11), .y(output_11_58));
wire output_13_58, output_13_11, output_12_58;
mixer gate_output_12_58(.a(output_13_58), .b(output_13_11), .y(output_12_58));
wire output_14_58, output_14_11, output_13_58;
mixer gate_output_13_58(.a(output_14_58), .b(output_14_11), .y(output_13_58));
wire output_15_58, output_15_11, output_14_58;
mixer gate_output_14_58(.a(output_15_58), .b(output_15_11), .y(output_14_58));
wire output_16_58, output_16_11, output_15_58;
mixer gate_output_15_58(.a(output_16_58), .b(output_16_11), .y(output_15_58));
wire output_1_59, output_1_12, output_0_59;
mixer gate_output_0_59(.a(output_1_59), .b(output_1_12), .y(output_0_59));
wire output_2_59, output_2_12, output_1_59;
mixer gate_output_1_59(.a(output_2_59), .b(output_2_12), .y(output_1_59));
wire output_3_59, output_3_12, output_2_59;
mixer gate_output_2_59(.a(output_3_59), .b(output_3_12), .y(output_2_59));
wire output_4_59, output_4_12, output_3_59;
mixer gate_output_3_59(.a(output_4_59), .b(output_4_12), .y(output_3_59));
wire output_5_59, output_5_12, output_4_59;
mixer gate_output_4_59(.a(output_5_59), .b(output_5_12), .y(output_4_59));
wire output_6_59, output_6_12, output_5_59;
mixer gate_output_5_59(.a(output_6_59), .b(output_6_12), .y(output_5_59));
wire output_7_59, output_7_12, output_6_59;
mixer gate_output_6_59(.a(output_7_59), .b(output_7_12), .y(output_6_59));
wire output_8_59, output_8_12, output_7_59;
mixer gate_output_7_59(.a(output_8_59), .b(output_8_12), .y(output_7_59));
wire output_9_59, output_9_12, output_8_59;
mixer gate_output_8_59(.a(output_9_59), .b(output_9_12), .y(output_8_59));
wire output_10_59, output_10_12, output_9_59;
mixer gate_output_9_59(.a(output_10_59), .b(output_10_12), .y(output_9_59));
wire output_11_59, output_11_12, output_10_59;
mixer gate_output_10_59(.a(output_11_59), .b(output_11_12), .y(output_10_59));
wire output_12_59, output_12_12, output_11_59;
mixer gate_output_11_59(.a(output_12_59), .b(output_12_12), .y(output_11_59));
wire output_13_59, output_13_12, output_12_59;
mixer gate_output_12_59(.a(output_13_59), .b(output_13_12), .y(output_12_59));
wire output_14_59, output_14_12, output_13_59;
mixer gate_output_13_59(.a(output_14_59), .b(output_14_12), .y(output_13_59));
wire output_15_59, output_15_12, output_14_59;
mixer gate_output_14_59(.a(output_15_59), .b(output_15_12), .y(output_14_59));
wire output_16_59, output_16_12, output_15_59;
mixer gate_output_15_59(.a(output_16_59), .b(output_16_12), .y(output_15_59));
wire output_1_60, output_1_13, output_0_60;
mixer gate_output_0_60(.a(output_1_60), .b(output_1_13), .y(output_0_60));
wire output_2_60, output_2_13, output_1_60;
mixer gate_output_1_60(.a(output_2_60), .b(output_2_13), .y(output_1_60));
wire output_3_60, output_3_13, output_2_60;
mixer gate_output_2_60(.a(output_3_60), .b(output_3_13), .y(output_2_60));
wire output_4_60, output_4_13, output_3_60;
mixer gate_output_3_60(.a(output_4_60), .b(output_4_13), .y(output_3_60));
wire output_5_60, output_5_13, output_4_60;
mixer gate_output_4_60(.a(output_5_60), .b(output_5_13), .y(output_4_60));
wire output_6_60, output_6_13, output_5_60;
mixer gate_output_5_60(.a(output_6_60), .b(output_6_13), .y(output_5_60));
wire output_7_60, output_7_13, output_6_60;
mixer gate_output_6_60(.a(output_7_60), .b(output_7_13), .y(output_6_60));
wire output_8_60, output_8_13, output_7_60;
mixer gate_output_7_60(.a(output_8_60), .b(output_8_13), .y(output_7_60));
wire output_9_60, output_9_13, output_8_60;
mixer gate_output_8_60(.a(output_9_60), .b(output_9_13), .y(output_8_60));
wire output_10_60, output_10_13, output_9_60;
mixer gate_output_9_60(.a(output_10_60), .b(output_10_13), .y(output_9_60));
wire output_11_60, output_11_13, output_10_60;
mixer gate_output_10_60(.a(output_11_60), .b(output_11_13), .y(output_10_60));
wire output_12_60, output_12_13, output_11_60;
mixer gate_output_11_60(.a(output_12_60), .b(output_12_13), .y(output_11_60));
wire output_13_60, output_13_13, output_12_60;
mixer gate_output_12_60(.a(output_13_60), .b(output_13_13), .y(output_12_60));
wire output_14_60, output_14_13, output_13_60;
mixer gate_output_13_60(.a(output_14_60), .b(output_14_13), .y(output_13_60));
wire output_15_60, output_15_13, output_14_60;
mixer gate_output_14_60(.a(output_15_60), .b(output_15_13), .y(output_14_60));
wire output_16_60, output_16_13, output_15_60;
mixer gate_output_15_60(.a(output_16_60), .b(output_16_13), .y(output_15_60));
wire output_1_61, output_1_14, output_0_61;
mixer gate_output_0_61(.a(output_1_61), .b(output_1_14), .y(output_0_61));
wire output_2_61, output_2_14, output_1_61;
mixer gate_output_1_61(.a(output_2_61), .b(output_2_14), .y(output_1_61));
wire output_3_61, output_3_14, output_2_61;
mixer gate_output_2_61(.a(output_3_61), .b(output_3_14), .y(output_2_61));
wire output_4_61, output_4_14, output_3_61;
mixer gate_output_3_61(.a(output_4_61), .b(output_4_14), .y(output_3_61));
wire output_5_61, output_5_14, output_4_61;
mixer gate_output_4_61(.a(output_5_61), .b(output_5_14), .y(output_4_61));
wire output_6_61, output_6_14, output_5_61;
mixer gate_output_5_61(.a(output_6_61), .b(output_6_14), .y(output_5_61));
wire output_7_61, output_7_14, output_6_61;
mixer gate_output_6_61(.a(output_7_61), .b(output_7_14), .y(output_6_61));
wire output_8_61, output_8_14, output_7_61;
mixer gate_output_7_61(.a(output_8_61), .b(output_8_14), .y(output_7_61));
wire output_9_61, output_9_14, output_8_61;
mixer gate_output_8_61(.a(output_9_61), .b(output_9_14), .y(output_8_61));
wire output_10_61, output_10_14, output_9_61;
mixer gate_output_9_61(.a(output_10_61), .b(output_10_14), .y(output_9_61));
wire output_11_61, output_11_14, output_10_61;
mixer gate_output_10_61(.a(output_11_61), .b(output_11_14), .y(output_10_61));
wire output_12_61, output_12_14, output_11_61;
mixer gate_output_11_61(.a(output_12_61), .b(output_12_14), .y(output_11_61));
wire output_13_61, output_13_14, output_12_61;
mixer gate_output_12_61(.a(output_13_61), .b(output_13_14), .y(output_12_61));
wire output_14_61, output_14_14, output_13_61;
mixer gate_output_13_61(.a(output_14_61), .b(output_14_14), .y(output_13_61));
wire output_15_61, output_15_14, output_14_61;
mixer gate_output_14_61(.a(output_15_61), .b(output_15_14), .y(output_14_61));
wire output_16_61, output_16_14, output_15_61;
mixer gate_output_15_61(.a(output_16_61), .b(output_16_14), .y(output_15_61));
wire output_1_62, output_1_15, output_0_62;
mixer gate_output_0_62(.a(output_1_62), .b(output_1_15), .y(output_0_62));
wire output_2_62, output_2_15, output_1_62;
mixer gate_output_1_62(.a(output_2_62), .b(output_2_15), .y(output_1_62));
wire output_3_62, output_3_15, output_2_62;
mixer gate_output_2_62(.a(output_3_62), .b(output_3_15), .y(output_2_62));
wire output_4_62, output_4_15, output_3_62;
mixer gate_output_3_62(.a(output_4_62), .b(output_4_15), .y(output_3_62));
wire output_5_62, output_5_15, output_4_62;
mixer gate_output_4_62(.a(output_5_62), .b(output_5_15), .y(output_4_62));
wire output_6_62, output_6_15, output_5_62;
mixer gate_output_5_62(.a(output_6_62), .b(output_6_15), .y(output_5_62));
wire output_7_62, output_7_15, output_6_62;
mixer gate_output_6_62(.a(output_7_62), .b(output_7_15), .y(output_6_62));
wire output_8_62, output_8_15, output_7_62;
mixer gate_output_7_62(.a(output_8_62), .b(output_8_15), .y(output_7_62));
wire output_9_62, output_9_15, output_8_62;
mixer gate_output_8_62(.a(output_9_62), .b(output_9_15), .y(output_8_62));
wire output_10_62, output_10_15, output_9_62;
mixer gate_output_9_62(.a(output_10_62), .b(output_10_15), .y(output_9_62));
wire output_11_62, output_11_15, output_10_62;
mixer gate_output_10_62(.a(output_11_62), .b(output_11_15), .y(output_10_62));
wire output_12_62, output_12_15, output_11_62;
mixer gate_output_11_62(.a(output_12_62), .b(output_12_15), .y(output_11_62));
wire output_13_62, output_13_15, output_12_62;
mixer gate_output_12_62(.a(output_13_62), .b(output_13_15), .y(output_12_62));
wire output_14_62, output_14_15, output_13_62;
mixer gate_output_13_62(.a(output_14_62), .b(output_14_15), .y(output_13_62));
wire output_15_62, output_15_15, output_14_62;
mixer gate_output_14_62(.a(output_15_62), .b(output_15_15), .y(output_14_62));
wire output_16_62, output_16_15, output_15_62;
mixer gate_output_15_62(.a(output_16_62), .b(output_16_15), .y(output_15_62));
wire output_1_63, output_1_0, output_0_63;
mixer gate_output_0_63(.a(output_1_63), .b(output_1_0), .y(output_0_63));
wire output_2_63, output_2_0, output_1_63;
mixer gate_output_1_63(.a(output_2_63), .b(output_2_0), .y(output_1_63));
wire output_3_63, output_3_0, output_2_63;
mixer gate_output_2_63(.a(output_3_63), .b(output_3_0), .y(output_2_63));
wire output_4_63, output_4_0, output_3_63;
mixer gate_output_3_63(.a(output_4_63), .b(output_4_0), .y(output_3_63));
wire output_5_63, output_5_0, output_4_63;
mixer gate_output_4_63(.a(output_5_63), .b(output_5_0), .y(output_4_63));
wire output_6_63, output_6_0, output_5_63;
mixer gate_output_5_63(.a(output_6_63), .b(output_6_0), .y(output_5_63));
wire output_7_63, output_7_0, output_6_63;
mixer gate_output_6_63(.a(output_7_63), .b(output_7_0), .y(output_6_63));
wire output_8_63, output_8_0, output_7_63;
mixer gate_output_7_63(.a(output_8_63), .b(output_8_0), .y(output_7_63));
wire output_9_63, output_9_0, output_8_63;
mixer gate_output_8_63(.a(output_9_63), .b(output_9_0), .y(output_8_63));
wire output_10_63, output_10_0, output_9_63;
mixer gate_output_9_63(.a(output_10_63), .b(output_10_0), .y(output_9_63));
wire output_11_63, output_11_0, output_10_63;
mixer gate_output_10_63(.a(output_11_63), .b(output_11_0), .y(output_10_63));
wire output_12_63, output_12_0, output_11_63;
mixer gate_output_11_63(.a(output_12_63), .b(output_12_0), .y(output_11_63));
wire output_13_63, output_13_0, output_12_63;
mixer gate_output_12_63(.a(output_13_63), .b(output_13_0), .y(output_12_63));
wire output_14_63, output_14_0, output_13_63;
mixer gate_output_13_63(.a(output_14_63), .b(output_14_0), .y(output_13_63));
wire output_15_63, output_15_0, output_14_63;
mixer gate_output_14_63(.a(output_15_63), .b(output_15_0), .y(output_14_63));
wire output_16_63, output_16_0, output_15_63;
mixer gate_output_15_63(.a(output_16_63), .b(output_16_0), .y(output_15_63));
wire output_1_64, output_1_1, output_0_64;
mixer gate_output_0_64(.a(output_1_64), .b(output_1_1), .y(output_0_64));
wire output_2_64, output_2_1, output_1_64;
mixer gate_output_1_64(.a(output_2_64), .b(output_2_1), .y(output_1_64));
wire output_3_64, output_3_1, output_2_64;
mixer gate_output_2_64(.a(output_3_64), .b(output_3_1), .y(output_2_64));
wire output_4_64, output_4_1, output_3_64;
mixer gate_output_3_64(.a(output_4_64), .b(output_4_1), .y(output_3_64));
wire output_5_64, output_5_1, output_4_64;
mixer gate_output_4_64(.a(output_5_64), .b(output_5_1), .y(output_4_64));
wire output_6_64, output_6_1, output_5_64;
mixer gate_output_5_64(.a(output_6_64), .b(output_6_1), .y(output_5_64));
wire output_7_64, output_7_1, output_6_64;
mixer gate_output_6_64(.a(output_7_64), .b(output_7_1), .y(output_6_64));
wire output_8_64, output_8_1, output_7_64;
mixer gate_output_7_64(.a(output_8_64), .b(output_8_1), .y(output_7_64));
wire output_9_64, output_9_1, output_8_64;
mixer gate_output_8_64(.a(output_9_64), .b(output_9_1), .y(output_8_64));
wire output_10_64, output_10_1, output_9_64;
mixer gate_output_9_64(.a(output_10_64), .b(output_10_1), .y(output_9_64));
wire output_11_64, output_11_1, output_10_64;
mixer gate_output_10_64(.a(output_11_64), .b(output_11_1), .y(output_10_64));
wire output_12_64, output_12_1, output_11_64;
mixer gate_output_11_64(.a(output_12_64), .b(output_12_1), .y(output_11_64));
wire output_13_64, output_13_1, output_12_64;
mixer gate_output_12_64(.a(output_13_64), .b(output_13_1), .y(output_12_64));
wire output_14_64, output_14_1, output_13_64;
mixer gate_output_13_64(.a(output_14_64), .b(output_14_1), .y(output_13_64));
wire output_15_64, output_15_1, output_14_64;
mixer gate_output_14_64(.a(output_15_64), .b(output_15_1), .y(output_14_64));
wire output_16_64, output_16_1, output_15_64;
mixer gate_output_15_64(.a(output_16_64), .b(output_16_1), .y(output_15_64));
wire output_1_65, output_1_2, output_0_65;
mixer gate_output_0_65(.a(output_1_65), .b(output_1_2), .y(output_0_65));
wire output_2_65, output_2_2, output_1_65;
mixer gate_output_1_65(.a(output_2_65), .b(output_2_2), .y(output_1_65));
wire output_3_65, output_3_2, output_2_65;
mixer gate_output_2_65(.a(output_3_65), .b(output_3_2), .y(output_2_65));
wire output_4_65, output_4_2, output_3_65;
mixer gate_output_3_65(.a(output_4_65), .b(output_4_2), .y(output_3_65));
wire output_5_65, output_5_2, output_4_65;
mixer gate_output_4_65(.a(output_5_65), .b(output_5_2), .y(output_4_65));
wire output_6_65, output_6_2, output_5_65;
mixer gate_output_5_65(.a(output_6_65), .b(output_6_2), .y(output_5_65));
wire output_7_65, output_7_2, output_6_65;
mixer gate_output_6_65(.a(output_7_65), .b(output_7_2), .y(output_6_65));
wire output_8_65, output_8_2, output_7_65;
mixer gate_output_7_65(.a(output_8_65), .b(output_8_2), .y(output_7_65));
wire output_9_65, output_9_2, output_8_65;
mixer gate_output_8_65(.a(output_9_65), .b(output_9_2), .y(output_8_65));
wire output_10_65, output_10_2, output_9_65;
mixer gate_output_9_65(.a(output_10_65), .b(output_10_2), .y(output_9_65));
wire output_11_65, output_11_2, output_10_65;
mixer gate_output_10_65(.a(output_11_65), .b(output_11_2), .y(output_10_65));
wire output_12_65, output_12_2, output_11_65;
mixer gate_output_11_65(.a(output_12_65), .b(output_12_2), .y(output_11_65));
wire output_13_65, output_13_2, output_12_65;
mixer gate_output_12_65(.a(output_13_65), .b(output_13_2), .y(output_12_65));
wire output_14_65, output_14_2, output_13_65;
mixer gate_output_13_65(.a(output_14_65), .b(output_14_2), .y(output_13_65));
wire output_15_65, output_15_2, output_14_65;
mixer gate_output_14_65(.a(output_15_65), .b(output_15_2), .y(output_14_65));
wire output_16_65, output_16_2, output_15_65;
mixer gate_output_15_65(.a(output_16_65), .b(output_16_2), .y(output_15_65));
wire output_1_66, output_1_3, output_0_66;
mixer gate_output_0_66(.a(output_1_66), .b(output_1_3), .y(output_0_66));
wire output_2_66, output_2_3, output_1_66;
mixer gate_output_1_66(.a(output_2_66), .b(output_2_3), .y(output_1_66));
wire output_3_66, output_3_3, output_2_66;
mixer gate_output_2_66(.a(output_3_66), .b(output_3_3), .y(output_2_66));
wire output_4_66, output_4_3, output_3_66;
mixer gate_output_3_66(.a(output_4_66), .b(output_4_3), .y(output_3_66));
wire output_5_66, output_5_3, output_4_66;
mixer gate_output_4_66(.a(output_5_66), .b(output_5_3), .y(output_4_66));
wire output_6_66, output_6_3, output_5_66;
mixer gate_output_5_66(.a(output_6_66), .b(output_6_3), .y(output_5_66));
wire output_7_66, output_7_3, output_6_66;
mixer gate_output_6_66(.a(output_7_66), .b(output_7_3), .y(output_6_66));
wire output_8_66, output_8_3, output_7_66;
mixer gate_output_7_66(.a(output_8_66), .b(output_8_3), .y(output_7_66));
wire output_9_66, output_9_3, output_8_66;
mixer gate_output_8_66(.a(output_9_66), .b(output_9_3), .y(output_8_66));
wire output_10_66, output_10_3, output_9_66;
mixer gate_output_9_66(.a(output_10_66), .b(output_10_3), .y(output_9_66));
wire output_11_66, output_11_3, output_10_66;
mixer gate_output_10_66(.a(output_11_66), .b(output_11_3), .y(output_10_66));
wire output_12_66, output_12_3, output_11_66;
mixer gate_output_11_66(.a(output_12_66), .b(output_12_3), .y(output_11_66));
wire output_13_66, output_13_3, output_12_66;
mixer gate_output_12_66(.a(output_13_66), .b(output_13_3), .y(output_12_66));
wire output_14_66, output_14_3, output_13_66;
mixer gate_output_13_66(.a(output_14_66), .b(output_14_3), .y(output_13_66));
wire output_15_66, output_15_3, output_14_66;
mixer gate_output_14_66(.a(output_15_66), .b(output_15_3), .y(output_14_66));
wire output_16_66, output_16_3, output_15_66;
mixer gate_output_15_66(.a(output_16_66), .b(output_16_3), .y(output_15_66));
wire output_1_67, output_1_4, output_0_67;
mixer gate_output_0_67(.a(output_1_67), .b(output_1_4), .y(output_0_67));
wire output_2_67, output_2_4, output_1_67;
mixer gate_output_1_67(.a(output_2_67), .b(output_2_4), .y(output_1_67));
wire output_3_67, output_3_4, output_2_67;
mixer gate_output_2_67(.a(output_3_67), .b(output_3_4), .y(output_2_67));
wire output_4_67, output_4_4, output_3_67;
mixer gate_output_3_67(.a(output_4_67), .b(output_4_4), .y(output_3_67));
wire output_5_67, output_5_4, output_4_67;
mixer gate_output_4_67(.a(output_5_67), .b(output_5_4), .y(output_4_67));
wire output_6_67, output_6_4, output_5_67;
mixer gate_output_5_67(.a(output_6_67), .b(output_6_4), .y(output_5_67));
wire output_7_67, output_7_4, output_6_67;
mixer gate_output_6_67(.a(output_7_67), .b(output_7_4), .y(output_6_67));
wire output_8_67, output_8_4, output_7_67;
mixer gate_output_7_67(.a(output_8_67), .b(output_8_4), .y(output_7_67));
wire output_9_67, output_9_4, output_8_67;
mixer gate_output_8_67(.a(output_9_67), .b(output_9_4), .y(output_8_67));
wire output_10_67, output_10_4, output_9_67;
mixer gate_output_9_67(.a(output_10_67), .b(output_10_4), .y(output_9_67));
wire output_11_67, output_11_4, output_10_67;
mixer gate_output_10_67(.a(output_11_67), .b(output_11_4), .y(output_10_67));
wire output_12_67, output_12_4, output_11_67;
mixer gate_output_11_67(.a(output_12_67), .b(output_12_4), .y(output_11_67));
wire output_13_67, output_13_4, output_12_67;
mixer gate_output_12_67(.a(output_13_67), .b(output_13_4), .y(output_12_67));
wire output_14_67, output_14_4, output_13_67;
mixer gate_output_13_67(.a(output_14_67), .b(output_14_4), .y(output_13_67));
wire output_15_67, output_15_4, output_14_67;
mixer gate_output_14_67(.a(output_15_67), .b(output_15_4), .y(output_14_67));
wire output_16_67, output_16_4, output_15_67;
mixer gate_output_15_67(.a(output_16_67), .b(output_16_4), .y(output_15_67));
wire output_1_68, output_1_5, output_0_68;
mixer gate_output_0_68(.a(output_1_68), .b(output_1_5), .y(output_0_68));
wire output_2_68, output_2_5, output_1_68;
mixer gate_output_1_68(.a(output_2_68), .b(output_2_5), .y(output_1_68));
wire output_3_68, output_3_5, output_2_68;
mixer gate_output_2_68(.a(output_3_68), .b(output_3_5), .y(output_2_68));
wire output_4_68, output_4_5, output_3_68;
mixer gate_output_3_68(.a(output_4_68), .b(output_4_5), .y(output_3_68));
wire output_5_68, output_5_5, output_4_68;
mixer gate_output_4_68(.a(output_5_68), .b(output_5_5), .y(output_4_68));
wire output_6_68, output_6_5, output_5_68;
mixer gate_output_5_68(.a(output_6_68), .b(output_6_5), .y(output_5_68));
wire output_7_68, output_7_5, output_6_68;
mixer gate_output_6_68(.a(output_7_68), .b(output_7_5), .y(output_6_68));
wire output_8_68, output_8_5, output_7_68;
mixer gate_output_7_68(.a(output_8_68), .b(output_8_5), .y(output_7_68));
wire output_9_68, output_9_5, output_8_68;
mixer gate_output_8_68(.a(output_9_68), .b(output_9_5), .y(output_8_68));
wire output_10_68, output_10_5, output_9_68;
mixer gate_output_9_68(.a(output_10_68), .b(output_10_5), .y(output_9_68));
wire output_11_68, output_11_5, output_10_68;
mixer gate_output_10_68(.a(output_11_68), .b(output_11_5), .y(output_10_68));
wire output_12_68, output_12_5, output_11_68;
mixer gate_output_11_68(.a(output_12_68), .b(output_12_5), .y(output_11_68));
wire output_13_68, output_13_5, output_12_68;
mixer gate_output_12_68(.a(output_13_68), .b(output_13_5), .y(output_12_68));
wire output_14_68, output_14_5, output_13_68;
mixer gate_output_13_68(.a(output_14_68), .b(output_14_5), .y(output_13_68));
wire output_15_68, output_15_5, output_14_68;
mixer gate_output_14_68(.a(output_15_68), .b(output_15_5), .y(output_14_68));
wire output_16_68, output_16_5, output_15_68;
mixer gate_output_15_68(.a(output_16_68), .b(output_16_5), .y(output_15_68));
wire output_1_69, output_1_6, output_0_69;
mixer gate_output_0_69(.a(output_1_69), .b(output_1_6), .y(output_0_69));
wire output_2_69, output_2_6, output_1_69;
mixer gate_output_1_69(.a(output_2_69), .b(output_2_6), .y(output_1_69));
wire output_3_69, output_3_6, output_2_69;
mixer gate_output_2_69(.a(output_3_69), .b(output_3_6), .y(output_2_69));
wire output_4_69, output_4_6, output_3_69;
mixer gate_output_3_69(.a(output_4_69), .b(output_4_6), .y(output_3_69));
wire output_5_69, output_5_6, output_4_69;
mixer gate_output_4_69(.a(output_5_69), .b(output_5_6), .y(output_4_69));
wire output_6_69, output_6_6, output_5_69;
mixer gate_output_5_69(.a(output_6_69), .b(output_6_6), .y(output_5_69));
wire output_7_69, output_7_6, output_6_69;
mixer gate_output_6_69(.a(output_7_69), .b(output_7_6), .y(output_6_69));
wire output_8_69, output_8_6, output_7_69;
mixer gate_output_7_69(.a(output_8_69), .b(output_8_6), .y(output_7_69));
wire output_9_69, output_9_6, output_8_69;
mixer gate_output_8_69(.a(output_9_69), .b(output_9_6), .y(output_8_69));
wire output_10_69, output_10_6, output_9_69;
mixer gate_output_9_69(.a(output_10_69), .b(output_10_6), .y(output_9_69));
wire output_11_69, output_11_6, output_10_69;
mixer gate_output_10_69(.a(output_11_69), .b(output_11_6), .y(output_10_69));
wire output_12_69, output_12_6, output_11_69;
mixer gate_output_11_69(.a(output_12_69), .b(output_12_6), .y(output_11_69));
wire output_13_69, output_13_6, output_12_69;
mixer gate_output_12_69(.a(output_13_69), .b(output_13_6), .y(output_12_69));
wire output_14_69, output_14_6, output_13_69;
mixer gate_output_13_69(.a(output_14_69), .b(output_14_6), .y(output_13_69));
wire output_15_69, output_15_6, output_14_69;
mixer gate_output_14_69(.a(output_15_69), .b(output_15_6), .y(output_14_69));
wire output_16_69, output_16_6, output_15_69;
mixer gate_output_15_69(.a(output_16_69), .b(output_16_6), .y(output_15_69));
wire output_1_70, output_1_7, output_0_70;
mixer gate_output_0_70(.a(output_1_70), .b(output_1_7), .y(output_0_70));
wire output_2_70, output_2_7, output_1_70;
mixer gate_output_1_70(.a(output_2_70), .b(output_2_7), .y(output_1_70));
wire output_3_70, output_3_7, output_2_70;
mixer gate_output_2_70(.a(output_3_70), .b(output_3_7), .y(output_2_70));
wire output_4_70, output_4_7, output_3_70;
mixer gate_output_3_70(.a(output_4_70), .b(output_4_7), .y(output_3_70));
wire output_5_70, output_5_7, output_4_70;
mixer gate_output_4_70(.a(output_5_70), .b(output_5_7), .y(output_4_70));
wire output_6_70, output_6_7, output_5_70;
mixer gate_output_5_70(.a(output_6_70), .b(output_6_7), .y(output_5_70));
wire output_7_70, output_7_7, output_6_70;
mixer gate_output_6_70(.a(output_7_70), .b(output_7_7), .y(output_6_70));
wire output_8_70, output_8_7, output_7_70;
mixer gate_output_7_70(.a(output_8_70), .b(output_8_7), .y(output_7_70));
wire output_9_70, output_9_7, output_8_70;
mixer gate_output_8_70(.a(output_9_70), .b(output_9_7), .y(output_8_70));
wire output_10_70, output_10_7, output_9_70;
mixer gate_output_9_70(.a(output_10_70), .b(output_10_7), .y(output_9_70));
wire output_11_70, output_11_7, output_10_70;
mixer gate_output_10_70(.a(output_11_70), .b(output_11_7), .y(output_10_70));
wire output_12_70, output_12_7, output_11_70;
mixer gate_output_11_70(.a(output_12_70), .b(output_12_7), .y(output_11_70));
wire output_13_70, output_13_7, output_12_70;
mixer gate_output_12_70(.a(output_13_70), .b(output_13_7), .y(output_12_70));
wire output_14_70, output_14_7, output_13_70;
mixer gate_output_13_70(.a(output_14_70), .b(output_14_7), .y(output_13_70));
wire output_15_70, output_15_7, output_14_70;
mixer gate_output_14_70(.a(output_15_70), .b(output_15_7), .y(output_14_70));
wire output_16_70, output_16_7, output_15_70;
mixer gate_output_15_70(.a(output_16_70), .b(output_16_7), .y(output_15_70));
wire output_1_71, output_1_8, output_0_71;
mixer gate_output_0_71(.a(output_1_71), .b(output_1_8), .y(output_0_71));
wire output_2_71, output_2_8, output_1_71;
mixer gate_output_1_71(.a(output_2_71), .b(output_2_8), .y(output_1_71));
wire output_3_71, output_3_8, output_2_71;
mixer gate_output_2_71(.a(output_3_71), .b(output_3_8), .y(output_2_71));
wire output_4_71, output_4_8, output_3_71;
mixer gate_output_3_71(.a(output_4_71), .b(output_4_8), .y(output_3_71));
wire output_5_71, output_5_8, output_4_71;
mixer gate_output_4_71(.a(output_5_71), .b(output_5_8), .y(output_4_71));
wire output_6_71, output_6_8, output_5_71;
mixer gate_output_5_71(.a(output_6_71), .b(output_6_8), .y(output_5_71));
wire output_7_71, output_7_8, output_6_71;
mixer gate_output_6_71(.a(output_7_71), .b(output_7_8), .y(output_6_71));
wire output_8_71, output_8_8, output_7_71;
mixer gate_output_7_71(.a(output_8_71), .b(output_8_8), .y(output_7_71));
wire output_9_71, output_9_8, output_8_71;
mixer gate_output_8_71(.a(output_9_71), .b(output_9_8), .y(output_8_71));
wire output_10_71, output_10_8, output_9_71;
mixer gate_output_9_71(.a(output_10_71), .b(output_10_8), .y(output_9_71));
wire output_11_71, output_11_8, output_10_71;
mixer gate_output_10_71(.a(output_11_71), .b(output_11_8), .y(output_10_71));
wire output_12_71, output_12_8, output_11_71;
mixer gate_output_11_71(.a(output_12_71), .b(output_12_8), .y(output_11_71));
wire output_13_71, output_13_8, output_12_71;
mixer gate_output_12_71(.a(output_13_71), .b(output_13_8), .y(output_12_71));
wire output_14_71, output_14_8, output_13_71;
mixer gate_output_13_71(.a(output_14_71), .b(output_14_8), .y(output_13_71));
wire output_15_71, output_15_8, output_14_71;
mixer gate_output_14_71(.a(output_15_71), .b(output_15_8), .y(output_14_71));
wire output_16_71, output_16_8, output_15_71;
mixer gate_output_15_71(.a(output_16_71), .b(output_16_8), .y(output_15_71));
wire output_1_72, output_1_9, output_0_72;
mixer gate_output_0_72(.a(output_1_72), .b(output_1_9), .y(output_0_72));
wire output_2_72, output_2_9, output_1_72;
mixer gate_output_1_72(.a(output_2_72), .b(output_2_9), .y(output_1_72));
wire output_3_72, output_3_9, output_2_72;
mixer gate_output_2_72(.a(output_3_72), .b(output_3_9), .y(output_2_72));
wire output_4_72, output_4_9, output_3_72;
mixer gate_output_3_72(.a(output_4_72), .b(output_4_9), .y(output_3_72));
wire output_5_72, output_5_9, output_4_72;
mixer gate_output_4_72(.a(output_5_72), .b(output_5_9), .y(output_4_72));
wire output_6_72, output_6_9, output_5_72;
mixer gate_output_5_72(.a(output_6_72), .b(output_6_9), .y(output_5_72));
wire output_7_72, output_7_9, output_6_72;
mixer gate_output_6_72(.a(output_7_72), .b(output_7_9), .y(output_6_72));
wire output_8_72, output_8_9, output_7_72;
mixer gate_output_7_72(.a(output_8_72), .b(output_8_9), .y(output_7_72));
wire output_9_72, output_9_9, output_8_72;
mixer gate_output_8_72(.a(output_9_72), .b(output_9_9), .y(output_8_72));
wire output_10_72, output_10_9, output_9_72;
mixer gate_output_9_72(.a(output_10_72), .b(output_10_9), .y(output_9_72));
wire output_11_72, output_11_9, output_10_72;
mixer gate_output_10_72(.a(output_11_72), .b(output_11_9), .y(output_10_72));
wire output_12_72, output_12_9, output_11_72;
mixer gate_output_11_72(.a(output_12_72), .b(output_12_9), .y(output_11_72));
wire output_13_72, output_13_9, output_12_72;
mixer gate_output_12_72(.a(output_13_72), .b(output_13_9), .y(output_12_72));
wire output_14_72, output_14_9, output_13_72;
mixer gate_output_13_72(.a(output_14_72), .b(output_14_9), .y(output_13_72));
wire output_15_72, output_15_9, output_14_72;
mixer gate_output_14_72(.a(output_15_72), .b(output_15_9), .y(output_14_72));
wire output_16_72, output_16_9, output_15_72;
mixer gate_output_15_72(.a(output_16_72), .b(output_16_9), .y(output_15_72));
wire output_1_73, output_1_10, output_0_73;
mixer gate_output_0_73(.a(output_1_73), .b(output_1_10), .y(output_0_73));
wire output_2_73, output_2_10, output_1_73;
mixer gate_output_1_73(.a(output_2_73), .b(output_2_10), .y(output_1_73));
wire output_3_73, output_3_10, output_2_73;
mixer gate_output_2_73(.a(output_3_73), .b(output_3_10), .y(output_2_73));
wire output_4_73, output_4_10, output_3_73;
mixer gate_output_3_73(.a(output_4_73), .b(output_4_10), .y(output_3_73));
wire output_5_73, output_5_10, output_4_73;
mixer gate_output_4_73(.a(output_5_73), .b(output_5_10), .y(output_4_73));
wire output_6_73, output_6_10, output_5_73;
mixer gate_output_5_73(.a(output_6_73), .b(output_6_10), .y(output_5_73));
wire output_7_73, output_7_10, output_6_73;
mixer gate_output_6_73(.a(output_7_73), .b(output_7_10), .y(output_6_73));
wire output_8_73, output_8_10, output_7_73;
mixer gate_output_7_73(.a(output_8_73), .b(output_8_10), .y(output_7_73));
wire output_9_73, output_9_10, output_8_73;
mixer gate_output_8_73(.a(output_9_73), .b(output_9_10), .y(output_8_73));
wire output_10_73, output_10_10, output_9_73;
mixer gate_output_9_73(.a(output_10_73), .b(output_10_10), .y(output_9_73));
wire output_11_73, output_11_10, output_10_73;
mixer gate_output_10_73(.a(output_11_73), .b(output_11_10), .y(output_10_73));
wire output_12_73, output_12_10, output_11_73;
mixer gate_output_11_73(.a(output_12_73), .b(output_12_10), .y(output_11_73));
wire output_13_73, output_13_10, output_12_73;
mixer gate_output_12_73(.a(output_13_73), .b(output_13_10), .y(output_12_73));
wire output_14_73, output_14_10, output_13_73;
mixer gate_output_13_73(.a(output_14_73), .b(output_14_10), .y(output_13_73));
wire output_15_73, output_15_10, output_14_73;
mixer gate_output_14_73(.a(output_15_73), .b(output_15_10), .y(output_14_73));
wire output_16_73, output_16_10, output_15_73;
mixer gate_output_15_73(.a(output_16_73), .b(output_16_10), .y(output_15_73));
wire output_1_74, output_1_11, output_0_74;
mixer gate_output_0_74(.a(output_1_74), .b(output_1_11), .y(output_0_74));
wire output_2_74, output_2_11, output_1_74;
mixer gate_output_1_74(.a(output_2_74), .b(output_2_11), .y(output_1_74));
wire output_3_74, output_3_11, output_2_74;
mixer gate_output_2_74(.a(output_3_74), .b(output_3_11), .y(output_2_74));
wire output_4_74, output_4_11, output_3_74;
mixer gate_output_3_74(.a(output_4_74), .b(output_4_11), .y(output_3_74));
wire output_5_74, output_5_11, output_4_74;
mixer gate_output_4_74(.a(output_5_74), .b(output_5_11), .y(output_4_74));
wire output_6_74, output_6_11, output_5_74;
mixer gate_output_5_74(.a(output_6_74), .b(output_6_11), .y(output_5_74));
wire output_7_74, output_7_11, output_6_74;
mixer gate_output_6_74(.a(output_7_74), .b(output_7_11), .y(output_6_74));
wire output_8_74, output_8_11, output_7_74;
mixer gate_output_7_74(.a(output_8_74), .b(output_8_11), .y(output_7_74));
wire output_9_74, output_9_11, output_8_74;
mixer gate_output_8_74(.a(output_9_74), .b(output_9_11), .y(output_8_74));
wire output_10_74, output_10_11, output_9_74;
mixer gate_output_9_74(.a(output_10_74), .b(output_10_11), .y(output_9_74));
wire output_11_74, output_11_11, output_10_74;
mixer gate_output_10_74(.a(output_11_74), .b(output_11_11), .y(output_10_74));
wire output_12_74, output_12_11, output_11_74;
mixer gate_output_11_74(.a(output_12_74), .b(output_12_11), .y(output_11_74));
wire output_13_74, output_13_11, output_12_74;
mixer gate_output_12_74(.a(output_13_74), .b(output_13_11), .y(output_12_74));
wire output_14_74, output_14_11, output_13_74;
mixer gate_output_13_74(.a(output_14_74), .b(output_14_11), .y(output_13_74));
wire output_15_74, output_15_11, output_14_74;
mixer gate_output_14_74(.a(output_15_74), .b(output_15_11), .y(output_14_74));
wire output_16_74, output_16_11, output_15_74;
mixer gate_output_15_74(.a(output_16_74), .b(output_16_11), .y(output_15_74));
wire output_1_75, output_1_12, output_0_75;
mixer gate_output_0_75(.a(output_1_75), .b(output_1_12), .y(output_0_75));
wire output_2_75, output_2_12, output_1_75;
mixer gate_output_1_75(.a(output_2_75), .b(output_2_12), .y(output_1_75));
wire output_3_75, output_3_12, output_2_75;
mixer gate_output_2_75(.a(output_3_75), .b(output_3_12), .y(output_2_75));
wire output_4_75, output_4_12, output_3_75;
mixer gate_output_3_75(.a(output_4_75), .b(output_4_12), .y(output_3_75));
wire output_5_75, output_5_12, output_4_75;
mixer gate_output_4_75(.a(output_5_75), .b(output_5_12), .y(output_4_75));
wire output_6_75, output_6_12, output_5_75;
mixer gate_output_5_75(.a(output_6_75), .b(output_6_12), .y(output_5_75));
wire output_7_75, output_7_12, output_6_75;
mixer gate_output_6_75(.a(output_7_75), .b(output_7_12), .y(output_6_75));
wire output_8_75, output_8_12, output_7_75;
mixer gate_output_7_75(.a(output_8_75), .b(output_8_12), .y(output_7_75));
wire output_9_75, output_9_12, output_8_75;
mixer gate_output_8_75(.a(output_9_75), .b(output_9_12), .y(output_8_75));
wire output_10_75, output_10_12, output_9_75;
mixer gate_output_9_75(.a(output_10_75), .b(output_10_12), .y(output_9_75));
wire output_11_75, output_11_12, output_10_75;
mixer gate_output_10_75(.a(output_11_75), .b(output_11_12), .y(output_10_75));
wire output_12_75, output_12_12, output_11_75;
mixer gate_output_11_75(.a(output_12_75), .b(output_12_12), .y(output_11_75));
wire output_13_75, output_13_12, output_12_75;
mixer gate_output_12_75(.a(output_13_75), .b(output_13_12), .y(output_12_75));
wire output_14_75, output_14_12, output_13_75;
mixer gate_output_13_75(.a(output_14_75), .b(output_14_12), .y(output_13_75));
wire output_15_75, output_15_12, output_14_75;
mixer gate_output_14_75(.a(output_15_75), .b(output_15_12), .y(output_14_75));
wire output_16_75, output_16_12, output_15_75;
mixer gate_output_15_75(.a(output_16_75), .b(output_16_12), .y(output_15_75));
wire output_1_76, output_1_13, output_0_76;
mixer gate_output_0_76(.a(output_1_76), .b(output_1_13), .y(output_0_76));
wire output_2_76, output_2_13, output_1_76;
mixer gate_output_1_76(.a(output_2_76), .b(output_2_13), .y(output_1_76));
wire output_3_76, output_3_13, output_2_76;
mixer gate_output_2_76(.a(output_3_76), .b(output_3_13), .y(output_2_76));
wire output_4_76, output_4_13, output_3_76;
mixer gate_output_3_76(.a(output_4_76), .b(output_4_13), .y(output_3_76));
wire output_5_76, output_5_13, output_4_76;
mixer gate_output_4_76(.a(output_5_76), .b(output_5_13), .y(output_4_76));
wire output_6_76, output_6_13, output_5_76;
mixer gate_output_5_76(.a(output_6_76), .b(output_6_13), .y(output_5_76));
wire output_7_76, output_7_13, output_6_76;
mixer gate_output_6_76(.a(output_7_76), .b(output_7_13), .y(output_6_76));
wire output_8_76, output_8_13, output_7_76;
mixer gate_output_7_76(.a(output_8_76), .b(output_8_13), .y(output_7_76));
wire output_9_76, output_9_13, output_8_76;
mixer gate_output_8_76(.a(output_9_76), .b(output_9_13), .y(output_8_76));
wire output_10_76, output_10_13, output_9_76;
mixer gate_output_9_76(.a(output_10_76), .b(output_10_13), .y(output_9_76));
wire output_11_76, output_11_13, output_10_76;
mixer gate_output_10_76(.a(output_11_76), .b(output_11_13), .y(output_10_76));
wire output_12_76, output_12_13, output_11_76;
mixer gate_output_11_76(.a(output_12_76), .b(output_12_13), .y(output_11_76));
wire output_13_76, output_13_13, output_12_76;
mixer gate_output_12_76(.a(output_13_76), .b(output_13_13), .y(output_12_76));
wire output_14_76, output_14_13, output_13_76;
mixer gate_output_13_76(.a(output_14_76), .b(output_14_13), .y(output_13_76));
wire output_15_76, output_15_13, output_14_76;
mixer gate_output_14_76(.a(output_15_76), .b(output_15_13), .y(output_14_76));
wire output_16_76, output_16_13, output_15_76;
mixer gate_output_15_76(.a(output_16_76), .b(output_16_13), .y(output_15_76));
wire output_1_77, output_1_14, output_0_77;
mixer gate_output_0_77(.a(output_1_77), .b(output_1_14), .y(output_0_77));
wire output_2_77, output_2_14, output_1_77;
mixer gate_output_1_77(.a(output_2_77), .b(output_2_14), .y(output_1_77));
wire output_3_77, output_3_14, output_2_77;
mixer gate_output_2_77(.a(output_3_77), .b(output_3_14), .y(output_2_77));
wire output_4_77, output_4_14, output_3_77;
mixer gate_output_3_77(.a(output_4_77), .b(output_4_14), .y(output_3_77));
wire output_5_77, output_5_14, output_4_77;
mixer gate_output_4_77(.a(output_5_77), .b(output_5_14), .y(output_4_77));
wire output_6_77, output_6_14, output_5_77;
mixer gate_output_5_77(.a(output_6_77), .b(output_6_14), .y(output_5_77));
wire output_7_77, output_7_14, output_6_77;
mixer gate_output_6_77(.a(output_7_77), .b(output_7_14), .y(output_6_77));
wire output_8_77, output_8_14, output_7_77;
mixer gate_output_7_77(.a(output_8_77), .b(output_8_14), .y(output_7_77));
wire output_9_77, output_9_14, output_8_77;
mixer gate_output_8_77(.a(output_9_77), .b(output_9_14), .y(output_8_77));
wire output_10_77, output_10_14, output_9_77;
mixer gate_output_9_77(.a(output_10_77), .b(output_10_14), .y(output_9_77));
wire output_11_77, output_11_14, output_10_77;
mixer gate_output_10_77(.a(output_11_77), .b(output_11_14), .y(output_10_77));
wire output_12_77, output_12_14, output_11_77;
mixer gate_output_11_77(.a(output_12_77), .b(output_12_14), .y(output_11_77));
wire output_13_77, output_13_14, output_12_77;
mixer gate_output_12_77(.a(output_13_77), .b(output_13_14), .y(output_12_77));
wire output_14_77, output_14_14, output_13_77;
mixer gate_output_13_77(.a(output_14_77), .b(output_14_14), .y(output_13_77));
wire output_15_77, output_15_14, output_14_77;
mixer gate_output_14_77(.a(output_15_77), .b(output_15_14), .y(output_14_77));
wire output_16_77, output_16_14, output_15_77;
mixer gate_output_15_77(.a(output_16_77), .b(output_16_14), .y(output_15_77));
wire output_1_78, output_1_15, output_0_78;
mixer gate_output_0_78(.a(output_1_78), .b(output_1_15), .y(output_0_78));
wire output_2_78, output_2_15, output_1_78;
mixer gate_output_1_78(.a(output_2_78), .b(output_2_15), .y(output_1_78));
wire output_3_78, output_3_15, output_2_78;
mixer gate_output_2_78(.a(output_3_78), .b(output_3_15), .y(output_2_78));
wire output_4_78, output_4_15, output_3_78;
mixer gate_output_3_78(.a(output_4_78), .b(output_4_15), .y(output_3_78));
wire output_5_78, output_5_15, output_4_78;
mixer gate_output_4_78(.a(output_5_78), .b(output_5_15), .y(output_4_78));
wire output_6_78, output_6_15, output_5_78;
mixer gate_output_5_78(.a(output_6_78), .b(output_6_15), .y(output_5_78));
wire output_7_78, output_7_15, output_6_78;
mixer gate_output_6_78(.a(output_7_78), .b(output_7_15), .y(output_6_78));
wire output_8_78, output_8_15, output_7_78;
mixer gate_output_7_78(.a(output_8_78), .b(output_8_15), .y(output_7_78));
wire output_9_78, output_9_15, output_8_78;
mixer gate_output_8_78(.a(output_9_78), .b(output_9_15), .y(output_8_78));
wire output_10_78, output_10_15, output_9_78;
mixer gate_output_9_78(.a(output_10_78), .b(output_10_15), .y(output_9_78));
wire output_11_78, output_11_15, output_10_78;
mixer gate_output_10_78(.a(output_11_78), .b(output_11_15), .y(output_10_78));
wire output_12_78, output_12_15, output_11_78;
mixer gate_output_11_78(.a(output_12_78), .b(output_12_15), .y(output_11_78));
wire output_13_78, output_13_15, output_12_78;
mixer gate_output_12_78(.a(output_13_78), .b(output_13_15), .y(output_12_78));
wire output_14_78, output_14_15, output_13_78;
mixer gate_output_13_78(.a(output_14_78), .b(output_14_15), .y(output_13_78));
wire output_15_78, output_15_15, output_14_78;
mixer gate_output_14_78(.a(output_15_78), .b(output_15_15), .y(output_14_78));
wire output_16_78, output_16_15, output_15_78;
mixer gate_output_15_78(.a(output_16_78), .b(output_16_15), .y(output_15_78));
wire output_1_79, output_1_0, output_0_79;
mixer gate_output_0_79(.a(output_1_79), .b(output_1_0), .y(output_0_79));
wire output_2_79, output_2_0, output_1_79;
mixer gate_output_1_79(.a(output_2_79), .b(output_2_0), .y(output_1_79));
wire output_3_79, output_3_0, output_2_79;
mixer gate_output_2_79(.a(output_3_79), .b(output_3_0), .y(output_2_79));
wire output_4_79, output_4_0, output_3_79;
mixer gate_output_3_79(.a(output_4_79), .b(output_4_0), .y(output_3_79));
wire output_5_79, output_5_0, output_4_79;
mixer gate_output_4_79(.a(output_5_79), .b(output_5_0), .y(output_4_79));
wire output_6_79, output_6_0, output_5_79;
mixer gate_output_5_79(.a(output_6_79), .b(output_6_0), .y(output_5_79));
wire output_7_79, output_7_0, output_6_79;
mixer gate_output_6_79(.a(output_7_79), .b(output_7_0), .y(output_6_79));
wire output_8_79, output_8_0, output_7_79;
mixer gate_output_7_79(.a(output_8_79), .b(output_8_0), .y(output_7_79));
wire output_9_79, output_9_0, output_8_79;
mixer gate_output_8_79(.a(output_9_79), .b(output_9_0), .y(output_8_79));
wire output_10_79, output_10_0, output_9_79;
mixer gate_output_9_79(.a(output_10_79), .b(output_10_0), .y(output_9_79));
wire output_11_79, output_11_0, output_10_79;
mixer gate_output_10_79(.a(output_11_79), .b(output_11_0), .y(output_10_79));
wire output_12_79, output_12_0, output_11_79;
mixer gate_output_11_79(.a(output_12_79), .b(output_12_0), .y(output_11_79));
wire output_13_79, output_13_0, output_12_79;
mixer gate_output_12_79(.a(output_13_79), .b(output_13_0), .y(output_12_79));
wire output_14_79, output_14_0, output_13_79;
mixer gate_output_13_79(.a(output_14_79), .b(output_14_0), .y(output_13_79));
wire output_15_79, output_15_0, output_14_79;
mixer gate_output_14_79(.a(output_15_79), .b(output_15_0), .y(output_14_79));
wire output_16_79, output_16_0, output_15_79;
mixer gate_output_15_79(.a(output_16_79), .b(output_16_0), .y(output_15_79));
wire output_1_80, output_1_1, output_0_80;
mixer gate_output_0_80(.a(output_1_80), .b(output_1_1), .y(output_0_80));
wire output_2_80, output_2_1, output_1_80;
mixer gate_output_1_80(.a(output_2_80), .b(output_2_1), .y(output_1_80));
wire output_3_80, output_3_1, output_2_80;
mixer gate_output_2_80(.a(output_3_80), .b(output_3_1), .y(output_2_80));
wire output_4_80, output_4_1, output_3_80;
mixer gate_output_3_80(.a(output_4_80), .b(output_4_1), .y(output_3_80));
wire output_5_80, output_5_1, output_4_80;
mixer gate_output_4_80(.a(output_5_80), .b(output_5_1), .y(output_4_80));
wire output_6_80, output_6_1, output_5_80;
mixer gate_output_5_80(.a(output_6_80), .b(output_6_1), .y(output_5_80));
wire output_7_80, output_7_1, output_6_80;
mixer gate_output_6_80(.a(output_7_80), .b(output_7_1), .y(output_6_80));
wire output_8_80, output_8_1, output_7_80;
mixer gate_output_7_80(.a(output_8_80), .b(output_8_1), .y(output_7_80));
wire output_9_80, output_9_1, output_8_80;
mixer gate_output_8_80(.a(output_9_80), .b(output_9_1), .y(output_8_80));
wire output_10_80, output_10_1, output_9_80;
mixer gate_output_9_80(.a(output_10_80), .b(output_10_1), .y(output_9_80));
wire output_11_80, output_11_1, output_10_80;
mixer gate_output_10_80(.a(output_11_80), .b(output_11_1), .y(output_10_80));
wire output_12_80, output_12_1, output_11_80;
mixer gate_output_11_80(.a(output_12_80), .b(output_12_1), .y(output_11_80));
wire output_13_80, output_13_1, output_12_80;
mixer gate_output_12_80(.a(output_13_80), .b(output_13_1), .y(output_12_80));
wire output_14_80, output_14_1, output_13_80;
mixer gate_output_13_80(.a(output_14_80), .b(output_14_1), .y(output_13_80));
wire output_15_80, output_15_1, output_14_80;
mixer gate_output_14_80(.a(output_15_80), .b(output_15_1), .y(output_14_80));
wire output_16_80, output_16_1, output_15_80;
mixer gate_output_15_80(.a(output_16_80), .b(output_16_1), .y(output_15_80));
wire output_1_81, output_1_2, output_0_81;
mixer gate_output_0_81(.a(output_1_81), .b(output_1_2), .y(output_0_81));
wire output_2_81, output_2_2, output_1_81;
mixer gate_output_1_81(.a(output_2_81), .b(output_2_2), .y(output_1_81));
wire output_3_81, output_3_2, output_2_81;
mixer gate_output_2_81(.a(output_3_81), .b(output_3_2), .y(output_2_81));
wire output_4_81, output_4_2, output_3_81;
mixer gate_output_3_81(.a(output_4_81), .b(output_4_2), .y(output_3_81));
wire output_5_81, output_5_2, output_4_81;
mixer gate_output_4_81(.a(output_5_81), .b(output_5_2), .y(output_4_81));
wire output_6_81, output_6_2, output_5_81;
mixer gate_output_5_81(.a(output_6_81), .b(output_6_2), .y(output_5_81));
wire output_7_81, output_7_2, output_6_81;
mixer gate_output_6_81(.a(output_7_81), .b(output_7_2), .y(output_6_81));
wire output_8_81, output_8_2, output_7_81;
mixer gate_output_7_81(.a(output_8_81), .b(output_8_2), .y(output_7_81));
wire output_9_81, output_9_2, output_8_81;
mixer gate_output_8_81(.a(output_9_81), .b(output_9_2), .y(output_8_81));
wire output_10_81, output_10_2, output_9_81;
mixer gate_output_9_81(.a(output_10_81), .b(output_10_2), .y(output_9_81));
wire output_11_81, output_11_2, output_10_81;
mixer gate_output_10_81(.a(output_11_81), .b(output_11_2), .y(output_10_81));
wire output_12_81, output_12_2, output_11_81;
mixer gate_output_11_81(.a(output_12_81), .b(output_12_2), .y(output_11_81));
wire output_13_81, output_13_2, output_12_81;
mixer gate_output_12_81(.a(output_13_81), .b(output_13_2), .y(output_12_81));
wire output_14_81, output_14_2, output_13_81;
mixer gate_output_13_81(.a(output_14_81), .b(output_14_2), .y(output_13_81));
wire output_15_81, output_15_2, output_14_81;
mixer gate_output_14_81(.a(output_15_81), .b(output_15_2), .y(output_14_81));
wire output_16_81, output_16_2, output_15_81;
mixer gate_output_15_81(.a(output_16_81), .b(output_16_2), .y(output_15_81));
wire output_1_82, output_1_3, output_0_82;
mixer gate_output_0_82(.a(output_1_82), .b(output_1_3), .y(output_0_82));
wire output_2_82, output_2_3, output_1_82;
mixer gate_output_1_82(.a(output_2_82), .b(output_2_3), .y(output_1_82));
wire output_3_82, output_3_3, output_2_82;
mixer gate_output_2_82(.a(output_3_82), .b(output_3_3), .y(output_2_82));
wire output_4_82, output_4_3, output_3_82;
mixer gate_output_3_82(.a(output_4_82), .b(output_4_3), .y(output_3_82));
wire output_5_82, output_5_3, output_4_82;
mixer gate_output_4_82(.a(output_5_82), .b(output_5_3), .y(output_4_82));
wire output_6_82, output_6_3, output_5_82;
mixer gate_output_5_82(.a(output_6_82), .b(output_6_3), .y(output_5_82));
wire output_7_82, output_7_3, output_6_82;
mixer gate_output_6_82(.a(output_7_82), .b(output_7_3), .y(output_6_82));
wire output_8_82, output_8_3, output_7_82;
mixer gate_output_7_82(.a(output_8_82), .b(output_8_3), .y(output_7_82));
wire output_9_82, output_9_3, output_8_82;
mixer gate_output_8_82(.a(output_9_82), .b(output_9_3), .y(output_8_82));
wire output_10_82, output_10_3, output_9_82;
mixer gate_output_9_82(.a(output_10_82), .b(output_10_3), .y(output_9_82));
wire output_11_82, output_11_3, output_10_82;
mixer gate_output_10_82(.a(output_11_82), .b(output_11_3), .y(output_10_82));
wire output_12_82, output_12_3, output_11_82;
mixer gate_output_11_82(.a(output_12_82), .b(output_12_3), .y(output_11_82));
wire output_13_82, output_13_3, output_12_82;
mixer gate_output_12_82(.a(output_13_82), .b(output_13_3), .y(output_12_82));
wire output_14_82, output_14_3, output_13_82;
mixer gate_output_13_82(.a(output_14_82), .b(output_14_3), .y(output_13_82));
wire output_15_82, output_15_3, output_14_82;
mixer gate_output_14_82(.a(output_15_82), .b(output_15_3), .y(output_14_82));
wire output_16_82, output_16_3, output_15_82;
mixer gate_output_15_82(.a(output_16_82), .b(output_16_3), .y(output_15_82));
wire output_1_83, output_1_4, output_0_83;
mixer gate_output_0_83(.a(output_1_83), .b(output_1_4), .y(output_0_83));
wire output_2_83, output_2_4, output_1_83;
mixer gate_output_1_83(.a(output_2_83), .b(output_2_4), .y(output_1_83));
wire output_3_83, output_3_4, output_2_83;
mixer gate_output_2_83(.a(output_3_83), .b(output_3_4), .y(output_2_83));
wire output_4_83, output_4_4, output_3_83;
mixer gate_output_3_83(.a(output_4_83), .b(output_4_4), .y(output_3_83));
wire output_5_83, output_5_4, output_4_83;
mixer gate_output_4_83(.a(output_5_83), .b(output_5_4), .y(output_4_83));
wire output_6_83, output_6_4, output_5_83;
mixer gate_output_5_83(.a(output_6_83), .b(output_6_4), .y(output_5_83));
wire output_7_83, output_7_4, output_6_83;
mixer gate_output_6_83(.a(output_7_83), .b(output_7_4), .y(output_6_83));
wire output_8_83, output_8_4, output_7_83;
mixer gate_output_7_83(.a(output_8_83), .b(output_8_4), .y(output_7_83));
wire output_9_83, output_9_4, output_8_83;
mixer gate_output_8_83(.a(output_9_83), .b(output_9_4), .y(output_8_83));
wire output_10_83, output_10_4, output_9_83;
mixer gate_output_9_83(.a(output_10_83), .b(output_10_4), .y(output_9_83));
wire output_11_83, output_11_4, output_10_83;
mixer gate_output_10_83(.a(output_11_83), .b(output_11_4), .y(output_10_83));
wire output_12_83, output_12_4, output_11_83;
mixer gate_output_11_83(.a(output_12_83), .b(output_12_4), .y(output_11_83));
wire output_13_83, output_13_4, output_12_83;
mixer gate_output_12_83(.a(output_13_83), .b(output_13_4), .y(output_12_83));
wire output_14_83, output_14_4, output_13_83;
mixer gate_output_13_83(.a(output_14_83), .b(output_14_4), .y(output_13_83));
wire output_15_83, output_15_4, output_14_83;
mixer gate_output_14_83(.a(output_15_83), .b(output_15_4), .y(output_14_83));
wire output_16_83, output_16_4, output_15_83;
mixer gate_output_15_83(.a(output_16_83), .b(output_16_4), .y(output_15_83));
wire output_1_84, output_1_5, output_0_84;
mixer gate_output_0_84(.a(output_1_84), .b(output_1_5), .y(output_0_84));
wire output_2_84, output_2_5, output_1_84;
mixer gate_output_1_84(.a(output_2_84), .b(output_2_5), .y(output_1_84));
wire output_3_84, output_3_5, output_2_84;
mixer gate_output_2_84(.a(output_3_84), .b(output_3_5), .y(output_2_84));
wire output_4_84, output_4_5, output_3_84;
mixer gate_output_3_84(.a(output_4_84), .b(output_4_5), .y(output_3_84));
wire output_5_84, output_5_5, output_4_84;
mixer gate_output_4_84(.a(output_5_84), .b(output_5_5), .y(output_4_84));
wire output_6_84, output_6_5, output_5_84;
mixer gate_output_5_84(.a(output_6_84), .b(output_6_5), .y(output_5_84));
wire output_7_84, output_7_5, output_6_84;
mixer gate_output_6_84(.a(output_7_84), .b(output_7_5), .y(output_6_84));
wire output_8_84, output_8_5, output_7_84;
mixer gate_output_7_84(.a(output_8_84), .b(output_8_5), .y(output_7_84));
wire output_9_84, output_9_5, output_8_84;
mixer gate_output_8_84(.a(output_9_84), .b(output_9_5), .y(output_8_84));
wire output_10_84, output_10_5, output_9_84;
mixer gate_output_9_84(.a(output_10_84), .b(output_10_5), .y(output_9_84));
wire output_11_84, output_11_5, output_10_84;
mixer gate_output_10_84(.a(output_11_84), .b(output_11_5), .y(output_10_84));
wire output_12_84, output_12_5, output_11_84;
mixer gate_output_11_84(.a(output_12_84), .b(output_12_5), .y(output_11_84));
wire output_13_84, output_13_5, output_12_84;
mixer gate_output_12_84(.a(output_13_84), .b(output_13_5), .y(output_12_84));
wire output_14_84, output_14_5, output_13_84;
mixer gate_output_13_84(.a(output_14_84), .b(output_14_5), .y(output_13_84));
wire output_15_84, output_15_5, output_14_84;
mixer gate_output_14_84(.a(output_15_84), .b(output_15_5), .y(output_14_84));
wire output_16_84, output_16_5, output_15_84;
mixer gate_output_15_84(.a(output_16_84), .b(output_16_5), .y(output_15_84));
wire output_1_85, output_1_6, output_0_85;
mixer gate_output_0_85(.a(output_1_85), .b(output_1_6), .y(output_0_85));
wire output_2_85, output_2_6, output_1_85;
mixer gate_output_1_85(.a(output_2_85), .b(output_2_6), .y(output_1_85));
wire output_3_85, output_3_6, output_2_85;
mixer gate_output_2_85(.a(output_3_85), .b(output_3_6), .y(output_2_85));
wire output_4_85, output_4_6, output_3_85;
mixer gate_output_3_85(.a(output_4_85), .b(output_4_6), .y(output_3_85));
wire output_5_85, output_5_6, output_4_85;
mixer gate_output_4_85(.a(output_5_85), .b(output_5_6), .y(output_4_85));
wire output_6_85, output_6_6, output_5_85;
mixer gate_output_5_85(.a(output_6_85), .b(output_6_6), .y(output_5_85));
wire output_7_85, output_7_6, output_6_85;
mixer gate_output_6_85(.a(output_7_85), .b(output_7_6), .y(output_6_85));
wire output_8_85, output_8_6, output_7_85;
mixer gate_output_7_85(.a(output_8_85), .b(output_8_6), .y(output_7_85));
wire output_9_85, output_9_6, output_8_85;
mixer gate_output_8_85(.a(output_9_85), .b(output_9_6), .y(output_8_85));
wire output_10_85, output_10_6, output_9_85;
mixer gate_output_9_85(.a(output_10_85), .b(output_10_6), .y(output_9_85));
wire output_11_85, output_11_6, output_10_85;
mixer gate_output_10_85(.a(output_11_85), .b(output_11_6), .y(output_10_85));
wire output_12_85, output_12_6, output_11_85;
mixer gate_output_11_85(.a(output_12_85), .b(output_12_6), .y(output_11_85));
wire output_13_85, output_13_6, output_12_85;
mixer gate_output_12_85(.a(output_13_85), .b(output_13_6), .y(output_12_85));
wire output_14_85, output_14_6, output_13_85;
mixer gate_output_13_85(.a(output_14_85), .b(output_14_6), .y(output_13_85));
wire output_15_85, output_15_6, output_14_85;
mixer gate_output_14_85(.a(output_15_85), .b(output_15_6), .y(output_14_85));
wire output_16_85, output_16_6, output_15_85;
mixer gate_output_15_85(.a(output_16_85), .b(output_16_6), .y(output_15_85));
wire output_1_86, output_1_7, output_0_86;
mixer gate_output_0_86(.a(output_1_86), .b(output_1_7), .y(output_0_86));
wire output_2_86, output_2_7, output_1_86;
mixer gate_output_1_86(.a(output_2_86), .b(output_2_7), .y(output_1_86));
wire output_3_86, output_3_7, output_2_86;
mixer gate_output_2_86(.a(output_3_86), .b(output_3_7), .y(output_2_86));
wire output_4_86, output_4_7, output_3_86;
mixer gate_output_3_86(.a(output_4_86), .b(output_4_7), .y(output_3_86));
wire output_5_86, output_5_7, output_4_86;
mixer gate_output_4_86(.a(output_5_86), .b(output_5_7), .y(output_4_86));
wire output_6_86, output_6_7, output_5_86;
mixer gate_output_5_86(.a(output_6_86), .b(output_6_7), .y(output_5_86));
wire output_7_86, output_7_7, output_6_86;
mixer gate_output_6_86(.a(output_7_86), .b(output_7_7), .y(output_6_86));
wire output_8_86, output_8_7, output_7_86;
mixer gate_output_7_86(.a(output_8_86), .b(output_8_7), .y(output_7_86));
wire output_9_86, output_9_7, output_8_86;
mixer gate_output_8_86(.a(output_9_86), .b(output_9_7), .y(output_8_86));
wire output_10_86, output_10_7, output_9_86;
mixer gate_output_9_86(.a(output_10_86), .b(output_10_7), .y(output_9_86));
wire output_11_86, output_11_7, output_10_86;
mixer gate_output_10_86(.a(output_11_86), .b(output_11_7), .y(output_10_86));
wire output_12_86, output_12_7, output_11_86;
mixer gate_output_11_86(.a(output_12_86), .b(output_12_7), .y(output_11_86));
wire output_13_86, output_13_7, output_12_86;
mixer gate_output_12_86(.a(output_13_86), .b(output_13_7), .y(output_12_86));
wire output_14_86, output_14_7, output_13_86;
mixer gate_output_13_86(.a(output_14_86), .b(output_14_7), .y(output_13_86));
wire output_15_86, output_15_7, output_14_86;
mixer gate_output_14_86(.a(output_15_86), .b(output_15_7), .y(output_14_86));
wire output_16_86, output_16_7, output_15_86;
mixer gate_output_15_86(.a(output_16_86), .b(output_16_7), .y(output_15_86));
wire output_1_87, output_1_8, output_0_87;
mixer gate_output_0_87(.a(output_1_87), .b(output_1_8), .y(output_0_87));
wire output_2_87, output_2_8, output_1_87;
mixer gate_output_1_87(.a(output_2_87), .b(output_2_8), .y(output_1_87));
wire output_3_87, output_3_8, output_2_87;
mixer gate_output_2_87(.a(output_3_87), .b(output_3_8), .y(output_2_87));
wire output_4_87, output_4_8, output_3_87;
mixer gate_output_3_87(.a(output_4_87), .b(output_4_8), .y(output_3_87));
wire output_5_87, output_5_8, output_4_87;
mixer gate_output_4_87(.a(output_5_87), .b(output_5_8), .y(output_4_87));
wire output_6_87, output_6_8, output_5_87;
mixer gate_output_5_87(.a(output_6_87), .b(output_6_8), .y(output_5_87));
wire output_7_87, output_7_8, output_6_87;
mixer gate_output_6_87(.a(output_7_87), .b(output_7_8), .y(output_6_87));
wire output_8_87, output_8_8, output_7_87;
mixer gate_output_7_87(.a(output_8_87), .b(output_8_8), .y(output_7_87));
wire output_9_87, output_9_8, output_8_87;
mixer gate_output_8_87(.a(output_9_87), .b(output_9_8), .y(output_8_87));
wire output_10_87, output_10_8, output_9_87;
mixer gate_output_9_87(.a(output_10_87), .b(output_10_8), .y(output_9_87));
wire output_11_87, output_11_8, output_10_87;
mixer gate_output_10_87(.a(output_11_87), .b(output_11_8), .y(output_10_87));
wire output_12_87, output_12_8, output_11_87;
mixer gate_output_11_87(.a(output_12_87), .b(output_12_8), .y(output_11_87));
wire output_13_87, output_13_8, output_12_87;
mixer gate_output_12_87(.a(output_13_87), .b(output_13_8), .y(output_12_87));
wire output_14_87, output_14_8, output_13_87;
mixer gate_output_13_87(.a(output_14_87), .b(output_14_8), .y(output_13_87));
wire output_15_87, output_15_8, output_14_87;
mixer gate_output_14_87(.a(output_15_87), .b(output_15_8), .y(output_14_87));
wire output_16_87, output_16_8, output_15_87;
mixer gate_output_15_87(.a(output_16_87), .b(output_16_8), .y(output_15_87));
wire output_1_88, output_1_9, output_0_88;
mixer gate_output_0_88(.a(output_1_88), .b(output_1_9), .y(output_0_88));
wire output_2_88, output_2_9, output_1_88;
mixer gate_output_1_88(.a(output_2_88), .b(output_2_9), .y(output_1_88));
wire output_3_88, output_3_9, output_2_88;
mixer gate_output_2_88(.a(output_3_88), .b(output_3_9), .y(output_2_88));
wire output_4_88, output_4_9, output_3_88;
mixer gate_output_3_88(.a(output_4_88), .b(output_4_9), .y(output_3_88));
wire output_5_88, output_5_9, output_4_88;
mixer gate_output_4_88(.a(output_5_88), .b(output_5_9), .y(output_4_88));
wire output_6_88, output_6_9, output_5_88;
mixer gate_output_5_88(.a(output_6_88), .b(output_6_9), .y(output_5_88));
wire output_7_88, output_7_9, output_6_88;
mixer gate_output_6_88(.a(output_7_88), .b(output_7_9), .y(output_6_88));
wire output_8_88, output_8_9, output_7_88;
mixer gate_output_7_88(.a(output_8_88), .b(output_8_9), .y(output_7_88));
wire output_9_88, output_9_9, output_8_88;
mixer gate_output_8_88(.a(output_9_88), .b(output_9_9), .y(output_8_88));
wire output_10_88, output_10_9, output_9_88;
mixer gate_output_9_88(.a(output_10_88), .b(output_10_9), .y(output_9_88));
wire output_11_88, output_11_9, output_10_88;
mixer gate_output_10_88(.a(output_11_88), .b(output_11_9), .y(output_10_88));
wire output_12_88, output_12_9, output_11_88;
mixer gate_output_11_88(.a(output_12_88), .b(output_12_9), .y(output_11_88));
wire output_13_88, output_13_9, output_12_88;
mixer gate_output_12_88(.a(output_13_88), .b(output_13_9), .y(output_12_88));
wire output_14_88, output_14_9, output_13_88;
mixer gate_output_13_88(.a(output_14_88), .b(output_14_9), .y(output_13_88));
wire output_15_88, output_15_9, output_14_88;
mixer gate_output_14_88(.a(output_15_88), .b(output_15_9), .y(output_14_88));
wire output_16_88, output_16_9, output_15_88;
mixer gate_output_15_88(.a(output_16_88), .b(output_16_9), .y(output_15_88));
wire output_1_89, output_1_10, output_0_89;
mixer gate_output_0_89(.a(output_1_89), .b(output_1_10), .y(output_0_89));
wire output_2_89, output_2_10, output_1_89;
mixer gate_output_1_89(.a(output_2_89), .b(output_2_10), .y(output_1_89));
wire output_3_89, output_3_10, output_2_89;
mixer gate_output_2_89(.a(output_3_89), .b(output_3_10), .y(output_2_89));
wire output_4_89, output_4_10, output_3_89;
mixer gate_output_3_89(.a(output_4_89), .b(output_4_10), .y(output_3_89));
wire output_5_89, output_5_10, output_4_89;
mixer gate_output_4_89(.a(output_5_89), .b(output_5_10), .y(output_4_89));
wire output_6_89, output_6_10, output_5_89;
mixer gate_output_5_89(.a(output_6_89), .b(output_6_10), .y(output_5_89));
wire output_7_89, output_7_10, output_6_89;
mixer gate_output_6_89(.a(output_7_89), .b(output_7_10), .y(output_6_89));
wire output_8_89, output_8_10, output_7_89;
mixer gate_output_7_89(.a(output_8_89), .b(output_8_10), .y(output_7_89));
wire output_9_89, output_9_10, output_8_89;
mixer gate_output_8_89(.a(output_9_89), .b(output_9_10), .y(output_8_89));
wire output_10_89, output_10_10, output_9_89;
mixer gate_output_9_89(.a(output_10_89), .b(output_10_10), .y(output_9_89));
wire output_11_89, output_11_10, output_10_89;
mixer gate_output_10_89(.a(output_11_89), .b(output_11_10), .y(output_10_89));
wire output_12_89, output_12_10, output_11_89;
mixer gate_output_11_89(.a(output_12_89), .b(output_12_10), .y(output_11_89));
wire output_13_89, output_13_10, output_12_89;
mixer gate_output_12_89(.a(output_13_89), .b(output_13_10), .y(output_12_89));
wire output_14_89, output_14_10, output_13_89;
mixer gate_output_13_89(.a(output_14_89), .b(output_14_10), .y(output_13_89));
wire output_15_89, output_15_10, output_14_89;
mixer gate_output_14_89(.a(output_15_89), .b(output_15_10), .y(output_14_89));
wire output_16_89, output_16_10, output_15_89;
mixer gate_output_15_89(.a(output_16_89), .b(output_16_10), .y(output_15_89));
wire output_1_90, output_1_11, output_0_90;
mixer gate_output_0_90(.a(output_1_90), .b(output_1_11), .y(output_0_90));
wire output_2_90, output_2_11, output_1_90;
mixer gate_output_1_90(.a(output_2_90), .b(output_2_11), .y(output_1_90));
wire output_3_90, output_3_11, output_2_90;
mixer gate_output_2_90(.a(output_3_90), .b(output_3_11), .y(output_2_90));
wire output_4_90, output_4_11, output_3_90;
mixer gate_output_3_90(.a(output_4_90), .b(output_4_11), .y(output_3_90));
wire output_5_90, output_5_11, output_4_90;
mixer gate_output_4_90(.a(output_5_90), .b(output_5_11), .y(output_4_90));
wire output_6_90, output_6_11, output_5_90;
mixer gate_output_5_90(.a(output_6_90), .b(output_6_11), .y(output_5_90));
wire output_7_90, output_7_11, output_6_90;
mixer gate_output_6_90(.a(output_7_90), .b(output_7_11), .y(output_6_90));
wire output_8_90, output_8_11, output_7_90;
mixer gate_output_7_90(.a(output_8_90), .b(output_8_11), .y(output_7_90));
wire output_9_90, output_9_11, output_8_90;
mixer gate_output_8_90(.a(output_9_90), .b(output_9_11), .y(output_8_90));
wire output_10_90, output_10_11, output_9_90;
mixer gate_output_9_90(.a(output_10_90), .b(output_10_11), .y(output_9_90));
wire output_11_90, output_11_11, output_10_90;
mixer gate_output_10_90(.a(output_11_90), .b(output_11_11), .y(output_10_90));
wire output_12_90, output_12_11, output_11_90;
mixer gate_output_11_90(.a(output_12_90), .b(output_12_11), .y(output_11_90));
wire output_13_90, output_13_11, output_12_90;
mixer gate_output_12_90(.a(output_13_90), .b(output_13_11), .y(output_12_90));
wire output_14_90, output_14_11, output_13_90;
mixer gate_output_13_90(.a(output_14_90), .b(output_14_11), .y(output_13_90));
wire output_15_90, output_15_11, output_14_90;
mixer gate_output_14_90(.a(output_15_90), .b(output_15_11), .y(output_14_90));
wire output_16_90, output_16_11, output_15_90;
mixer gate_output_15_90(.a(output_16_90), .b(output_16_11), .y(output_15_90));
wire output_1_91, output_1_12, output_0_91;
mixer gate_output_0_91(.a(output_1_91), .b(output_1_12), .y(output_0_91));
wire output_2_91, output_2_12, output_1_91;
mixer gate_output_1_91(.a(output_2_91), .b(output_2_12), .y(output_1_91));
wire output_3_91, output_3_12, output_2_91;
mixer gate_output_2_91(.a(output_3_91), .b(output_3_12), .y(output_2_91));
wire output_4_91, output_4_12, output_3_91;
mixer gate_output_3_91(.a(output_4_91), .b(output_4_12), .y(output_3_91));
wire output_5_91, output_5_12, output_4_91;
mixer gate_output_4_91(.a(output_5_91), .b(output_5_12), .y(output_4_91));
wire output_6_91, output_6_12, output_5_91;
mixer gate_output_5_91(.a(output_6_91), .b(output_6_12), .y(output_5_91));
wire output_7_91, output_7_12, output_6_91;
mixer gate_output_6_91(.a(output_7_91), .b(output_7_12), .y(output_6_91));
wire output_8_91, output_8_12, output_7_91;
mixer gate_output_7_91(.a(output_8_91), .b(output_8_12), .y(output_7_91));
wire output_9_91, output_9_12, output_8_91;
mixer gate_output_8_91(.a(output_9_91), .b(output_9_12), .y(output_8_91));
wire output_10_91, output_10_12, output_9_91;
mixer gate_output_9_91(.a(output_10_91), .b(output_10_12), .y(output_9_91));
wire output_11_91, output_11_12, output_10_91;
mixer gate_output_10_91(.a(output_11_91), .b(output_11_12), .y(output_10_91));
wire output_12_91, output_12_12, output_11_91;
mixer gate_output_11_91(.a(output_12_91), .b(output_12_12), .y(output_11_91));
wire output_13_91, output_13_12, output_12_91;
mixer gate_output_12_91(.a(output_13_91), .b(output_13_12), .y(output_12_91));
wire output_14_91, output_14_12, output_13_91;
mixer gate_output_13_91(.a(output_14_91), .b(output_14_12), .y(output_13_91));
wire output_15_91, output_15_12, output_14_91;
mixer gate_output_14_91(.a(output_15_91), .b(output_15_12), .y(output_14_91));
wire output_16_91, output_16_12, output_15_91;
mixer gate_output_15_91(.a(output_16_91), .b(output_16_12), .y(output_15_91));
wire output_1_92, output_1_13, output_0_92;
mixer gate_output_0_92(.a(output_1_92), .b(output_1_13), .y(output_0_92));
wire output_2_92, output_2_13, output_1_92;
mixer gate_output_1_92(.a(output_2_92), .b(output_2_13), .y(output_1_92));
wire output_3_92, output_3_13, output_2_92;
mixer gate_output_2_92(.a(output_3_92), .b(output_3_13), .y(output_2_92));
wire output_4_92, output_4_13, output_3_92;
mixer gate_output_3_92(.a(output_4_92), .b(output_4_13), .y(output_3_92));
wire output_5_92, output_5_13, output_4_92;
mixer gate_output_4_92(.a(output_5_92), .b(output_5_13), .y(output_4_92));
wire output_6_92, output_6_13, output_5_92;
mixer gate_output_5_92(.a(output_6_92), .b(output_6_13), .y(output_5_92));
wire output_7_92, output_7_13, output_6_92;
mixer gate_output_6_92(.a(output_7_92), .b(output_7_13), .y(output_6_92));
wire output_8_92, output_8_13, output_7_92;
mixer gate_output_7_92(.a(output_8_92), .b(output_8_13), .y(output_7_92));
wire output_9_92, output_9_13, output_8_92;
mixer gate_output_8_92(.a(output_9_92), .b(output_9_13), .y(output_8_92));
wire output_10_92, output_10_13, output_9_92;
mixer gate_output_9_92(.a(output_10_92), .b(output_10_13), .y(output_9_92));
wire output_11_92, output_11_13, output_10_92;
mixer gate_output_10_92(.a(output_11_92), .b(output_11_13), .y(output_10_92));
wire output_12_92, output_12_13, output_11_92;
mixer gate_output_11_92(.a(output_12_92), .b(output_12_13), .y(output_11_92));
wire output_13_92, output_13_13, output_12_92;
mixer gate_output_12_92(.a(output_13_92), .b(output_13_13), .y(output_12_92));
wire output_14_92, output_14_13, output_13_92;
mixer gate_output_13_92(.a(output_14_92), .b(output_14_13), .y(output_13_92));
wire output_15_92, output_15_13, output_14_92;
mixer gate_output_14_92(.a(output_15_92), .b(output_15_13), .y(output_14_92));
wire output_16_92, output_16_13, output_15_92;
mixer gate_output_15_92(.a(output_16_92), .b(output_16_13), .y(output_15_92));
wire output_1_93, output_1_14, output_0_93;
mixer gate_output_0_93(.a(output_1_93), .b(output_1_14), .y(output_0_93));
wire output_2_93, output_2_14, output_1_93;
mixer gate_output_1_93(.a(output_2_93), .b(output_2_14), .y(output_1_93));
wire output_3_93, output_3_14, output_2_93;
mixer gate_output_2_93(.a(output_3_93), .b(output_3_14), .y(output_2_93));
wire output_4_93, output_4_14, output_3_93;
mixer gate_output_3_93(.a(output_4_93), .b(output_4_14), .y(output_3_93));
wire output_5_93, output_5_14, output_4_93;
mixer gate_output_4_93(.a(output_5_93), .b(output_5_14), .y(output_4_93));
wire output_6_93, output_6_14, output_5_93;
mixer gate_output_5_93(.a(output_6_93), .b(output_6_14), .y(output_5_93));
wire output_7_93, output_7_14, output_6_93;
mixer gate_output_6_93(.a(output_7_93), .b(output_7_14), .y(output_6_93));
wire output_8_93, output_8_14, output_7_93;
mixer gate_output_7_93(.a(output_8_93), .b(output_8_14), .y(output_7_93));
wire output_9_93, output_9_14, output_8_93;
mixer gate_output_8_93(.a(output_9_93), .b(output_9_14), .y(output_8_93));
wire output_10_93, output_10_14, output_9_93;
mixer gate_output_9_93(.a(output_10_93), .b(output_10_14), .y(output_9_93));
wire output_11_93, output_11_14, output_10_93;
mixer gate_output_10_93(.a(output_11_93), .b(output_11_14), .y(output_10_93));
wire output_12_93, output_12_14, output_11_93;
mixer gate_output_11_93(.a(output_12_93), .b(output_12_14), .y(output_11_93));
wire output_13_93, output_13_14, output_12_93;
mixer gate_output_12_93(.a(output_13_93), .b(output_13_14), .y(output_12_93));
wire output_14_93, output_14_14, output_13_93;
mixer gate_output_13_93(.a(output_14_93), .b(output_14_14), .y(output_13_93));
wire output_15_93, output_15_14, output_14_93;
mixer gate_output_14_93(.a(output_15_93), .b(output_15_14), .y(output_14_93));
wire output_16_93, output_16_14, output_15_93;
mixer gate_output_15_93(.a(output_16_93), .b(output_16_14), .y(output_15_93));
wire output_1_94, output_1_15, output_0_94;
mixer gate_output_0_94(.a(output_1_94), .b(output_1_15), .y(output_0_94));
wire output_2_94, output_2_15, output_1_94;
mixer gate_output_1_94(.a(output_2_94), .b(output_2_15), .y(output_1_94));
wire output_3_94, output_3_15, output_2_94;
mixer gate_output_2_94(.a(output_3_94), .b(output_3_15), .y(output_2_94));
wire output_4_94, output_4_15, output_3_94;
mixer gate_output_3_94(.a(output_4_94), .b(output_4_15), .y(output_3_94));
wire output_5_94, output_5_15, output_4_94;
mixer gate_output_4_94(.a(output_5_94), .b(output_5_15), .y(output_4_94));
wire output_6_94, output_6_15, output_5_94;
mixer gate_output_5_94(.a(output_6_94), .b(output_6_15), .y(output_5_94));
wire output_7_94, output_7_15, output_6_94;
mixer gate_output_6_94(.a(output_7_94), .b(output_7_15), .y(output_6_94));
wire output_8_94, output_8_15, output_7_94;
mixer gate_output_7_94(.a(output_8_94), .b(output_8_15), .y(output_7_94));
wire output_9_94, output_9_15, output_8_94;
mixer gate_output_8_94(.a(output_9_94), .b(output_9_15), .y(output_8_94));
wire output_10_94, output_10_15, output_9_94;
mixer gate_output_9_94(.a(output_10_94), .b(output_10_15), .y(output_9_94));
wire output_11_94, output_11_15, output_10_94;
mixer gate_output_10_94(.a(output_11_94), .b(output_11_15), .y(output_10_94));
wire output_12_94, output_12_15, output_11_94;
mixer gate_output_11_94(.a(output_12_94), .b(output_12_15), .y(output_11_94));
wire output_13_94, output_13_15, output_12_94;
mixer gate_output_12_94(.a(output_13_94), .b(output_13_15), .y(output_12_94));
wire output_14_94, output_14_15, output_13_94;
mixer gate_output_13_94(.a(output_14_94), .b(output_14_15), .y(output_13_94));
wire output_15_94, output_15_15, output_14_94;
mixer gate_output_14_94(.a(output_15_94), .b(output_15_15), .y(output_14_94));
wire output_16_94, output_16_15, output_15_94;
mixer gate_output_15_94(.a(output_16_94), .b(output_16_15), .y(output_15_94));
wire output_1_95, output_1_0, output_0_95;
mixer gate_output_0_95(.a(output_1_95), .b(output_1_0), .y(output_0_95));
wire output_2_95, output_2_0, output_1_95;
mixer gate_output_1_95(.a(output_2_95), .b(output_2_0), .y(output_1_95));
wire output_3_95, output_3_0, output_2_95;
mixer gate_output_2_95(.a(output_3_95), .b(output_3_0), .y(output_2_95));
wire output_4_95, output_4_0, output_3_95;
mixer gate_output_3_95(.a(output_4_95), .b(output_4_0), .y(output_3_95));
wire output_5_95, output_5_0, output_4_95;
mixer gate_output_4_95(.a(output_5_95), .b(output_5_0), .y(output_4_95));
wire output_6_95, output_6_0, output_5_95;
mixer gate_output_5_95(.a(output_6_95), .b(output_6_0), .y(output_5_95));
wire output_7_95, output_7_0, output_6_95;
mixer gate_output_6_95(.a(output_7_95), .b(output_7_0), .y(output_6_95));
wire output_8_95, output_8_0, output_7_95;
mixer gate_output_7_95(.a(output_8_95), .b(output_8_0), .y(output_7_95));
wire output_9_95, output_9_0, output_8_95;
mixer gate_output_8_95(.a(output_9_95), .b(output_9_0), .y(output_8_95));
wire output_10_95, output_10_0, output_9_95;
mixer gate_output_9_95(.a(output_10_95), .b(output_10_0), .y(output_9_95));
wire output_11_95, output_11_0, output_10_95;
mixer gate_output_10_95(.a(output_11_95), .b(output_11_0), .y(output_10_95));
wire output_12_95, output_12_0, output_11_95;
mixer gate_output_11_95(.a(output_12_95), .b(output_12_0), .y(output_11_95));
wire output_13_95, output_13_0, output_12_95;
mixer gate_output_12_95(.a(output_13_95), .b(output_13_0), .y(output_12_95));
wire output_14_95, output_14_0, output_13_95;
mixer gate_output_13_95(.a(output_14_95), .b(output_14_0), .y(output_13_95));
wire output_15_95, output_15_0, output_14_95;
mixer gate_output_14_95(.a(output_15_95), .b(output_15_0), .y(output_14_95));
wire output_16_95, output_16_0, output_15_95;
mixer gate_output_15_95(.a(output_16_95), .b(output_16_0), .y(output_15_95));
assign output_0 = output_0_0;
wire output_0_96;
assign output_0_96 = input_0;
assign output_1 = output_1_0;
wire output_1_96;
assign output_1_96 = input_1;
assign output_2 = output_2_0;
wire output_2_96;
assign output_2_96 = input_2;
assign output_3 = output_3_0;
wire output_3_96;
assign output_3_96 = input_3;
assign output_4 = output_4_0;
wire output_4_96;
assign output_4_96 = input_4;
assign output_5 = output_5_0;
wire output_5_96;
assign output_5_96 = input_5;
assign output_6 = output_6_0;
wire output_6_96;
assign output_6_96 = input_6;
assign output_7 = output_7_0;
wire output_7_96;
assign output_7_96 = input_7;
assign output_8 = output_8_0;
wire output_8_96;
assign output_8_96 = input_8;
assign output_9 = output_9_0;
wire output_9_96;
assign output_9_96 = input_9;
assign output_10 = output_10_0;
wire output_10_96;
assign output_10_96 = input_10;
assign output_11 = output_11_0;
wire output_11_96;
assign output_11_96 = input_11;
assign output_12 = output_12_0;
wire output_12_96;
assign output_12_96 = input_12;
assign output_13 = output_13_0;
wire output_13_96;
assign output_13_96 = input_13;
assign output_14 = output_14_0;
wire output_14_96;
assign output_14_96 = input_14;
assign output_15 = output_15_0;
wire output_15_96;
assign output_15_96 = input_15;
endmodule
