  module protein_assay(input DsS,
                       DsB1, DsB2, DsB3, DsB4, DsB5, DsB6, DsB7, DsB8, DsB9, DsB10, DsB11, DsB12, DsB13, DsB14, DsB15, DsB16, DsB17, DsB18, DsB19, DsB20, DsB21, DsB22, DsB23, DsB24, DsB25, DsB26, DsB27, DsB28, DsB29, DsB30, DsB31, DsB32, DsB33, DsB34, DsB35, DsB36, DsB37, DsB38, DsB39,
                       output Opt1, Opt2, Opt3, Opt4, Opt5, Opt6, Opt7, Opt8);
